module multiplier_256bits_version11(product, A, B);

    output [511:0] product;
    input [255:0] A, B;

    wire [255:0] pp0;
    wire [255:0] pp1;
    wire [255:0] pp2;
    wire [255:0] pp3;
    wire [255:0] pp4;
    wire [255:0] pp5;
    wire [255:0] pp6;
    wire [255:0] pp7;
    wire [255:0] pp8;
    wire [255:0] pp9;
    wire [255:0] pp10;
    wire [255:0] pp11;
    wire [255:0] pp12;
    wire [255:0] pp13;
    wire [255:0] pp14;
    wire [255:0] pp15;
    wire [255:0] pp16;
    wire [255:0] pp17;
    wire [255:0] pp18;
    wire [255:0] pp19;
    wire [255:0] pp20;
    wire [255:0] pp21;
    wire [255:0] pp22;
    wire [255:0] pp23;
    wire [255:0] pp24;
    wire [255:0] pp25;
    wire [255:0] pp26;
    wire [255:0] pp27;
    wire [255:0] pp28;
    wire [255:0] pp29;
    wire [255:0] pp30;
    wire [255:0] pp31;
    wire [255:0] pp32;
    wire [255:0] pp33;
    wire [255:0] pp34;
    wire [255:0] pp35;
    wire [255:0] pp36;
    wire [255:0] pp37;
    wire [255:0] pp38;
    wire [255:0] pp39;
    wire [255:0] pp40;
    wire [255:0] pp41;
    wire [255:0] pp42;
    wire [255:0] pp43;
    wire [255:0] pp44;
    wire [255:0] pp45;
    wire [255:0] pp46;
    wire [255:0] pp47;
    wire [255:0] pp48;
    wire [255:0] pp49;
    wire [255:0] pp50;
    wire [255:0] pp51;
    wire [255:0] pp52;
    wire [255:0] pp53;
    wire [255:0] pp54;
    wire [255:0] pp55;
    wire [255:0] pp56;
    wire [255:0] pp57;
    wire [255:0] pp58;
    wire [255:0] pp59;
    wire [255:0] pp60;
    wire [255:0] pp61;
    wire [255:0] pp62;
    wire [255:0] pp63;
    wire [255:0] pp64;
    wire [255:0] pp65;
    wire [255:0] pp66;
    wire [255:0] pp67;
    wire [255:0] pp68;
    wire [255:0] pp69;
    wire [255:0] pp70;
    wire [255:0] pp71;
    wire [255:0] pp72;
    wire [255:0] pp73;
    wire [255:0] pp74;
    wire [255:0] pp75;
    wire [255:0] pp76;
    wire [255:0] pp77;
    wire [255:0] pp78;
    wire [255:0] pp79;
    wire [255:0] pp80;
    wire [255:0] pp81;
    wire [255:0] pp82;
    wire [255:0] pp83;
    wire [255:0] pp84;
    wire [255:0] pp85;
    wire [255:0] pp86;
    wire [255:0] pp87;
    wire [255:0] pp88;
    wire [255:0] pp89;
    wire [255:0] pp90;
    wire [255:0] pp91;
    wire [255:0] pp92;
    wire [255:0] pp93;
    wire [255:0] pp94;
    wire [255:0] pp95;
    wire [255:0] pp96;
    wire [255:0] pp97;
    wire [255:0] pp98;
    wire [255:0] pp99;
    wire [255:0] pp100;
    wire [255:0] pp101;
    wire [255:0] pp102;
    wire [255:0] pp103;
    wire [255:0] pp104;
    wire [255:0] pp105;
    wire [255:0] pp106;
    wire [255:0] pp107;
    wire [255:0] pp108;
    wire [255:0] pp109;
    wire [255:0] pp110;
    wire [255:0] pp111;
    wire [255:0] pp112;
    wire [255:0] pp113;
    wire [255:0] pp114;
    wire [255:0] pp115;
    wire [255:0] pp116;
    wire [255:0] pp117;
    wire [255:0] pp118;
    wire [255:0] pp119;
    wire [255:0] pp120;
    wire [255:0] pp121;
    wire [255:0] pp122;
    wire [255:0] pp123;
    wire [255:0] pp124;
    wire [255:0] pp125;
    wire [255:0] pp126;
    wire [255:0] pp127;
    wire [255:0] pp128;
    wire [255:0] pp129;
    wire [255:0] pp130;
    wire [255:0] pp131;
    wire [255:0] pp132;
    wire [255:0] pp133;
    wire [255:0] pp134;
    wire [255:0] pp135;
    wire [255:0] pp136;
    wire [255:0] pp137;
    wire [255:0] pp138;
    wire [255:0] pp139;
    wire [255:0] pp140;
    wire [255:0] pp141;
    wire [255:0] pp142;
    wire [255:0] pp143;
    wire [255:0] pp144;
    wire [255:0] pp145;
    wire [255:0] pp146;
    wire [255:0] pp147;
    wire [255:0] pp148;
    wire [255:0] pp149;
    wire [255:0] pp150;
    wire [255:0] pp151;
    wire [255:0] pp152;
    wire [255:0] pp153;
    wire [255:0] pp154;
    wire [255:0] pp155;
    wire [255:0] pp156;
    wire [255:0] pp157;
    wire [255:0] pp158;
    wire [255:0] pp159;
    wire [255:0] pp160;
    wire [255:0] pp161;
    wire [255:0] pp162;
    wire [255:0] pp163;
    wire [255:0] pp164;
    wire [255:0] pp165;
    wire [255:0] pp166;
    wire [255:0] pp167;
    wire [255:0] pp168;
    wire [255:0] pp169;
    wire [255:0] pp170;
    wire [255:0] pp171;
    wire [255:0] pp172;
    wire [255:0] pp173;
    wire [255:0] pp174;
    wire [255:0] pp175;
    wire [255:0] pp176;
    wire [255:0] pp177;
    wire [255:0] pp178;
    wire [255:0] pp179;
    wire [255:0] pp180;
    wire [255:0] pp181;
    wire [255:0] pp182;
    wire [255:0] pp183;
    wire [255:0] pp184;
    wire [255:0] pp185;
    wire [255:0] pp186;
    wire [255:0] pp187;
    wire [255:0] pp188;
    wire [255:0] pp189;
    wire [255:0] pp190;
    wire [255:0] pp191;
    wire [255:0] pp192;
    wire [255:0] pp193;
    wire [255:0] pp194;
    wire [255:0] pp195;
    wire [255:0] pp196;
    wire [255:0] pp197;
    wire [255:0] pp198;
    wire [255:0] pp199;
    wire [255:0] pp200;
    wire [255:0] pp201;
    wire [255:0] pp202;
    wire [255:0] pp203;
    wire [255:0] pp204;
    wire [255:0] pp205;
    wire [255:0] pp206;
    wire [255:0] pp207;
    wire [255:0] pp208;
    wire [255:0] pp209;
    wire [255:0] pp210;
    wire [255:0] pp211;
    wire [255:0] pp212;
    wire [255:0] pp213;
    wire [255:0] pp214;
    wire [255:0] pp215;
    wire [255:0] pp216;
    wire [255:0] pp217;
    wire [255:0] pp218;
    wire [255:0] pp219;
    wire [255:0] pp220;
    wire [255:0] pp221;
    wire [255:0] pp222;
    wire [255:0] pp223;
    wire [255:0] pp224;
    wire [255:0] pp225;
    wire [255:0] pp226;
    wire [255:0] pp227;
    wire [255:0] pp228;
    wire [255:0] pp229;
    wire [255:0] pp230;
    wire [255:0] pp231;
    wire [255:0] pp232;
    wire [255:0] pp233;
    wire [255:0] pp234;
    wire [255:0] pp235;
    wire [255:0] pp236;
    wire [255:0] pp237;
    wire [255:0] pp238;
    wire [255:0] pp239;
    wire [255:0] pp240;
    wire [255:0] pp241;
    wire [255:0] pp242;
    wire [255:0] pp243;
    wire [255:0] pp244;
    wire [255:0] pp245;
    wire [255:0] pp246;
    wire [255:0] pp247;
    wire [255:0] pp248;
    wire [255:0] pp249;
    wire [255:0] pp250;
    wire [255:0] pp251;
    wire [255:0] pp252;
    wire [255:0] pp253;
    wire [255:0] pp254;
    wire [255:0] pp255;


    assign pp0 = A[0] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp64 = A[64] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp65 = A[65] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp66 = A[66] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp67 = A[67] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp68 = A[68] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp69 = A[69] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp70 = A[70] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp71 = A[71] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp72 = A[72] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp73 = A[73] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp74 = A[74] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp75 = A[75] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp76 = A[76] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp77 = A[77] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp78 = A[78] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp79 = A[79] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp80 = A[80] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp81 = A[81] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp82 = A[82] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp83 = A[83] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp84 = A[84] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp85 = A[85] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp86 = A[86] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp87 = A[87] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp88 = A[88] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp89 = A[89] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp90 = A[90] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp91 = A[91] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp92 = A[92] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp93 = A[93] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp94 = A[94] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp95 = A[95] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp96 = A[96] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp97 = A[97] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp98 = A[98] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp99 = A[99] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp100 = A[100] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp101 = A[101] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp102 = A[102] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp103 = A[103] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp104 = A[104] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp105 = A[105] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp106 = A[106] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp107 = A[107] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp108 = A[108] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp109 = A[109] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp110 = A[110] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp111 = A[111] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp112 = A[112] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp113 = A[113] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp114 = A[114] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp115 = A[115] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp116 = A[116] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp117 = A[117] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp118 = A[118] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp119 = A[119] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp120 = A[120] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp121 = A[121] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp122 = A[122] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp123 = A[123] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp124 = A[124] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp125 = A[125] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp126 = A[126] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp127 = A[127] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp128 = A[128] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp129 = A[129] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp130 = A[130] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp131 = A[131] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp132 = A[132] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp133 = A[133] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp134 = A[134] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp135 = A[135] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp136 = A[136] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp137 = A[137] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp138 = A[138] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp139 = A[139] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp140 = A[140] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp141 = A[141] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp142 = A[142] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp143 = A[143] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp144 = A[144] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp145 = A[145] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp146 = A[146] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp147 = A[147] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp148 = A[148] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp149 = A[149] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp150 = A[150] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp151 = A[151] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp152 = A[152] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp153 = A[153] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp154 = A[154] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp155 = A[155] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp156 = A[156] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp157 = A[157] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp158 = A[158] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp159 = A[159] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp160 = A[160] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp161 = A[161] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp162 = A[162] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp163 = A[163] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp164 = A[164] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp165 = A[165] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp166 = A[166] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp167 = A[167] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp168 = A[168] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp169 = A[169] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp170 = A[170] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp171 = A[171] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp172 = A[172] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp173 = A[173] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp174 = A[174] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp175 = A[175] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp176 = A[176] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp177 = A[177] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp178 = A[178] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp179 = A[179] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp180 = A[180] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp181 = A[181] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp182 = A[182] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp183 = A[183] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp184 = A[184] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp185 = A[185] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp186 = A[186] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp187 = A[187] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp188 = A[188] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp189 = A[189] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp190 = A[190] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp191 = A[191] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp192 = A[192] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp193 = A[193] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp194 = A[194] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp195 = A[195] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp196 = A[196] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp197 = A[197] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp198 = A[198] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp199 = A[199] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp200 = A[200] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp201 = A[201] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp202 = A[202] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp203 = A[203] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp204 = A[204] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp205 = A[205] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp206 = A[206] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp207 = A[207] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp208 = A[208] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp209 = A[209] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp210 = A[210] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp211 = A[211] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp212 = A[212] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp213 = A[213] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp214 = A[214] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp215 = A[215] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp216 = A[216] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp217 = A[217] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp218 = A[218] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp219 = A[219] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp220 = A[220] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp221 = A[221] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp222 = A[222] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp223 = A[223] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp224 = A[224] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp225 = A[225] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp226 = A[226] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp227 = A[227] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp228 = A[228] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp229 = A[229] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp230 = A[230] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp231 = A[231] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp232 = A[232] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp233 = A[233] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp234 = A[234] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp235 = A[235] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp236 = A[236] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp237 = A[237] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp238 = A[238] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp239 = A[239] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp240 = A[240] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp241 = A[241] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp242 = A[242] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp243 = A[243] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp244 = A[244] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp245 = A[245] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp246 = A[246] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp247 = A[247] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp248 = A[248] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp249 = A[249] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp250 = A[250] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp251 = A[251] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp252 = A[252] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp253 = A[253] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp254 = A[254] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp255 = A[255] ? B: 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[255:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp10[118],pp10[119],pp10[120],pp10[121],pp10[122],pp10[123],pp10[124],pp10[125],pp10[126],pp10[127],pp10[128],pp10[129],pp10[130],pp10[131],pp10[132],pp10[133],pp10[134],pp10[135],pp10[136],pp10[137],pp10[138],pp10[139],pp10[140],pp10[141],pp10[142],pp10[143],pp10[144],pp10[145],pp10[146],pp10[147],pp10[148],pp10[149],pp10[150],pp10[151],pp10[152],pp10[153],pp10[154],pp10[155],pp10[156],pp10[157],pp10[158],pp10[159],pp10[160],pp10[161],pp10[162],pp10[163],pp10[164],pp10[165],pp10[166],pp10[167],pp10[168],pp10[169],pp10[170],pp10[171],pp10[172],pp10[173],pp10[174],pp10[175],pp10[176],pp10[177],pp10[178],pp10[179],pp10[180],pp10[181],pp10[182],pp10[183],pp10[184],pp10[185],pp10[186],pp10[187],pp10[188],pp10[189],pp100[100],pp100[101],pp100[102],pp100[103],pp100[104],pp100[105],pp100[106],pp100[107],pp100[108],pp100[109],pp100[110],pp100[111],pp100[112],pp100[113],pp100[114],pp100[115],pp100[116],pp100[117],pp100[118],pp100[119],pp100[120],pp100[121],pp100[122],pp100[123],pp100[124],pp100[125],pp100[126],pp100[127],pp100[128],pp100[129],pp100[130],pp100[131],pp100[132],pp100[133],pp100[134],pp100[135],pp100[136],pp100[137],pp100[138],pp100[139],pp100[140],pp100[141],pp100[142],pp100[143],pp100[144],pp100[145],pp100[146],pp100[147],pp100[148],pp100[149],pp100[150],pp100[151],pp100[152],pp100[153],pp100[154],pp100[155],pp100[156],pp100[157],pp100[158],pp100[159],pp100[160],pp100[161],pp100[162],pp100[163],pp100[164],pp100[165],pp100[166],pp100[167],pp100[168],pp100[169],pp100[170],pp100[171],pp100[172],pp100[173],pp100[174],pp100[175],pp100[176],pp100[177],pp100[178],pp100[179],pp100[180],pp100[181],pp100[182],pp100[183],pp100[184],pp100[185],pp100[186],pp100[187],pp100[188],pp100[189],pp100[190],pp100[191],pp100[192],pp100[193],pp100[194],pp100[195],pp100[196],pp100[197],pp100[198],pp100[199],pp100[200],pp100[201],pp100[202],pp100[203],pp100[204],pp100[205],pp100[206],pp100[207],pp100[208],pp100[209],pp100[210],pp100[211],pp100[212],pp100[213],pp100[214],pp100[215],pp100[216],pp100[217],pp100[218],pp100[219],pp100[220],pp100[221],pp100[222],pp100[223],pp100[224],pp100[225],pp100[226],pp100[227],pp100[228],pp100[229],pp100[230],pp100[231],pp100[232],pp100[233],pp100[234],pp100[235],pp100[236],pp100[237],pp100[238],pp100[239],pp100[240],pp100[241],pp100[242],pp100[243],pp100[244],pp100[245],pp100[246],pp100[247],pp100[248],pp100[249],pp100[250],pp100[251],pp100[252],pp100[253],pp100[254],pp100[255],pp101[255],pp102[255],pp103[255],pp104[255],pp105[255],pp106[255],pp107[255],pp108[255],pp109[255],pp110[255],pp111[255],pp112[255],pp113[255],pp114[255],pp115[255],pp116[255],pp117[255],pp118[255],pp119[255],pp120[255],pp121[255],pp122[255],pp123[255],pp124[255],pp125[255],pp126[255],pp127[255],pp128[255]};
    assign in1_2 = {pp11[117],pp11[118],pp11[119],pp11[120],pp11[121],pp11[122],pp11[123],pp11[124],pp11[125],pp11[126],pp11[127],pp11[128],pp11[129],pp11[130],pp11[131],pp11[132],pp11[133],pp11[134],pp11[135],pp11[136],pp11[137],pp11[138],pp11[139],pp11[140],pp11[141],pp11[142],pp11[143],pp11[144],pp11[145],pp11[146],pp11[147],pp11[148],pp11[149],pp11[150],pp11[151],pp11[152],pp11[153],pp11[154],pp11[155],pp11[156],pp11[157],pp11[158],pp11[159],pp11[160],pp11[161],pp11[162],pp11[163],pp11[164],pp11[165],pp11[166],pp11[167],pp11[168],pp11[169],pp11[170],pp11[171],pp11[172],pp11[173],pp11[174],pp11[175],pp11[176],pp11[177],pp11[178],pp11[179],pp11[180],pp11[181],pp11[182],pp11[183],pp11[184],pp11[185],pp11[186],pp11[187],pp11[188],pp10[190],pp101[100],pp101[101],pp101[102],pp101[103],pp101[104],pp101[105],pp101[106],pp101[107],pp101[108],pp101[109],pp101[110],pp101[111],pp101[112],pp101[113],pp101[114],pp101[115],pp101[116],pp101[117],pp101[118],pp101[119],pp101[120],pp101[121],pp101[122],pp101[123],pp101[124],pp101[125],pp101[126],pp101[127],pp101[128],pp101[129],pp101[130],pp101[131],pp101[132],pp101[133],pp101[134],pp101[135],pp101[136],pp101[137],pp101[138],pp101[139],pp101[140],pp101[141],pp101[142],pp101[143],pp101[144],pp101[145],pp101[146],pp101[147],pp101[148],pp101[149],pp101[150],pp101[151],pp101[152],pp101[153],pp101[154],pp101[155],pp101[156],pp101[157],pp101[158],pp101[159],pp101[160],pp101[161],pp101[162],pp101[163],pp101[164],pp101[165],pp101[166],pp101[167],pp101[168],pp101[169],pp101[170],pp101[171],pp101[172],pp101[173],pp101[174],pp101[175],pp101[176],pp101[177],pp101[178],pp101[179],pp101[180],pp101[181],pp101[182],pp101[183],pp101[184],pp101[185],pp101[186],pp101[187],pp101[188],pp101[189],pp101[190],pp101[191],pp101[192],pp101[193],pp101[194],pp101[195],pp101[196],pp101[197],pp101[198],pp101[199],pp101[200],pp101[201],pp101[202],pp101[203],pp101[204],pp101[205],pp101[206],pp101[207],pp101[208],pp101[209],pp101[210],pp101[211],pp101[212],pp101[213],pp101[214],pp101[215],pp101[216],pp101[217],pp101[218],pp101[219],pp101[220],pp101[221],pp101[222],pp101[223],pp101[224],pp101[225],pp101[226],pp101[227],pp101[228],pp101[229],pp101[230],pp101[231],pp101[232],pp101[233],pp101[234],pp101[235],pp101[236],pp101[237],pp101[238],pp101[239],pp101[240],pp101[241],pp101[242],pp101[243],pp101[244],pp101[245],pp101[246],pp101[247],pp101[248],pp101[249],pp101[250],pp101[251],pp101[252],pp101[253],pp101[254],pp102[254],pp103[254],pp104[254],pp105[254],pp106[254],pp107[254],pp108[254],pp109[254],pp110[254],pp111[254],pp112[254],pp113[254],pp114[254],pp115[254],pp116[254],pp117[254],pp118[254],pp119[254],pp120[254],pp121[254],pp122[254],pp123[254],pp124[254],pp125[254],pp126[254],pp127[254],pp128[254],pp129[254]};
    CLA_256 KS_1(s1, c1, in1_1, in1_2);
    wire[253:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp12[117],pp12[118],pp12[119],pp12[120],pp12[121],pp12[122],pp12[123],pp12[124],pp12[125],pp12[126],pp12[127],pp12[128],pp12[129],pp12[130],pp12[131],pp12[132],pp12[133],pp12[134],pp12[135],pp12[136],pp12[137],pp12[138],pp12[139],pp12[140],pp12[141],pp12[142],pp12[143],pp12[144],pp12[145],pp12[146],pp12[147],pp12[148],pp12[149],pp12[150],pp12[151],pp12[152],pp12[153],pp12[154],pp12[155],pp12[156],pp12[157],pp12[158],pp12[159],pp12[160],pp12[161],pp12[162],pp12[163],pp12[164],pp12[165],pp12[166],pp12[167],pp12[168],pp12[169],pp12[170],pp12[171],pp12[172],pp12[173],pp12[174],pp12[175],pp12[176],pp12[177],pp12[178],pp12[179],pp12[180],pp12[181],pp12[182],pp12[183],pp12[184],pp12[185],pp12[186],pp12[187],pp11[189],pp10[191],pp102[100],pp102[101],pp102[102],pp102[103],pp102[104],pp102[105],pp102[106],pp102[107],pp102[108],pp102[109],pp102[110],pp102[111],pp102[112],pp102[113],pp102[114],pp102[115],pp102[116],pp102[117],pp102[118],pp102[119],pp102[120],pp102[121],pp102[122],pp102[123],pp102[124],pp102[125],pp102[126],pp102[127],pp102[128],pp102[129],pp102[130],pp102[131],pp102[132],pp102[133],pp102[134],pp102[135],pp102[136],pp102[137],pp102[138],pp102[139],pp102[140],pp102[141],pp102[142],pp102[143],pp102[144],pp102[145],pp102[146],pp102[147],pp102[148],pp102[149],pp102[150],pp102[151],pp102[152],pp102[153],pp102[154],pp102[155],pp102[156],pp102[157],pp102[158],pp102[159],pp102[160],pp102[161],pp102[162],pp102[163],pp102[164],pp102[165],pp102[166],pp102[167],pp102[168],pp102[169],pp102[170],pp102[171],pp102[172],pp102[173],pp102[174],pp102[175],pp102[176],pp102[177],pp102[178],pp102[179],pp102[180],pp102[181],pp102[182],pp102[183],pp102[184],pp102[185],pp102[186],pp102[187],pp102[188],pp102[189],pp102[190],pp102[191],pp102[192],pp102[193],pp102[194],pp102[195],pp102[196],pp102[197],pp102[198],pp102[199],pp102[200],pp102[201],pp102[202],pp102[203],pp102[204],pp102[205],pp102[206],pp102[207],pp102[208],pp102[209],pp102[210],pp102[211],pp102[212],pp102[213],pp102[214],pp102[215],pp102[216],pp102[217],pp102[218],pp102[219],pp102[220],pp102[221],pp102[222],pp102[223],pp102[224],pp102[225],pp102[226],pp102[227],pp102[228],pp102[229],pp102[230],pp102[231],pp102[232],pp102[233],pp102[234],pp102[235],pp102[236],pp102[237],pp102[238],pp102[239],pp102[240],pp102[241],pp102[242],pp102[243],pp102[244],pp102[245],pp102[246],pp102[247],pp102[248],pp102[249],pp102[250],pp102[251],pp102[252],pp102[253],pp103[253],pp104[253],pp105[253],pp106[253],pp107[253],pp108[253],pp109[253],pp110[253],pp111[253],pp112[253],pp113[253],pp114[253],pp115[253],pp116[253],pp117[253],pp118[253],pp119[253],pp120[253],pp121[253],pp122[253],pp123[253],pp124[253],pp125[253],pp126[253],pp127[253],pp128[253],pp129[253]};
    assign in2_2 = {pp13[116],pp13[117],pp13[118],pp13[119],pp13[120],pp13[121],pp13[122],pp13[123],pp13[124],pp13[125],pp13[126],pp13[127],pp13[128],pp13[129],pp13[130],pp13[131],pp13[132],pp13[133],pp13[134],pp13[135],pp13[136],pp13[137],pp13[138],pp13[139],pp13[140],pp13[141],pp13[142],pp13[143],pp13[144],pp13[145],pp13[146],pp13[147],pp13[148],pp13[149],pp13[150],pp13[151],pp13[152],pp13[153],pp13[154],pp13[155],pp13[156],pp13[157],pp13[158],pp13[159],pp13[160],pp13[161],pp13[162],pp13[163],pp13[164],pp13[165],pp13[166],pp13[167],pp13[168],pp13[169],pp13[170],pp13[171],pp13[172],pp13[173],pp13[174],pp13[175],pp13[176],pp13[177],pp13[178],pp13[179],pp13[180],pp13[181],pp13[182],pp13[183],pp13[184],pp13[185],pp13[186],pp12[188],pp11[190],pp10[192],pp103[100],pp103[101],pp103[102],pp103[103],pp103[104],pp103[105],pp103[106],pp103[107],pp103[108],pp103[109],pp103[110],pp103[111],pp103[112],pp103[113],pp103[114],pp103[115],pp103[116],pp103[117],pp103[118],pp103[119],pp103[120],pp103[121],pp103[122],pp103[123],pp103[124],pp103[125],pp103[126],pp103[127],pp103[128],pp103[129],pp103[130],pp103[131],pp103[132],pp103[133],pp103[134],pp103[135],pp103[136],pp103[137],pp103[138],pp103[139],pp103[140],pp103[141],pp103[142],pp103[143],pp103[144],pp103[145],pp103[146],pp103[147],pp103[148],pp103[149],pp103[150],pp103[151],pp103[152],pp103[153],pp103[154],pp103[155],pp103[156],pp103[157],pp103[158],pp103[159],pp103[160],pp103[161],pp103[162],pp103[163],pp103[164],pp103[165],pp103[166],pp103[167],pp103[168],pp103[169],pp103[170],pp103[171],pp103[172],pp103[173],pp103[174],pp103[175],pp103[176],pp103[177],pp103[178],pp103[179],pp103[180],pp103[181],pp103[182],pp103[183],pp103[184],pp103[185],pp103[186],pp103[187],pp103[188],pp103[189],pp103[190],pp103[191],pp103[192],pp103[193],pp103[194],pp103[195],pp103[196],pp103[197],pp103[198],pp103[199],pp103[200],pp103[201],pp103[202],pp103[203],pp103[204],pp103[205],pp103[206],pp103[207],pp103[208],pp103[209],pp103[210],pp103[211],pp103[212],pp103[213],pp103[214],pp103[215],pp103[216],pp103[217],pp103[218],pp103[219],pp103[220],pp103[221],pp103[222],pp103[223],pp103[224],pp103[225],pp103[226],pp103[227],pp103[228],pp103[229],pp103[230],pp103[231],pp103[232],pp103[233],pp103[234],pp103[235],pp103[236],pp103[237],pp103[238],pp103[239],pp103[240],pp103[241],pp103[242],pp103[243],pp103[244],pp103[245],pp103[246],pp103[247],pp103[248],pp103[249],pp103[250],pp103[251],pp103[252],pp104[252],pp105[252],pp106[252],pp107[252],pp108[252],pp109[252],pp110[252],pp111[252],pp112[252],pp113[252],pp114[252],pp115[252],pp116[252],pp117[252],pp118[252],pp119[252],pp120[252],pp121[252],pp122[252],pp123[252],pp124[252],pp125[252],pp126[252],pp127[252],pp128[252],pp129[252],pp130[252]};
    CLA_254 KS_2(s2, c2, in2_1, in2_2);
    wire[251:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp14[116],pp14[117],pp14[118],pp14[119],pp14[120],pp14[121],pp14[122],pp14[123],pp14[124],pp14[125],pp14[126],pp14[127],pp14[128],pp14[129],pp14[130],pp14[131],pp14[132],pp14[133],pp14[134],pp14[135],pp14[136],pp14[137],pp14[138],pp14[139],pp14[140],pp14[141],pp14[142],pp14[143],pp14[144],pp14[145],pp14[146],pp14[147],pp14[148],pp14[149],pp14[150],pp14[151],pp14[152],pp14[153],pp14[154],pp14[155],pp14[156],pp14[157],pp14[158],pp14[159],pp14[160],pp14[161],pp14[162],pp14[163],pp14[164],pp14[165],pp14[166],pp14[167],pp14[168],pp14[169],pp14[170],pp14[171],pp14[172],pp14[173],pp14[174],pp14[175],pp14[176],pp14[177],pp14[178],pp14[179],pp14[180],pp14[181],pp14[182],pp14[183],pp14[184],pp14[185],pp13[187],pp12[189],pp11[191],pp10[193],pp104[100],pp104[101],pp104[102],pp104[103],pp104[104],pp104[105],pp104[106],pp104[107],pp104[108],pp104[109],pp104[110],pp104[111],pp104[112],pp104[113],pp104[114],pp104[115],pp104[116],pp104[117],pp104[118],pp104[119],pp104[120],pp104[121],pp104[122],pp104[123],pp104[124],pp104[125],pp104[126],pp104[127],pp104[128],pp104[129],pp104[130],pp104[131],pp104[132],pp104[133],pp104[134],pp104[135],pp104[136],pp104[137],pp104[138],pp104[139],pp104[140],pp104[141],pp104[142],pp104[143],pp104[144],pp104[145],pp104[146],pp104[147],pp104[148],pp104[149],pp104[150],pp104[151],pp104[152],pp104[153],pp104[154],pp104[155],pp104[156],pp104[157],pp104[158],pp104[159],pp104[160],pp104[161],pp104[162],pp104[163],pp104[164],pp104[165],pp104[166],pp104[167],pp104[168],pp104[169],pp104[170],pp104[171],pp104[172],pp104[173],pp104[174],pp104[175],pp104[176],pp104[177],pp104[178],pp104[179],pp104[180],pp104[181],pp104[182],pp104[183],pp104[184],pp104[185],pp104[186],pp104[187],pp104[188],pp104[189],pp104[190],pp104[191],pp104[192],pp104[193],pp104[194],pp104[195],pp104[196],pp104[197],pp104[198],pp104[199],pp104[200],pp104[201],pp104[202],pp104[203],pp104[204],pp104[205],pp104[206],pp104[207],pp104[208],pp104[209],pp104[210],pp104[211],pp104[212],pp104[213],pp104[214],pp104[215],pp104[216],pp104[217],pp104[218],pp104[219],pp104[220],pp104[221],pp104[222],pp104[223],pp104[224],pp104[225],pp104[226],pp104[227],pp104[228],pp104[229],pp104[230],pp104[231],pp104[232],pp104[233],pp104[234],pp104[235],pp104[236],pp104[237],pp104[238],pp104[239],pp104[240],pp104[241],pp104[242],pp104[243],pp104[244],pp104[245],pp104[246],pp104[247],pp104[248],pp104[249],pp104[250],pp104[251],pp105[251],pp106[251],pp107[251],pp108[251],pp109[251],pp110[251],pp111[251],pp112[251],pp113[251],pp114[251],pp115[251],pp116[251],pp117[251],pp118[251],pp119[251],pp120[251],pp121[251],pp122[251],pp123[251],pp124[251],pp125[251],pp126[251],pp127[251],pp128[251],pp129[251],pp130[251]};
    assign in3_2 = {pp15[115],pp15[116],pp15[117],pp15[118],pp15[119],pp15[120],pp15[121],pp15[122],pp15[123],pp15[124],pp15[125],pp15[126],pp15[127],pp15[128],pp15[129],pp15[130],pp15[131],pp15[132],pp15[133],pp15[134],pp15[135],pp15[136],pp15[137],pp15[138],pp15[139],pp15[140],pp15[141],pp15[142],pp15[143],pp15[144],pp15[145],pp15[146],pp15[147],pp15[148],pp15[149],pp15[150],pp15[151],pp15[152],pp15[153],pp15[154],pp15[155],pp15[156],pp15[157],pp15[158],pp15[159],pp15[160],pp15[161],pp15[162],pp15[163],pp15[164],pp15[165],pp15[166],pp15[167],pp15[168],pp15[169],pp15[170],pp15[171],pp15[172],pp15[173],pp15[174],pp15[175],pp15[176],pp15[177],pp15[178],pp15[179],pp15[180],pp15[181],pp15[182],pp15[183],pp15[184],pp14[186],pp13[188],pp12[190],pp11[192],pp10[194],pp105[100],pp105[101],pp105[102],pp105[103],pp105[104],pp105[105],pp105[106],pp105[107],pp105[108],pp105[109],pp105[110],pp105[111],pp105[112],pp105[113],pp105[114],pp105[115],pp105[116],pp105[117],pp105[118],pp105[119],pp105[120],pp105[121],pp105[122],pp105[123],pp105[124],pp105[125],pp105[126],pp105[127],pp105[128],pp105[129],pp105[130],pp105[131],pp105[132],pp105[133],pp105[134],pp105[135],pp105[136],pp105[137],pp105[138],pp105[139],pp105[140],pp105[141],pp105[142],pp105[143],pp105[144],pp105[145],pp105[146],pp105[147],pp105[148],pp105[149],pp105[150],pp105[151],pp105[152],pp105[153],pp105[154],pp105[155],pp105[156],pp105[157],pp105[158],pp105[159],pp105[160],pp105[161],pp105[162],pp105[163],pp105[164],pp105[165],pp105[166],pp105[167],pp105[168],pp105[169],pp105[170],pp105[171],pp105[172],pp105[173],pp105[174],pp105[175],pp105[176],pp105[177],pp105[178],pp105[179],pp105[180],pp105[181],pp105[182],pp105[183],pp105[184],pp105[185],pp105[186],pp105[187],pp105[188],pp105[189],pp105[190],pp105[191],pp105[192],pp105[193],pp105[194],pp105[195],pp105[196],pp105[197],pp105[198],pp105[199],pp105[200],pp105[201],pp105[202],pp105[203],pp105[204],pp105[205],pp105[206],pp105[207],pp105[208],pp105[209],pp105[210],pp105[211],pp105[212],pp105[213],pp105[214],pp105[215],pp105[216],pp105[217],pp105[218],pp105[219],pp105[220],pp105[221],pp105[222],pp105[223],pp105[224],pp105[225],pp105[226],pp105[227],pp105[228],pp105[229],pp105[230],pp105[231],pp105[232],pp105[233],pp105[234],pp105[235],pp105[236],pp105[237],pp105[238],pp105[239],pp105[240],pp105[241],pp105[242],pp105[243],pp105[244],pp105[245],pp105[246],pp105[247],pp105[248],pp105[249],pp105[250],pp106[250],pp107[250],pp108[250],pp109[250],pp110[250],pp111[250],pp112[250],pp113[250],pp114[250],pp115[250],pp116[250],pp117[250],pp118[250],pp119[250],pp120[250],pp121[250],pp122[250],pp123[250],pp124[250],pp125[250],pp126[250],pp127[250],pp128[250],pp129[250],pp130[250],pp131[250]};
    CLA_252 KS_3(s3, c3, in3_1, in3_2);
    wire[249:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp16[115],pp16[116],pp16[117],pp16[118],pp16[119],pp16[120],pp16[121],pp16[122],pp16[123],pp16[124],pp16[125],pp16[126],pp16[127],pp16[128],pp16[129],pp16[130],pp16[131],pp16[132],pp16[133],pp16[134],pp16[135],pp16[136],pp16[137],pp16[138],pp16[139],pp16[140],pp16[141],pp16[142],pp16[143],pp16[144],pp16[145],pp16[146],pp16[147],pp16[148],pp16[149],pp16[150],pp16[151],pp16[152],pp16[153],pp16[154],pp16[155],pp16[156],pp16[157],pp16[158],pp16[159],pp16[160],pp16[161],pp16[162],pp16[163],pp16[164],pp16[165],pp16[166],pp16[167],pp16[168],pp16[169],pp16[170],pp16[171],pp16[172],pp16[173],pp16[174],pp16[175],pp16[176],pp16[177],pp16[178],pp16[179],pp16[180],pp16[181],pp16[182],pp16[183],pp15[185],pp14[187],pp13[189],pp12[191],pp11[193],pp10[195],pp106[100],pp106[101],pp106[102],pp106[103],pp106[104],pp106[105],pp106[106],pp106[107],pp106[108],pp106[109],pp106[110],pp106[111],pp106[112],pp106[113],pp106[114],pp106[115],pp106[116],pp106[117],pp106[118],pp106[119],pp106[120],pp106[121],pp106[122],pp106[123],pp106[124],pp106[125],pp106[126],pp106[127],pp106[128],pp106[129],pp106[130],pp106[131],pp106[132],pp106[133],pp106[134],pp106[135],pp106[136],pp106[137],pp106[138],pp106[139],pp106[140],pp106[141],pp106[142],pp106[143],pp106[144],pp106[145],pp106[146],pp106[147],pp106[148],pp106[149],pp106[150],pp106[151],pp106[152],pp106[153],pp106[154],pp106[155],pp106[156],pp106[157],pp106[158],pp106[159],pp106[160],pp106[161],pp106[162],pp106[163],pp106[164],pp106[165],pp106[166],pp106[167],pp106[168],pp106[169],pp106[170],pp106[171],pp106[172],pp106[173],pp106[174],pp106[175],pp106[176],pp106[177],pp106[178],pp106[179],pp106[180],pp106[181],pp106[182],pp106[183],pp106[184],pp106[185],pp106[186],pp106[187],pp106[188],pp106[189],pp106[190],pp106[191],pp106[192],pp106[193],pp106[194],pp106[195],pp106[196],pp106[197],pp106[198],pp106[199],pp106[200],pp106[201],pp106[202],pp106[203],pp106[204],pp106[205],pp106[206],pp106[207],pp106[208],pp106[209],pp106[210],pp106[211],pp106[212],pp106[213],pp106[214],pp106[215],pp106[216],pp106[217],pp106[218],pp106[219],pp106[220],pp106[221],pp106[222],pp106[223],pp106[224],pp106[225],pp106[226],pp106[227],pp106[228],pp106[229],pp106[230],pp106[231],pp106[232],pp106[233],pp106[234],pp106[235],pp106[236],pp106[237],pp106[238],pp106[239],pp106[240],pp106[241],pp106[242],pp106[243],pp106[244],pp106[245],pp106[246],pp106[247],pp106[248],pp106[249],pp107[249],pp108[249],pp109[249],pp110[249],pp111[249],pp112[249],pp113[249],pp114[249],pp115[249],pp116[249],pp117[249],pp118[249],pp119[249],pp120[249],pp121[249],pp122[249],pp123[249],pp124[249],pp125[249],pp126[249],pp127[249],pp128[249],pp129[249],pp130[249],pp131[249]};
    assign in4_2 = {pp17[114],pp17[115],pp17[116],pp17[117],pp17[118],pp17[119],pp17[120],pp17[121],pp17[122],pp17[123],pp17[124],pp17[125],pp17[126],pp17[127],pp17[128],pp17[129],pp17[130],pp17[131],pp17[132],pp17[133],pp17[134],pp17[135],pp17[136],pp17[137],pp17[138],pp17[139],pp17[140],pp17[141],pp17[142],pp17[143],pp17[144],pp17[145],pp17[146],pp17[147],pp17[148],pp17[149],pp17[150],pp17[151],pp17[152],pp17[153],pp17[154],pp17[155],pp17[156],pp17[157],pp17[158],pp17[159],pp17[160],pp17[161],pp17[162],pp17[163],pp17[164],pp17[165],pp17[166],pp17[167],pp17[168],pp17[169],pp17[170],pp17[171],pp17[172],pp17[173],pp17[174],pp17[175],pp17[176],pp17[177],pp17[178],pp17[179],pp17[180],pp17[181],pp17[182],pp16[184],pp15[186],pp14[188],pp13[190],pp12[192],pp11[194],pp10[196],pp107[100],pp107[101],pp107[102],pp107[103],pp107[104],pp107[105],pp107[106],pp107[107],pp107[108],pp107[109],pp107[110],pp107[111],pp107[112],pp107[113],pp107[114],pp107[115],pp107[116],pp107[117],pp107[118],pp107[119],pp107[120],pp107[121],pp107[122],pp107[123],pp107[124],pp107[125],pp107[126],pp107[127],pp107[128],pp107[129],pp107[130],pp107[131],pp107[132],pp107[133],pp107[134],pp107[135],pp107[136],pp107[137],pp107[138],pp107[139],pp107[140],pp107[141],pp107[142],pp107[143],pp107[144],pp107[145],pp107[146],pp107[147],pp107[148],pp107[149],pp107[150],pp107[151],pp107[152],pp107[153],pp107[154],pp107[155],pp107[156],pp107[157],pp107[158],pp107[159],pp107[160],pp107[161],pp107[162],pp107[163],pp107[164],pp107[165],pp107[166],pp107[167],pp107[168],pp107[169],pp107[170],pp107[171],pp107[172],pp107[173],pp107[174],pp107[175],pp107[176],pp107[177],pp107[178],pp107[179],pp107[180],pp107[181],pp107[182],pp107[183],pp107[184],pp107[185],pp107[186],pp107[187],pp107[188],pp107[189],pp107[190],pp107[191],pp107[192],pp107[193],pp107[194],pp107[195],pp107[196],pp107[197],pp107[198],pp107[199],pp107[200],pp107[201],pp107[202],pp107[203],pp107[204],pp107[205],pp107[206],pp107[207],pp107[208],pp107[209],pp107[210],pp107[211],pp107[212],pp107[213],pp107[214],pp107[215],pp107[216],pp107[217],pp107[218],pp107[219],pp107[220],pp107[221],pp107[222],pp107[223],pp107[224],pp107[225],pp107[226],pp107[227],pp107[228],pp107[229],pp107[230],pp107[231],pp107[232],pp107[233],pp107[234],pp107[235],pp107[236],pp107[237],pp107[238],pp107[239],pp107[240],pp107[241],pp107[242],pp107[243],pp107[244],pp107[245],pp107[246],pp107[247],pp107[248],pp108[248],pp109[248],pp110[248],pp111[248],pp112[248],pp113[248],pp114[248],pp115[248],pp116[248],pp117[248],pp118[248],pp119[248],pp120[248],pp121[248],pp122[248],pp123[248],pp124[248],pp125[248],pp126[248],pp127[248],pp128[248],pp129[248],pp130[248],pp131[248],pp132[248]};
    CLA_250 KS_4(s4, c4, in4_1, in4_2);
    wire[247:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp18[114],pp18[115],pp18[116],pp18[117],pp18[118],pp18[119],pp18[120],pp18[121],pp18[122],pp18[123],pp18[124],pp18[125],pp18[126],pp18[127],pp18[128],pp18[129],pp18[130],pp18[131],pp18[132],pp18[133],pp18[134],pp18[135],pp18[136],pp18[137],pp18[138],pp18[139],pp18[140],pp18[141],pp18[142],pp18[143],pp18[144],pp18[145],pp18[146],pp18[147],pp18[148],pp18[149],pp18[150],pp18[151],pp18[152],pp18[153],pp18[154],pp18[155],pp18[156],pp18[157],pp18[158],pp18[159],pp18[160],pp18[161],pp18[162],pp18[163],pp18[164],pp18[165],pp18[166],pp18[167],pp18[168],pp18[169],pp18[170],pp18[171],pp18[172],pp18[173],pp18[174],pp18[175],pp18[176],pp18[177],pp18[178],pp18[179],pp18[180],pp18[181],pp17[183],pp16[185],pp15[187],pp14[189],pp13[191],pp12[193],pp11[195],pp10[197],pp108[100],pp108[101],pp108[102],pp108[103],pp108[104],pp108[105],pp108[106],pp108[107],pp108[108],pp108[109],pp108[110],pp108[111],pp108[112],pp108[113],pp108[114],pp108[115],pp108[116],pp108[117],pp108[118],pp108[119],pp108[120],pp108[121],pp108[122],pp108[123],pp108[124],pp108[125],pp108[126],pp108[127],pp108[128],pp108[129],pp108[130],pp108[131],pp108[132],pp108[133],pp108[134],pp108[135],pp108[136],pp108[137],pp108[138],pp108[139],pp108[140],pp108[141],pp108[142],pp108[143],pp108[144],pp108[145],pp108[146],pp108[147],pp108[148],pp108[149],pp108[150],pp108[151],pp108[152],pp108[153],pp108[154],pp108[155],pp108[156],pp108[157],pp108[158],pp108[159],pp108[160],pp108[161],pp108[162],pp108[163],pp108[164],pp108[165],pp108[166],pp108[167],pp108[168],pp108[169],pp108[170],pp108[171],pp108[172],pp108[173],pp108[174],pp108[175],pp108[176],pp108[177],pp108[178],pp108[179],pp108[180],pp108[181],pp108[182],pp108[183],pp108[184],pp108[185],pp108[186],pp108[187],pp108[188],pp108[189],pp108[190],pp108[191],pp108[192],pp108[193],pp108[194],pp108[195],pp108[196],pp108[197],pp108[198],pp108[199],pp108[200],pp108[201],pp108[202],pp108[203],pp108[204],pp108[205],pp108[206],pp108[207],pp108[208],pp108[209],pp108[210],pp108[211],pp108[212],pp108[213],pp108[214],pp108[215],pp108[216],pp108[217],pp108[218],pp108[219],pp108[220],pp108[221],pp108[222],pp108[223],pp108[224],pp108[225],pp108[226],pp108[227],pp108[228],pp108[229],pp108[230],pp108[231],pp108[232],pp108[233],pp108[234],pp108[235],pp108[236],pp108[237],pp108[238],pp108[239],pp108[240],pp108[241],pp108[242],pp108[243],pp108[244],pp108[245],pp108[246],pp108[247],pp109[247],pp110[247],pp111[247],pp112[247],pp113[247],pp114[247],pp115[247],pp116[247],pp117[247],pp118[247],pp119[247],pp120[247],pp121[247],pp122[247],pp123[247],pp124[247],pp125[247],pp126[247],pp127[247],pp128[247],pp129[247],pp130[247],pp131[247],pp132[247]};
    assign in5_2 = {pp19[113],pp19[114],pp19[115],pp19[116],pp19[117],pp19[118],pp19[119],pp19[120],pp19[121],pp19[122],pp19[123],pp19[124],pp19[125],pp19[126],pp19[127],pp19[128],pp19[129],pp19[130],pp19[131],pp19[132],pp19[133],pp19[134],pp19[135],pp19[136],pp19[137],pp19[138],pp19[139],pp19[140],pp19[141],pp19[142],pp19[143],pp19[144],pp19[145],pp19[146],pp19[147],pp19[148],pp19[149],pp19[150],pp19[151],pp19[152],pp19[153],pp19[154],pp19[155],pp19[156],pp19[157],pp19[158],pp19[159],pp19[160],pp19[161],pp19[162],pp19[163],pp19[164],pp19[165],pp19[166],pp19[167],pp19[168],pp19[169],pp19[170],pp19[171],pp19[172],pp19[173],pp19[174],pp19[175],pp19[176],pp19[177],pp19[178],pp19[179],pp19[180],pp18[182],pp17[184],pp16[186],pp15[188],pp14[190],pp13[192],pp12[194],pp11[196],pp10[198],pp109[100],pp109[101],pp109[102],pp109[103],pp109[104],pp109[105],pp109[106],pp109[107],pp109[108],pp109[109],pp109[110],pp109[111],pp109[112],pp109[113],pp109[114],pp109[115],pp109[116],pp109[117],pp109[118],pp109[119],pp109[120],pp109[121],pp109[122],pp109[123],pp109[124],pp109[125],pp109[126],pp109[127],pp109[128],pp109[129],pp109[130],pp109[131],pp109[132],pp109[133],pp109[134],pp109[135],pp109[136],pp109[137],pp109[138],pp109[139],pp109[140],pp109[141],pp109[142],pp109[143],pp109[144],pp109[145],pp109[146],pp109[147],pp109[148],pp109[149],pp109[150],pp109[151],pp109[152],pp109[153],pp109[154],pp109[155],pp109[156],pp109[157],pp109[158],pp109[159],pp109[160],pp109[161],pp109[162],pp109[163],pp109[164],pp109[165],pp109[166],pp109[167],pp109[168],pp109[169],pp109[170],pp109[171],pp109[172],pp109[173],pp109[174],pp109[175],pp109[176],pp109[177],pp109[178],pp109[179],pp109[180],pp109[181],pp109[182],pp109[183],pp109[184],pp109[185],pp109[186],pp109[187],pp109[188],pp109[189],pp109[190],pp109[191],pp109[192],pp109[193],pp109[194],pp109[195],pp109[196],pp109[197],pp109[198],pp109[199],pp109[200],pp109[201],pp109[202],pp109[203],pp109[204],pp109[205],pp109[206],pp109[207],pp109[208],pp109[209],pp109[210],pp109[211],pp109[212],pp109[213],pp109[214],pp109[215],pp109[216],pp109[217],pp109[218],pp109[219],pp109[220],pp109[221],pp109[222],pp109[223],pp109[224],pp109[225],pp109[226],pp109[227],pp109[228],pp109[229],pp109[230],pp109[231],pp109[232],pp109[233],pp109[234],pp109[235],pp109[236],pp109[237],pp109[238],pp109[239],pp109[240],pp109[241],pp109[242],pp109[243],pp109[244],pp109[245],pp109[246],pp110[246],pp111[246],pp112[246],pp113[246],pp114[246],pp115[246],pp116[246],pp117[246],pp118[246],pp119[246],pp120[246],pp121[246],pp122[246],pp123[246],pp124[246],pp125[246],pp126[246],pp127[246],pp128[246],pp129[246],pp130[246],pp131[246],pp132[246],pp133[246]};
    CLA_248 KS_5(s5, c5, in5_1, in5_2);
    wire[245:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp20[113],pp20[114],pp20[115],pp20[116],pp20[117],pp20[118],pp20[119],pp20[120],pp20[121],pp20[122],pp20[123],pp20[124],pp20[125],pp20[126],pp20[127],pp20[128],pp20[129],pp20[130],pp20[131],pp20[132],pp20[133],pp20[134],pp20[135],pp20[136],pp20[137],pp20[138],pp20[139],pp20[140],pp20[141],pp20[142],pp20[143],pp20[144],pp20[145],pp20[146],pp20[147],pp20[148],pp20[149],pp20[150],pp20[151],pp20[152],pp20[153],pp20[154],pp20[155],pp20[156],pp20[157],pp20[158],pp20[159],pp20[160],pp20[161],pp20[162],pp20[163],pp20[164],pp20[165],pp20[166],pp20[167],pp20[168],pp20[169],pp20[170],pp20[171],pp20[172],pp20[173],pp20[174],pp20[175],pp20[176],pp20[177],pp20[178],pp20[179],pp19[181],pp18[183],pp17[185],pp16[187],pp15[189],pp14[191],pp13[193],pp12[195],pp11[197],pp10[199],pp110[100],pp110[101],pp110[102],pp110[103],pp110[104],pp110[105],pp110[106],pp110[107],pp110[108],pp110[109],pp110[110],pp110[111],pp110[112],pp110[113],pp110[114],pp110[115],pp110[116],pp110[117],pp110[118],pp110[119],pp110[120],pp110[121],pp110[122],pp110[123],pp110[124],pp110[125],pp110[126],pp110[127],pp110[128],pp110[129],pp110[130],pp110[131],pp110[132],pp110[133],pp110[134],pp110[135],pp110[136],pp110[137],pp110[138],pp110[139],pp110[140],pp110[141],pp110[142],pp110[143],pp110[144],pp110[145],pp110[146],pp110[147],pp110[148],pp110[149],pp110[150],pp110[151],pp110[152],pp110[153],pp110[154],pp110[155],pp110[156],pp110[157],pp110[158],pp110[159],pp110[160],pp110[161],pp110[162],pp110[163],pp110[164],pp110[165],pp110[166],pp110[167],pp110[168],pp110[169],pp110[170],pp110[171],pp110[172],pp110[173],pp110[174],pp110[175],pp110[176],pp110[177],pp110[178],pp110[179],pp110[180],pp110[181],pp110[182],pp110[183],pp110[184],pp110[185],pp110[186],pp110[187],pp110[188],pp110[189],pp110[190],pp110[191],pp110[192],pp110[193],pp110[194],pp110[195],pp110[196],pp110[197],pp110[198],pp110[199],pp110[200],pp110[201],pp110[202],pp110[203],pp110[204],pp110[205],pp110[206],pp110[207],pp110[208],pp110[209],pp110[210],pp110[211],pp110[212],pp110[213],pp110[214],pp110[215],pp110[216],pp110[217],pp110[218],pp110[219],pp110[220],pp110[221],pp110[222],pp110[223],pp110[224],pp110[225],pp110[226],pp110[227],pp110[228],pp110[229],pp110[230],pp110[231],pp110[232],pp110[233],pp110[234],pp110[235],pp110[236],pp110[237],pp110[238],pp110[239],pp110[240],pp110[241],pp110[242],pp110[243],pp110[244],pp110[245],pp111[245],pp112[245],pp113[245],pp114[245],pp115[245],pp116[245],pp117[245],pp118[245],pp119[245],pp120[245],pp121[245],pp122[245],pp123[245],pp124[245],pp125[245],pp126[245],pp127[245],pp128[245],pp129[245],pp130[245],pp131[245],pp132[245],pp133[245]};
    assign in6_2 = {pp21[112],pp21[113],pp21[114],pp21[115],pp21[116],pp21[117],pp21[118],pp21[119],pp21[120],pp21[121],pp21[122],pp21[123],pp21[124],pp21[125],pp21[126],pp21[127],pp21[128],pp21[129],pp21[130],pp21[131],pp21[132],pp21[133],pp21[134],pp21[135],pp21[136],pp21[137],pp21[138],pp21[139],pp21[140],pp21[141],pp21[142],pp21[143],pp21[144],pp21[145],pp21[146],pp21[147],pp21[148],pp21[149],pp21[150],pp21[151],pp21[152],pp21[153],pp21[154],pp21[155],pp21[156],pp21[157],pp21[158],pp21[159],pp21[160],pp21[161],pp21[162],pp21[163],pp21[164],pp21[165],pp21[166],pp21[167],pp21[168],pp21[169],pp21[170],pp21[171],pp21[172],pp21[173],pp21[174],pp21[175],pp21[176],pp21[177],pp21[178],pp20[180],pp19[182],pp18[184],pp17[186],pp16[188],pp15[190],pp14[192],pp13[194],pp12[196],pp11[198],pp10[200],pp111[100],pp111[101],pp111[102],pp111[103],pp111[104],pp111[105],pp111[106],pp111[107],pp111[108],pp111[109],pp111[110],pp111[111],pp111[112],pp111[113],pp111[114],pp111[115],pp111[116],pp111[117],pp111[118],pp111[119],pp111[120],pp111[121],pp111[122],pp111[123],pp111[124],pp111[125],pp111[126],pp111[127],pp111[128],pp111[129],pp111[130],pp111[131],pp111[132],pp111[133],pp111[134],pp111[135],pp111[136],pp111[137],pp111[138],pp111[139],pp111[140],pp111[141],pp111[142],pp111[143],pp111[144],pp111[145],pp111[146],pp111[147],pp111[148],pp111[149],pp111[150],pp111[151],pp111[152],pp111[153],pp111[154],pp111[155],pp111[156],pp111[157],pp111[158],pp111[159],pp111[160],pp111[161],pp111[162],pp111[163],pp111[164],pp111[165],pp111[166],pp111[167],pp111[168],pp111[169],pp111[170],pp111[171],pp111[172],pp111[173],pp111[174],pp111[175],pp111[176],pp111[177],pp111[178],pp111[179],pp111[180],pp111[181],pp111[182],pp111[183],pp111[184],pp111[185],pp111[186],pp111[187],pp111[188],pp111[189],pp111[190],pp111[191],pp111[192],pp111[193],pp111[194],pp111[195],pp111[196],pp111[197],pp111[198],pp111[199],pp111[200],pp111[201],pp111[202],pp111[203],pp111[204],pp111[205],pp111[206],pp111[207],pp111[208],pp111[209],pp111[210],pp111[211],pp111[212],pp111[213],pp111[214],pp111[215],pp111[216],pp111[217],pp111[218],pp111[219],pp111[220],pp111[221],pp111[222],pp111[223],pp111[224],pp111[225],pp111[226],pp111[227],pp111[228],pp111[229],pp111[230],pp111[231],pp111[232],pp111[233],pp111[234],pp111[235],pp111[236],pp111[237],pp111[238],pp111[239],pp111[240],pp111[241],pp111[242],pp111[243],pp111[244],pp112[244],pp113[244],pp114[244],pp115[244],pp116[244],pp117[244],pp118[244],pp119[244],pp120[244],pp121[244],pp122[244],pp123[244],pp124[244],pp125[244],pp126[244],pp127[244],pp128[244],pp129[244],pp130[244],pp131[244],pp132[244],pp133[244],pp134[244]};
    CLA_246 KS_6(s6, c6, in6_1, in6_2);
    wire[243:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp22[112],pp22[113],pp22[114],pp22[115],pp22[116],pp22[117],pp22[118],pp22[119],pp22[120],pp22[121],pp22[122],pp22[123],pp22[124],pp22[125],pp22[126],pp22[127],pp22[128],pp22[129],pp22[130],pp22[131],pp22[132],pp22[133],pp22[134],pp22[135],pp22[136],pp22[137],pp22[138],pp22[139],pp22[140],pp22[141],pp22[142],pp22[143],pp22[144],pp22[145],pp22[146],pp22[147],pp22[148],pp22[149],pp22[150],pp22[151],pp22[152],pp22[153],pp22[154],pp22[155],pp22[156],pp22[157],pp22[158],pp22[159],pp22[160],pp22[161],pp22[162],pp22[163],pp22[164],pp22[165],pp22[166],pp22[167],pp22[168],pp22[169],pp22[170],pp22[171],pp22[172],pp22[173],pp22[174],pp22[175],pp22[176],pp22[177],pp21[179],pp20[181],pp19[183],pp18[185],pp17[187],pp16[189],pp15[191],pp14[193],pp13[195],pp12[197],pp11[199],pp10[201],pp112[100],pp112[101],pp112[102],pp112[103],pp112[104],pp112[105],pp112[106],pp112[107],pp112[108],pp112[109],pp112[110],pp112[111],pp112[112],pp112[113],pp112[114],pp112[115],pp112[116],pp112[117],pp112[118],pp112[119],pp112[120],pp112[121],pp112[122],pp112[123],pp112[124],pp112[125],pp112[126],pp112[127],pp112[128],pp112[129],pp112[130],pp112[131],pp112[132],pp112[133],pp112[134],pp112[135],pp112[136],pp112[137],pp112[138],pp112[139],pp112[140],pp112[141],pp112[142],pp112[143],pp112[144],pp112[145],pp112[146],pp112[147],pp112[148],pp112[149],pp112[150],pp112[151],pp112[152],pp112[153],pp112[154],pp112[155],pp112[156],pp112[157],pp112[158],pp112[159],pp112[160],pp112[161],pp112[162],pp112[163],pp112[164],pp112[165],pp112[166],pp112[167],pp112[168],pp112[169],pp112[170],pp112[171],pp112[172],pp112[173],pp112[174],pp112[175],pp112[176],pp112[177],pp112[178],pp112[179],pp112[180],pp112[181],pp112[182],pp112[183],pp112[184],pp112[185],pp112[186],pp112[187],pp112[188],pp112[189],pp112[190],pp112[191],pp112[192],pp112[193],pp112[194],pp112[195],pp112[196],pp112[197],pp112[198],pp112[199],pp112[200],pp112[201],pp112[202],pp112[203],pp112[204],pp112[205],pp112[206],pp112[207],pp112[208],pp112[209],pp112[210],pp112[211],pp112[212],pp112[213],pp112[214],pp112[215],pp112[216],pp112[217],pp112[218],pp112[219],pp112[220],pp112[221],pp112[222],pp112[223],pp112[224],pp112[225],pp112[226],pp112[227],pp112[228],pp112[229],pp112[230],pp112[231],pp112[232],pp112[233],pp112[234],pp112[235],pp112[236],pp112[237],pp112[238],pp112[239],pp112[240],pp112[241],pp112[242],pp112[243],pp113[243],pp114[243],pp115[243],pp116[243],pp117[243],pp118[243],pp119[243],pp120[243],pp121[243],pp122[243],pp123[243],pp124[243],pp125[243],pp126[243],pp127[243],pp128[243],pp129[243],pp130[243],pp131[243],pp132[243],pp133[243],pp134[243]};
    assign in7_2 = {pp23[111],pp23[112],pp23[113],pp23[114],pp23[115],pp23[116],pp23[117],pp23[118],pp23[119],pp23[120],pp23[121],pp23[122],pp23[123],pp23[124],pp23[125],pp23[126],pp23[127],pp23[128],pp23[129],pp23[130],pp23[131],pp23[132],pp23[133],pp23[134],pp23[135],pp23[136],pp23[137],pp23[138],pp23[139],pp23[140],pp23[141],pp23[142],pp23[143],pp23[144],pp23[145],pp23[146],pp23[147],pp23[148],pp23[149],pp23[150],pp23[151],pp23[152],pp23[153],pp23[154],pp23[155],pp23[156],pp23[157],pp23[158],pp23[159],pp23[160],pp23[161],pp23[162],pp23[163],pp23[164],pp23[165],pp23[166],pp23[167],pp23[168],pp23[169],pp23[170],pp23[171],pp23[172],pp23[173],pp23[174],pp23[175],pp23[176],pp22[178],pp21[180],pp20[182],pp19[184],pp18[186],pp17[188],pp16[190],pp15[192],pp14[194],pp13[196],pp12[198],pp11[200],pp10[202],pp113[100],pp113[101],pp113[102],pp113[103],pp113[104],pp113[105],pp113[106],pp113[107],pp113[108],pp113[109],pp113[110],pp113[111],pp113[112],pp113[113],pp113[114],pp113[115],pp113[116],pp113[117],pp113[118],pp113[119],pp113[120],pp113[121],pp113[122],pp113[123],pp113[124],pp113[125],pp113[126],pp113[127],pp113[128],pp113[129],pp113[130],pp113[131],pp113[132],pp113[133],pp113[134],pp113[135],pp113[136],pp113[137],pp113[138],pp113[139],pp113[140],pp113[141],pp113[142],pp113[143],pp113[144],pp113[145],pp113[146],pp113[147],pp113[148],pp113[149],pp113[150],pp113[151],pp113[152],pp113[153],pp113[154],pp113[155],pp113[156],pp113[157],pp113[158],pp113[159],pp113[160],pp113[161],pp113[162],pp113[163],pp113[164],pp113[165],pp113[166],pp113[167],pp113[168],pp113[169],pp113[170],pp113[171],pp113[172],pp113[173],pp113[174],pp113[175],pp113[176],pp113[177],pp113[178],pp113[179],pp113[180],pp113[181],pp113[182],pp113[183],pp113[184],pp113[185],pp113[186],pp113[187],pp113[188],pp113[189],pp113[190],pp113[191],pp113[192],pp113[193],pp113[194],pp113[195],pp113[196],pp113[197],pp113[198],pp113[199],pp113[200],pp113[201],pp113[202],pp113[203],pp113[204],pp113[205],pp113[206],pp113[207],pp113[208],pp113[209],pp113[210],pp113[211],pp113[212],pp113[213],pp113[214],pp113[215],pp113[216],pp113[217],pp113[218],pp113[219],pp113[220],pp113[221],pp113[222],pp113[223],pp113[224],pp113[225],pp113[226],pp113[227],pp113[228],pp113[229],pp113[230],pp113[231],pp113[232],pp113[233],pp113[234],pp113[235],pp113[236],pp113[237],pp113[238],pp113[239],pp113[240],pp113[241],pp113[242],pp114[242],pp115[242],pp116[242],pp117[242],pp118[242],pp119[242],pp120[242],pp121[242],pp122[242],pp123[242],pp124[242],pp125[242],pp126[242],pp127[242],pp128[242],pp129[242],pp130[242],pp131[242],pp132[242],pp133[242],pp134[242],pp135[242]};
    CLA_244 KS_7(s7, c7, in7_1, in7_2);
    wire[241:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp24[111],pp24[112],pp24[113],pp24[114],pp24[115],pp24[116],pp24[117],pp24[118],pp24[119],pp24[120],pp24[121],pp24[122],pp24[123],pp24[124],pp24[125],pp24[126],pp24[127],pp24[128],pp24[129],pp24[130],pp24[131],pp24[132],pp24[133],pp24[134],pp24[135],pp24[136],pp24[137],pp24[138],pp24[139],pp24[140],pp24[141],pp24[142],pp24[143],pp24[144],pp24[145],pp24[146],pp24[147],pp24[148],pp24[149],pp24[150],pp24[151],pp24[152],pp24[153],pp24[154],pp24[155],pp24[156],pp24[157],pp24[158],pp24[159],pp24[160],pp24[161],pp24[162],pp24[163],pp24[164],pp24[165],pp24[166],pp24[167],pp24[168],pp24[169],pp24[170],pp24[171],pp24[172],pp24[173],pp24[174],pp24[175],pp23[177],pp22[179],pp21[181],pp20[183],pp19[185],pp18[187],pp17[189],pp16[191],pp15[193],pp14[195],pp13[197],pp12[199],pp11[201],pp10[203],pp114[100],pp114[101],pp114[102],pp114[103],pp114[104],pp114[105],pp114[106],pp114[107],pp114[108],pp114[109],pp114[110],pp114[111],pp114[112],pp114[113],pp114[114],pp114[115],pp114[116],pp114[117],pp114[118],pp114[119],pp114[120],pp114[121],pp114[122],pp114[123],pp114[124],pp114[125],pp114[126],pp114[127],pp114[128],pp114[129],pp114[130],pp114[131],pp114[132],pp114[133],pp114[134],pp114[135],pp114[136],pp114[137],pp114[138],pp114[139],pp114[140],pp114[141],pp114[142],pp114[143],pp114[144],pp114[145],pp114[146],pp114[147],pp114[148],pp114[149],pp114[150],pp114[151],pp114[152],pp114[153],pp114[154],pp114[155],pp114[156],pp114[157],pp114[158],pp114[159],pp114[160],pp114[161],pp114[162],pp114[163],pp114[164],pp114[165],pp114[166],pp114[167],pp114[168],pp114[169],pp114[170],pp114[171],pp114[172],pp114[173],pp114[174],pp114[175],pp114[176],pp114[177],pp114[178],pp114[179],pp114[180],pp114[181],pp114[182],pp114[183],pp114[184],pp114[185],pp114[186],pp114[187],pp114[188],pp114[189],pp114[190],pp114[191],pp114[192],pp114[193],pp114[194],pp114[195],pp114[196],pp114[197],pp114[198],pp114[199],pp114[200],pp114[201],pp114[202],pp114[203],pp114[204],pp114[205],pp114[206],pp114[207],pp114[208],pp114[209],pp114[210],pp114[211],pp114[212],pp114[213],pp114[214],pp114[215],pp114[216],pp114[217],pp114[218],pp114[219],pp114[220],pp114[221],pp114[222],pp114[223],pp114[224],pp114[225],pp114[226],pp114[227],pp114[228],pp114[229],pp114[230],pp114[231],pp114[232],pp114[233],pp114[234],pp114[235],pp114[236],pp114[237],pp114[238],pp114[239],pp114[240],pp114[241],pp115[241],pp116[241],pp117[241],pp118[241],pp119[241],pp120[241],pp121[241],pp122[241],pp123[241],pp124[241],pp125[241],pp126[241],pp127[241],pp128[241],pp129[241],pp130[241],pp131[241],pp132[241],pp133[241],pp134[241],pp135[241]};
    assign in8_2 = {pp25[110],pp25[111],pp25[112],pp25[113],pp25[114],pp25[115],pp25[116],pp25[117],pp25[118],pp25[119],pp25[120],pp25[121],pp25[122],pp25[123],pp25[124],pp25[125],pp25[126],pp25[127],pp25[128],pp25[129],pp25[130],pp25[131],pp25[132],pp25[133],pp25[134],pp25[135],pp25[136],pp25[137],pp25[138],pp25[139],pp25[140],pp25[141],pp25[142],pp25[143],pp25[144],pp25[145],pp25[146],pp25[147],pp25[148],pp25[149],pp25[150],pp25[151],pp25[152],pp25[153],pp25[154],pp25[155],pp25[156],pp25[157],pp25[158],pp25[159],pp25[160],pp25[161],pp25[162],pp25[163],pp25[164],pp25[165],pp25[166],pp25[167],pp25[168],pp25[169],pp25[170],pp25[171],pp25[172],pp25[173],pp25[174],pp24[176],pp23[178],pp22[180],pp21[182],pp20[184],pp19[186],pp18[188],pp17[190],pp16[192],pp15[194],pp14[196],pp13[198],pp12[200],pp11[202],pp10[204],pp115[100],pp115[101],pp115[102],pp115[103],pp115[104],pp115[105],pp115[106],pp115[107],pp115[108],pp115[109],pp115[110],pp115[111],pp115[112],pp115[113],pp115[114],pp115[115],pp115[116],pp115[117],pp115[118],pp115[119],pp115[120],pp115[121],pp115[122],pp115[123],pp115[124],pp115[125],pp115[126],pp115[127],pp115[128],pp115[129],pp115[130],pp115[131],pp115[132],pp115[133],pp115[134],pp115[135],pp115[136],pp115[137],pp115[138],pp115[139],pp115[140],pp115[141],pp115[142],pp115[143],pp115[144],pp115[145],pp115[146],pp115[147],pp115[148],pp115[149],pp115[150],pp115[151],pp115[152],pp115[153],pp115[154],pp115[155],pp115[156],pp115[157],pp115[158],pp115[159],pp115[160],pp115[161],pp115[162],pp115[163],pp115[164],pp115[165],pp115[166],pp115[167],pp115[168],pp115[169],pp115[170],pp115[171],pp115[172],pp115[173],pp115[174],pp115[175],pp115[176],pp115[177],pp115[178],pp115[179],pp115[180],pp115[181],pp115[182],pp115[183],pp115[184],pp115[185],pp115[186],pp115[187],pp115[188],pp115[189],pp115[190],pp115[191],pp115[192],pp115[193],pp115[194],pp115[195],pp115[196],pp115[197],pp115[198],pp115[199],pp115[200],pp115[201],pp115[202],pp115[203],pp115[204],pp115[205],pp115[206],pp115[207],pp115[208],pp115[209],pp115[210],pp115[211],pp115[212],pp115[213],pp115[214],pp115[215],pp115[216],pp115[217],pp115[218],pp115[219],pp115[220],pp115[221],pp115[222],pp115[223],pp115[224],pp115[225],pp115[226],pp115[227],pp115[228],pp115[229],pp115[230],pp115[231],pp115[232],pp115[233],pp115[234],pp115[235],pp115[236],pp115[237],pp115[238],pp115[239],pp115[240],pp116[240],pp117[240],pp118[240],pp119[240],pp120[240],pp121[240],pp122[240],pp123[240],pp124[240],pp125[240],pp126[240],pp127[240],pp128[240],pp129[240],pp130[240],pp131[240],pp132[240],pp133[240],pp134[240],pp135[240],pp136[240]};
    CLA_242 KS_8(s8, c8, in8_1, in8_2);
    wire[239:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp26[110],pp26[111],pp26[112],pp26[113],pp26[114],pp26[115],pp26[116],pp26[117],pp26[118],pp26[119],pp26[120],pp26[121],pp26[122],pp26[123],pp26[124],pp26[125],pp26[126],pp26[127],pp26[128],pp26[129],pp26[130],pp26[131],pp26[132],pp26[133],pp26[134],pp26[135],pp26[136],pp26[137],pp26[138],pp26[139],pp26[140],pp26[141],pp26[142],pp26[143],pp26[144],pp26[145],pp26[146],pp26[147],pp26[148],pp26[149],pp26[150],pp26[151],pp26[152],pp26[153],pp26[154],pp26[155],pp26[156],pp26[157],pp26[158],pp26[159],pp26[160],pp26[161],pp26[162],pp26[163],pp26[164],pp26[165],pp26[166],pp26[167],pp26[168],pp26[169],pp26[170],pp26[171],pp26[172],pp26[173],pp25[175],pp24[177],pp23[179],pp22[181],pp21[183],pp20[185],pp19[187],pp18[189],pp17[191],pp16[193],pp15[195],pp14[197],pp13[199],pp12[201],pp11[203],pp10[205],pp116[100],pp116[101],pp116[102],pp116[103],pp116[104],pp116[105],pp116[106],pp116[107],pp116[108],pp116[109],pp116[110],pp116[111],pp116[112],pp116[113],pp116[114],pp116[115],pp116[116],pp116[117],pp116[118],pp116[119],pp116[120],pp116[121],pp116[122],pp116[123],pp116[124],pp116[125],pp116[126],pp116[127],pp116[128],pp116[129],pp116[130],pp116[131],pp116[132],pp116[133],pp116[134],pp116[135],pp116[136],pp116[137],pp116[138],pp116[139],pp116[140],pp116[141],pp116[142],pp116[143],pp116[144],pp116[145],pp116[146],pp116[147],pp116[148],pp116[149],pp116[150],pp116[151],pp116[152],pp116[153],pp116[154],pp116[155],pp116[156],pp116[157],pp116[158],pp116[159],pp116[160],pp116[161],pp116[162],pp116[163],pp116[164],pp116[165],pp116[166],pp116[167],pp116[168],pp116[169],pp116[170],pp116[171],pp116[172],pp116[173],pp116[174],pp116[175],pp116[176],pp116[177],pp116[178],pp116[179],pp116[180],pp116[181],pp116[182],pp116[183],pp116[184],pp116[185],pp116[186],pp116[187],pp116[188],pp116[189],pp116[190],pp116[191],pp116[192],pp116[193],pp116[194],pp116[195],pp116[196],pp116[197],pp116[198],pp116[199],pp116[200],pp116[201],pp116[202],pp116[203],pp116[204],pp116[205],pp116[206],pp116[207],pp116[208],pp116[209],pp116[210],pp116[211],pp116[212],pp116[213],pp116[214],pp116[215],pp116[216],pp116[217],pp116[218],pp116[219],pp116[220],pp116[221],pp116[222],pp116[223],pp116[224],pp116[225],pp116[226],pp116[227],pp116[228],pp116[229],pp116[230],pp116[231],pp116[232],pp116[233],pp116[234],pp116[235],pp116[236],pp116[237],pp116[238],pp116[239],pp117[239],pp118[239],pp119[239],pp120[239],pp121[239],pp122[239],pp123[239],pp124[239],pp125[239],pp126[239],pp127[239],pp128[239],pp129[239],pp130[239],pp131[239],pp132[239],pp133[239],pp134[239],pp135[239],pp136[239]};
    assign in9_2 = {pp27[109],pp27[110],pp27[111],pp27[112],pp27[113],pp27[114],pp27[115],pp27[116],pp27[117],pp27[118],pp27[119],pp27[120],pp27[121],pp27[122],pp27[123],pp27[124],pp27[125],pp27[126],pp27[127],pp27[128],pp27[129],pp27[130],pp27[131],pp27[132],pp27[133],pp27[134],pp27[135],pp27[136],pp27[137],pp27[138],pp27[139],pp27[140],pp27[141],pp27[142],pp27[143],pp27[144],pp27[145],pp27[146],pp27[147],pp27[148],pp27[149],pp27[150],pp27[151],pp27[152],pp27[153],pp27[154],pp27[155],pp27[156],pp27[157],pp27[158],pp27[159],pp27[160],pp27[161],pp27[162],pp27[163],pp27[164],pp27[165],pp27[166],pp27[167],pp27[168],pp27[169],pp27[170],pp27[171],pp27[172],pp26[174],pp25[176],pp24[178],pp23[180],pp22[182],pp21[184],pp20[186],pp19[188],pp18[190],pp17[192],pp16[194],pp15[196],pp14[198],pp13[200],pp12[202],pp11[204],pp10[206],pp117[100],pp117[101],pp117[102],pp117[103],pp117[104],pp117[105],pp117[106],pp117[107],pp117[108],pp117[109],pp117[110],pp117[111],pp117[112],pp117[113],pp117[114],pp117[115],pp117[116],pp117[117],pp117[118],pp117[119],pp117[120],pp117[121],pp117[122],pp117[123],pp117[124],pp117[125],pp117[126],pp117[127],pp117[128],pp117[129],pp117[130],pp117[131],pp117[132],pp117[133],pp117[134],pp117[135],pp117[136],pp117[137],pp117[138],pp117[139],pp117[140],pp117[141],pp117[142],pp117[143],pp117[144],pp117[145],pp117[146],pp117[147],pp117[148],pp117[149],pp117[150],pp117[151],pp117[152],pp117[153],pp117[154],pp117[155],pp117[156],pp117[157],pp117[158],pp117[159],pp117[160],pp117[161],pp117[162],pp117[163],pp117[164],pp117[165],pp117[166],pp117[167],pp117[168],pp117[169],pp117[170],pp117[171],pp117[172],pp117[173],pp117[174],pp117[175],pp117[176],pp117[177],pp117[178],pp117[179],pp117[180],pp117[181],pp117[182],pp117[183],pp117[184],pp117[185],pp117[186],pp117[187],pp117[188],pp117[189],pp117[190],pp117[191],pp117[192],pp117[193],pp117[194],pp117[195],pp117[196],pp117[197],pp117[198],pp117[199],pp117[200],pp117[201],pp117[202],pp117[203],pp117[204],pp117[205],pp117[206],pp117[207],pp117[208],pp117[209],pp117[210],pp117[211],pp117[212],pp117[213],pp117[214],pp117[215],pp117[216],pp117[217],pp117[218],pp117[219],pp117[220],pp117[221],pp117[222],pp117[223],pp117[224],pp117[225],pp117[226],pp117[227],pp117[228],pp117[229],pp117[230],pp117[231],pp117[232],pp117[233],pp117[234],pp117[235],pp117[236],pp117[237],pp117[238],pp118[238],pp119[238],pp120[238],pp121[238],pp122[238],pp123[238],pp124[238],pp125[238],pp126[238],pp127[238],pp128[238],pp129[238],pp130[238],pp131[238],pp132[238],pp133[238],pp134[238],pp135[238],pp136[238],pp137[238]};
    CLA_240 KS_9(s9, c9, in9_1, in9_2);
    wire[237:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp28[109],pp28[110],pp28[111],pp28[112],pp28[113],pp28[114],pp28[115],pp28[116],pp28[117],pp28[118],pp28[119],pp28[120],pp28[121],pp28[122],pp28[123],pp28[124],pp28[125],pp28[126],pp28[127],pp28[128],pp28[129],pp28[130],pp28[131],pp28[132],pp28[133],pp28[134],pp28[135],pp28[136],pp28[137],pp28[138],pp28[139],pp28[140],pp28[141],pp28[142],pp28[143],pp28[144],pp28[145],pp28[146],pp28[147],pp28[148],pp28[149],pp28[150],pp28[151],pp28[152],pp28[153],pp28[154],pp28[155],pp28[156],pp28[157],pp28[158],pp28[159],pp28[160],pp28[161],pp28[162],pp28[163],pp28[164],pp28[165],pp28[166],pp28[167],pp28[168],pp28[169],pp28[170],pp28[171],pp27[173],pp26[175],pp25[177],pp24[179],pp23[181],pp22[183],pp21[185],pp20[187],pp19[189],pp18[191],pp17[193],pp16[195],pp15[197],pp14[199],pp13[201],pp12[203],pp11[205],pp10[207],pp118[100],pp118[101],pp118[102],pp118[103],pp118[104],pp118[105],pp118[106],pp118[107],pp118[108],pp118[109],pp118[110],pp118[111],pp118[112],pp118[113],pp118[114],pp118[115],pp118[116],pp118[117],pp118[118],pp118[119],pp118[120],pp118[121],pp118[122],pp118[123],pp118[124],pp118[125],pp118[126],pp118[127],pp118[128],pp118[129],pp118[130],pp118[131],pp118[132],pp118[133],pp118[134],pp118[135],pp118[136],pp118[137],pp118[138],pp118[139],pp118[140],pp118[141],pp118[142],pp118[143],pp118[144],pp118[145],pp118[146],pp118[147],pp118[148],pp118[149],pp118[150],pp118[151],pp118[152],pp118[153],pp118[154],pp118[155],pp118[156],pp118[157],pp118[158],pp118[159],pp118[160],pp118[161],pp118[162],pp118[163],pp118[164],pp118[165],pp118[166],pp118[167],pp118[168],pp118[169],pp118[170],pp118[171],pp118[172],pp118[173],pp118[174],pp118[175],pp118[176],pp118[177],pp118[178],pp118[179],pp118[180],pp118[181],pp118[182],pp118[183],pp118[184],pp118[185],pp118[186],pp118[187],pp118[188],pp118[189],pp118[190],pp118[191],pp118[192],pp118[193],pp118[194],pp118[195],pp118[196],pp118[197],pp118[198],pp118[199],pp118[200],pp118[201],pp118[202],pp118[203],pp118[204],pp118[205],pp118[206],pp118[207],pp118[208],pp118[209],pp118[210],pp118[211],pp118[212],pp118[213],pp118[214],pp118[215],pp118[216],pp118[217],pp118[218],pp118[219],pp118[220],pp118[221],pp118[222],pp118[223],pp118[224],pp118[225],pp118[226],pp118[227],pp118[228],pp118[229],pp118[230],pp118[231],pp118[232],pp118[233],pp118[234],pp118[235],pp118[236],pp118[237],pp119[237],pp120[237],pp121[237],pp122[237],pp123[237],pp124[237],pp125[237],pp126[237],pp127[237],pp128[237],pp129[237],pp130[237],pp131[237],pp132[237],pp133[237],pp134[237],pp135[237],pp136[237],pp137[237]};
    assign in10_2 = {pp29[108],pp29[109],pp29[110],pp29[111],pp29[112],pp29[113],pp29[114],pp29[115],pp29[116],pp29[117],pp29[118],pp29[119],pp29[120],pp29[121],pp29[122],pp29[123],pp29[124],pp29[125],pp29[126],pp29[127],pp29[128],pp29[129],pp29[130],pp29[131],pp29[132],pp29[133],pp29[134],pp29[135],pp29[136],pp29[137],pp29[138],pp29[139],pp29[140],pp29[141],pp29[142],pp29[143],pp29[144],pp29[145],pp29[146],pp29[147],pp29[148],pp29[149],pp29[150],pp29[151],pp29[152],pp29[153],pp29[154],pp29[155],pp29[156],pp29[157],pp29[158],pp29[159],pp29[160],pp29[161],pp29[162],pp29[163],pp29[164],pp29[165],pp29[166],pp29[167],pp29[168],pp29[169],pp29[170],pp28[172],pp27[174],pp26[176],pp25[178],pp24[180],pp23[182],pp22[184],pp21[186],pp20[188],pp19[190],pp18[192],pp17[194],pp16[196],pp15[198],pp14[200],pp13[202],pp12[204],pp11[206],pp10[208],pp119[100],pp119[101],pp119[102],pp119[103],pp119[104],pp119[105],pp119[106],pp119[107],pp119[108],pp119[109],pp119[110],pp119[111],pp119[112],pp119[113],pp119[114],pp119[115],pp119[116],pp119[117],pp119[118],pp119[119],pp119[120],pp119[121],pp119[122],pp119[123],pp119[124],pp119[125],pp119[126],pp119[127],pp119[128],pp119[129],pp119[130],pp119[131],pp119[132],pp119[133],pp119[134],pp119[135],pp119[136],pp119[137],pp119[138],pp119[139],pp119[140],pp119[141],pp119[142],pp119[143],pp119[144],pp119[145],pp119[146],pp119[147],pp119[148],pp119[149],pp119[150],pp119[151],pp119[152],pp119[153],pp119[154],pp119[155],pp119[156],pp119[157],pp119[158],pp119[159],pp119[160],pp119[161],pp119[162],pp119[163],pp119[164],pp119[165],pp119[166],pp119[167],pp119[168],pp119[169],pp119[170],pp119[171],pp119[172],pp119[173],pp119[174],pp119[175],pp119[176],pp119[177],pp119[178],pp119[179],pp119[180],pp119[181],pp119[182],pp119[183],pp119[184],pp119[185],pp119[186],pp119[187],pp119[188],pp119[189],pp119[190],pp119[191],pp119[192],pp119[193],pp119[194],pp119[195],pp119[196],pp119[197],pp119[198],pp119[199],pp119[200],pp119[201],pp119[202],pp119[203],pp119[204],pp119[205],pp119[206],pp119[207],pp119[208],pp119[209],pp119[210],pp119[211],pp119[212],pp119[213],pp119[214],pp119[215],pp119[216],pp119[217],pp119[218],pp119[219],pp119[220],pp119[221],pp119[222],pp119[223],pp119[224],pp119[225],pp119[226],pp119[227],pp119[228],pp119[229],pp119[230],pp119[231],pp119[232],pp119[233],pp119[234],pp119[235],pp119[236],pp120[236],pp121[236],pp122[236],pp123[236],pp124[236],pp125[236],pp126[236],pp127[236],pp128[236],pp129[236],pp130[236],pp131[236],pp132[236],pp133[236],pp134[236],pp135[236],pp136[236],pp137[236],pp138[236]};
    CLA_238 KS_10(s10, c10, in10_1, in10_2);
    wire[235:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp30[108],pp30[109],pp30[110],pp30[111],pp30[112],pp30[113],pp30[114],pp30[115],pp30[116],pp30[117],pp30[118],pp30[119],pp30[120],pp30[121],pp30[122],pp30[123],pp30[124],pp30[125],pp30[126],pp30[127],pp30[128],pp30[129],pp30[130],pp30[131],pp30[132],pp30[133],pp30[134],pp30[135],pp30[136],pp30[137],pp30[138],pp30[139],pp30[140],pp30[141],pp30[142],pp30[143],pp30[144],pp30[145],pp30[146],pp30[147],pp30[148],pp30[149],pp30[150],pp30[151],pp30[152],pp30[153],pp30[154],pp30[155],pp30[156],pp30[157],pp30[158],pp30[159],pp30[160],pp30[161],pp30[162],pp30[163],pp30[164],pp30[165],pp30[166],pp30[167],pp30[168],pp30[169],pp29[171],pp28[173],pp27[175],pp26[177],pp25[179],pp24[181],pp23[183],pp22[185],pp21[187],pp20[189],pp19[191],pp18[193],pp17[195],pp16[197],pp15[199],pp14[201],pp13[203],pp12[205],pp11[207],pp10[209],pp120[100],pp120[101],pp120[102],pp120[103],pp120[104],pp120[105],pp120[106],pp120[107],pp120[108],pp120[109],pp120[110],pp120[111],pp120[112],pp120[113],pp120[114],pp120[115],pp120[116],pp120[117],pp120[118],pp120[119],pp120[120],pp120[121],pp120[122],pp120[123],pp120[124],pp120[125],pp120[126],pp120[127],pp120[128],pp120[129],pp120[130],pp120[131],pp120[132],pp120[133],pp120[134],pp120[135],pp120[136],pp120[137],pp120[138],pp120[139],pp120[140],pp120[141],pp120[142],pp120[143],pp120[144],pp120[145],pp120[146],pp120[147],pp120[148],pp120[149],pp120[150],pp120[151],pp120[152],pp120[153],pp120[154],pp120[155],pp120[156],pp120[157],pp120[158],pp120[159],pp120[160],pp120[161],pp120[162],pp120[163],pp120[164],pp120[165],pp120[166],pp120[167],pp120[168],pp120[169],pp120[170],pp120[171],pp120[172],pp120[173],pp120[174],pp120[175],pp120[176],pp120[177],pp120[178],pp120[179],pp120[180],pp120[181],pp120[182],pp120[183],pp120[184],pp120[185],pp120[186],pp120[187],pp120[188],pp120[189],pp120[190],pp120[191],pp120[192],pp120[193],pp120[194],pp120[195],pp120[196],pp120[197],pp120[198],pp120[199],pp120[200],pp120[201],pp120[202],pp120[203],pp120[204],pp120[205],pp120[206],pp120[207],pp120[208],pp120[209],pp120[210],pp120[211],pp120[212],pp120[213],pp120[214],pp120[215],pp120[216],pp120[217],pp120[218],pp120[219],pp120[220],pp120[221],pp120[222],pp120[223],pp120[224],pp120[225],pp120[226],pp120[227],pp120[228],pp120[229],pp120[230],pp120[231],pp120[232],pp120[233],pp120[234],pp120[235],pp121[235],pp122[235],pp123[235],pp124[235],pp125[235],pp126[235],pp127[235],pp128[235],pp129[235],pp130[235],pp131[235],pp132[235],pp133[235],pp134[235],pp135[235],pp136[235],pp137[235],pp138[235]};
    assign in11_2 = {pp31[107],pp31[108],pp31[109],pp31[110],pp31[111],pp31[112],pp31[113],pp31[114],pp31[115],pp31[116],pp31[117],pp31[118],pp31[119],pp31[120],pp31[121],pp31[122],pp31[123],pp31[124],pp31[125],pp31[126],pp31[127],pp31[128],pp31[129],pp31[130],pp31[131],pp31[132],pp31[133],pp31[134],pp31[135],pp31[136],pp31[137],pp31[138],pp31[139],pp31[140],pp31[141],pp31[142],pp31[143],pp31[144],pp31[145],pp31[146],pp31[147],pp31[148],pp31[149],pp31[150],pp31[151],pp31[152],pp31[153],pp31[154],pp31[155],pp31[156],pp31[157],pp31[158],pp31[159],pp31[160],pp31[161],pp31[162],pp31[163],pp31[164],pp31[165],pp31[166],pp31[167],pp31[168],pp30[170],pp29[172],pp28[174],pp27[176],pp26[178],pp25[180],pp24[182],pp23[184],pp22[186],pp21[188],pp20[190],pp19[192],pp18[194],pp17[196],pp16[198],pp15[200],pp14[202],pp13[204],pp12[206],pp11[208],pp10[210],pp121[100],pp121[101],pp121[102],pp121[103],pp121[104],pp121[105],pp121[106],pp121[107],pp121[108],pp121[109],pp121[110],pp121[111],pp121[112],pp121[113],pp121[114],pp121[115],pp121[116],pp121[117],pp121[118],pp121[119],pp121[120],pp121[121],pp121[122],pp121[123],pp121[124],pp121[125],pp121[126],pp121[127],pp121[128],pp121[129],pp121[130],pp121[131],pp121[132],pp121[133],pp121[134],pp121[135],pp121[136],pp121[137],pp121[138],pp121[139],pp121[140],pp121[141],pp121[142],pp121[143],pp121[144],pp121[145],pp121[146],pp121[147],pp121[148],pp121[149],pp121[150],pp121[151],pp121[152],pp121[153],pp121[154],pp121[155],pp121[156],pp121[157],pp121[158],pp121[159],pp121[160],pp121[161],pp121[162],pp121[163],pp121[164],pp121[165],pp121[166],pp121[167],pp121[168],pp121[169],pp121[170],pp121[171],pp121[172],pp121[173],pp121[174],pp121[175],pp121[176],pp121[177],pp121[178],pp121[179],pp121[180],pp121[181],pp121[182],pp121[183],pp121[184],pp121[185],pp121[186],pp121[187],pp121[188],pp121[189],pp121[190],pp121[191],pp121[192],pp121[193],pp121[194],pp121[195],pp121[196],pp121[197],pp121[198],pp121[199],pp121[200],pp121[201],pp121[202],pp121[203],pp121[204],pp121[205],pp121[206],pp121[207],pp121[208],pp121[209],pp121[210],pp121[211],pp121[212],pp121[213],pp121[214],pp121[215],pp121[216],pp121[217],pp121[218],pp121[219],pp121[220],pp121[221],pp121[222],pp121[223],pp121[224],pp121[225],pp121[226],pp121[227],pp121[228],pp121[229],pp121[230],pp121[231],pp121[232],pp121[233],pp121[234],pp122[234],pp123[234],pp124[234],pp125[234],pp126[234],pp127[234],pp128[234],pp129[234],pp130[234],pp131[234],pp132[234],pp133[234],pp134[234],pp135[234],pp136[234],pp137[234],pp138[234],pp139[234]};
    CLA_236 KS_11(s11, c11, in11_1, in11_2);
    wire[233:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp32[107],pp32[108],pp32[109],pp32[110],pp32[111],pp32[112],pp32[113],pp32[114],pp32[115],pp32[116],pp32[117],pp32[118],pp32[119],pp32[120],pp32[121],pp32[122],pp32[123],pp32[124],pp32[125],pp32[126],pp32[127],pp32[128],pp32[129],pp32[130],pp32[131],pp32[132],pp32[133],pp32[134],pp32[135],pp32[136],pp32[137],pp32[138],pp32[139],pp32[140],pp32[141],pp32[142],pp32[143],pp32[144],pp32[145],pp32[146],pp32[147],pp32[148],pp32[149],pp32[150],pp32[151],pp32[152],pp32[153],pp32[154],pp32[155],pp32[156],pp32[157],pp32[158],pp32[159],pp32[160],pp32[161],pp32[162],pp32[163],pp32[164],pp32[165],pp32[166],pp32[167],pp31[169],pp30[171],pp29[173],pp28[175],pp27[177],pp26[179],pp25[181],pp24[183],pp23[185],pp22[187],pp21[189],pp20[191],pp19[193],pp18[195],pp17[197],pp16[199],pp15[201],pp14[203],pp13[205],pp12[207],pp11[209],pp10[211],pp122[100],pp122[101],pp122[102],pp122[103],pp122[104],pp122[105],pp122[106],pp122[107],pp122[108],pp122[109],pp122[110],pp122[111],pp122[112],pp122[113],pp122[114],pp122[115],pp122[116],pp122[117],pp122[118],pp122[119],pp122[120],pp122[121],pp122[122],pp122[123],pp122[124],pp122[125],pp122[126],pp122[127],pp122[128],pp122[129],pp122[130],pp122[131],pp122[132],pp122[133],pp122[134],pp122[135],pp122[136],pp122[137],pp122[138],pp122[139],pp122[140],pp122[141],pp122[142],pp122[143],pp122[144],pp122[145],pp122[146],pp122[147],pp122[148],pp122[149],pp122[150],pp122[151],pp122[152],pp122[153],pp122[154],pp122[155],pp122[156],pp122[157],pp122[158],pp122[159],pp122[160],pp122[161],pp122[162],pp122[163],pp122[164],pp122[165],pp122[166],pp122[167],pp122[168],pp122[169],pp122[170],pp122[171],pp122[172],pp122[173],pp122[174],pp122[175],pp122[176],pp122[177],pp122[178],pp122[179],pp122[180],pp122[181],pp122[182],pp122[183],pp122[184],pp122[185],pp122[186],pp122[187],pp122[188],pp122[189],pp122[190],pp122[191],pp122[192],pp122[193],pp122[194],pp122[195],pp122[196],pp122[197],pp122[198],pp122[199],pp122[200],pp122[201],pp122[202],pp122[203],pp122[204],pp122[205],pp122[206],pp122[207],pp122[208],pp122[209],pp122[210],pp122[211],pp122[212],pp122[213],pp122[214],pp122[215],pp122[216],pp122[217],pp122[218],pp122[219],pp122[220],pp122[221],pp122[222],pp122[223],pp122[224],pp122[225],pp122[226],pp122[227],pp122[228],pp122[229],pp122[230],pp122[231],pp122[232],pp122[233],pp123[233],pp124[233],pp125[233],pp126[233],pp127[233],pp128[233],pp129[233],pp130[233],pp131[233],pp132[233],pp133[233],pp134[233],pp135[233],pp136[233],pp137[233],pp138[233],pp139[233]};
    assign in12_2 = {pp33[106],pp33[107],pp33[108],pp33[109],pp33[110],pp33[111],pp33[112],pp33[113],pp33[114],pp33[115],pp33[116],pp33[117],pp33[118],pp33[119],pp33[120],pp33[121],pp33[122],pp33[123],pp33[124],pp33[125],pp33[126],pp33[127],pp33[128],pp33[129],pp33[130],pp33[131],pp33[132],pp33[133],pp33[134],pp33[135],pp33[136],pp33[137],pp33[138],pp33[139],pp33[140],pp33[141],pp33[142],pp33[143],pp33[144],pp33[145],pp33[146],pp33[147],pp33[148],pp33[149],pp33[150],pp33[151],pp33[152],pp33[153],pp33[154],pp33[155],pp33[156],pp33[157],pp33[158],pp33[159],pp33[160],pp33[161],pp33[162],pp33[163],pp33[164],pp33[165],pp33[166],pp32[168],pp31[170],pp30[172],pp29[174],pp28[176],pp27[178],pp26[180],pp25[182],pp24[184],pp23[186],pp22[188],pp21[190],pp20[192],pp19[194],pp18[196],pp17[198],pp16[200],pp15[202],pp14[204],pp13[206],pp12[208],pp11[210],pp10[212],pp123[100],pp123[101],pp123[102],pp123[103],pp123[104],pp123[105],pp123[106],pp123[107],pp123[108],pp123[109],pp123[110],pp123[111],pp123[112],pp123[113],pp123[114],pp123[115],pp123[116],pp123[117],pp123[118],pp123[119],pp123[120],pp123[121],pp123[122],pp123[123],pp123[124],pp123[125],pp123[126],pp123[127],pp123[128],pp123[129],pp123[130],pp123[131],pp123[132],pp123[133],pp123[134],pp123[135],pp123[136],pp123[137],pp123[138],pp123[139],pp123[140],pp123[141],pp123[142],pp123[143],pp123[144],pp123[145],pp123[146],pp123[147],pp123[148],pp123[149],pp123[150],pp123[151],pp123[152],pp123[153],pp123[154],pp123[155],pp123[156],pp123[157],pp123[158],pp123[159],pp123[160],pp123[161],pp123[162],pp123[163],pp123[164],pp123[165],pp123[166],pp123[167],pp123[168],pp123[169],pp123[170],pp123[171],pp123[172],pp123[173],pp123[174],pp123[175],pp123[176],pp123[177],pp123[178],pp123[179],pp123[180],pp123[181],pp123[182],pp123[183],pp123[184],pp123[185],pp123[186],pp123[187],pp123[188],pp123[189],pp123[190],pp123[191],pp123[192],pp123[193],pp123[194],pp123[195],pp123[196],pp123[197],pp123[198],pp123[199],pp123[200],pp123[201],pp123[202],pp123[203],pp123[204],pp123[205],pp123[206],pp123[207],pp123[208],pp123[209],pp123[210],pp123[211],pp123[212],pp123[213],pp123[214],pp123[215],pp123[216],pp123[217],pp123[218],pp123[219],pp123[220],pp123[221],pp123[222],pp123[223],pp123[224],pp123[225],pp123[226],pp123[227],pp123[228],pp123[229],pp123[230],pp123[231],pp123[232],pp124[232],pp125[232],pp126[232],pp127[232],pp128[232],pp129[232],pp130[232],pp131[232],pp132[232],pp133[232],pp134[232],pp135[232],pp136[232],pp137[232],pp138[232],pp139[232],pp140[232]};
    CLA_234 KS_12(s12, c12, in12_1, in12_2);
    wire[231:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp34[106],pp34[107],pp34[108],pp34[109],pp34[110],pp34[111],pp34[112],pp34[113],pp34[114],pp34[115],pp34[116],pp34[117],pp34[118],pp34[119],pp34[120],pp34[121],pp34[122],pp34[123],pp34[124],pp34[125],pp34[126],pp34[127],pp34[128],pp34[129],pp34[130],pp34[131],pp34[132],pp34[133],pp34[134],pp34[135],pp34[136],pp34[137],pp34[138],pp34[139],pp34[140],pp34[141],pp34[142],pp34[143],pp34[144],pp34[145],pp34[146],pp34[147],pp34[148],pp34[149],pp34[150],pp34[151],pp34[152],pp34[153],pp34[154],pp34[155],pp34[156],pp34[157],pp34[158],pp34[159],pp34[160],pp34[161],pp34[162],pp34[163],pp34[164],pp34[165],pp33[167],pp32[169],pp31[171],pp30[173],pp29[175],pp28[177],pp27[179],pp26[181],pp25[183],pp24[185],pp23[187],pp22[189],pp21[191],pp20[193],pp19[195],pp18[197],pp17[199],pp16[201],pp15[203],pp14[205],pp13[207],pp12[209],pp11[211],pp10[213],pp124[100],pp124[101],pp124[102],pp124[103],pp124[104],pp124[105],pp124[106],pp124[107],pp124[108],pp124[109],pp124[110],pp124[111],pp124[112],pp124[113],pp124[114],pp124[115],pp124[116],pp124[117],pp124[118],pp124[119],pp124[120],pp124[121],pp124[122],pp124[123],pp124[124],pp124[125],pp124[126],pp124[127],pp124[128],pp124[129],pp124[130],pp124[131],pp124[132],pp124[133],pp124[134],pp124[135],pp124[136],pp124[137],pp124[138],pp124[139],pp124[140],pp124[141],pp124[142],pp124[143],pp124[144],pp124[145],pp124[146],pp124[147],pp124[148],pp124[149],pp124[150],pp124[151],pp124[152],pp124[153],pp124[154],pp124[155],pp124[156],pp124[157],pp124[158],pp124[159],pp124[160],pp124[161],pp124[162],pp124[163],pp124[164],pp124[165],pp124[166],pp124[167],pp124[168],pp124[169],pp124[170],pp124[171],pp124[172],pp124[173],pp124[174],pp124[175],pp124[176],pp124[177],pp124[178],pp124[179],pp124[180],pp124[181],pp124[182],pp124[183],pp124[184],pp124[185],pp124[186],pp124[187],pp124[188],pp124[189],pp124[190],pp124[191],pp124[192],pp124[193],pp124[194],pp124[195],pp124[196],pp124[197],pp124[198],pp124[199],pp124[200],pp124[201],pp124[202],pp124[203],pp124[204],pp124[205],pp124[206],pp124[207],pp124[208],pp124[209],pp124[210],pp124[211],pp124[212],pp124[213],pp124[214],pp124[215],pp124[216],pp124[217],pp124[218],pp124[219],pp124[220],pp124[221],pp124[222],pp124[223],pp124[224],pp124[225],pp124[226],pp124[227],pp124[228],pp124[229],pp124[230],pp124[231],pp125[231],pp126[231],pp127[231],pp128[231],pp129[231],pp130[231],pp131[231],pp132[231],pp133[231],pp134[231],pp135[231],pp136[231],pp137[231],pp138[231],pp139[231],pp140[231]};
    assign in13_2 = {pp35[105],pp35[106],pp35[107],pp35[108],pp35[109],pp35[110],pp35[111],pp35[112],pp35[113],pp35[114],pp35[115],pp35[116],pp35[117],pp35[118],pp35[119],pp35[120],pp35[121],pp35[122],pp35[123],pp35[124],pp35[125],pp35[126],pp35[127],pp35[128],pp35[129],pp35[130],pp35[131],pp35[132],pp35[133],pp35[134],pp35[135],pp35[136],pp35[137],pp35[138],pp35[139],pp35[140],pp35[141],pp35[142],pp35[143],pp35[144],pp35[145],pp35[146],pp35[147],pp35[148],pp35[149],pp35[150],pp35[151],pp35[152],pp35[153],pp35[154],pp35[155],pp35[156],pp35[157],pp35[158],pp35[159],pp35[160],pp35[161],pp35[162],pp35[163],pp35[164],pp34[166],pp33[168],pp32[170],pp31[172],pp30[174],pp29[176],pp28[178],pp27[180],pp26[182],pp25[184],pp24[186],pp23[188],pp22[190],pp21[192],pp20[194],pp19[196],pp18[198],pp17[200],pp16[202],pp15[204],pp14[206],pp13[208],pp12[210],pp11[212],pp10[214],pp125[100],pp125[101],pp125[102],pp125[103],pp125[104],pp125[105],pp125[106],pp125[107],pp125[108],pp125[109],pp125[110],pp125[111],pp125[112],pp125[113],pp125[114],pp125[115],pp125[116],pp125[117],pp125[118],pp125[119],pp125[120],pp125[121],pp125[122],pp125[123],pp125[124],pp125[125],pp125[126],pp125[127],pp125[128],pp125[129],pp125[130],pp125[131],pp125[132],pp125[133],pp125[134],pp125[135],pp125[136],pp125[137],pp125[138],pp125[139],pp125[140],pp125[141],pp125[142],pp125[143],pp125[144],pp125[145],pp125[146],pp125[147],pp125[148],pp125[149],pp125[150],pp125[151],pp125[152],pp125[153],pp125[154],pp125[155],pp125[156],pp125[157],pp125[158],pp125[159],pp125[160],pp125[161],pp125[162],pp125[163],pp125[164],pp125[165],pp125[166],pp125[167],pp125[168],pp125[169],pp125[170],pp125[171],pp125[172],pp125[173],pp125[174],pp125[175],pp125[176],pp125[177],pp125[178],pp125[179],pp125[180],pp125[181],pp125[182],pp125[183],pp125[184],pp125[185],pp125[186],pp125[187],pp125[188],pp125[189],pp125[190],pp125[191],pp125[192],pp125[193],pp125[194],pp125[195],pp125[196],pp125[197],pp125[198],pp125[199],pp125[200],pp125[201],pp125[202],pp125[203],pp125[204],pp125[205],pp125[206],pp125[207],pp125[208],pp125[209],pp125[210],pp125[211],pp125[212],pp125[213],pp125[214],pp125[215],pp125[216],pp125[217],pp125[218],pp125[219],pp125[220],pp125[221],pp125[222],pp125[223],pp125[224],pp125[225],pp125[226],pp125[227],pp125[228],pp125[229],pp125[230],pp126[230],pp127[230],pp128[230],pp129[230],pp130[230],pp131[230],pp132[230],pp133[230],pp134[230],pp135[230],pp136[230],pp137[230],pp138[230],pp139[230],pp140[230],pp141[230]};
    CLA_232 KS_13(s13, c13, in13_1, in13_2);
    wire[229:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp36[105],pp36[106],pp36[107],pp36[108],pp36[109],pp36[110],pp36[111],pp36[112],pp36[113],pp36[114],pp36[115],pp36[116],pp36[117],pp36[118],pp36[119],pp36[120],pp36[121],pp36[122],pp36[123],pp36[124],pp36[125],pp36[126],pp36[127],pp36[128],pp36[129],pp36[130],pp36[131],pp36[132],pp36[133],pp36[134],pp36[135],pp36[136],pp36[137],pp36[138],pp36[139],pp36[140],pp36[141],pp36[142],pp36[143],pp36[144],pp36[145],pp36[146],pp36[147],pp36[148],pp36[149],pp36[150],pp36[151],pp36[152],pp36[153],pp36[154],pp36[155],pp36[156],pp36[157],pp36[158],pp36[159],pp36[160],pp36[161],pp36[162],pp36[163],pp35[165],pp34[167],pp33[169],pp32[171],pp31[173],pp30[175],pp29[177],pp28[179],pp27[181],pp26[183],pp25[185],pp24[187],pp23[189],pp22[191],pp21[193],pp20[195],pp19[197],pp18[199],pp17[201],pp16[203],pp15[205],pp14[207],pp13[209],pp12[211],pp11[213],pp10[215],pp126[100],pp126[101],pp126[102],pp126[103],pp126[104],pp126[105],pp126[106],pp126[107],pp126[108],pp126[109],pp126[110],pp126[111],pp126[112],pp126[113],pp126[114],pp126[115],pp126[116],pp126[117],pp126[118],pp126[119],pp126[120],pp126[121],pp126[122],pp126[123],pp126[124],pp126[125],pp126[126],pp126[127],pp126[128],pp126[129],pp126[130],pp126[131],pp126[132],pp126[133],pp126[134],pp126[135],pp126[136],pp126[137],pp126[138],pp126[139],pp126[140],pp126[141],pp126[142],pp126[143],pp126[144],pp126[145],pp126[146],pp126[147],pp126[148],pp126[149],pp126[150],pp126[151],pp126[152],pp126[153],pp126[154],pp126[155],pp126[156],pp126[157],pp126[158],pp126[159],pp126[160],pp126[161],pp126[162],pp126[163],pp126[164],pp126[165],pp126[166],pp126[167],pp126[168],pp126[169],pp126[170],pp126[171],pp126[172],pp126[173],pp126[174],pp126[175],pp126[176],pp126[177],pp126[178],pp126[179],pp126[180],pp126[181],pp126[182],pp126[183],pp126[184],pp126[185],pp126[186],pp126[187],pp126[188],pp126[189],pp126[190],pp126[191],pp126[192],pp126[193],pp126[194],pp126[195],pp126[196],pp126[197],pp126[198],pp126[199],pp126[200],pp126[201],pp126[202],pp126[203],pp126[204],pp126[205],pp126[206],pp126[207],pp126[208],pp126[209],pp126[210],pp126[211],pp126[212],pp126[213],pp126[214],pp126[215],pp126[216],pp126[217],pp126[218],pp126[219],pp126[220],pp126[221],pp126[222],pp126[223],pp126[224],pp126[225],pp126[226],pp126[227],pp126[228],pp126[229],pp127[229],pp128[229],pp129[229],pp130[229],pp131[229],pp132[229],pp133[229],pp134[229],pp135[229],pp136[229],pp137[229],pp138[229],pp139[229],pp140[229],pp141[229]};
    assign in14_2 = {pp37[104],pp37[105],pp37[106],pp37[107],pp37[108],pp37[109],pp37[110],pp37[111],pp37[112],pp37[113],pp37[114],pp37[115],pp37[116],pp37[117],pp37[118],pp37[119],pp37[120],pp37[121],pp37[122],pp37[123],pp37[124],pp37[125],pp37[126],pp37[127],pp37[128],pp37[129],pp37[130],pp37[131],pp37[132],pp37[133],pp37[134],pp37[135],pp37[136],pp37[137],pp37[138],pp37[139],pp37[140],pp37[141],pp37[142],pp37[143],pp37[144],pp37[145],pp37[146],pp37[147],pp37[148],pp37[149],pp37[150],pp37[151],pp37[152],pp37[153],pp37[154],pp37[155],pp37[156],pp37[157],pp37[158],pp37[159],pp37[160],pp37[161],pp37[162],pp36[164],pp35[166],pp34[168],pp33[170],pp32[172],pp31[174],pp30[176],pp29[178],pp28[180],pp27[182],pp26[184],pp25[186],pp24[188],pp23[190],pp22[192],pp21[194],pp20[196],pp19[198],pp18[200],pp17[202],pp16[204],pp15[206],pp14[208],pp13[210],pp12[212],pp11[214],pp10[216],pp127[100],pp127[101],pp127[102],pp127[103],pp127[104],pp127[105],pp127[106],pp127[107],pp127[108],pp127[109],pp127[110],pp127[111],pp127[112],pp127[113],pp127[114],pp127[115],pp127[116],pp127[117],pp127[118],pp127[119],pp127[120],pp127[121],pp127[122],pp127[123],pp127[124],pp127[125],pp127[126],pp127[127],pp127[128],pp127[129],pp127[130],pp127[131],pp127[132],pp127[133],pp127[134],pp127[135],pp127[136],pp127[137],pp127[138],pp127[139],pp127[140],pp127[141],pp127[142],pp127[143],pp127[144],pp127[145],pp127[146],pp127[147],pp127[148],pp127[149],pp127[150],pp127[151],pp127[152],pp127[153],pp127[154],pp127[155],pp127[156],pp127[157],pp127[158],pp127[159],pp127[160],pp127[161],pp127[162],pp127[163],pp127[164],pp127[165],pp127[166],pp127[167],pp127[168],pp127[169],pp127[170],pp127[171],pp127[172],pp127[173],pp127[174],pp127[175],pp127[176],pp127[177],pp127[178],pp127[179],pp127[180],pp127[181],pp127[182],pp127[183],pp127[184],pp127[185],pp127[186],pp127[187],pp127[188],pp127[189],pp127[190],pp127[191],pp127[192],pp127[193],pp127[194],pp127[195],pp127[196],pp127[197],pp127[198],pp127[199],pp127[200],pp127[201],pp127[202],pp127[203],pp127[204],pp127[205],pp127[206],pp127[207],pp127[208],pp127[209],pp127[210],pp127[211],pp127[212],pp127[213],pp127[214],pp127[215],pp127[216],pp127[217],pp127[218],pp127[219],pp127[220],pp127[221],pp127[222],pp127[223],pp127[224],pp127[225],pp127[226],pp127[227],pp127[228],pp128[228],pp129[228],pp130[228],pp131[228],pp132[228],pp133[228],pp134[228],pp135[228],pp136[228],pp137[228],pp138[228],pp139[228],pp140[228],pp141[228],pp142[228]};
    CLA_230 KS_14(s14, c14, in14_1, in14_2);
    wire[227:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp38[104],pp38[105],pp38[106],pp38[107],pp38[108],pp38[109],pp38[110],pp38[111],pp38[112],pp38[113],pp38[114],pp38[115],pp38[116],pp38[117],pp38[118],pp38[119],pp38[120],pp38[121],pp38[122],pp38[123],pp38[124],pp38[125],pp38[126],pp38[127],pp38[128],pp38[129],pp38[130],pp38[131],pp38[132],pp38[133],pp38[134],pp38[135],pp38[136],pp38[137],pp38[138],pp38[139],pp38[140],pp38[141],pp38[142],pp38[143],pp38[144],pp38[145],pp38[146],pp38[147],pp38[148],pp38[149],pp38[150],pp38[151],pp38[152],pp38[153],pp38[154],pp38[155],pp38[156],pp38[157],pp38[158],pp38[159],pp38[160],pp38[161],pp37[163],pp36[165],pp35[167],pp34[169],pp33[171],pp32[173],pp31[175],pp30[177],pp29[179],pp28[181],pp27[183],pp26[185],pp25[187],pp24[189],pp23[191],pp22[193],pp21[195],pp20[197],pp19[199],pp18[201],pp17[203],pp16[205],pp15[207],pp14[209],pp13[211],pp12[213],pp11[215],pp10[217],pp128[100],pp128[101],pp128[102],pp128[103],pp128[104],pp128[105],pp128[106],pp128[107],pp128[108],pp128[109],pp128[110],pp128[111],pp128[112],pp128[113],pp128[114],pp128[115],pp128[116],pp128[117],pp128[118],pp128[119],pp128[120],pp128[121],pp128[122],pp128[123],pp128[124],pp128[125],pp128[126],pp128[127],pp128[128],pp128[129],pp128[130],pp128[131],pp128[132],pp128[133],pp128[134],pp128[135],pp128[136],pp128[137],pp128[138],pp128[139],pp128[140],pp128[141],pp128[142],pp128[143],pp128[144],pp128[145],pp128[146],pp128[147],pp128[148],pp128[149],pp128[150],pp128[151],pp128[152],pp128[153],pp128[154],pp128[155],pp128[156],pp128[157],pp128[158],pp128[159],pp128[160],pp128[161],pp128[162],pp128[163],pp128[164],pp128[165],pp128[166],pp128[167],pp128[168],pp128[169],pp128[170],pp128[171],pp128[172],pp128[173],pp128[174],pp128[175],pp128[176],pp128[177],pp128[178],pp128[179],pp128[180],pp128[181],pp128[182],pp128[183],pp128[184],pp128[185],pp128[186],pp128[187],pp128[188],pp128[189],pp128[190],pp128[191],pp128[192],pp128[193],pp128[194],pp128[195],pp128[196],pp128[197],pp128[198],pp128[199],pp128[200],pp128[201],pp128[202],pp128[203],pp128[204],pp128[205],pp128[206],pp128[207],pp128[208],pp128[209],pp128[210],pp128[211],pp128[212],pp128[213],pp128[214],pp128[215],pp128[216],pp128[217],pp128[218],pp128[219],pp128[220],pp128[221],pp128[222],pp128[223],pp128[224],pp128[225],pp128[226],pp128[227],pp129[227],pp130[227],pp131[227],pp132[227],pp133[227],pp134[227],pp135[227],pp136[227],pp137[227],pp138[227],pp139[227],pp140[227],pp141[227],pp142[227]};
    assign in15_2 = {pp39[103],pp39[104],pp39[105],pp39[106],pp39[107],pp39[108],pp39[109],pp39[110],pp39[111],pp39[112],pp39[113],pp39[114],pp39[115],pp39[116],pp39[117],pp39[118],pp39[119],pp39[120],pp39[121],pp39[122],pp39[123],pp39[124],pp39[125],pp39[126],pp39[127],pp39[128],pp39[129],pp39[130],pp39[131],pp39[132],pp39[133],pp39[134],pp39[135],pp39[136],pp39[137],pp39[138],pp39[139],pp39[140],pp39[141],pp39[142],pp39[143],pp39[144],pp39[145],pp39[146],pp39[147],pp39[148],pp39[149],pp39[150],pp39[151],pp39[152],pp39[153],pp39[154],pp39[155],pp39[156],pp39[157],pp39[158],pp39[159],pp39[160],pp38[162],pp37[164],pp36[166],pp35[168],pp34[170],pp33[172],pp32[174],pp31[176],pp30[178],pp29[180],pp28[182],pp27[184],pp26[186],pp25[188],pp24[190],pp23[192],pp22[194],pp21[196],pp20[198],pp19[200],pp18[202],pp17[204],pp16[206],pp15[208],pp14[210],pp13[212],pp12[214],pp11[216],pp10[218],pp129[100],pp129[101],pp129[102],pp129[103],pp129[104],pp129[105],pp129[106],pp129[107],pp129[108],pp129[109],pp129[110],pp129[111],pp129[112],pp129[113],pp129[114],pp129[115],pp129[116],pp129[117],pp129[118],pp129[119],pp129[120],pp129[121],pp129[122],pp129[123],pp129[124],pp129[125],pp129[126],pp129[127],pp129[128],pp129[129],pp129[130],pp129[131],pp129[132],pp129[133],pp129[134],pp129[135],pp129[136],pp129[137],pp129[138],pp129[139],pp129[140],pp129[141],pp129[142],pp129[143],pp129[144],pp129[145],pp129[146],pp129[147],pp129[148],pp129[149],pp129[150],pp129[151],pp129[152],pp129[153],pp129[154],pp129[155],pp129[156],pp129[157],pp129[158],pp129[159],pp129[160],pp129[161],pp129[162],pp129[163],pp129[164],pp129[165],pp129[166],pp129[167],pp129[168],pp129[169],pp129[170],pp129[171],pp129[172],pp129[173],pp129[174],pp129[175],pp129[176],pp129[177],pp129[178],pp129[179],pp129[180],pp129[181],pp129[182],pp129[183],pp129[184],pp129[185],pp129[186],pp129[187],pp129[188],pp129[189],pp129[190],pp129[191],pp129[192],pp129[193],pp129[194],pp129[195],pp129[196],pp129[197],pp129[198],pp129[199],pp129[200],pp129[201],pp129[202],pp129[203],pp129[204],pp129[205],pp129[206],pp129[207],pp129[208],pp129[209],pp129[210],pp129[211],pp129[212],pp129[213],pp129[214],pp129[215],pp129[216],pp129[217],pp129[218],pp129[219],pp129[220],pp129[221],pp129[222],pp129[223],pp129[224],pp129[225],pp129[226],pp130[226],pp131[226],pp132[226],pp133[226],pp134[226],pp135[226],pp136[226],pp137[226],pp138[226],pp139[226],pp140[226],pp141[226],pp142[226],pp143[226]};
    CLA_228 KS_15(s15, c15, in15_1, in15_2);
    wire[225:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp40[103],pp40[104],pp40[105],pp40[106],pp40[107],pp40[108],pp40[109],pp40[110],pp40[111],pp40[112],pp40[113],pp40[114],pp40[115],pp40[116],pp40[117],pp40[118],pp40[119],pp40[120],pp40[121],pp40[122],pp40[123],pp40[124],pp40[125],pp40[126],pp40[127],pp40[128],pp40[129],pp40[130],pp40[131],pp40[132],pp40[133],pp40[134],pp40[135],pp40[136],pp40[137],pp40[138],pp40[139],pp40[140],pp40[141],pp40[142],pp40[143],pp40[144],pp40[145],pp40[146],pp40[147],pp40[148],pp40[149],pp40[150],pp40[151],pp40[152],pp40[153],pp40[154],pp40[155],pp40[156],pp40[157],pp40[158],pp40[159],pp39[161],pp38[163],pp37[165],pp36[167],pp35[169],pp34[171],pp33[173],pp32[175],pp31[177],pp30[179],pp29[181],pp28[183],pp27[185],pp26[187],pp25[189],pp24[191],pp23[193],pp22[195],pp21[197],pp20[199],pp19[201],pp18[203],pp17[205],pp16[207],pp15[209],pp14[211],pp13[213],pp12[215],pp11[217],pp10[219],pp130[100],pp130[101],pp130[102],pp130[103],pp130[104],pp130[105],pp130[106],pp130[107],pp130[108],pp130[109],pp130[110],pp130[111],pp130[112],pp130[113],pp130[114],pp130[115],pp130[116],pp130[117],pp130[118],pp130[119],pp130[120],pp130[121],pp130[122],pp130[123],pp130[124],pp130[125],pp130[126],pp130[127],pp130[128],pp130[129],pp130[130],pp130[131],pp130[132],pp130[133],pp130[134],pp130[135],pp130[136],pp130[137],pp130[138],pp130[139],pp130[140],pp130[141],pp130[142],pp130[143],pp130[144],pp130[145],pp130[146],pp130[147],pp130[148],pp130[149],pp130[150],pp130[151],pp130[152],pp130[153],pp130[154],pp130[155],pp130[156],pp130[157],pp130[158],pp130[159],pp130[160],pp130[161],pp130[162],pp130[163],pp130[164],pp130[165],pp130[166],pp130[167],pp130[168],pp130[169],pp130[170],pp130[171],pp130[172],pp130[173],pp130[174],pp130[175],pp130[176],pp130[177],pp130[178],pp130[179],pp130[180],pp130[181],pp130[182],pp130[183],pp130[184],pp130[185],pp130[186],pp130[187],pp130[188],pp130[189],pp130[190],pp130[191],pp130[192],pp130[193],pp130[194],pp130[195],pp130[196],pp130[197],pp130[198],pp130[199],pp130[200],pp130[201],pp130[202],pp130[203],pp130[204],pp130[205],pp130[206],pp130[207],pp130[208],pp130[209],pp130[210],pp130[211],pp130[212],pp130[213],pp130[214],pp130[215],pp130[216],pp130[217],pp130[218],pp130[219],pp130[220],pp130[221],pp130[222],pp130[223],pp130[224],pp130[225],pp131[225],pp132[225],pp133[225],pp134[225],pp135[225],pp136[225],pp137[225],pp138[225],pp139[225],pp140[225],pp141[225],pp142[225],pp143[225]};
    assign in16_2 = {pp41[102],pp41[103],pp41[104],pp41[105],pp41[106],pp41[107],pp41[108],pp41[109],pp41[110],pp41[111],pp41[112],pp41[113],pp41[114],pp41[115],pp41[116],pp41[117],pp41[118],pp41[119],pp41[120],pp41[121],pp41[122],pp41[123],pp41[124],pp41[125],pp41[126],pp41[127],pp41[128],pp41[129],pp41[130],pp41[131],pp41[132],pp41[133],pp41[134],pp41[135],pp41[136],pp41[137],pp41[138],pp41[139],pp41[140],pp41[141],pp41[142],pp41[143],pp41[144],pp41[145],pp41[146],pp41[147],pp41[148],pp41[149],pp41[150],pp41[151],pp41[152],pp41[153],pp41[154],pp41[155],pp41[156],pp41[157],pp41[158],pp40[160],pp39[162],pp38[164],pp37[166],pp36[168],pp35[170],pp34[172],pp33[174],pp32[176],pp31[178],pp30[180],pp29[182],pp28[184],pp27[186],pp26[188],pp25[190],pp24[192],pp23[194],pp22[196],pp21[198],pp20[200],pp19[202],pp18[204],pp17[206],pp16[208],pp15[210],pp14[212],pp13[214],pp12[216],pp11[218],pp10[220],pp131[100],pp131[101],pp131[102],pp131[103],pp131[104],pp131[105],pp131[106],pp131[107],pp131[108],pp131[109],pp131[110],pp131[111],pp131[112],pp131[113],pp131[114],pp131[115],pp131[116],pp131[117],pp131[118],pp131[119],pp131[120],pp131[121],pp131[122],pp131[123],pp131[124],pp131[125],pp131[126],pp131[127],pp131[128],pp131[129],pp131[130],pp131[131],pp131[132],pp131[133],pp131[134],pp131[135],pp131[136],pp131[137],pp131[138],pp131[139],pp131[140],pp131[141],pp131[142],pp131[143],pp131[144],pp131[145],pp131[146],pp131[147],pp131[148],pp131[149],pp131[150],pp131[151],pp131[152],pp131[153],pp131[154],pp131[155],pp131[156],pp131[157],pp131[158],pp131[159],pp131[160],pp131[161],pp131[162],pp131[163],pp131[164],pp131[165],pp131[166],pp131[167],pp131[168],pp131[169],pp131[170],pp131[171],pp131[172],pp131[173],pp131[174],pp131[175],pp131[176],pp131[177],pp131[178],pp131[179],pp131[180],pp131[181],pp131[182],pp131[183],pp131[184],pp131[185],pp131[186],pp131[187],pp131[188],pp131[189],pp131[190],pp131[191],pp131[192],pp131[193],pp131[194],pp131[195],pp131[196],pp131[197],pp131[198],pp131[199],pp131[200],pp131[201],pp131[202],pp131[203],pp131[204],pp131[205],pp131[206],pp131[207],pp131[208],pp131[209],pp131[210],pp131[211],pp131[212],pp131[213],pp131[214],pp131[215],pp131[216],pp131[217],pp131[218],pp131[219],pp131[220],pp131[221],pp131[222],pp131[223],pp131[224],pp132[224],pp133[224],pp134[224],pp135[224],pp136[224],pp137[224],pp138[224],pp139[224],pp140[224],pp141[224],pp142[224],pp143[224],pp144[224]};
    CLA_226 KS_16(s16, c16, in16_1, in16_2);
    wire[223:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp42[102],pp42[103],pp42[104],pp42[105],pp42[106],pp42[107],pp42[108],pp42[109],pp42[110],pp42[111],pp42[112],pp42[113],pp42[114],pp42[115],pp42[116],pp42[117],pp42[118],pp42[119],pp42[120],pp42[121],pp42[122],pp42[123],pp42[124],pp42[125],pp42[126],pp42[127],pp42[128],pp42[129],pp42[130],pp42[131],pp42[132],pp42[133],pp42[134],pp42[135],pp42[136],pp42[137],pp42[138],pp42[139],pp42[140],pp42[141],pp42[142],pp42[143],pp42[144],pp42[145],pp42[146],pp42[147],pp42[148],pp42[149],pp42[150],pp42[151],pp42[152],pp42[153],pp42[154],pp42[155],pp42[156],pp42[157],pp41[159],pp40[161],pp39[163],pp38[165],pp37[167],pp36[169],pp35[171],pp34[173],pp33[175],pp32[177],pp31[179],pp30[181],pp29[183],pp28[185],pp27[187],pp26[189],pp25[191],pp24[193],pp23[195],pp22[197],pp21[199],pp20[201],pp19[203],pp18[205],pp17[207],pp16[209],pp15[211],pp14[213],pp13[215],pp12[217],pp11[219],pp10[221],pp132[100],pp132[101],pp132[102],pp132[103],pp132[104],pp132[105],pp132[106],pp132[107],pp132[108],pp132[109],pp132[110],pp132[111],pp132[112],pp132[113],pp132[114],pp132[115],pp132[116],pp132[117],pp132[118],pp132[119],pp132[120],pp132[121],pp132[122],pp132[123],pp132[124],pp132[125],pp132[126],pp132[127],pp132[128],pp132[129],pp132[130],pp132[131],pp132[132],pp132[133],pp132[134],pp132[135],pp132[136],pp132[137],pp132[138],pp132[139],pp132[140],pp132[141],pp132[142],pp132[143],pp132[144],pp132[145],pp132[146],pp132[147],pp132[148],pp132[149],pp132[150],pp132[151],pp132[152],pp132[153],pp132[154],pp132[155],pp132[156],pp132[157],pp132[158],pp132[159],pp132[160],pp132[161],pp132[162],pp132[163],pp132[164],pp132[165],pp132[166],pp132[167],pp132[168],pp132[169],pp132[170],pp132[171],pp132[172],pp132[173],pp132[174],pp132[175],pp132[176],pp132[177],pp132[178],pp132[179],pp132[180],pp132[181],pp132[182],pp132[183],pp132[184],pp132[185],pp132[186],pp132[187],pp132[188],pp132[189],pp132[190],pp132[191],pp132[192],pp132[193],pp132[194],pp132[195],pp132[196],pp132[197],pp132[198],pp132[199],pp132[200],pp132[201],pp132[202],pp132[203],pp132[204],pp132[205],pp132[206],pp132[207],pp132[208],pp132[209],pp132[210],pp132[211],pp132[212],pp132[213],pp132[214],pp132[215],pp132[216],pp132[217],pp132[218],pp132[219],pp132[220],pp132[221],pp132[222],pp132[223],pp133[223],pp134[223],pp135[223],pp136[223],pp137[223],pp138[223],pp139[223],pp140[223],pp141[223],pp142[223],pp143[223],pp144[223]};
    assign in17_2 = {pp43[101],pp43[102],pp43[103],pp43[104],pp43[105],pp43[106],pp43[107],pp43[108],pp43[109],pp43[110],pp43[111],pp43[112],pp43[113],pp43[114],pp43[115],pp43[116],pp43[117],pp43[118],pp43[119],pp43[120],pp43[121],pp43[122],pp43[123],pp43[124],pp43[125],pp43[126],pp43[127],pp43[128],pp43[129],pp43[130],pp43[131],pp43[132],pp43[133],pp43[134],pp43[135],pp43[136],pp43[137],pp43[138],pp43[139],pp43[140],pp43[141],pp43[142],pp43[143],pp43[144],pp43[145],pp43[146],pp43[147],pp43[148],pp43[149],pp43[150],pp43[151],pp43[152],pp43[153],pp43[154],pp43[155],pp43[156],pp42[158],pp41[160],pp40[162],pp39[164],pp38[166],pp37[168],pp36[170],pp35[172],pp34[174],pp33[176],pp32[178],pp31[180],pp30[182],pp29[184],pp28[186],pp27[188],pp26[190],pp25[192],pp24[194],pp23[196],pp22[198],pp21[200],pp20[202],pp19[204],pp18[206],pp17[208],pp16[210],pp15[212],pp14[214],pp13[216],pp12[218],pp11[220],pp10[222],pp133[100],pp133[101],pp133[102],pp133[103],pp133[104],pp133[105],pp133[106],pp133[107],pp133[108],pp133[109],pp133[110],pp133[111],pp133[112],pp133[113],pp133[114],pp133[115],pp133[116],pp133[117],pp133[118],pp133[119],pp133[120],pp133[121],pp133[122],pp133[123],pp133[124],pp133[125],pp133[126],pp133[127],pp133[128],pp133[129],pp133[130],pp133[131],pp133[132],pp133[133],pp133[134],pp133[135],pp133[136],pp133[137],pp133[138],pp133[139],pp133[140],pp133[141],pp133[142],pp133[143],pp133[144],pp133[145],pp133[146],pp133[147],pp133[148],pp133[149],pp133[150],pp133[151],pp133[152],pp133[153],pp133[154],pp133[155],pp133[156],pp133[157],pp133[158],pp133[159],pp133[160],pp133[161],pp133[162],pp133[163],pp133[164],pp133[165],pp133[166],pp133[167],pp133[168],pp133[169],pp133[170],pp133[171],pp133[172],pp133[173],pp133[174],pp133[175],pp133[176],pp133[177],pp133[178],pp133[179],pp133[180],pp133[181],pp133[182],pp133[183],pp133[184],pp133[185],pp133[186],pp133[187],pp133[188],pp133[189],pp133[190],pp133[191],pp133[192],pp133[193],pp133[194],pp133[195],pp133[196],pp133[197],pp133[198],pp133[199],pp133[200],pp133[201],pp133[202],pp133[203],pp133[204],pp133[205],pp133[206],pp133[207],pp133[208],pp133[209],pp133[210],pp133[211],pp133[212],pp133[213],pp133[214],pp133[215],pp133[216],pp133[217],pp133[218],pp133[219],pp133[220],pp133[221],pp133[222],pp134[222],pp135[222],pp136[222],pp137[222],pp138[222],pp139[222],pp140[222],pp141[222],pp142[222],pp143[222],pp144[222],pp145[222]};
    CLA_224 KS_17(s17, c17, in17_1, in17_2);
    wire[221:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp44[101],pp44[102],pp44[103],pp44[104],pp44[105],pp44[106],pp44[107],pp44[108],pp44[109],pp44[110],pp44[111],pp44[112],pp44[113],pp44[114],pp44[115],pp44[116],pp44[117],pp44[118],pp44[119],pp44[120],pp44[121],pp44[122],pp44[123],pp44[124],pp44[125],pp44[126],pp44[127],pp44[128],pp44[129],pp44[130],pp44[131],pp44[132],pp44[133],pp44[134],pp44[135],pp44[136],pp44[137],pp44[138],pp44[139],pp44[140],pp44[141],pp44[142],pp44[143],pp44[144],pp44[145],pp44[146],pp44[147],pp44[148],pp44[149],pp44[150],pp44[151],pp44[152],pp44[153],pp44[154],pp44[155],pp43[157],pp42[159],pp41[161],pp40[163],pp39[165],pp38[167],pp37[169],pp36[171],pp35[173],pp34[175],pp33[177],pp32[179],pp31[181],pp30[183],pp29[185],pp28[187],pp27[189],pp26[191],pp25[193],pp24[195],pp23[197],pp22[199],pp21[201],pp20[203],pp19[205],pp18[207],pp17[209],pp16[211],pp15[213],pp14[215],pp13[217],pp12[219],pp11[221],pp10[223],pp134[100],pp134[101],pp134[102],pp134[103],pp134[104],pp134[105],pp134[106],pp134[107],pp134[108],pp134[109],pp134[110],pp134[111],pp134[112],pp134[113],pp134[114],pp134[115],pp134[116],pp134[117],pp134[118],pp134[119],pp134[120],pp134[121],pp134[122],pp134[123],pp134[124],pp134[125],pp134[126],pp134[127],pp134[128],pp134[129],pp134[130],pp134[131],pp134[132],pp134[133],pp134[134],pp134[135],pp134[136],pp134[137],pp134[138],pp134[139],pp134[140],pp134[141],pp134[142],pp134[143],pp134[144],pp134[145],pp134[146],pp134[147],pp134[148],pp134[149],pp134[150],pp134[151],pp134[152],pp134[153],pp134[154],pp134[155],pp134[156],pp134[157],pp134[158],pp134[159],pp134[160],pp134[161],pp134[162],pp134[163],pp134[164],pp134[165],pp134[166],pp134[167],pp134[168],pp134[169],pp134[170],pp134[171],pp134[172],pp134[173],pp134[174],pp134[175],pp134[176],pp134[177],pp134[178],pp134[179],pp134[180],pp134[181],pp134[182],pp134[183],pp134[184],pp134[185],pp134[186],pp134[187],pp134[188],pp134[189],pp134[190],pp134[191],pp134[192],pp134[193],pp134[194],pp134[195],pp134[196],pp134[197],pp134[198],pp134[199],pp134[200],pp134[201],pp134[202],pp134[203],pp134[204],pp134[205],pp134[206],pp134[207],pp134[208],pp134[209],pp134[210],pp134[211],pp134[212],pp134[213],pp134[214],pp134[215],pp134[216],pp134[217],pp134[218],pp134[219],pp134[220],pp134[221],pp135[221],pp136[221],pp137[221],pp138[221],pp139[221],pp140[221],pp141[221],pp142[221],pp143[221],pp144[221],pp145[221]};
    assign in18_2 = {pp45[100],pp45[101],pp45[102],pp45[103],pp45[104],pp45[105],pp45[106],pp45[107],pp45[108],pp45[109],pp45[110],pp45[111],pp45[112],pp45[113],pp45[114],pp45[115],pp45[116],pp45[117],pp45[118],pp45[119],pp45[120],pp45[121],pp45[122],pp45[123],pp45[124],pp45[125],pp45[126],pp45[127],pp45[128],pp45[129],pp45[130],pp45[131],pp45[132],pp45[133],pp45[134],pp45[135],pp45[136],pp45[137],pp45[138],pp45[139],pp45[140],pp45[141],pp45[142],pp45[143],pp45[144],pp45[145],pp45[146],pp45[147],pp45[148],pp45[149],pp45[150],pp45[151],pp45[152],pp45[153],pp45[154],pp44[156],pp43[158],pp42[160],pp41[162],pp40[164],pp39[166],pp38[168],pp37[170],pp36[172],pp35[174],pp34[176],pp33[178],pp32[180],pp31[182],pp30[184],pp29[186],pp28[188],pp27[190],pp26[192],pp25[194],pp24[196],pp23[198],pp22[200],pp21[202],pp20[204],pp19[206],pp18[208],pp17[210],pp16[212],pp15[214],pp14[216],pp13[218],pp12[220],pp11[222],pp10[224],pp135[100],pp135[101],pp135[102],pp135[103],pp135[104],pp135[105],pp135[106],pp135[107],pp135[108],pp135[109],pp135[110],pp135[111],pp135[112],pp135[113],pp135[114],pp135[115],pp135[116],pp135[117],pp135[118],pp135[119],pp135[120],pp135[121],pp135[122],pp135[123],pp135[124],pp135[125],pp135[126],pp135[127],pp135[128],pp135[129],pp135[130],pp135[131],pp135[132],pp135[133],pp135[134],pp135[135],pp135[136],pp135[137],pp135[138],pp135[139],pp135[140],pp135[141],pp135[142],pp135[143],pp135[144],pp135[145],pp135[146],pp135[147],pp135[148],pp135[149],pp135[150],pp135[151],pp135[152],pp135[153],pp135[154],pp135[155],pp135[156],pp135[157],pp135[158],pp135[159],pp135[160],pp135[161],pp135[162],pp135[163],pp135[164],pp135[165],pp135[166],pp135[167],pp135[168],pp135[169],pp135[170],pp135[171],pp135[172],pp135[173],pp135[174],pp135[175],pp135[176],pp135[177],pp135[178],pp135[179],pp135[180],pp135[181],pp135[182],pp135[183],pp135[184],pp135[185],pp135[186],pp135[187],pp135[188],pp135[189],pp135[190],pp135[191],pp135[192],pp135[193],pp135[194],pp135[195],pp135[196],pp135[197],pp135[198],pp135[199],pp135[200],pp135[201],pp135[202],pp135[203],pp135[204],pp135[205],pp135[206],pp135[207],pp135[208],pp135[209],pp135[210],pp135[211],pp135[212],pp135[213],pp135[214],pp135[215],pp135[216],pp135[217],pp135[218],pp135[219],pp135[220],pp136[220],pp137[220],pp138[220],pp139[220],pp140[220],pp141[220],pp142[220],pp143[220],pp144[220],pp145[220],pp146[220]};
    CLA_222 KS_18(s18, c18, in18_1, in18_2);
    wire[219:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp46[100],pp46[101],pp46[102],pp46[103],pp46[104],pp46[105],pp46[106],pp46[107],pp46[108],pp46[109],pp46[110],pp46[111],pp46[112],pp46[113],pp46[114],pp46[115],pp46[116],pp46[117],pp46[118],pp46[119],pp46[120],pp46[121],pp46[122],pp46[123],pp46[124],pp46[125],pp46[126],pp46[127],pp46[128],pp46[129],pp46[130],pp46[131],pp46[132],pp46[133],pp46[134],pp46[135],pp46[136],pp46[137],pp46[138],pp46[139],pp46[140],pp46[141],pp46[142],pp46[143],pp46[144],pp46[145],pp46[146],pp46[147],pp46[148],pp46[149],pp46[150],pp46[151],pp46[152],pp46[153],pp45[155],pp44[157],pp43[159],pp42[161],pp41[163],pp40[165],pp39[167],pp38[169],pp37[171],pp36[173],pp35[175],pp34[177],pp33[179],pp32[181],pp31[183],pp30[185],pp29[187],pp28[189],pp27[191],pp26[193],pp25[195],pp24[197],pp23[199],pp22[201],pp21[203],pp20[205],pp19[207],pp18[209],pp17[211],pp16[213],pp15[215],pp14[217],pp13[219],pp12[221],pp11[223],pp10[225],pp136[100],pp136[101],pp136[102],pp136[103],pp136[104],pp136[105],pp136[106],pp136[107],pp136[108],pp136[109],pp136[110],pp136[111],pp136[112],pp136[113],pp136[114],pp136[115],pp136[116],pp136[117],pp136[118],pp136[119],pp136[120],pp136[121],pp136[122],pp136[123],pp136[124],pp136[125],pp136[126],pp136[127],pp136[128],pp136[129],pp136[130],pp136[131],pp136[132],pp136[133],pp136[134],pp136[135],pp136[136],pp136[137],pp136[138],pp136[139],pp136[140],pp136[141],pp136[142],pp136[143],pp136[144],pp136[145],pp136[146],pp136[147],pp136[148],pp136[149],pp136[150],pp136[151],pp136[152],pp136[153],pp136[154],pp136[155],pp136[156],pp136[157],pp136[158],pp136[159],pp136[160],pp136[161],pp136[162],pp136[163],pp136[164],pp136[165],pp136[166],pp136[167],pp136[168],pp136[169],pp136[170],pp136[171],pp136[172],pp136[173],pp136[174],pp136[175],pp136[176],pp136[177],pp136[178],pp136[179],pp136[180],pp136[181],pp136[182],pp136[183],pp136[184],pp136[185],pp136[186],pp136[187],pp136[188],pp136[189],pp136[190],pp136[191],pp136[192],pp136[193],pp136[194],pp136[195],pp136[196],pp136[197],pp136[198],pp136[199],pp136[200],pp136[201],pp136[202],pp136[203],pp136[204],pp136[205],pp136[206],pp136[207],pp136[208],pp136[209],pp136[210],pp136[211],pp136[212],pp136[213],pp136[214],pp136[215],pp136[216],pp136[217],pp136[218],pp136[219],pp137[219],pp138[219],pp139[219],pp140[219],pp141[219],pp142[219],pp143[219],pp144[219],pp145[219],pp146[219]};
    assign in19_2 = {pp100[46],pp47[100],pp47[101],pp47[102],pp47[103],pp47[104],pp47[105],pp47[106],pp47[107],pp47[108],pp47[109],pp47[110],pp47[111],pp47[112],pp47[113],pp47[114],pp47[115],pp47[116],pp47[117],pp47[118],pp47[119],pp47[120],pp47[121],pp47[122],pp47[123],pp47[124],pp47[125],pp47[126],pp47[127],pp47[128],pp47[129],pp47[130],pp47[131],pp47[132],pp47[133],pp47[134],pp47[135],pp47[136],pp47[137],pp47[138],pp47[139],pp47[140],pp47[141],pp47[142],pp47[143],pp47[144],pp47[145],pp47[146],pp47[147],pp47[148],pp47[149],pp47[150],pp47[151],pp47[152],pp46[154],pp45[156],pp44[158],pp43[160],pp42[162],pp41[164],pp40[166],pp39[168],pp38[170],pp37[172],pp36[174],pp35[176],pp34[178],pp33[180],pp32[182],pp31[184],pp30[186],pp29[188],pp28[190],pp27[192],pp26[194],pp25[196],pp24[198],pp23[200],pp22[202],pp21[204],pp20[206],pp19[208],pp18[210],pp17[212],pp16[214],pp15[216],pp14[218],pp13[220],pp12[222],pp11[224],pp10[226],pp137[100],pp137[101],pp137[102],pp137[103],pp137[104],pp137[105],pp137[106],pp137[107],pp137[108],pp137[109],pp137[110],pp137[111],pp137[112],pp137[113],pp137[114],pp137[115],pp137[116],pp137[117],pp137[118],pp137[119],pp137[120],pp137[121],pp137[122],pp137[123],pp137[124],pp137[125],pp137[126],pp137[127],pp137[128],pp137[129],pp137[130],pp137[131],pp137[132],pp137[133],pp137[134],pp137[135],pp137[136],pp137[137],pp137[138],pp137[139],pp137[140],pp137[141],pp137[142],pp137[143],pp137[144],pp137[145],pp137[146],pp137[147],pp137[148],pp137[149],pp137[150],pp137[151],pp137[152],pp137[153],pp137[154],pp137[155],pp137[156],pp137[157],pp137[158],pp137[159],pp137[160],pp137[161],pp137[162],pp137[163],pp137[164],pp137[165],pp137[166],pp137[167],pp137[168],pp137[169],pp137[170],pp137[171],pp137[172],pp137[173],pp137[174],pp137[175],pp137[176],pp137[177],pp137[178],pp137[179],pp137[180],pp137[181],pp137[182],pp137[183],pp137[184],pp137[185],pp137[186],pp137[187],pp137[188],pp137[189],pp137[190],pp137[191],pp137[192],pp137[193],pp137[194],pp137[195],pp137[196],pp137[197],pp137[198],pp137[199],pp137[200],pp137[201],pp137[202],pp137[203],pp137[204],pp137[205],pp137[206],pp137[207],pp137[208],pp137[209],pp137[210],pp137[211],pp137[212],pp137[213],pp137[214],pp137[215],pp137[216],pp137[217],pp137[218],pp138[218],pp139[218],pp140[218],pp141[218],pp142[218],pp143[218],pp144[218],pp145[218],pp146[218],pp147[218]};
    CLA_220 KS_19(s19, c19, in19_1, in19_2);
    wire[217:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp100[47],pp48[100],pp48[101],pp48[102],pp48[103],pp48[104],pp48[105],pp48[106],pp48[107],pp48[108],pp48[109],pp48[110],pp48[111],pp48[112],pp48[113],pp48[114],pp48[115],pp48[116],pp48[117],pp48[118],pp48[119],pp48[120],pp48[121],pp48[122],pp48[123],pp48[124],pp48[125],pp48[126],pp48[127],pp48[128],pp48[129],pp48[130],pp48[131],pp48[132],pp48[133],pp48[134],pp48[135],pp48[136],pp48[137],pp48[138],pp48[139],pp48[140],pp48[141],pp48[142],pp48[143],pp48[144],pp48[145],pp48[146],pp48[147],pp48[148],pp48[149],pp48[150],pp48[151],pp47[153],pp46[155],pp45[157],pp44[159],pp43[161],pp42[163],pp41[165],pp40[167],pp39[169],pp38[171],pp37[173],pp36[175],pp35[177],pp34[179],pp33[181],pp32[183],pp31[185],pp30[187],pp29[189],pp28[191],pp27[193],pp26[195],pp25[197],pp24[199],pp23[201],pp22[203],pp21[205],pp20[207],pp19[209],pp18[211],pp17[213],pp16[215],pp15[217],pp14[219],pp13[221],pp12[223],pp11[225],pp10[227],pp138[100],pp138[101],pp138[102],pp138[103],pp138[104],pp138[105],pp138[106],pp138[107],pp138[108],pp138[109],pp138[110],pp138[111],pp138[112],pp138[113],pp138[114],pp138[115],pp138[116],pp138[117],pp138[118],pp138[119],pp138[120],pp138[121],pp138[122],pp138[123],pp138[124],pp138[125],pp138[126],pp138[127],pp138[128],pp138[129],pp138[130],pp138[131],pp138[132],pp138[133],pp138[134],pp138[135],pp138[136],pp138[137],pp138[138],pp138[139],pp138[140],pp138[141],pp138[142],pp138[143],pp138[144],pp138[145],pp138[146],pp138[147],pp138[148],pp138[149],pp138[150],pp138[151],pp138[152],pp138[153],pp138[154],pp138[155],pp138[156],pp138[157],pp138[158],pp138[159],pp138[160],pp138[161],pp138[162],pp138[163],pp138[164],pp138[165],pp138[166],pp138[167],pp138[168],pp138[169],pp138[170],pp138[171],pp138[172],pp138[173],pp138[174],pp138[175],pp138[176],pp138[177],pp138[178],pp138[179],pp138[180],pp138[181],pp138[182],pp138[183],pp138[184],pp138[185],pp138[186],pp138[187],pp138[188],pp138[189],pp138[190],pp138[191],pp138[192],pp138[193],pp138[194],pp138[195],pp138[196],pp138[197],pp138[198],pp138[199],pp138[200],pp138[201],pp138[202],pp138[203],pp138[204],pp138[205],pp138[206],pp138[207],pp138[208],pp138[209],pp138[210],pp138[211],pp138[212],pp138[213],pp138[214],pp138[215],pp138[216],pp138[217],pp139[217],pp140[217],pp141[217],pp142[217],pp143[217],pp144[217],pp145[217],pp146[217],pp147[217]};
    assign in20_2 = {pp101[46],pp100[48],pp49[100],pp49[101],pp49[102],pp49[103],pp49[104],pp49[105],pp49[106],pp49[107],pp49[108],pp49[109],pp49[110],pp49[111],pp49[112],pp49[113],pp49[114],pp49[115],pp49[116],pp49[117],pp49[118],pp49[119],pp49[120],pp49[121],pp49[122],pp49[123],pp49[124],pp49[125],pp49[126],pp49[127],pp49[128],pp49[129],pp49[130],pp49[131],pp49[132],pp49[133],pp49[134],pp49[135],pp49[136],pp49[137],pp49[138],pp49[139],pp49[140],pp49[141],pp49[142],pp49[143],pp49[144],pp49[145],pp49[146],pp49[147],pp49[148],pp49[149],pp49[150],pp48[152],pp47[154],pp46[156],pp45[158],pp44[160],pp43[162],pp42[164],pp41[166],pp40[168],pp39[170],pp38[172],pp37[174],pp36[176],pp35[178],pp34[180],pp33[182],pp32[184],pp31[186],pp30[188],pp29[190],pp28[192],pp27[194],pp26[196],pp25[198],pp24[200],pp23[202],pp22[204],pp21[206],pp20[208],pp19[210],pp18[212],pp17[214],pp16[216],pp15[218],pp14[220],pp13[222],pp12[224],pp11[226],pp10[228],pp139[100],pp139[101],pp139[102],pp139[103],pp139[104],pp139[105],pp139[106],pp139[107],pp139[108],pp139[109],pp139[110],pp139[111],pp139[112],pp139[113],pp139[114],pp139[115],pp139[116],pp139[117],pp139[118],pp139[119],pp139[120],pp139[121],pp139[122],pp139[123],pp139[124],pp139[125],pp139[126],pp139[127],pp139[128],pp139[129],pp139[130],pp139[131],pp139[132],pp139[133],pp139[134],pp139[135],pp139[136],pp139[137],pp139[138],pp139[139],pp139[140],pp139[141],pp139[142],pp139[143],pp139[144],pp139[145],pp139[146],pp139[147],pp139[148],pp139[149],pp139[150],pp139[151],pp139[152],pp139[153],pp139[154],pp139[155],pp139[156],pp139[157],pp139[158],pp139[159],pp139[160],pp139[161],pp139[162],pp139[163],pp139[164],pp139[165],pp139[166],pp139[167],pp139[168],pp139[169],pp139[170],pp139[171],pp139[172],pp139[173],pp139[174],pp139[175],pp139[176],pp139[177],pp139[178],pp139[179],pp139[180],pp139[181],pp139[182],pp139[183],pp139[184],pp139[185],pp139[186],pp139[187],pp139[188],pp139[189],pp139[190],pp139[191],pp139[192],pp139[193],pp139[194],pp139[195],pp139[196],pp139[197],pp139[198],pp139[199],pp139[200],pp139[201],pp139[202],pp139[203],pp139[204],pp139[205],pp139[206],pp139[207],pp139[208],pp139[209],pp139[210],pp139[211],pp139[212],pp139[213],pp139[214],pp139[215],pp139[216],pp140[216],pp141[216],pp142[216],pp143[216],pp144[216],pp145[216],pp146[216],pp147[216],pp148[216]};
    CLA_218 KS_20(s20, c20, in20_1, in20_2);
    wire[215:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp101[47],pp100[49],pp50[100],pp50[101],pp50[102],pp50[103],pp50[104],pp50[105],pp50[106],pp50[107],pp50[108],pp50[109],pp50[110],pp50[111],pp50[112],pp50[113],pp50[114],pp50[115],pp50[116],pp50[117],pp50[118],pp50[119],pp50[120],pp50[121],pp50[122],pp50[123],pp50[124],pp50[125],pp50[126],pp50[127],pp50[128],pp50[129],pp50[130],pp50[131],pp50[132],pp50[133],pp50[134],pp50[135],pp50[136],pp50[137],pp50[138],pp50[139],pp50[140],pp50[141],pp50[142],pp50[143],pp50[144],pp50[145],pp50[146],pp50[147],pp50[148],pp50[149],pp49[151],pp48[153],pp47[155],pp46[157],pp45[159],pp44[161],pp43[163],pp42[165],pp41[167],pp40[169],pp39[171],pp38[173],pp37[175],pp36[177],pp35[179],pp34[181],pp33[183],pp32[185],pp31[187],pp30[189],pp29[191],pp28[193],pp27[195],pp26[197],pp25[199],pp24[201],pp23[203],pp22[205],pp21[207],pp20[209],pp19[211],pp18[213],pp17[215],pp16[217],pp15[219],pp14[221],pp13[223],pp12[225],pp11[227],pp10[229],pp140[100],pp140[101],pp140[102],pp140[103],pp140[104],pp140[105],pp140[106],pp140[107],pp140[108],pp140[109],pp140[110],pp140[111],pp140[112],pp140[113],pp140[114],pp140[115],pp140[116],pp140[117],pp140[118],pp140[119],pp140[120],pp140[121],pp140[122],pp140[123],pp140[124],pp140[125],pp140[126],pp140[127],pp140[128],pp140[129],pp140[130],pp140[131],pp140[132],pp140[133],pp140[134],pp140[135],pp140[136],pp140[137],pp140[138],pp140[139],pp140[140],pp140[141],pp140[142],pp140[143],pp140[144],pp140[145],pp140[146],pp140[147],pp140[148],pp140[149],pp140[150],pp140[151],pp140[152],pp140[153],pp140[154],pp140[155],pp140[156],pp140[157],pp140[158],pp140[159],pp140[160],pp140[161],pp140[162],pp140[163],pp140[164],pp140[165],pp140[166],pp140[167],pp140[168],pp140[169],pp140[170],pp140[171],pp140[172],pp140[173],pp140[174],pp140[175],pp140[176],pp140[177],pp140[178],pp140[179],pp140[180],pp140[181],pp140[182],pp140[183],pp140[184],pp140[185],pp140[186],pp140[187],pp140[188],pp140[189],pp140[190],pp140[191],pp140[192],pp140[193],pp140[194],pp140[195],pp140[196],pp140[197],pp140[198],pp140[199],pp140[200],pp140[201],pp140[202],pp140[203],pp140[204],pp140[205],pp140[206],pp140[207],pp140[208],pp140[209],pp140[210],pp140[211],pp140[212],pp140[213],pp140[214],pp140[215],pp141[215],pp142[215],pp143[215],pp144[215],pp145[215],pp146[215],pp147[215],pp148[215]};
    assign in21_2 = {pp102[46],pp101[48],pp100[50],pp51[100],pp51[101],pp51[102],pp51[103],pp51[104],pp51[105],pp51[106],pp51[107],pp51[108],pp51[109],pp51[110],pp51[111],pp51[112],pp51[113],pp51[114],pp51[115],pp51[116],pp51[117],pp51[118],pp51[119],pp51[120],pp51[121],pp51[122],pp51[123],pp51[124],pp51[125],pp51[126],pp51[127],pp51[128],pp51[129],pp51[130],pp51[131],pp51[132],pp51[133],pp51[134],pp51[135],pp51[136],pp51[137],pp51[138],pp51[139],pp51[140],pp51[141],pp51[142],pp51[143],pp51[144],pp51[145],pp51[146],pp51[147],pp51[148],pp50[150],pp49[152],pp48[154],pp47[156],pp46[158],pp45[160],pp44[162],pp43[164],pp42[166],pp41[168],pp40[170],pp39[172],pp38[174],pp37[176],pp36[178],pp35[180],pp34[182],pp33[184],pp32[186],pp31[188],pp30[190],pp29[192],pp28[194],pp27[196],pp26[198],pp25[200],pp24[202],pp23[204],pp22[206],pp21[208],pp20[210],pp19[212],pp18[214],pp17[216],pp16[218],pp15[220],pp14[222],pp13[224],pp12[226],pp11[228],pp10[230],pp141[100],pp141[101],pp141[102],pp141[103],pp141[104],pp141[105],pp141[106],pp141[107],pp141[108],pp141[109],pp141[110],pp141[111],pp141[112],pp141[113],pp141[114],pp141[115],pp141[116],pp141[117],pp141[118],pp141[119],pp141[120],pp141[121],pp141[122],pp141[123],pp141[124],pp141[125],pp141[126],pp141[127],pp141[128],pp141[129],pp141[130],pp141[131],pp141[132],pp141[133],pp141[134],pp141[135],pp141[136],pp141[137],pp141[138],pp141[139],pp141[140],pp141[141],pp141[142],pp141[143],pp141[144],pp141[145],pp141[146],pp141[147],pp141[148],pp141[149],pp141[150],pp141[151],pp141[152],pp141[153],pp141[154],pp141[155],pp141[156],pp141[157],pp141[158],pp141[159],pp141[160],pp141[161],pp141[162],pp141[163],pp141[164],pp141[165],pp141[166],pp141[167],pp141[168],pp141[169],pp141[170],pp141[171],pp141[172],pp141[173],pp141[174],pp141[175],pp141[176],pp141[177],pp141[178],pp141[179],pp141[180],pp141[181],pp141[182],pp141[183],pp141[184],pp141[185],pp141[186],pp141[187],pp141[188],pp141[189],pp141[190],pp141[191],pp141[192],pp141[193],pp141[194],pp141[195],pp141[196],pp141[197],pp141[198],pp141[199],pp141[200],pp141[201],pp141[202],pp141[203],pp141[204],pp141[205],pp141[206],pp141[207],pp141[208],pp141[209],pp141[210],pp141[211],pp141[212],pp141[213],pp141[214],pp142[214],pp143[214],pp144[214],pp145[214],pp146[214],pp147[214],pp148[214],pp149[214]};
    CLA_216 KS_21(s21, c21, in21_1, in21_2);
    wire[213:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp102[47],pp101[49],pp100[51],pp52[100],pp52[101],pp52[102],pp52[103],pp52[104],pp52[105],pp52[106],pp52[107],pp52[108],pp52[109],pp52[110],pp52[111],pp52[112],pp52[113],pp52[114],pp52[115],pp52[116],pp52[117],pp52[118],pp52[119],pp52[120],pp52[121],pp52[122],pp52[123],pp52[124],pp52[125],pp52[126],pp52[127],pp52[128],pp52[129],pp52[130],pp52[131],pp52[132],pp52[133],pp52[134],pp52[135],pp52[136],pp52[137],pp52[138],pp52[139],pp52[140],pp52[141],pp52[142],pp52[143],pp52[144],pp52[145],pp52[146],pp52[147],pp51[149],pp50[151],pp49[153],pp48[155],pp47[157],pp46[159],pp45[161],pp44[163],pp43[165],pp42[167],pp41[169],pp40[171],pp39[173],pp38[175],pp37[177],pp36[179],pp35[181],pp34[183],pp33[185],pp32[187],pp31[189],pp30[191],pp29[193],pp28[195],pp27[197],pp26[199],pp25[201],pp24[203],pp23[205],pp22[207],pp21[209],pp20[211],pp19[213],pp18[215],pp17[217],pp16[219],pp15[221],pp14[223],pp13[225],pp12[227],pp11[229],pp10[231],pp142[100],pp142[101],pp142[102],pp142[103],pp142[104],pp142[105],pp142[106],pp142[107],pp142[108],pp142[109],pp142[110],pp142[111],pp142[112],pp142[113],pp142[114],pp142[115],pp142[116],pp142[117],pp142[118],pp142[119],pp142[120],pp142[121],pp142[122],pp142[123],pp142[124],pp142[125],pp142[126],pp142[127],pp142[128],pp142[129],pp142[130],pp142[131],pp142[132],pp142[133],pp142[134],pp142[135],pp142[136],pp142[137],pp142[138],pp142[139],pp142[140],pp142[141],pp142[142],pp142[143],pp142[144],pp142[145],pp142[146],pp142[147],pp142[148],pp142[149],pp142[150],pp142[151],pp142[152],pp142[153],pp142[154],pp142[155],pp142[156],pp142[157],pp142[158],pp142[159],pp142[160],pp142[161],pp142[162],pp142[163],pp142[164],pp142[165],pp142[166],pp142[167],pp142[168],pp142[169],pp142[170],pp142[171],pp142[172],pp142[173],pp142[174],pp142[175],pp142[176],pp142[177],pp142[178],pp142[179],pp142[180],pp142[181],pp142[182],pp142[183],pp142[184],pp142[185],pp142[186],pp142[187],pp142[188],pp142[189],pp142[190],pp142[191],pp142[192],pp142[193],pp142[194],pp142[195],pp142[196],pp142[197],pp142[198],pp142[199],pp142[200],pp142[201],pp142[202],pp142[203],pp142[204],pp142[205],pp142[206],pp142[207],pp142[208],pp142[209],pp142[210],pp142[211],pp142[212],pp142[213],pp143[213],pp144[213],pp145[213],pp146[213],pp147[213],pp148[213],pp149[213]};
    assign in22_2 = {pp103[46],pp102[48],pp101[50],pp100[52],pp53[100],pp53[101],pp53[102],pp53[103],pp53[104],pp53[105],pp53[106],pp53[107],pp53[108],pp53[109],pp53[110],pp53[111],pp53[112],pp53[113],pp53[114],pp53[115],pp53[116],pp53[117],pp53[118],pp53[119],pp53[120],pp53[121],pp53[122],pp53[123],pp53[124],pp53[125],pp53[126],pp53[127],pp53[128],pp53[129],pp53[130],pp53[131],pp53[132],pp53[133],pp53[134],pp53[135],pp53[136],pp53[137],pp53[138],pp53[139],pp53[140],pp53[141],pp53[142],pp53[143],pp53[144],pp53[145],pp53[146],pp52[148],pp51[150],pp50[152],pp49[154],pp48[156],pp47[158],pp46[160],pp45[162],pp44[164],pp43[166],pp42[168],pp41[170],pp40[172],pp39[174],pp38[176],pp37[178],pp36[180],pp35[182],pp34[184],pp33[186],pp32[188],pp31[190],pp30[192],pp29[194],pp28[196],pp27[198],pp26[200],pp25[202],pp24[204],pp23[206],pp22[208],pp21[210],pp20[212],pp19[214],pp18[216],pp17[218],pp16[220],pp15[222],pp14[224],pp13[226],pp12[228],pp11[230],pp10[232],pp143[100],pp143[101],pp143[102],pp143[103],pp143[104],pp143[105],pp143[106],pp143[107],pp143[108],pp143[109],pp143[110],pp143[111],pp143[112],pp143[113],pp143[114],pp143[115],pp143[116],pp143[117],pp143[118],pp143[119],pp143[120],pp143[121],pp143[122],pp143[123],pp143[124],pp143[125],pp143[126],pp143[127],pp143[128],pp143[129],pp143[130],pp143[131],pp143[132],pp143[133],pp143[134],pp143[135],pp143[136],pp143[137],pp143[138],pp143[139],pp143[140],pp143[141],pp143[142],pp143[143],pp143[144],pp143[145],pp143[146],pp143[147],pp143[148],pp143[149],pp143[150],pp143[151],pp143[152],pp143[153],pp143[154],pp143[155],pp143[156],pp143[157],pp143[158],pp143[159],pp143[160],pp143[161],pp143[162],pp143[163],pp143[164],pp143[165],pp143[166],pp143[167],pp143[168],pp143[169],pp143[170],pp143[171],pp143[172],pp143[173],pp143[174],pp143[175],pp143[176],pp143[177],pp143[178],pp143[179],pp143[180],pp143[181],pp143[182],pp143[183],pp143[184],pp143[185],pp143[186],pp143[187],pp143[188],pp143[189],pp143[190],pp143[191],pp143[192],pp143[193],pp143[194],pp143[195],pp143[196],pp143[197],pp143[198],pp143[199],pp143[200],pp143[201],pp143[202],pp143[203],pp143[204],pp143[205],pp143[206],pp143[207],pp143[208],pp143[209],pp143[210],pp143[211],pp143[212],pp144[212],pp145[212],pp146[212],pp147[212],pp148[212],pp149[212],pp150[212]};
    CLA_214 KS_22(s22, c22, in22_1, in22_2);
    wire[211:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp103[47],pp102[49],pp101[51],pp100[53],pp54[100],pp54[101],pp54[102],pp54[103],pp54[104],pp54[105],pp54[106],pp54[107],pp54[108],pp54[109],pp54[110],pp54[111],pp54[112],pp54[113],pp54[114],pp54[115],pp54[116],pp54[117],pp54[118],pp54[119],pp54[120],pp54[121],pp54[122],pp54[123],pp54[124],pp54[125],pp54[126],pp54[127],pp54[128],pp54[129],pp54[130],pp54[131],pp54[132],pp54[133],pp54[134],pp54[135],pp54[136],pp54[137],pp54[138],pp54[139],pp54[140],pp54[141],pp54[142],pp54[143],pp54[144],pp54[145],pp53[147],pp52[149],pp51[151],pp50[153],pp49[155],pp48[157],pp47[159],pp46[161],pp45[163],pp44[165],pp43[167],pp42[169],pp41[171],pp40[173],pp39[175],pp38[177],pp37[179],pp36[181],pp35[183],pp34[185],pp33[187],pp32[189],pp31[191],pp30[193],pp29[195],pp28[197],pp27[199],pp26[201],pp25[203],pp24[205],pp23[207],pp22[209],pp21[211],pp20[213],pp19[215],pp18[217],pp17[219],pp16[221],pp15[223],pp14[225],pp13[227],pp12[229],pp11[231],pp10[233],pp144[100],pp144[101],pp144[102],pp144[103],pp144[104],pp144[105],pp144[106],pp144[107],pp144[108],pp144[109],pp144[110],pp144[111],pp144[112],pp144[113],pp144[114],pp144[115],pp144[116],pp144[117],pp144[118],pp144[119],pp144[120],pp144[121],pp144[122],pp144[123],pp144[124],pp144[125],pp144[126],pp144[127],pp144[128],pp144[129],pp144[130],pp144[131],pp144[132],pp144[133],pp144[134],pp144[135],pp144[136],pp144[137],pp144[138],pp144[139],pp144[140],pp144[141],pp144[142],pp144[143],pp144[144],pp144[145],pp144[146],pp144[147],pp144[148],pp144[149],pp144[150],pp144[151],pp144[152],pp144[153],pp144[154],pp144[155],pp144[156],pp144[157],pp144[158],pp144[159],pp144[160],pp144[161],pp144[162],pp144[163],pp144[164],pp144[165],pp144[166],pp144[167],pp144[168],pp144[169],pp144[170],pp144[171],pp144[172],pp144[173],pp144[174],pp144[175],pp144[176],pp144[177],pp144[178],pp144[179],pp144[180],pp144[181],pp144[182],pp144[183],pp144[184],pp144[185],pp144[186],pp144[187],pp144[188],pp144[189],pp144[190],pp144[191],pp144[192],pp144[193],pp144[194],pp144[195],pp144[196],pp144[197],pp144[198],pp144[199],pp144[200],pp144[201],pp144[202],pp144[203],pp144[204],pp144[205],pp144[206],pp144[207],pp144[208],pp144[209],pp144[210],pp144[211],pp145[211],pp146[211],pp147[211],pp148[211],pp149[211],pp150[211]};
    assign in23_2 = {pp104[46],pp103[48],pp102[50],pp101[52],pp100[54],pp55[100],pp55[101],pp55[102],pp55[103],pp55[104],pp55[105],pp55[106],pp55[107],pp55[108],pp55[109],pp55[110],pp55[111],pp55[112],pp55[113],pp55[114],pp55[115],pp55[116],pp55[117],pp55[118],pp55[119],pp55[120],pp55[121],pp55[122],pp55[123],pp55[124],pp55[125],pp55[126],pp55[127],pp55[128],pp55[129],pp55[130],pp55[131],pp55[132],pp55[133],pp55[134],pp55[135],pp55[136],pp55[137],pp55[138],pp55[139],pp55[140],pp55[141],pp55[142],pp55[143],pp55[144],pp54[146],pp53[148],pp52[150],pp51[152],pp50[154],pp49[156],pp48[158],pp47[160],pp46[162],pp45[164],pp44[166],pp43[168],pp42[170],pp41[172],pp40[174],pp39[176],pp38[178],pp37[180],pp36[182],pp35[184],pp34[186],pp33[188],pp32[190],pp31[192],pp30[194],pp29[196],pp28[198],pp27[200],pp26[202],pp25[204],pp24[206],pp23[208],pp22[210],pp21[212],pp20[214],pp19[216],pp18[218],pp17[220],pp16[222],pp15[224],pp14[226],pp13[228],pp12[230],pp11[232],pp10[234],pp145[100],pp145[101],pp145[102],pp145[103],pp145[104],pp145[105],pp145[106],pp145[107],pp145[108],pp145[109],pp145[110],pp145[111],pp145[112],pp145[113],pp145[114],pp145[115],pp145[116],pp145[117],pp145[118],pp145[119],pp145[120],pp145[121],pp145[122],pp145[123],pp145[124],pp145[125],pp145[126],pp145[127],pp145[128],pp145[129],pp145[130],pp145[131],pp145[132],pp145[133],pp145[134],pp145[135],pp145[136],pp145[137],pp145[138],pp145[139],pp145[140],pp145[141],pp145[142],pp145[143],pp145[144],pp145[145],pp145[146],pp145[147],pp145[148],pp145[149],pp145[150],pp145[151],pp145[152],pp145[153],pp145[154],pp145[155],pp145[156],pp145[157],pp145[158],pp145[159],pp145[160],pp145[161],pp145[162],pp145[163],pp145[164],pp145[165],pp145[166],pp145[167],pp145[168],pp145[169],pp145[170],pp145[171],pp145[172],pp145[173],pp145[174],pp145[175],pp145[176],pp145[177],pp145[178],pp145[179],pp145[180],pp145[181],pp145[182],pp145[183],pp145[184],pp145[185],pp145[186],pp145[187],pp145[188],pp145[189],pp145[190],pp145[191],pp145[192],pp145[193],pp145[194],pp145[195],pp145[196],pp145[197],pp145[198],pp145[199],pp145[200],pp145[201],pp145[202],pp145[203],pp145[204],pp145[205],pp145[206],pp145[207],pp145[208],pp145[209],pp145[210],pp146[210],pp147[210],pp148[210],pp149[210],pp150[210],pp151[210]};
    CLA_212 KS_23(s23, c23, in23_1, in23_2);
    wire[209:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp104[47],pp103[49],pp102[51],pp101[53],pp100[55],pp56[100],pp56[101],pp56[102],pp56[103],pp56[104],pp56[105],pp56[106],pp56[107],pp56[108],pp56[109],pp56[110],pp56[111],pp56[112],pp56[113],pp56[114],pp56[115],pp56[116],pp56[117],pp56[118],pp56[119],pp56[120],pp56[121],pp56[122],pp56[123],pp56[124],pp56[125],pp56[126],pp56[127],pp56[128],pp56[129],pp56[130],pp56[131],pp56[132],pp56[133],pp56[134],pp56[135],pp56[136],pp56[137],pp56[138],pp56[139],pp56[140],pp56[141],pp56[142],pp56[143],pp55[145],pp54[147],pp53[149],pp52[151],pp51[153],pp50[155],pp49[157],pp48[159],pp47[161],pp46[163],pp45[165],pp44[167],pp43[169],pp42[171],pp41[173],pp40[175],pp39[177],pp38[179],pp37[181],pp36[183],pp35[185],pp34[187],pp33[189],pp32[191],pp31[193],pp30[195],pp29[197],pp28[199],pp27[201],pp26[203],pp25[205],pp24[207],pp23[209],pp22[211],pp21[213],pp20[215],pp19[217],pp18[219],pp17[221],pp16[223],pp15[225],pp14[227],pp13[229],pp12[231],pp11[233],pp10[235],pp146[100],pp146[101],pp146[102],pp146[103],pp146[104],pp146[105],pp146[106],pp146[107],pp146[108],pp146[109],pp146[110],pp146[111],pp146[112],pp146[113],pp146[114],pp146[115],pp146[116],pp146[117],pp146[118],pp146[119],pp146[120],pp146[121],pp146[122],pp146[123],pp146[124],pp146[125],pp146[126],pp146[127],pp146[128],pp146[129],pp146[130],pp146[131],pp146[132],pp146[133],pp146[134],pp146[135],pp146[136],pp146[137],pp146[138],pp146[139],pp146[140],pp146[141],pp146[142],pp146[143],pp146[144],pp146[145],pp146[146],pp146[147],pp146[148],pp146[149],pp146[150],pp146[151],pp146[152],pp146[153],pp146[154],pp146[155],pp146[156],pp146[157],pp146[158],pp146[159],pp146[160],pp146[161],pp146[162],pp146[163],pp146[164],pp146[165],pp146[166],pp146[167],pp146[168],pp146[169],pp146[170],pp146[171],pp146[172],pp146[173],pp146[174],pp146[175],pp146[176],pp146[177],pp146[178],pp146[179],pp146[180],pp146[181],pp146[182],pp146[183],pp146[184],pp146[185],pp146[186],pp146[187],pp146[188],pp146[189],pp146[190],pp146[191],pp146[192],pp146[193],pp146[194],pp146[195],pp146[196],pp146[197],pp146[198],pp146[199],pp146[200],pp146[201],pp146[202],pp146[203],pp146[204],pp146[205],pp146[206],pp146[207],pp146[208],pp146[209],pp147[209],pp148[209],pp149[209],pp150[209],pp151[209]};
    assign in24_2 = {pp105[46],pp104[48],pp103[50],pp102[52],pp101[54],pp100[56],pp57[100],pp57[101],pp57[102],pp57[103],pp57[104],pp57[105],pp57[106],pp57[107],pp57[108],pp57[109],pp57[110],pp57[111],pp57[112],pp57[113],pp57[114],pp57[115],pp57[116],pp57[117],pp57[118],pp57[119],pp57[120],pp57[121],pp57[122],pp57[123],pp57[124],pp57[125],pp57[126],pp57[127],pp57[128],pp57[129],pp57[130],pp57[131],pp57[132],pp57[133],pp57[134],pp57[135],pp57[136],pp57[137],pp57[138],pp57[139],pp57[140],pp57[141],pp57[142],pp56[144],pp55[146],pp54[148],pp53[150],pp52[152],pp51[154],pp50[156],pp49[158],pp48[160],pp47[162],pp46[164],pp45[166],pp44[168],pp43[170],pp42[172],pp41[174],pp40[176],pp39[178],pp38[180],pp37[182],pp36[184],pp35[186],pp34[188],pp33[190],pp32[192],pp31[194],pp30[196],pp29[198],pp28[200],pp27[202],pp26[204],pp25[206],pp24[208],pp23[210],pp22[212],pp21[214],pp20[216],pp19[218],pp18[220],pp17[222],pp16[224],pp15[226],pp14[228],pp13[230],pp12[232],pp11[234],pp10[236],pp147[100],pp147[101],pp147[102],pp147[103],pp147[104],pp147[105],pp147[106],pp147[107],pp147[108],pp147[109],pp147[110],pp147[111],pp147[112],pp147[113],pp147[114],pp147[115],pp147[116],pp147[117],pp147[118],pp147[119],pp147[120],pp147[121],pp147[122],pp147[123],pp147[124],pp147[125],pp147[126],pp147[127],pp147[128],pp147[129],pp147[130],pp147[131],pp147[132],pp147[133],pp147[134],pp147[135],pp147[136],pp147[137],pp147[138],pp147[139],pp147[140],pp147[141],pp147[142],pp147[143],pp147[144],pp147[145],pp147[146],pp147[147],pp147[148],pp147[149],pp147[150],pp147[151],pp147[152],pp147[153],pp147[154],pp147[155],pp147[156],pp147[157],pp147[158],pp147[159],pp147[160],pp147[161],pp147[162],pp147[163],pp147[164],pp147[165],pp147[166],pp147[167],pp147[168],pp147[169],pp147[170],pp147[171],pp147[172],pp147[173],pp147[174],pp147[175],pp147[176],pp147[177],pp147[178],pp147[179],pp147[180],pp147[181],pp147[182],pp147[183],pp147[184],pp147[185],pp147[186],pp147[187],pp147[188],pp147[189],pp147[190],pp147[191],pp147[192],pp147[193],pp147[194],pp147[195],pp147[196],pp147[197],pp147[198],pp147[199],pp147[200],pp147[201],pp147[202],pp147[203],pp147[204],pp147[205],pp147[206],pp147[207],pp147[208],pp148[208],pp149[208],pp150[208],pp151[208],pp152[208]};
    CLA_210 KS_24(s24, c24, in24_1, in24_2);
    wire[207:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp105[47],pp104[49],pp103[51],pp102[53],pp101[55],pp100[57],pp58[100],pp58[101],pp58[102],pp58[103],pp58[104],pp58[105],pp58[106],pp58[107],pp58[108],pp58[109],pp58[110],pp58[111],pp58[112],pp58[113],pp58[114],pp58[115],pp58[116],pp58[117],pp58[118],pp58[119],pp58[120],pp58[121],pp58[122],pp58[123],pp58[124],pp58[125],pp58[126],pp58[127],pp58[128],pp58[129],pp58[130],pp58[131],pp58[132],pp58[133],pp58[134],pp58[135],pp58[136],pp58[137],pp58[138],pp58[139],pp58[140],pp58[141],pp57[143],pp56[145],pp55[147],pp54[149],pp53[151],pp52[153],pp51[155],pp50[157],pp49[159],pp48[161],pp47[163],pp46[165],pp45[167],pp44[169],pp43[171],pp42[173],pp41[175],pp40[177],pp39[179],pp38[181],pp37[183],pp36[185],pp35[187],pp34[189],pp33[191],pp32[193],pp31[195],pp30[197],pp29[199],pp28[201],pp27[203],pp26[205],pp25[207],pp24[209],pp23[211],pp22[213],pp21[215],pp20[217],pp19[219],pp18[221],pp17[223],pp16[225],pp15[227],pp14[229],pp13[231],pp12[233],pp11[235],pp10[237],pp148[100],pp148[101],pp148[102],pp148[103],pp148[104],pp148[105],pp148[106],pp148[107],pp148[108],pp148[109],pp148[110],pp148[111],pp148[112],pp148[113],pp148[114],pp148[115],pp148[116],pp148[117],pp148[118],pp148[119],pp148[120],pp148[121],pp148[122],pp148[123],pp148[124],pp148[125],pp148[126],pp148[127],pp148[128],pp148[129],pp148[130],pp148[131],pp148[132],pp148[133],pp148[134],pp148[135],pp148[136],pp148[137],pp148[138],pp148[139],pp148[140],pp148[141],pp148[142],pp148[143],pp148[144],pp148[145],pp148[146],pp148[147],pp148[148],pp148[149],pp148[150],pp148[151],pp148[152],pp148[153],pp148[154],pp148[155],pp148[156],pp148[157],pp148[158],pp148[159],pp148[160],pp148[161],pp148[162],pp148[163],pp148[164],pp148[165],pp148[166],pp148[167],pp148[168],pp148[169],pp148[170],pp148[171],pp148[172],pp148[173],pp148[174],pp148[175],pp148[176],pp148[177],pp148[178],pp148[179],pp148[180],pp148[181],pp148[182],pp148[183],pp148[184],pp148[185],pp148[186],pp148[187],pp148[188],pp148[189],pp148[190],pp148[191],pp148[192],pp148[193],pp148[194],pp148[195],pp148[196],pp148[197],pp148[198],pp148[199],pp148[200],pp148[201],pp148[202],pp148[203],pp148[204],pp148[205],pp148[206],pp148[207],pp149[207],pp150[207],pp151[207],pp152[207]};
    assign in25_2 = {pp106[46],pp105[48],pp104[50],pp103[52],pp102[54],pp101[56],pp100[58],pp59[100],pp59[101],pp59[102],pp59[103],pp59[104],pp59[105],pp59[106],pp59[107],pp59[108],pp59[109],pp59[110],pp59[111],pp59[112],pp59[113],pp59[114],pp59[115],pp59[116],pp59[117],pp59[118],pp59[119],pp59[120],pp59[121],pp59[122],pp59[123],pp59[124],pp59[125],pp59[126],pp59[127],pp59[128],pp59[129],pp59[130],pp59[131],pp59[132],pp59[133],pp59[134],pp59[135],pp59[136],pp59[137],pp59[138],pp59[139],pp59[140],pp58[142],pp57[144],pp56[146],pp55[148],pp54[150],pp53[152],pp52[154],pp51[156],pp50[158],pp49[160],pp48[162],pp47[164],pp46[166],pp45[168],pp44[170],pp43[172],pp42[174],pp41[176],pp40[178],pp39[180],pp38[182],pp37[184],pp36[186],pp35[188],pp34[190],pp33[192],pp32[194],pp31[196],pp30[198],pp29[200],pp28[202],pp27[204],pp26[206],pp25[208],pp24[210],pp23[212],pp22[214],pp21[216],pp20[218],pp19[220],pp18[222],pp17[224],pp16[226],pp15[228],pp14[230],pp13[232],pp12[234],pp11[236],pp10[238],pp149[100],pp149[101],pp149[102],pp149[103],pp149[104],pp149[105],pp149[106],pp149[107],pp149[108],pp149[109],pp149[110],pp149[111],pp149[112],pp149[113],pp149[114],pp149[115],pp149[116],pp149[117],pp149[118],pp149[119],pp149[120],pp149[121],pp149[122],pp149[123],pp149[124],pp149[125],pp149[126],pp149[127],pp149[128],pp149[129],pp149[130],pp149[131],pp149[132],pp149[133],pp149[134],pp149[135],pp149[136],pp149[137],pp149[138],pp149[139],pp149[140],pp149[141],pp149[142],pp149[143],pp149[144],pp149[145],pp149[146],pp149[147],pp149[148],pp149[149],pp149[150],pp149[151],pp149[152],pp149[153],pp149[154],pp149[155],pp149[156],pp149[157],pp149[158],pp149[159],pp149[160],pp149[161],pp149[162],pp149[163],pp149[164],pp149[165],pp149[166],pp149[167],pp149[168],pp149[169],pp149[170],pp149[171],pp149[172],pp149[173],pp149[174],pp149[175],pp149[176],pp149[177],pp149[178],pp149[179],pp149[180],pp149[181],pp149[182],pp149[183],pp149[184],pp149[185],pp149[186],pp149[187],pp149[188],pp149[189],pp149[190],pp149[191],pp149[192],pp149[193],pp149[194],pp149[195],pp149[196],pp149[197],pp149[198],pp149[199],pp149[200],pp149[201],pp149[202],pp149[203],pp149[204],pp149[205],pp149[206],pp150[206],pp151[206],pp152[206],pp153[206]};
    CLA_208 KS_25(s25, c25, in25_1, in25_2);
    wire[205:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp106[47],pp105[49],pp104[51],pp103[53],pp102[55],pp101[57],pp100[59],pp60[100],pp60[101],pp60[102],pp60[103],pp60[104],pp60[105],pp60[106],pp60[107],pp60[108],pp60[109],pp60[110],pp60[111],pp60[112],pp60[113],pp60[114],pp60[115],pp60[116],pp60[117],pp60[118],pp60[119],pp60[120],pp60[121],pp60[122],pp60[123],pp60[124],pp60[125],pp60[126],pp60[127],pp60[128],pp60[129],pp60[130],pp60[131],pp60[132],pp60[133],pp60[134],pp60[135],pp60[136],pp60[137],pp60[138],pp60[139],pp59[141],pp58[143],pp57[145],pp56[147],pp55[149],pp54[151],pp53[153],pp52[155],pp51[157],pp50[159],pp49[161],pp48[163],pp47[165],pp46[167],pp45[169],pp44[171],pp43[173],pp42[175],pp41[177],pp40[179],pp39[181],pp38[183],pp37[185],pp36[187],pp35[189],pp34[191],pp33[193],pp32[195],pp31[197],pp30[199],pp29[201],pp28[203],pp27[205],pp26[207],pp25[209],pp24[211],pp23[213],pp22[215],pp21[217],pp20[219],pp19[221],pp18[223],pp17[225],pp16[227],pp15[229],pp14[231],pp13[233],pp12[235],pp11[237],pp10[239],pp150[100],pp150[101],pp150[102],pp150[103],pp150[104],pp150[105],pp150[106],pp150[107],pp150[108],pp150[109],pp150[110],pp150[111],pp150[112],pp150[113],pp150[114],pp150[115],pp150[116],pp150[117],pp150[118],pp150[119],pp150[120],pp150[121],pp150[122],pp150[123],pp150[124],pp150[125],pp150[126],pp150[127],pp150[128],pp150[129],pp150[130],pp150[131],pp150[132],pp150[133],pp150[134],pp150[135],pp150[136],pp150[137],pp150[138],pp150[139],pp150[140],pp150[141],pp150[142],pp150[143],pp150[144],pp150[145],pp150[146],pp150[147],pp150[148],pp150[149],pp150[150],pp150[151],pp150[152],pp150[153],pp150[154],pp150[155],pp150[156],pp150[157],pp150[158],pp150[159],pp150[160],pp150[161],pp150[162],pp150[163],pp150[164],pp150[165],pp150[166],pp150[167],pp150[168],pp150[169],pp150[170],pp150[171],pp150[172],pp150[173],pp150[174],pp150[175],pp150[176],pp150[177],pp150[178],pp150[179],pp150[180],pp150[181],pp150[182],pp150[183],pp150[184],pp150[185],pp150[186],pp150[187],pp150[188],pp150[189],pp150[190],pp150[191],pp150[192],pp150[193],pp150[194],pp150[195],pp150[196],pp150[197],pp150[198],pp150[199],pp150[200],pp150[201],pp150[202],pp150[203],pp150[204],pp150[205],pp151[205],pp152[205],pp153[205]};
    assign in26_2 = {pp107[46],pp106[48],pp105[50],pp104[52],pp103[54],pp102[56],pp101[58],pp100[60],pp61[100],pp61[101],pp61[102],pp61[103],pp61[104],pp61[105],pp61[106],pp61[107],pp61[108],pp61[109],pp61[110],pp61[111],pp61[112],pp61[113],pp61[114],pp61[115],pp61[116],pp61[117],pp61[118],pp61[119],pp61[120],pp61[121],pp61[122],pp61[123],pp61[124],pp61[125],pp61[126],pp61[127],pp61[128],pp61[129],pp61[130],pp61[131],pp61[132],pp61[133],pp61[134],pp61[135],pp61[136],pp61[137],pp61[138],pp60[140],pp59[142],pp58[144],pp57[146],pp56[148],pp55[150],pp54[152],pp53[154],pp52[156],pp51[158],pp50[160],pp49[162],pp48[164],pp47[166],pp46[168],pp45[170],pp44[172],pp43[174],pp42[176],pp41[178],pp40[180],pp39[182],pp38[184],pp37[186],pp36[188],pp35[190],pp34[192],pp33[194],pp32[196],pp31[198],pp30[200],pp29[202],pp28[204],pp27[206],pp26[208],pp25[210],pp24[212],pp23[214],pp22[216],pp21[218],pp20[220],pp19[222],pp18[224],pp17[226],pp16[228],pp15[230],pp14[232],pp13[234],pp12[236],pp11[238],pp10[240],pp151[100],pp151[101],pp151[102],pp151[103],pp151[104],pp151[105],pp151[106],pp151[107],pp151[108],pp151[109],pp151[110],pp151[111],pp151[112],pp151[113],pp151[114],pp151[115],pp151[116],pp151[117],pp151[118],pp151[119],pp151[120],pp151[121],pp151[122],pp151[123],pp151[124],pp151[125],pp151[126],pp151[127],pp151[128],pp151[129],pp151[130],pp151[131],pp151[132],pp151[133],pp151[134],pp151[135],pp151[136],pp151[137],pp151[138],pp151[139],pp151[140],pp151[141],pp151[142],pp151[143],pp151[144],pp151[145],pp151[146],pp151[147],pp151[148],pp151[149],pp151[150],pp151[151],pp151[152],pp151[153],pp151[154],pp151[155],pp151[156],pp151[157],pp151[158],pp151[159],pp151[160],pp151[161],pp151[162],pp151[163],pp151[164],pp151[165],pp151[166],pp151[167],pp151[168],pp151[169],pp151[170],pp151[171],pp151[172],pp151[173],pp151[174],pp151[175],pp151[176],pp151[177],pp151[178],pp151[179],pp151[180],pp151[181],pp151[182],pp151[183],pp151[184],pp151[185],pp151[186],pp151[187],pp151[188],pp151[189],pp151[190],pp151[191],pp151[192],pp151[193],pp151[194],pp151[195],pp151[196],pp151[197],pp151[198],pp151[199],pp151[200],pp151[201],pp151[202],pp151[203],pp151[204],pp152[204],pp153[204],pp154[204]};
    CLA_206 KS_26(s26, c26, in26_1, in26_2);
    wire[203:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp107[47],pp106[49],pp105[51],pp104[53],pp103[55],pp102[57],pp101[59],pp100[61],pp62[100],pp62[101],pp62[102],pp62[103],pp62[104],pp62[105],pp62[106],pp62[107],pp62[108],pp62[109],pp62[110],pp62[111],pp62[112],pp62[113],pp62[114],pp62[115],pp62[116],pp62[117],pp62[118],pp62[119],pp62[120],pp62[121],pp62[122],pp62[123],pp62[124],pp62[125],pp62[126],pp62[127],pp62[128],pp62[129],pp62[130],pp62[131],pp62[132],pp62[133],pp62[134],pp62[135],pp62[136],pp62[137],pp61[139],pp60[141],pp59[143],pp58[145],pp57[147],pp56[149],pp55[151],pp54[153],pp53[155],pp52[157],pp51[159],pp50[161],pp49[163],pp48[165],pp47[167],pp46[169],pp45[171],pp44[173],pp43[175],pp42[177],pp41[179],pp40[181],pp39[183],pp38[185],pp37[187],pp36[189],pp35[191],pp34[193],pp33[195],pp32[197],pp31[199],pp30[201],pp29[203],pp28[205],pp27[207],pp26[209],pp25[211],pp24[213],pp23[215],pp22[217],pp21[219],pp20[221],pp19[223],pp18[225],pp17[227],pp16[229],pp15[231],pp14[233],pp13[235],pp12[237],pp11[239],pp10[241],pp152[100],pp152[101],pp152[102],pp152[103],pp152[104],pp152[105],pp152[106],pp152[107],pp152[108],pp152[109],pp152[110],pp152[111],pp152[112],pp152[113],pp152[114],pp152[115],pp152[116],pp152[117],pp152[118],pp152[119],pp152[120],pp152[121],pp152[122],pp152[123],pp152[124],pp152[125],pp152[126],pp152[127],pp152[128],pp152[129],pp152[130],pp152[131],pp152[132],pp152[133],pp152[134],pp152[135],pp152[136],pp152[137],pp152[138],pp152[139],pp152[140],pp152[141],pp152[142],pp152[143],pp152[144],pp152[145],pp152[146],pp152[147],pp152[148],pp152[149],pp152[150],pp152[151],pp152[152],pp152[153],pp152[154],pp152[155],pp152[156],pp152[157],pp152[158],pp152[159],pp152[160],pp152[161],pp152[162],pp152[163],pp152[164],pp152[165],pp152[166],pp152[167],pp152[168],pp152[169],pp152[170],pp152[171],pp152[172],pp152[173],pp152[174],pp152[175],pp152[176],pp152[177],pp152[178],pp152[179],pp152[180],pp152[181],pp152[182],pp152[183],pp152[184],pp152[185],pp152[186],pp152[187],pp152[188],pp152[189],pp152[190],pp152[191],pp152[192],pp152[193],pp152[194],pp152[195],pp152[196],pp152[197],pp152[198],pp152[199],pp152[200],pp152[201],pp152[202],pp152[203],pp153[203],pp154[203]};
    assign in27_2 = {pp108[46],pp107[48],pp106[50],pp105[52],pp104[54],pp103[56],pp102[58],pp101[60],pp100[62],pp63[100],pp63[101],pp63[102],pp63[103],pp63[104],pp63[105],pp63[106],pp63[107],pp63[108],pp63[109],pp63[110],pp63[111],pp63[112],pp63[113],pp63[114],pp63[115],pp63[116],pp63[117],pp63[118],pp63[119],pp63[120],pp63[121],pp63[122],pp63[123],pp63[124],pp63[125],pp63[126],pp63[127],pp63[128],pp63[129],pp63[130],pp63[131],pp63[132],pp63[133],pp63[134],pp63[135],pp63[136],pp62[138],pp61[140],pp60[142],pp59[144],pp58[146],pp57[148],pp56[150],pp55[152],pp54[154],pp53[156],pp52[158],pp51[160],pp50[162],pp49[164],pp48[166],pp47[168],pp46[170],pp45[172],pp44[174],pp43[176],pp42[178],pp41[180],pp40[182],pp39[184],pp38[186],pp37[188],pp36[190],pp35[192],pp34[194],pp33[196],pp32[198],pp31[200],pp30[202],pp29[204],pp28[206],pp27[208],pp26[210],pp25[212],pp24[214],pp23[216],pp22[218],pp21[220],pp20[222],pp19[224],pp18[226],pp17[228],pp16[230],pp15[232],pp14[234],pp13[236],pp12[238],pp11[240],pp10[242],pp153[100],pp153[101],pp153[102],pp153[103],pp153[104],pp153[105],pp153[106],pp153[107],pp153[108],pp153[109],pp153[110],pp153[111],pp153[112],pp153[113],pp153[114],pp153[115],pp153[116],pp153[117],pp153[118],pp153[119],pp153[120],pp153[121],pp153[122],pp153[123],pp153[124],pp153[125],pp153[126],pp153[127],pp153[128],pp153[129],pp153[130],pp153[131],pp153[132],pp153[133],pp153[134],pp153[135],pp153[136],pp153[137],pp153[138],pp153[139],pp153[140],pp153[141],pp153[142],pp153[143],pp153[144],pp153[145],pp153[146],pp153[147],pp153[148],pp153[149],pp153[150],pp153[151],pp153[152],pp153[153],pp153[154],pp153[155],pp153[156],pp153[157],pp153[158],pp153[159],pp153[160],pp153[161],pp153[162],pp153[163],pp153[164],pp153[165],pp153[166],pp153[167],pp153[168],pp153[169],pp153[170],pp153[171],pp153[172],pp153[173],pp153[174],pp153[175],pp153[176],pp153[177],pp153[178],pp153[179],pp153[180],pp153[181],pp153[182],pp153[183],pp153[184],pp153[185],pp153[186],pp153[187],pp153[188],pp153[189],pp153[190],pp153[191],pp153[192],pp153[193],pp153[194],pp153[195],pp153[196],pp153[197],pp153[198],pp153[199],pp153[200],pp153[201],pp153[202],pp154[202],pp155[202]};
    CLA_204 KS_27(s27, c27, in27_1, in27_2);
    wire[201:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp108[47],pp107[49],pp106[51],pp105[53],pp104[55],pp103[57],pp102[59],pp101[61],pp100[63],pp64[100],pp64[101],pp64[102],pp64[103],pp64[104],pp64[105],pp64[106],pp64[107],pp64[108],pp64[109],pp64[110],pp64[111],pp64[112],pp64[113],pp64[114],pp64[115],pp64[116],pp64[117],pp64[118],pp64[119],pp64[120],pp64[121],pp64[122],pp64[123],pp64[124],pp64[125],pp64[126],pp64[127],pp64[128],pp64[129],pp64[130],pp64[131],pp64[132],pp64[133],pp64[134],pp64[135],pp63[137],pp62[139],pp61[141],pp60[143],pp59[145],pp58[147],pp57[149],pp56[151],pp55[153],pp54[155],pp53[157],pp52[159],pp51[161],pp50[163],pp49[165],pp48[167],pp47[169],pp46[171],pp45[173],pp44[175],pp43[177],pp42[179],pp41[181],pp40[183],pp39[185],pp38[187],pp37[189],pp36[191],pp35[193],pp34[195],pp33[197],pp32[199],pp31[201],pp30[203],pp29[205],pp28[207],pp27[209],pp26[211],pp25[213],pp24[215],pp23[217],pp22[219],pp21[221],pp20[223],pp19[225],pp18[227],pp17[229],pp16[231],pp15[233],pp14[235],pp13[237],pp12[239],pp11[241],pp10[243],pp154[100],pp154[101],pp154[102],pp154[103],pp154[104],pp154[105],pp154[106],pp154[107],pp154[108],pp154[109],pp154[110],pp154[111],pp154[112],pp154[113],pp154[114],pp154[115],pp154[116],pp154[117],pp154[118],pp154[119],pp154[120],pp154[121],pp154[122],pp154[123],pp154[124],pp154[125],pp154[126],pp154[127],pp154[128],pp154[129],pp154[130],pp154[131],pp154[132],pp154[133],pp154[134],pp154[135],pp154[136],pp154[137],pp154[138],pp154[139],pp154[140],pp154[141],pp154[142],pp154[143],pp154[144],pp154[145],pp154[146],pp154[147],pp154[148],pp154[149],pp154[150],pp154[151],pp154[152],pp154[153],pp154[154],pp154[155],pp154[156],pp154[157],pp154[158],pp154[159],pp154[160],pp154[161],pp154[162],pp154[163],pp154[164],pp154[165],pp154[166],pp154[167],pp154[168],pp154[169],pp154[170],pp154[171],pp154[172],pp154[173],pp154[174],pp154[175],pp154[176],pp154[177],pp154[178],pp154[179],pp154[180],pp154[181],pp154[182],pp154[183],pp154[184],pp154[185],pp154[186],pp154[187],pp154[188],pp154[189],pp154[190],pp154[191],pp154[192],pp154[193],pp154[194],pp154[195],pp154[196],pp154[197],pp154[198],pp154[199],pp154[200],pp154[201],pp155[201]};
    assign in28_2 = {pp109[46],pp108[48],pp107[50],pp106[52],pp105[54],pp104[56],pp103[58],pp102[60],pp101[62],pp100[64],pp65[100],pp65[101],pp65[102],pp65[103],pp65[104],pp65[105],pp65[106],pp65[107],pp65[108],pp65[109],pp65[110],pp65[111],pp65[112],pp65[113],pp65[114],pp65[115],pp65[116],pp65[117],pp65[118],pp65[119],pp65[120],pp65[121],pp65[122],pp65[123],pp65[124],pp65[125],pp65[126],pp65[127],pp65[128],pp65[129],pp65[130],pp65[131],pp65[132],pp65[133],pp65[134],pp64[136],pp63[138],pp62[140],pp61[142],pp60[144],pp59[146],pp58[148],pp57[150],pp56[152],pp55[154],pp54[156],pp53[158],pp52[160],pp51[162],pp50[164],pp49[166],pp48[168],pp47[170],pp46[172],pp45[174],pp44[176],pp43[178],pp42[180],pp41[182],pp40[184],pp39[186],pp38[188],pp37[190],pp36[192],pp35[194],pp34[196],pp33[198],pp32[200],pp31[202],pp30[204],pp29[206],pp28[208],pp27[210],pp26[212],pp25[214],pp24[216],pp23[218],pp22[220],pp21[222],pp20[224],pp19[226],pp18[228],pp17[230],pp16[232],pp15[234],pp14[236],pp13[238],pp12[240],pp11[242],pp10[244],pp155[100],pp155[101],pp155[102],pp155[103],pp155[104],pp155[105],pp155[106],pp155[107],pp155[108],pp155[109],pp155[110],pp155[111],pp155[112],pp155[113],pp155[114],pp155[115],pp155[116],pp155[117],pp155[118],pp155[119],pp155[120],pp155[121],pp155[122],pp155[123],pp155[124],pp155[125],pp155[126],pp155[127],pp155[128],pp155[129],pp155[130],pp155[131],pp155[132],pp155[133],pp155[134],pp155[135],pp155[136],pp155[137],pp155[138],pp155[139],pp155[140],pp155[141],pp155[142],pp155[143],pp155[144],pp155[145],pp155[146],pp155[147],pp155[148],pp155[149],pp155[150],pp155[151],pp155[152],pp155[153],pp155[154],pp155[155],pp155[156],pp155[157],pp155[158],pp155[159],pp155[160],pp155[161],pp155[162],pp155[163],pp155[164],pp155[165],pp155[166],pp155[167],pp155[168],pp155[169],pp155[170],pp155[171],pp155[172],pp155[173],pp155[174],pp155[175],pp155[176],pp155[177],pp155[178],pp155[179],pp155[180],pp155[181],pp155[182],pp155[183],pp155[184],pp155[185],pp155[186],pp155[187],pp155[188],pp155[189],pp155[190],pp155[191],pp155[192],pp155[193],pp155[194],pp155[195],pp155[196],pp155[197],pp155[198],pp155[199],pp155[200],pp156[200]};
    CLA_202 KS_28(s28, c28, in28_1, in28_2);
    wire[199:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp109[47],pp108[49],pp107[51],pp106[53],pp105[55],pp104[57],pp103[59],pp102[61],pp101[63],pp100[65],pp66[100],pp66[101],pp66[102],pp66[103],pp66[104],pp66[105],pp66[106],pp66[107],pp66[108],pp66[109],pp66[110],pp66[111],pp66[112],pp66[113],pp66[114],pp66[115],pp66[116],pp66[117],pp66[118],pp66[119],pp66[120],pp66[121],pp66[122],pp66[123],pp66[124],pp66[125],pp66[126],pp66[127],pp66[128],pp66[129],pp66[130],pp66[131],pp66[132],pp66[133],pp65[135],pp64[137],pp63[139],pp62[141],pp61[143],pp60[145],pp59[147],pp58[149],pp57[151],pp56[153],pp55[155],pp54[157],pp53[159],pp52[161],pp51[163],pp50[165],pp49[167],pp48[169],pp47[171],pp46[173],pp45[175],pp44[177],pp43[179],pp42[181],pp41[183],pp40[185],pp39[187],pp38[189],pp37[191],pp36[193],pp35[195],pp34[197],pp33[199],pp32[201],pp31[203],pp30[205],pp29[207],pp28[209],pp27[211],pp26[213],pp25[215],pp24[217],pp23[219],pp22[221],pp21[223],pp20[225],pp19[227],pp18[229],pp17[231],pp16[233],pp15[235],pp14[237],pp13[239],pp12[241],pp11[243],pp10[245],pp156[100],pp156[101],pp156[102],pp156[103],pp156[104],pp156[105],pp156[106],pp156[107],pp156[108],pp156[109],pp156[110],pp156[111],pp156[112],pp156[113],pp156[114],pp156[115],pp156[116],pp156[117],pp156[118],pp156[119],pp156[120],pp156[121],pp156[122],pp156[123],pp156[124],pp156[125],pp156[126],pp156[127],pp156[128],pp156[129],pp156[130],pp156[131],pp156[132],pp156[133],pp156[134],pp156[135],pp156[136],pp156[137],pp156[138],pp156[139],pp156[140],pp156[141],pp156[142],pp156[143],pp156[144],pp156[145],pp156[146],pp156[147],pp156[148],pp156[149],pp156[150],pp156[151],pp156[152],pp156[153],pp156[154],pp156[155],pp156[156],pp156[157],pp156[158],pp156[159],pp156[160],pp156[161],pp156[162],pp156[163],pp156[164],pp156[165],pp156[166],pp156[167],pp156[168],pp156[169],pp156[170],pp156[171],pp156[172],pp156[173],pp156[174],pp156[175],pp156[176],pp156[177],pp156[178],pp156[179],pp156[180],pp156[181],pp156[182],pp156[183],pp156[184],pp156[185],pp156[186],pp156[187],pp156[188],pp156[189],pp156[190],pp156[191],pp156[192],pp156[193],pp156[194],pp156[195],pp156[196],pp156[197],pp156[198],pp156[199]};
    assign in29_2 = {pp110[46],pp109[48],pp108[50],pp107[52],pp106[54],pp105[56],pp104[58],pp103[60],pp102[62],pp101[64],pp100[66],pp67[100],pp67[101],pp67[102],pp67[103],pp67[104],pp67[105],pp67[106],pp67[107],pp67[108],pp67[109],pp67[110],pp67[111],pp67[112],pp67[113],pp67[114],pp67[115],pp67[116],pp67[117],pp67[118],pp67[119],pp67[120],pp67[121],pp67[122],pp67[123],pp67[124],pp67[125],pp67[126],pp67[127],pp67[128],pp67[129],pp67[130],pp67[131],pp67[132],pp66[134],pp65[136],pp64[138],pp63[140],pp62[142],pp61[144],pp60[146],pp59[148],pp58[150],pp57[152],pp56[154],pp55[156],pp54[158],pp53[160],pp52[162],pp51[164],pp50[166],pp49[168],pp48[170],pp47[172],pp46[174],pp45[176],pp44[178],pp43[180],pp42[182],pp41[184],pp40[186],pp39[188],pp38[190],pp37[192],pp36[194],pp35[196],pp34[198],pp33[200],pp32[202],pp31[204],pp30[206],pp29[208],pp28[210],pp27[212],pp26[214],pp25[216],pp24[218],pp23[220],pp22[222],pp21[224],pp20[226],pp19[228],pp18[230],pp17[232],pp16[234],pp15[236],pp14[238],pp13[240],pp12[242],pp11[244],pp10[246],pp157[100],pp157[101],pp157[102],pp157[103],pp157[104],pp157[105],pp157[106],pp157[107],pp157[108],pp157[109],pp157[110],pp157[111],pp157[112],pp157[113],pp157[114],pp157[115],pp157[116],pp157[117],pp157[118],pp157[119],pp157[120],pp157[121],pp157[122],pp157[123],pp157[124],pp157[125],pp157[126],pp157[127],pp157[128],pp157[129],pp157[130],pp157[131],pp157[132],pp157[133],pp157[134],pp157[135],pp157[136],pp157[137],pp157[138],pp157[139],pp157[140],pp157[141],pp157[142],pp157[143],pp157[144],pp157[145],pp157[146],pp157[147],pp157[148],pp157[149],pp157[150],pp157[151],pp157[152],pp157[153],pp157[154],pp157[155],pp157[156],pp157[157],pp157[158],pp157[159],pp157[160],pp157[161],pp157[162],pp157[163],pp157[164],pp157[165],pp157[166],pp157[167],pp157[168],pp157[169],pp157[170],pp157[171],pp157[172],pp157[173],pp157[174],pp157[175],pp157[176],pp157[177],pp157[178],pp157[179],pp157[180],pp157[181],pp157[182],pp157[183],pp157[184],pp157[185],pp157[186],pp157[187],pp157[188],pp157[189],pp157[190],pp157[191],pp157[192],pp157[193],pp157[194],pp157[195],pp157[196],pp157[197],pp157[198]};
    CLA_200 KS_29(s29, c29, in29_1, in29_2);
    wire[197:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp110[47],pp109[49],pp108[51],pp107[53],pp106[55],pp105[57],pp104[59],pp103[61],pp102[63],pp101[65],pp100[67],pp68[100],pp68[101],pp68[102],pp68[103],pp68[104],pp68[105],pp68[106],pp68[107],pp68[108],pp68[109],pp68[110],pp68[111],pp68[112],pp68[113],pp68[114],pp68[115],pp68[116],pp68[117],pp68[118],pp68[119],pp68[120],pp68[121],pp68[122],pp68[123],pp68[124],pp68[125],pp68[126],pp68[127],pp68[128],pp68[129],pp68[130],pp68[131],pp67[133],pp66[135],pp65[137],pp64[139],pp63[141],pp62[143],pp61[145],pp60[147],pp59[149],pp58[151],pp57[153],pp56[155],pp55[157],pp54[159],pp53[161],pp52[163],pp51[165],pp50[167],pp49[169],pp48[171],pp47[173],pp46[175],pp45[177],pp44[179],pp43[181],pp42[183],pp41[185],pp40[187],pp39[189],pp38[191],pp37[193],pp36[195],pp35[197],pp34[199],pp33[201],pp32[203],pp31[205],pp30[207],pp29[209],pp28[211],pp27[213],pp26[215],pp25[217],pp24[219],pp23[221],pp22[223],pp21[225],pp20[227],pp19[229],pp18[231],pp17[233],pp16[235],pp15[237],pp14[239],pp13[241],pp12[243],pp11[245],pp10[247],pp158[100],pp158[101],pp158[102],pp158[103],pp158[104],pp158[105],pp158[106],pp158[107],pp158[108],pp158[109],pp158[110],pp158[111],pp158[112],pp158[113],pp158[114],pp158[115],pp158[116],pp158[117],pp158[118],pp158[119],pp158[120],pp158[121],pp158[122],pp158[123],pp158[124],pp158[125],pp158[126],pp158[127],pp158[128],pp158[129],pp158[130],pp158[131],pp158[132],pp158[133],pp158[134],pp158[135],pp158[136],pp158[137],pp158[138],pp158[139],pp158[140],pp158[141],pp158[142],pp158[143],pp158[144],pp158[145],pp158[146],pp158[147],pp158[148],pp158[149],pp158[150],pp158[151],pp158[152],pp158[153],pp158[154],pp158[155],pp158[156],pp158[157],pp158[158],pp158[159],pp158[160],pp158[161],pp158[162],pp158[163],pp158[164],pp158[165],pp158[166],pp158[167],pp158[168],pp158[169],pp158[170],pp158[171],pp158[172],pp158[173],pp158[174],pp158[175],pp158[176],pp158[177],pp158[178],pp158[179],pp158[180],pp158[181],pp158[182],pp158[183],pp158[184],pp158[185],pp158[186],pp158[187],pp158[188],pp158[189],pp158[190],pp158[191],pp158[192],pp158[193],pp158[194],pp158[195],pp158[196]};
    assign in30_2 = {pp111[46],pp110[48],pp109[50],pp108[52],pp107[54],pp106[56],pp105[58],pp104[60],pp103[62],pp102[64],pp101[66],pp100[68],pp69[100],pp69[101],pp69[102],pp69[103],pp69[104],pp69[105],pp69[106],pp69[107],pp69[108],pp69[109],pp69[110],pp69[111],pp69[112],pp69[113],pp69[114],pp69[115],pp69[116],pp69[117],pp69[118],pp69[119],pp69[120],pp69[121],pp69[122],pp69[123],pp69[124],pp69[125],pp69[126],pp69[127],pp69[128],pp69[129],pp69[130],pp68[132],pp67[134],pp66[136],pp65[138],pp64[140],pp63[142],pp62[144],pp61[146],pp60[148],pp59[150],pp58[152],pp57[154],pp56[156],pp55[158],pp54[160],pp53[162],pp52[164],pp51[166],pp50[168],pp49[170],pp48[172],pp47[174],pp46[176],pp45[178],pp44[180],pp43[182],pp42[184],pp41[186],pp40[188],pp39[190],pp38[192],pp37[194],pp36[196],pp35[198],pp34[200],pp33[202],pp32[204],pp31[206],pp30[208],pp29[210],pp28[212],pp27[214],pp26[216],pp25[218],pp24[220],pp23[222],pp22[224],pp21[226],pp20[228],pp19[230],pp18[232],pp17[234],pp16[236],pp15[238],pp14[240],pp13[242],pp12[244],pp11[246],pp10[248],pp159[100],pp159[101],pp159[102],pp159[103],pp159[104],pp159[105],pp159[106],pp159[107],pp159[108],pp159[109],pp159[110],pp159[111],pp159[112],pp159[113],pp159[114],pp159[115],pp159[116],pp159[117],pp159[118],pp159[119],pp159[120],pp159[121],pp159[122],pp159[123],pp159[124],pp159[125],pp159[126],pp159[127],pp159[128],pp159[129],pp159[130],pp159[131],pp159[132],pp159[133],pp159[134],pp159[135],pp159[136],pp159[137],pp159[138],pp159[139],pp159[140],pp159[141],pp159[142],pp159[143],pp159[144],pp159[145],pp159[146],pp159[147],pp159[148],pp159[149],pp159[150],pp159[151],pp159[152],pp159[153],pp159[154],pp159[155],pp159[156],pp159[157],pp159[158],pp159[159],pp159[160],pp159[161],pp159[162],pp159[163],pp159[164],pp159[165],pp159[166],pp159[167],pp159[168],pp159[169],pp159[170],pp159[171],pp159[172],pp159[173],pp159[174],pp159[175],pp159[176],pp159[177],pp159[178],pp159[179],pp159[180],pp159[181],pp159[182],pp159[183],pp159[184],pp159[185],pp159[186],pp159[187],pp159[188],pp159[189],pp159[190],pp159[191],pp159[192],pp159[193],pp159[194],pp159[195]};
    CLA_198 KS_30(s30, c30, in30_1, in30_2);
    wire[195:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp111[47],pp110[49],pp109[51],pp108[53],pp107[55],pp106[57],pp105[59],pp104[61],pp103[63],pp102[65],pp101[67],pp100[69],pp70[100],pp70[101],pp70[102],pp70[103],pp70[104],pp70[105],pp70[106],pp70[107],pp70[108],pp70[109],pp70[110],pp70[111],pp70[112],pp70[113],pp70[114],pp70[115],pp70[116],pp70[117],pp70[118],pp70[119],pp70[120],pp70[121],pp70[122],pp70[123],pp70[124],pp70[125],pp70[126],pp70[127],pp70[128],pp70[129],pp69[131],pp68[133],pp67[135],pp66[137],pp65[139],pp64[141],pp63[143],pp62[145],pp61[147],pp60[149],pp59[151],pp58[153],pp57[155],pp56[157],pp55[159],pp54[161],pp53[163],pp52[165],pp51[167],pp50[169],pp49[171],pp48[173],pp47[175],pp46[177],pp45[179],pp44[181],pp43[183],pp42[185],pp41[187],pp40[189],pp39[191],pp38[193],pp37[195],pp36[197],pp35[199],pp34[201],pp33[203],pp32[205],pp31[207],pp30[209],pp29[211],pp28[213],pp27[215],pp26[217],pp25[219],pp24[221],pp23[223],pp22[225],pp21[227],pp20[229],pp19[231],pp18[233],pp17[235],pp16[237],pp15[239],pp14[241],pp13[243],pp12[245],pp11[247],pp10[249],pp160[100],pp160[101],pp160[102],pp160[103],pp160[104],pp160[105],pp160[106],pp160[107],pp160[108],pp160[109],pp160[110],pp160[111],pp160[112],pp160[113],pp160[114],pp160[115],pp160[116],pp160[117],pp160[118],pp160[119],pp160[120],pp160[121],pp160[122],pp160[123],pp160[124],pp160[125],pp160[126],pp160[127],pp160[128],pp160[129],pp160[130],pp160[131],pp160[132],pp160[133],pp160[134],pp160[135],pp160[136],pp160[137],pp160[138],pp160[139],pp160[140],pp160[141],pp160[142],pp160[143],pp160[144],pp160[145],pp160[146],pp160[147],pp160[148],pp160[149],pp160[150],pp160[151],pp160[152],pp160[153],pp160[154],pp160[155],pp160[156],pp160[157],pp160[158],pp160[159],pp160[160],pp160[161],pp160[162],pp160[163],pp160[164],pp160[165],pp160[166],pp160[167],pp160[168],pp160[169],pp160[170],pp160[171],pp160[172],pp160[173],pp160[174],pp160[175],pp160[176],pp160[177],pp160[178],pp160[179],pp160[180],pp160[181],pp160[182],pp160[183],pp160[184],pp160[185],pp160[186],pp160[187],pp160[188],pp160[189],pp160[190],pp160[191],pp160[192],pp160[193]};
    assign in31_2 = {pp112[46],pp111[48],pp110[50],pp109[52],pp108[54],pp107[56],pp106[58],pp105[60],pp104[62],pp103[64],pp102[66],pp101[68],pp100[70],pp71[100],pp71[101],pp71[102],pp71[103],pp71[104],pp71[105],pp71[106],pp71[107],pp71[108],pp71[109],pp71[110],pp71[111],pp71[112],pp71[113],pp71[114],pp71[115],pp71[116],pp71[117],pp71[118],pp71[119],pp71[120],pp71[121],pp71[122],pp71[123],pp71[124],pp71[125],pp71[126],pp71[127],pp71[128],pp70[130],pp69[132],pp68[134],pp67[136],pp66[138],pp65[140],pp64[142],pp63[144],pp62[146],pp61[148],pp60[150],pp59[152],pp58[154],pp57[156],pp56[158],pp55[160],pp54[162],pp53[164],pp52[166],pp51[168],pp50[170],pp49[172],pp48[174],pp47[176],pp46[178],pp45[180],pp44[182],pp43[184],pp42[186],pp41[188],pp40[190],pp39[192],pp38[194],pp37[196],pp36[198],pp35[200],pp34[202],pp33[204],pp32[206],pp31[208],pp30[210],pp29[212],pp28[214],pp27[216],pp26[218],pp25[220],pp24[222],pp23[224],pp22[226],pp21[228],pp20[230],pp19[232],pp18[234],pp17[236],pp16[238],pp15[240],pp14[242],pp13[244],pp12[246],pp11[248],pp10[250],pp161[100],pp161[101],pp161[102],pp161[103],pp161[104],pp161[105],pp161[106],pp161[107],pp161[108],pp161[109],pp161[110],pp161[111],pp161[112],pp161[113],pp161[114],pp161[115],pp161[116],pp161[117],pp161[118],pp161[119],pp161[120],pp161[121],pp161[122],pp161[123],pp161[124],pp161[125],pp161[126],pp161[127],pp161[128],pp161[129],pp161[130],pp161[131],pp161[132],pp161[133],pp161[134],pp161[135],pp161[136],pp161[137],pp161[138],pp161[139],pp161[140],pp161[141],pp161[142],pp161[143],pp161[144],pp161[145],pp161[146],pp161[147],pp161[148],pp161[149],pp161[150],pp161[151],pp161[152],pp161[153],pp161[154],pp161[155],pp161[156],pp161[157],pp161[158],pp161[159],pp161[160],pp161[161],pp161[162],pp161[163],pp161[164],pp161[165],pp161[166],pp161[167],pp161[168],pp161[169],pp161[170],pp161[171],pp161[172],pp161[173],pp161[174],pp161[175],pp161[176],pp161[177],pp161[178],pp161[179],pp161[180],pp161[181],pp161[182],pp161[183],pp161[184],pp161[185],pp161[186],pp161[187],pp161[188],pp161[189],pp161[190],pp161[191],pp161[192]};
    CLA_196 KS_31(s31, c31, in31_1, in31_2);
    wire[193:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp112[47],pp111[49],pp110[51],pp109[53],pp108[55],pp107[57],pp106[59],pp105[61],pp104[63],pp103[65],pp102[67],pp101[69],pp100[71],pp72[100],pp72[101],pp72[102],pp72[103],pp72[104],pp72[105],pp72[106],pp72[107],pp72[108],pp72[109],pp72[110],pp72[111],pp72[112],pp72[113],pp72[114],pp72[115],pp72[116],pp72[117],pp72[118],pp72[119],pp72[120],pp72[121],pp72[122],pp72[123],pp72[124],pp72[125],pp72[126],pp72[127],pp71[129],pp70[131],pp69[133],pp68[135],pp67[137],pp66[139],pp65[141],pp64[143],pp63[145],pp62[147],pp61[149],pp60[151],pp59[153],pp58[155],pp57[157],pp56[159],pp55[161],pp54[163],pp53[165],pp52[167],pp51[169],pp50[171],pp49[173],pp48[175],pp47[177],pp46[179],pp45[181],pp44[183],pp43[185],pp42[187],pp41[189],pp40[191],pp39[193],pp38[195],pp37[197],pp36[199],pp35[201],pp34[203],pp33[205],pp32[207],pp31[209],pp30[211],pp29[213],pp28[215],pp27[217],pp26[219],pp25[221],pp24[223],pp23[225],pp22[227],pp21[229],pp20[231],pp19[233],pp18[235],pp17[237],pp16[239],pp15[241],pp14[243],pp13[245],pp12[247],pp11[249],pp10[251],pp162[100],pp162[101],pp162[102],pp162[103],pp162[104],pp162[105],pp162[106],pp162[107],pp162[108],pp162[109],pp162[110],pp162[111],pp162[112],pp162[113],pp162[114],pp162[115],pp162[116],pp162[117],pp162[118],pp162[119],pp162[120],pp162[121],pp162[122],pp162[123],pp162[124],pp162[125],pp162[126],pp162[127],pp162[128],pp162[129],pp162[130],pp162[131],pp162[132],pp162[133],pp162[134],pp162[135],pp162[136],pp162[137],pp162[138],pp162[139],pp162[140],pp162[141],pp162[142],pp162[143],pp162[144],pp162[145],pp162[146],pp162[147],pp162[148],pp162[149],pp162[150],pp162[151],pp162[152],pp162[153],pp162[154],pp162[155],pp162[156],pp162[157],pp162[158],pp162[159],pp162[160],pp162[161],pp162[162],pp162[163],pp162[164],pp162[165],pp162[166],pp162[167],pp162[168],pp162[169],pp162[170],pp162[171],pp162[172],pp162[173],pp162[174],pp162[175],pp162[176],pp162[177],pp162[178],pp162[179],pp162[180],pp162[181],pp162[182],pp162[183],pp162[184],pp162[185],pp162[186],pp162[187],pp162[188],pp162[189],pp162[190]};
    assign in32_2 = {pp113[46],pp112[48],pp111[50],pp110[52],pp109[54],pp108[56],pp107[58],pp106[60],pp105[62],pp104[64],pp103[66],pp102[68],pp101[70],pp100[72],pp73[100],pp73[101],pp73[102],pp73[103],pp73[104],pp73[105],pp73[106],pp73[107],pp73[108],pp73[109],pp73[110],pp73[111],pp73[112],pp73[113],pp73[114],pp73[115],pp73[116],pp73[117],pp73[118],pp73[119],pp73[120],pp73[121],pp73[122],pp73[123],pp73[124],pp73[125],pp73[126],pp72[128],pp71[130],pp70[132],pp69[134],pp68[136],pp67[138],pp66[140],pp65[142],pp64[144],pp63[146],pp62[148],pp61[150],pp60[152],pp59[154],pp58[156],pp57[158],pp56[160],pp55[162],pp54[164],pp53[166],pp52[168],pp51[170],pp50[172],pp49[174],pp48[176],pp47[178],pp46[180],pp45[182],pp44[184],pp43[186],pp42[188],pp41[190],pp40[192],pp39[194],pp38[196],pp37[198],pp36[200],pp35[202],pp34[204],pp33[206],pp32[208],pp31[210],pp30[212],pp29[214],pp28[216],pp27[218],pp26[220],pp25[222],pp24[224],pp23[226],pp22[228],pp21[230],pp20[232],pp19[234],pp18[236],pp17[238],pp16[240],pp15[242],pp14[244],pp13[246],pp12[248],pp11[250],pp10[252],pp163[100],pp163[101],pp163[102],pp163[103],pp163[104],pp163[105],pp163[106],pp163[107],pp163[108],pp163[109],pp163[110],pp163[111],pp163[112],pp163[113],pp163[114],pp163[115],pp163[116],pp163[117],pp163[118],pp163[119],pp163[120],pp163[121],pp163[122],pp163[123],pp163[124],pp163[125],pp163[126],pp163[127],pp163[128],pp163[129],pp163[130],pp163[131],pp163[132],pp163[133],pp163[134],pp163[135],pp163[136],pp163[137],pp163[138],pp163[139],pp163[140],pp163[141],pp163[142],pp163[143],pp163[144],pp163[145],pp163[146],pp163[147],pp163[148],pp163[149],pp163[150],pp163[151],pp163[152],pp163[153],pp163[154],pp163[155],pp163[156],pp163[157],pp163[158],pp163[159],pp163[160],pp163[161],pp163[162],pp163[163],pp163[164],pp163[165],pp163[166],pp163[167],pp163[168],pp163[169],pp163[170],pp163[171],pp163[172],pp163[173],pp163[174],pp163[175],pp163[176],pp163[177],pp163[178],pp163[179],pp163[180],pp163[181],pp163[182],pp163[183],pp163[184],pp163[185],pp163[186],pp163[187],pp163[188],pp163[189]};
    CLA_194 KS_32(s32, c32, in32_1, in32_2);
    wire[191:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp113[47],pp112[49],pp111[51],pp110[53],pp109[55],pp108[57],pp107[59],pp106[61],pp105[63],pp104[65],pp103[67],pp102[69],pp101[71],pp100[73],pp74[100],pp74[101],pp74[102],pp74[103],pp74[104],pp74[105],pp74[106],pp74[107],pp74[108],pp74[109],pp74[110],pp74[111],pp74[112],pp74[113],pp74[114],pp74[115],pp74[116],pp74[117],pp74[118],pp74[119],pp74[120],pp74[121],pp74[122],pp74[123],pp74[124],pp74[125],pp73[127],pp72[129],pp71[131],pp70[133],pp69[135],pp68[137],pp67[139],pp66[141],pp65[143],pp64[145],pp63[147],pp62[149],pp61[151],pp60[153],pp59[155],pp58[157],pp57[159],pp56[161],pp55[163],pp54[165],pp53[167],pp52[169],pp51[171],pp50[173],pp49[175],pp48[177],pp47[179],pp46[181],pp45[183],pp44[185],pp43[187],pp42[189],pp41[191],pp40[193],pp39[195],pp38[197],pp37[199],pp36[201],pp35[203],pp34[205],pp33[207],pp32[209],pp31[211],pp30[213],pp29[215],pp28[217],pp27[219],pp26[221],pp25[223],pp24[225],pp23[227],pp22[229],pp21[231],pp20[233],pp19[235],pp18[237],pp17[239],pp16[241],pp15[243],pp14[245],pp13[247],pp12[249],pp11[251],pp10[253],pp164[100],pp164[101],pp164[102],pp164[103],pp164[104],pp164[105],pp164[106],pp164[107],pp164[108],pp164[109],pp164[110],pp164[111],pp164[112],pp164[113],pp164[114],pp164[115],pp164[116],pp164[117],pp164[118],pp164[119],pp164[120],pp164[121],pp164[122],pp164[123],pp164[124],pp164[125],pp164[126],pp164[127],pp164[128],pp164[129],pp164[130],pp164[131],pp164[132],pp164[133],pp164[134],pp164[135],pp164[136],pp164[137],pp164[138],pp164[139],pp164[140],pp164[141],pp164[142],pp164[143],pp164[144],pp164[145],pp164[146],pp164[147],pp164[148],pp164[149],pp164[150],pp164[151],pp164[152],pp164[153],pp164[154],pp164[155],pp164[156],pp164[157],pp164[158],pp164[159],pp164[160],pp164[161],pp164[162],pp164[163],pp164[164],pp164[165],pp164[166],pp164[167],pp164[168],pp164[169],pp164[170],pp164[171],pp164[172],pp164[173],pp164[174],pp164[175],pp164[176],pp164[177],pp164[178],pp164[179],pp164[180],pp164[181],pp164[182],pp164[183],pp164[184],pp164[185],pp164[186],pp164[187]};
    assign in33_2 = {pp114[46],pp113[48],pp112[50],pp111[52],pp110[54],pp109[56],pp108[58],pp107[60],pp106[62],pp105[64],pp104[66],pp103[68],pp102[70],pp101[72],pp100[74],pp75[100],pp75[101],pp75[102],pp75[103],pp75[104],pp75[105],pp75[106],pp75[107],pp75[108],pp75[109],pp75[110],pp75[111],pp75[112],pp75[113],pp75[114],pp75[115],pp75[116],pp75[117],pp75[118],pp75[119],pp75[120],pp75[121],pp75[122],pp75[123],pp75[124],pp74[126],pp73[128],pp72[130],pp71[132],pp70[134],pp69[136],pp68[138],pp67[140],pp66[142],pp65[144],pp64[146],pp63[148],pp62[150],pp61[152],pp60[154],pp59[156],pp58[158],pp57[160],pp56[162],pp55[164],pp54[166],pp53[168],pp52[170],pp51[172],pp50[174],pp49[176],pp48[178],pp47[180],pp46[182],pp45[184],pp44[186],pp43[188],pp42[190],pp41[192],pp40[194],pp39[196],pp38[198],pp37[200],pp36[202],pp35[204],pp34[206],pp33[208],pp32[210],pp31[212],pp30[214],pp29[216],pp28[218],pp27[220],pp26[222],pp25[224],pp24[226],pp23[228],pp22[230],pp21[232],pp20[234],pp19[236],pp18[238],pp17[240],pp16[242],pp15[244],pp14[246],pp13[248],pp12[250],pp11[252],pp10[254],pp165[100],pp165[101],pp165[102],pp165[103],pp165[104],pp165[105],pp165[106],pp165[107],pp165[108],pp165[109],pp165[110],pp165[111],pp165[112],pp165[113],pp165[114],pp165[115],pp165[116],pp165[117],pp165[118],pp165[119],pp165[120],pp165[121],pp165[122],pp165[123],pp165[124],pp165[125],pp165[126],pp165[127],pp165[128],pp165[129],pp165[130],pp165[131],pp165[132],pp165[133],pp165[134],pp165[135],pp165[136],pp165[137],pp165[138],pp165[139],pp165[140],pp165[141],pp165[142],pp165[143],pp165[144],pp165[145],pp165[146],pp165[147],pp165[148],pp165[149],pp165[150],pp165[151],pp165[152],pp165[153],pp165[154],pp165[155],pp165[156],pp165[157],pp165[158],pp165[159],pp165[160],pp165[161],pp165[162],pp165[163],pp165[164],pp165[165],pp165[166],pp165[167],pp165[168],pp165[169],pp165[170],pp165[171],pp165[172],pp165[173],pp165[174],pp165[175],pp165[176],pp165[177],pp165[178],pp165[179],pp165[180],pp165[181],pp165[182],pp165[183],pp165[184],pp165[185],pp165[186]};
    CLA_192 KS_33(s33, c33, in33_1, in33_2);
    wire[189:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp114[47],pp113[49],pp112[51],pp111[53],pp110[55],pp109[57],pp108[59],pp107[61],pp106[63],pp105[65],pp104[67],pp103[69],pp102[71],pp101[73],pp100[75],pp76[100],pp76[101],pp76[102],pp76[103],pp76[104],pp76[105],pp76[106],pp76[107],pp76[108],pp76[109],pp76[110],pp76[111],pp76[112],pp76[113],pp76[114],pp76[115],pp76[116],pp76[117],pp76[118],pp76[119],pp76[120],pp76[121],pp76[122],pp76[123],pp75[125],pp74[127],pp73[129],pp72[131],pp71[133],pp70[135],pp69[137],pp68[139],pp67[141],pp66[143],pp65[145],pp64[147],pp63[149],pp62[151],pp61[153],pp60[155],pp59[157],pp58[159],pp57[161],pp56[163],pp55[165],pp54[167],pp53[169],pp52[171],pp51[173],pp50[175],pp49[177],pp48[179],pp47[181],pp46[183],pp45[185],pp44[187],pp43[189],pp42[191],pp41[193],pp40[195],pp39[197],pp38[199],pp37[201],pp36[203],pp35[205],pp34[207],pp33[209],pp32[211],pp31[213],pp30[215],pp29[217],pp28[219],pp27[221],pp26[223],pp25[225],pp24[227],pp23[229],pp22[231],pp21[233],pp20[235],pp19[237],pp18[239],pp17[241],pp16[243],pp15[245],pp14[247],pp13[249],pp12[251],pp11[253],pp10[255],pp166[100],pp166[101],pp166[102],pp166[103],pp166[104],pp166[105],pp166[106],pp166[107],pp166[108],pp166[109],pp166[110],pp166[111],pp166[112],pp166[113],pp166[114],pp166[115],pp166[116],pp166[117],pp166[118],pp166[119],pp166[120],pp166[121],pp166[122],pp166[123],pp166[124],pp166[125],pp166[126],pp166[127],pp166[128],pp166[129],pp166[130],pp166[131],pp166[132],pp166[133],pp166[134],pp166[135],pp166[136],pp166[137],pp166[138],pp166[139],pp166[140],pp166[141],pp166[142],pp166[143],pp166[144],pp166[145],pp166[146],pp166[147],pp166[148],pp166[149],pp166[150],pp166[151],pp166[152],pp166[153],pp166[154],pp166[155],pp166[156],pp166[157],pp166[158],pp166[159],pp166[160],pp166[161],pp166[162],pp166[163],pp166[164],pp166[165],pp166[166],pp166[167],pp166[168],pp166[169],pp166[170],pp166[171],pp166[172],pp166[173],pp166[174],pp166[175],pp166[176],pp166[177],pp166[178],pp166[179],pp166[180],pp166[181],pp166[182],pp166[183],pp166[184]};
    assign in34_2 = {pp115[46],pp114[48],pp113[50],pp112[52],pp111[54],pp110[56],pp109[58],pp108[60],pp107[62],pp106[64],pp105[66],pp104[68],pp103[70],pp102[72],pp101[74],pp100[76],pp77[100],pp77[101],pp77[102],pp77[103],pp77[104],pp77[105],pp77[106],pp77[107],pp77[108],pp77[109],pp77[110],pp77[111],pp77[112],pp77[113],pp77[114],pp77[115],pp77[116],pp77[117],pp77[118],pp77[119],pp77[120],pp77[121],pp77[122],pp76[124],pp75[126],pp74[128],pp73[130],pp72[132],pp71[134],pp70[136],pp69[138],pp68[140],pp67[142],pp66[144],pp65[146],pp64[148],pp63[150],pp62[152],pp61[154],pp60[156],pp59[158],pp58[160],pp57[162],pp56[164],pp55[166],pp54[168],pp53[170],pp52[172],pp51[174],pp50[176],pp49[178],pp48[180],pp47[182],pp46[184],pp45[186],pp44[188],pp43[190],pp42[192],pp41[194],pp40[196],pp39[198],pp38[200],pp37[202],pp36[204],pp35[206],pp34[208],pp33[210],pp32[212],pp31[214],pp30[216],pp29[218],pp28[220],pp27[222],pp26[224],pp25[226],pp24[228],pp23[230],pp22[232],pp21[234],pp20[236],pp19[238],pp18[240],pp17[242],pp16[244],pp15[246],pp14[248],pp13[250],pp12[252],pp11[254],pp11[255],pp167[100],pp167[101],pp167[102],pp167[103],pp167[104],pp167[105],pp167[106],pp167[107],pp167[108],pp167[109],pp167[110],pp167[111],pp167[112],pp167[113],pp167[114],pp167[115],pp167[116],pp167[117],pp167[118],pp167[119],pp167[120],pp167[121],pp167[122],pp167[123],pp167[124],pp167[125],pp167[126],pp167[127],pp167[128],pp167[129],pp167[130],pp167[131],pp167[132],pp167[133],pp167[134],pp167[135],pp167[136],pp167[137],pp167[138],pp167[139],pp167[140],pp167[141],pp167[142],pp167[143],pp167[144],pp167[145],pp167[146],pp167[147],pp167[148],pp167[149],pp167[150],pp167[151],pp167[152],pp167[153],pp167[154],pp167[155],pp167[156],pp167[157],pp167[158],pp167[159],pp167[160],pp167[161],pp167[162],pp167[163],pp167[164],pp167[165],pp167[166],pp167[167],pp167[168],pp167[169],pp167[170],pp167[171],pp167[172],pp167[173],pp167[174],pp167[175],pp167[176],pp167[177],pp167[178],pp167[179],pp167[180],pp167[181],pp167[182],pp167[183]};
    CLA_190 KS_34(s34, c34, in34_1, in34_2);
    wire[187:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp115[47],pp114[49],pp113[51],pp112[53],pp111[55],pp110[57],pp109[59],pp108[61],pp107[63],pp106[65],pp105[67],pp104[69],pp103[71],pp102[73],pp101[75],pp100[77],pp78[100],pp78[101],pp78[102],pp78[103],pp78[104],pp78[105],pp78[106],pp78[107],pp78[108],pp78[109],pp78[110],pp78[111],pp78[112],pp78[113],pp78[114],pp78[115],pp78[116],pp78[117],pp78[118],pp78[119],pp78[120],pp78[121],pp77[123],pp76[125],pp75[127],pp74[129],pp73[131],pp72[133],pp71[135],pp70[137],pp69[139],pp68[141],pp67[143],pp66[145],pp65[147],pp64[149],pp63[151],pp62[153],pp61[155],pp60[157],pp59[159],pp58[161],pp57[163],pp56[165],pp55[167],pp54[169],pp53[171],pp52[173],pp51[175],pp50[177],pp49[179],pp48[181],pp47[183],pp46[185],pp45[187],pp44[189],pp43[191],pp42[193],pp41[195],pp40[197],pp39[199],pp38[201],pp37[203],pp36[205],pp35[207],pp34[209],pp33[211],pp32[213],pp31[215],pp30[217],pp29[219],pp28[221],pp27[223],pp26[225],pp25[227],pp24[229],pp23[231],pp22[233],pp21[235],pp20[237],pp19[239],pp18[241],pp17[243],pp16[245],pp15[247],pp14[249],pp13[251],pp12[253],pp12[254],pp12[255],pp168[100],pp168[101],pp168[102],pp168[103],pp168[104],pp168[105],pp168[106],pp168[107],pp168[108],pp168[109],pp168[110],pp168[111],pp168[112],pp168[113],pp168[114],pp168[115],pp168[116],pp168[117],pp168[118],pp168[119],pp168[120],pp168[121],pp168[122],pp168[123],pp168[124],pp168[125],pp168[126],pp168[127],pp168[128],pp168[129],pp168[130],pp168[131],pp168[132],pp168[133],pp168[134],pp168[135],pp168[136],pp168[137],pp168[138],pp168[139],pp168[140],pp168[141],pp168[142],pp168[143],pp168[144],pp168[145],pp168[146],pp168[147],pp168[148],pp168[149],pp168[150],pp168[151],pp168[152],pp168[153],pp168[154],pp168[155],pp168[156],pp168[157],pp168[158],pp168[159],pp168[160],pp168[161],pp168[162],pp168[163],pp168[164],pp168[165],pp168[166],pp168[167],pp168[168],pp168[169],pp168[170],pp168[171],pp168[172],pp168[173],pp168[174],pp168[175],pp168[176],pp168[177],pp168[178],pp168[179],pp168[180],pp168[181]};
    assign in35_2 = {pp116[46],pp115[48],pp114[50],pp113[52],pp112[54],pp111[56],pp110[58],pp109[60],pp108[62],pp107[64],pp106[66],pp105[68],pp104[70],pp103[72],pp102[74],pp101[76],pp100[78],pp79[100],pp79[101],pp79[102],pp79[103],pp79[104],pp79[105],pp79[106],pp79[107],pp79[108],pp79[109],pp79[110],pp79[111],pp79[112],pp79[113],pp79[114],pp79[115],pp79[116],pp79[117],pp79[118],pp79[119],pp79[120],pp78[122],pp77[124],pp76[126],pp75[128],pp74[130],pp73[132],pp72[134],pp71[136],pp70[138],pp69[140],pp68[142],pp67[144],pp66[146],pp65[148],pp64[150],pp63[152],pp62[154],pp61[156],pp60[158],pp59[160],pp58[162],pp57[164],pp56[166],pp55[168],pp54[170],pp53[172],pp52[174],pp51[176],pp50[178],pp49[180],pp48[182],pp47[184],pp46[186],pp45[188],pp44[190],pp43[192],pp42[194],pp41[196],pp40[198],pp39[200],pp38[202],pp37[204],pp36[206],pp35[208],pp34[210],pp33[212],pp32[214],pp31[216],pp30[218],pp29[220],pp28[222],pp27[224],pp26[226],pp25[228],pp24[230],pp23[232],pp22[234],pp21[236],pp20[238],pp19[240],pp18[242],pp17[244],pp16[246],pp15[248],pp14[250],pp13[252],pp13[253],pp13[254],pp13[255],pp169[100],pp169[101],pp169[102],pp169[103],pp169[104],pp169[105],pp169[106],pp169[107],pp169[108],pp169[109],pp169[110],pp169[111],pp169[112],pp169[113],pp169[114],pp169[115],pp169[116],pp169[117],pp169[118],pp169[119],pp169[120],pp169[121],pp169[122],pp169[123],pp169[124],pp169[125],pp169[126],pp169[127],pp169[128],pp169[129],pp169[130],pp169[131],pp169[132],pp169[133],pp169[134],pp169[135],pp169[136],pp169[137],pp169[138],pp169[139],pp169[140],pp169[141],pp169[142],pp169[143],pp169[144],pp169[145],pp169[146],pp169[147],pp169[148],pp169[149],pp169[150],pp169[151],pp169[152],pp169[153],pp169[154],pp169[155],pp169[156],pp169[157],pp169[158],pp169[159],pp169[160],pp169[161],pp169[162],pp169[163],pp169[164],pp169[165],pp169[166],pp169[167],pp169[168],pp169[169],pp169[170],pp169[171],pp169[172],pp169[173],pp169[174],pp169[175],pp169[176],pp169[177],pp169[178],pp169[179],pp169[180]};
    CLA_188 KS_35(s35, c35, in35_1, in35_2);
    wire[185:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp116[47],pp115[49],pp114[51],pp113[53],pp112[55],pp111[57],pp110[59],pp109[61],pp108[63],pp107[65],pp106[67],pp105[69],pp104[71],pp103[73],pp102[75],pp101[77],pp100[79],pp80[100],pp80[101],pp80[102],pp80[103],pp80[104],pp80[105],pp80[106],pp80[107],pp80[108],pp80[109],pp80[110],pp80[111],pp80[112],pp80[113],pp80[114],pp80[115],pp80[116],pp80[117],pp80[118],pp80[119],pp79[121],pp78[123],pp77[125],pp76[127],pp75[129],pp74[131],pp73[133],pp72[135],pp71[137],pp70[139],pp69[141],pp68[143],pp67[145],pp66[147],pp65[149],pp64[151],pp63[153],pp62[155],pp61[157],pp60[159],pp59[161],pp58[163],pp57[165],pp56[167],pp55[169],pp54[171],pp53[173],pp52[175],pp51[177],pp50[179],pp49[181],pp48[183],pp47[185],pp46[187],pp45[189],pp44[191],pp43[193],pp42[195],pp41[197],pp40[199],pp39[201],pp38[203],pp37[205],pp36[207],pp35[209],pp34[211],pp33[213],pp32[215],pp31[217],pp30[219],pp29[221],pp28[223],pp27[225],pp26[227],pp25[229],pp24[231],pp23[233],pp22[235],pp21[237],pp20[239],pp19[241],pp18[243],pp17[245],pp16[247],pp15[249],pp14[251],pp14[252],pp14[253],pp14[254],pp14[255],pp170[100],pp170[101],pp170[102],pp170[103],pp170[104],pp170[105],pp170[106],pp170[107],pp170[108],pp170[109],pp170[110],pp170[111],pp170[112],pp170[113],pp170[114],pp170[115],pp170[116],pp170[117],pp170[118],pp170[119],pp170[120],pp170[121],pp170[122],pp170[123],pp170[124],pp170[125],pp170[126],pp170[127],pp170[128],pp170[129],pp170[130],pp170[131],pp170[132],pp170[133],pp170[134],pp170[135],pp170[136],pp170[137],pp170[138],pp170[139],pp170[140],pp170[141],pp170[142],pp170[143],pp170[144],pp170[145],pp170[146],pp170[147],pp170[148],pp170[149],pp170[150],pp170[151],pp170[152],pp170[153],pp170[154],pp170[155],pp170[156],pp170[157],pp170[158],pp170[159],pp170[160],pp170[161],pp170[162],pp170[163],pp170[164],pp170[165],pp170[166],pp170[167],pp170[168],pp170[169],pp170[170],pp170[171],pp170[172],pp170[173],pp170[174],pp170[175],pp170[176],pp170[177],pp170[178]};
    assign in36_2 = {pp117[46],pp116[48],pp115[50],pp114[52],pp113[54],pp112[56],pp111[58],pp110[60],pp109[62],pp108[64],pp107[66],pp106[68],pp105[70],pp104[72],pp103[74],pp102[76],pp101[78],pp100[80],pp81[100],pp81[101],pp81[102],pp81[103],pp81[104],pp81[105],pp81[106],pp81[107],pp81[108],pp81[109],pp81[110],pp81[111],pp81[112],pp81[113],pp81[114],pp81[115],pp81[116],pp81[117],pp81[118],pp80[120],pp79[122],pp78[124],pp77[126],pp76[128],pp75[130],pp74[132],pp73[134],pp72[136],pp71[138],pp70[140],pp69[142],pp68[144],pp67[146],pp66[148],pp65[150],pp64[152],pp63[154],pp62[156],pp61[158],pp60[160],pp59[162],pp58[164],pp57[166],pp56[168],pp55[170],pp54[172],pp53[174],pp52[176],pp51[178],pp50[180],pp49[182],pp48[184],pp47[186],pp46[188],pp45[190],pp44[192],pp43[194],pp42[196],pp41[198],pp40[200],pp39[202],pp38[204],pp37[206],pp36[208],pp35[210],pp34[212],pp33[214],pp32[216],pp31[218],pp30[220],pp29[222],pp28[224],pp27[226],pp26[228],pp25[230],pp24[232],pp23[234],pp22[236],pp21[238],pp20[240],pp19[242],pp18[244],pp17[246],pp16[248],pp15[250],pp15[251],pp15[252],pp15[253],pp15[254],pp15[255],pp171[100],pp171[101],pp171[102],pp171[103],pp171[104],pp171[105],pp171[106],pp171[107],pp171[108],pp171[109],pp171[110],pp171[111],pp171[112],pp171[113],pp171[114],pp171[115],pp171[116],pp171[117],pp171[118],pp171[119],pp171[120],pp171[121],pp171[122],pp171[123],pp171[124],pp171[125],pp171[126],pp171[127],pp171[128],pp171[129],pp171[130],pp171[131],pp171[132],pp171[133],pp171[134],pp171[135],pp171[136],pp171[137],pp171[138],pp171[139],pp171[140],pp171[141],pp171[142],pp171[143],pp171[144],pp171[145],pp171[146],pp171[147],pp171[148],pp171[149],pp171[150],pp171[151],pp171[152],pp171[153],pp171[154],pp171[155],pp171[156],pp171[157],pp171[158],pp171[159],pp171[160],pp171[161],pp171[162],pp171[163],pp171[164],pp171[165],pp171[166],pp171[167],pp171[168],pp171[169],pp171[170],pp171[171],pp171[172],pp171[173],pp171[174],pp171[175],pp171[176],pp171[177]};
    CLA_186 KS_36(s36, c36, in36_1, in36_2);
    wire[183:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp117[47],pp116[49],pp115[51],pp114[53],pp113[55],pp112[57],pp111[59],pp110[61],pp109[63],pp108[65],pp107[67],pp106[69],pp105[71],pp104[73],pp103[75],pp102[77],pp101[79],pp100[81],pp82[100],pp82[101],pp82[102],pp82[103],pp82[104],pp82[105],pp82[106],pp82[107],pp82[108],pp82[109],pp82[110],pp82[111],pp82[112],pp82[113],pp82[114],pp82[115],pp82[116],pp82[117],pp81[119],pp80[121],pp79[123],pp78[125],pp77[127],pp76[129],pp75[131],pp74[133],pp73[135],pp72[137],pp71[139],pp70[141],pp69[143],pp68[145],pp67[147],pp66[149],pp65[151],pp64[153],pp63[155],pp62[157],pp61[159],pp60[161],pp59[163],pp58[165],pp57[167],pp56[169],pp55[171],pp54[173],pp53[175],pp52[177],pp51[179],pp50[181],pp49[183],pp48[185],pp47[187],pp46[189],pp45[191],pp44[193],pp43[195],pp42[197],pp41[199],pp40[201],pp39[203],pp38[205],pp37[207],pp36[209],pp35[211],pp34[213],pp33[215],pp32[217],pp31[219],pp30[221],pp29[223],pp28[225],pp27[227],pp26[229],pp25[231],pp24[233],pp23[235],pp22[237],pp21[239],pp20[241],pp19[243],pp18[245],pp17[247],pp16[249],pp16[250],pp16[251],pp16[252],pp16[253],pp16[254],pp16[255],pp172[100],pp172[101],pp172[102],pp172[103],pp172[104],pp172[105],pp172[106],pp172[107],pp172[108],pp172[109],pp172[110],pp172[111],pp172[112],pp172[113],pp172[114],pp172[115],pp172[116],pp172[117],pp172[118],pp172[119],pp172[120],pp172[121],pp172[122],pp172[123],pp172[124],pp172[125],pp172[126],pp172[127],pp172[128],pp172[129],pp172[130],pp172[131],pp172[132],pp172[133],pp172[134],pp172[135],pp172[136],pp172[137],pp172[138],pp172[139],pp172[140],pp172[141],pp172[142],pp172[143],pp172[144],pp172[145],pp172[146],pp172[147],pp172[148],pp172[149],pp172[150],pp172[151],pp172[152],pp172[153],pp172[154],pp172[155],pp172[156],pp172[157],pp172[158],pp172[159],pp172[160],pp172[161],pp172[162],pp172[163],pp172[164],pp172[165],pp172[166],pp172[167],pp172[168],pp172[169],pp172[170],pp172[171],pp172[172],pp172[173],pp172[174],pp172[175]};
    assign in37_2 = {pp118[46],pp117[48],pp116[50],pp115[52],pp114[54],pp113[56],pp112[58],pp111[60],pp110[62],pp109[64],pp108[66],pp107[68],pp106[70],pp105[72],pp104[74],pp103[76],pp102[78],pp101[80],pp100[82],pp83[100],pp83[101],pp83[102],pp83[103],pp83[104],pp83[105],pp83[106],pp83[107],pp83[108],pp83[109],pp83[110],pp83[111],pp83[112],pp83[113],pp83[114],pp83[115],pp83[116],pp82[118],pp81[120],pp80[122],pp79[124],pp78[126],pp77[128],pp76[130],pp75[132],pp74[134],pp73[136],pp72[138],pp71[140],pp70[142],pp69[144],pp68[146],pp67[148],pp66[150],pp65[152],pp64[154],pp63[156],pp62[158],pp61[160],pp60[162],pp59[164],pp58[166],pp57[168],pp56[170],pp55[172],pp54[174],pp53[176],pp52[178],pp51[180],pp50[182],pp49[184],pp48[186],pp47[188],pp46[190],pp45[192],pp44[194],pp43[196],pp42[198],pp41[200],pp40[202],pp39[204],pp38[206],pp37[208],pp36[210],pp35[212],pp34[214],pp33[216],pp32[218],pp31[220],pp30[222],pp29[224],pp28[226],pp27[228],pp26[230],pp25[232],pp24[234],pp23[236],pp22[238],pp21[240],pp20[242],pp19[244],pp18[246],pp17[248],pp17[249],pp17[250],pp17[251],pp17[252],pp17[253],pp17[254],pp17[255],pp173[100],pp173[101],pp173[102],pp173[103],pp173[104],pp173[105],pp173[106],pp173[107],pp173[108],pp173[109],pp173[110],pp173[111],pp173[112],pp173[113],pp173[114],pp173[115],pp173[116],pp173[117],pp173[118],pp173[119],pp173[120],pp173[121],pp173[122],pp173[123],pp173[124],pp173[125],pp173[126],pp173[127],pp173[128],pp173[129],pp173[130],pp173[131],pp173[132],pp173[133],pp173[134],pp173[135],pp173[136],pp173[137],pp173[138],pp173[139],pp173[140],pp173[141],pp173[142],pp173[143],pp173[144],pp173[145],pp173[146],pp173[147],pp173[148],pp173[149],pp173[150],pp173[151],pp173[152],pp173[153],pp173[154],pp173[155],pp173[156],pp173[157],pp173[158],pp173[159],pp173[160],pp173[161],pp173[162],pp173[163],pp173[164],pp173[165],pp173[166],pp173[167],pp173[168],pp173[169],pp173[170],pp173[171],pp173[172],pp173[173],pp173[174]};
    CLA_184 KS_37(s37, c37, in37_1, in37_2);
    wire[181:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp118[47],pp117[49],pp116[51],pp115[53],pp114[55],pp113[57],pp112[59],pp111[61],pp110[63],pp109[65],pp108[67],pp107[69],pp106[71],pp105[73],pp104[75],pp103[77],pp102[79],pp101[81],pp100[83],pp84[100],pp84[101],pp84[102],pp84[103],pp84[104],pp84[105],pp84[106],pp84[107],pp84[108],pp84[109],pp84[110],pp84[111],pp84[112],pp84[113],pp84[114],pp84[115],pp83[117],pp82[119],pp81[121],pp80[123],pp79[125],pp78[127],pp77[129],pp76[131],pp75[133],pp74[135],pp73[137],pp72[139],pp71[141],pp70[143],pp69[145],pp68[147],pp67[149],pp66[151],pp65[153],pp64[155],pp63[157],pp62[159],pp61[161],pp60[163],pp59[165],pp58[167],pp57[169],pp56[171],pp55[173],pp54[175],pp53[177],pp52[179],pp51[181],pp50[183],pp49[185],pp48[187],pp47[189],pp46[191],pp45[193],pp44[195],pp43[197],pp42[199],pp41[201],pp40[203],pp39[205],pp38[207],pp37[209],pp36[211],pp35[213],pp34[215],pp33[217],pp32[219],pp31[221],pp30[223],pp29[225],pp28[227],pp27[229],pp26[231],pp25[233],pp24[235],pp23[237],pp22[239],pp21[241],pp20[243],pp19[245],pp18[247],pp18[248],pp18[249],pp18[250],pp18[251],pp18[252],pp18[253],pp18[254],pp18[255],pp174[100],pp174[101],pp174[102],pp174[103],pp174[104],pp174[105],pp174[106],pp174[107],pp174[108],pp174[109],pp174[110],pp174[111],pp174[112],pp174[113],pp174[114],pp174[115],pp174[116],pp174[117],pp174[118],pp174[119],pp174[120],pp174[121],pp174[122],pp174[123],pp174[124],pp174[125],pp174[126],pp174[127],pp174[128],pp174[129],pp174[130],pp174[131],pp174[132],pp174[133],pp174[134],pp174[135],pp174[136],pp174[137],pp174[138],pp174[139],pp174[140],pp174[141],pp174[142],pp174[143],pp174[144],pp174[145],pp174[146],pp174[147],pp174[148],pp174[149],pp174[150],pp174[151],pp174[152],pp174[153],pp174[154],pp174[155],pp174[156],pp174[157],pp174[158],pp174[159],pp174[160],pp174[161],pp174[162],pp174[163],pp174[164],pp174[165],pp174[166],pp174[167],pp174[168],pp174[169],pp174[170],pp174[171],pp174[172]};
    assign in38_2 = {pp119[46],pp118[48],pp117[50],pp116[52],pp115[54],pp114[56],pp113[58],pp112[60],pp111[62],pp110[64],pp109[66],pp108[68],pp107[70],pp106[72],pp105[74],pp104[76],pp103[78],pp102[80],pp101[82],pp100[84],pp85[100],pp85[101],pp85[102],pp85[103],pp85[104],pp85[105],pp85[106],pp85[107],pp85[108],pp85[109],pp85[110],pp85[111],pp85[112],pp85[113],pp85[114],pp84[116],pp83[118],pp82[120],pp81[122],pp80[124],pp79[126],pp78[128],pp77[130],pp76[132],pp75[134],pp74[136],pp73[138],pp72[140],pp71[142],pp70[144],pp69[146],pp68[148],pp67[150],pp66[152],pp65[154],pp64[156],pp63[158],pp62[160],pp61[162],pp60[164],pp59[166],pp58[168],pp57[170],pp56[172],pp55[174],pp54[176],pp53[178],pp52[180],pp51[182],pp50[184],pp49[186],pp48[188],pp47[190],pp46[192],pp45[194],pp44[196],pp43[198],pp42[200],pp41[202],pp40[204],pp39[206],pp38[208],pp37[210],pp36[212],pp35[214],pp34[216],pp33[218],pp32[220],pp31[222],pp30[224],pp29[226],pp28[228],pp27[230],pp26[232],pp25[234],pp24[236],pp23[238],pp22[240],pp21[242],pp20[244],pp19[246],pp19[247],pp19[248],pp19[249],pp19[250],pp19[251],pp19[252],pp19[253],pp19[254],pp19[255],pp175[100],pp175[101],pp175[102],pp175[103],pp175[104],pp175[105],pp175[106],pp175[107],pp175[108],pp175[109],pp175[110],pp175[111],pp175[112],pp175[113],pp175[114],pp175[115],pp175[116],pp175[117],pp175[118],pp175[119],pp175[120],pp175[121],pp175[122],pp175[123],pp175[124],pp175[125],pp175[126],pp175[127],pp175[128],pp175[129],pp175[130],pp175[131],pp175[132],pp175[133],pp175[134],pp175[135],pp175[136],pp175[137],pp175[138],pp175[139],pp175[140],pp175[141],pp175[142],pp175[143],pp175[144],pp175[145],pp175[146],pp175[147],pp175[148],pp175[149],pp175[150],pp175[151],pp175[152],pp175[153],pp175[154],pp175[155],pp175[156],pp175[157],pp175[158],pp175[159],pp175[160],pp175[161],pp175[162],pp175[163],pp175[164],pp175[165],pp175[166],pp175[167],pp175[168],pp175[169],pp175[170],pp175[171]};
    CLA_182 KS_38(s38, c38, in38_1, in38_2);
    wire[179:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp119[47],pp118[49],pp117[51],pp116[53],pp115[55],pp114[57],pp113[59],pp112[61],pp111[63],pp110[65],pp109[67],pp108[69],pp107[71],pp106[73],pp105[75],pp104[77],pp103[79],pp102[81],pp101[83],pp100[85],pp86[100],pp86[101],pp86[102],pp86[103],pp86[104],pp86[105],pp86[106],pp86[107],pp86[108],pp86[109],pp86[110],pp86[111],pp86[112],pp86[113],pp85[115],pp84[117],pp83[119],pp82[121],pp81[123],pp80[125],pp79[127],pp78[129],pp77[131],pp76[133],pp75[135],pp74[137],pp73[139],pp72[141],pp71[143],pp70[145],pp69[147],pp68[149],pp67[151],pp66[153],pp65[155],pp64[157],pp63[159],pp62[161],pp61[163],pp60[165],pp59[167],pp58[169],pp57[171],pp56[173],pp55[175],pp54[177],pp53[179],pp52[181],pp51[183],pp50[185],pp49[187],pp48[189],pp47[191],pp46[193],pp45[195],pp44[197],pp43[199],pp42[201],pp41[203],pp40[205],pp39[207],pp38[209],pp37[211],pp36[213],pp35[215],pp34[217],pp33[219],pp32[221],pp31[223],pp30[225],pp29[227],pp28[229],pp27[231],pp26[233],pp25[235],pp24[237],pp23[239],pp22[241],pp21[243],pp20[245],pp20[246],pp20[247],pp20[248],pp20[249],pp20[250],pp20[251],pp20[252],pp20[253],pp20[254],pp20[255],pp176[100],pp176[101],pp176[102],pp176[103],pp176[104],pp176[105],pp176[106],pp176[107],pp176[108],pp176[109],pp176[110],pp176[111],pp176[112],pp176[113],pp176[114],pp176[115],pp176[116],pp176[117],pp176[118],pp176[119],pp176[120],pp176[121],pp176[122],pp176[123],pp176[124],pp176[125],pp176[126],pp176[127],pp176[128],pp176[129],pp176[130],pp176[131],pp176[132],pp176[133],pp176[134],pp176[135],pp176[136],pp176[137],pp176[138],pp176[139],pp176[140],pp176[141],pp176[142],pp176[143],pp176[144],pp176[145],pp176[146],pp176[147],pp176[148],pp176[149],pp176[150],pp176[151],pp176[152],pp176[153],pp176[154],pp176[155],pp176[156],pp176[157],pp176[158],pp176[159],pp176[160],pp176[161],pp176[162],pp176[163],pp176[164],pp176[165],pp176[166],pp176[167],pp176[168],pp176[169]};
    assign in39_2 = {pp120[46],pp119[48],pp118[50],pp117[52],pp116[54],pp115[56],pp114[58],pp113[60],pp112[62],pp111[64],pp110[66],pp109[68],pp108[70],pp107[72],pp106[74],pp105[76],pp104[78],pp103[80],pp102[82],pp101[84],pp100[86],pp87[100],pp87[101],pp87[102],pp87[103],pp87[104],pp87[105],pp87[106],pp87[107],pp87[108],pp87[109],pp87[110],pp87[111],pp87[112],pp86[114],pp85[116],pp84[118],pp83[120],pp82[122],pp81[124],pp80[126],pp79[128],pp78[130],pp77[132],pp76[134],pp75[136],pp74[138],pp73[140],pp72[142],pp71[144],pp70[146],pp69[148],pp68[150],pp67[152],pp66[154],pp65[156],pp64[158],pp63[160],pp62[162],pp61[164],pp60[166],pp59[168],pp58[170],pp57[172],pp56[174],pp55[176],pp54[178],pp53[180],pp52[182],pp51[184],pp50[186],pp49[188],pp48[190],pp47[192],pp46[194],pp45[196],pp44[198],pp43[200],pp42[202],pp41[204],pp40[206],pp39[208],pp38[210],pp37[212],pp36[214],pp35[216],pp34[218],pp33[220],pp32[222],pp31[224],pp30[226],pp29[228],pp28[230],pp27[232],pp26[234],pp25[236],pp24[238],pp23[240],pp22[242],pp21[244],pp21[245],pp21[246],pp21[247],pp21[248],pp21[249],pp21[250],pp21[251],pp21[252],pp21[253],pp21[254],pp21[255],pp177[100],pp177[101],pp177[102],pp177[103],pp177[104],pp177[105],pp177[106],pp177[107],pp177[108],pp177[109],pp177[110],pp177[111],pp177[112],pp177[113],pp177[114],pp177[115],pp177[116],pp177[117],pp177[118],pp177[119],pp177[120],pp177[121],pp177[122],pp177[123],pp177[124],pp177[125],pp177[126],pp177[127],pp177[128],pp177[129],pp177[130],pp177[131],pp177[132],pp177[133],pp177[134],pp177[135],pp177[136],pp177[137],pp177[138],pp177[139],pp177[140],pp177[141],pp177[142],pp177[143],pp177[144],pp177[145],pp177[146],pp177[147],pp177[148],pp177[149],pp177[150],pp177[151],pp177[152],pp177[153],pp177[154],pp177[155],pp177[156],pp177[157],pp177[158],pp177[159],pp177[160],pp177[161],pp177[162],pp177[163],pp177[164],pp177[165],pp177[166],pp177[167],pp177[168]};
    CLA_180 KS_39(s39, c39, in39_1, in39_2);
    wire[177:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp120[47],pp119[49],pp118[51],pp117[53],pp116[55],pp115[57],pp114[59],pp113[61],pp112[63],pp111[65],pp110[67],pp109[69],pp108[71],pp107[73],pp106[75],pp105[77],pp104[79],pp103[81],pp102[83],pp101[85],pp100[87],pp88[100],pp88[101],pp88[102],pp88[103],pp88[104],pp88[105],pp88[106],pp88[107],pp88[108],pp88[109],pp88[110],pp88[111],pp87[113],pp86[115],pp85[117],pp84[119],pp83[121],pp82[123],pp81[125],pp80[127],pp79[129],pp78[131],pp77[133],pp76[135],pp75[137],pp74[139],pp73[141],pp72[143],pp71[145],pp70[147],pp69[149],pp68[151],pp67[153],pp66[155],pp65[157],pp64[159],pp63[161],pp62[163],pp61[165],pp60[167],pp59[169],pp58[171],pp57[173],pp56[175],pp55[177],pp54[179],pp53[181],pp52[183],pp51[185],pp50[187],pp49[189],pp48[191],pp47[193],pp46[195],pp45[197],pp44[199],pp43[201],pp42[203],pp41[205],pp40[207],pp39[209],pp38[211],pp37[213],pp36[215],pp35[217],pp34[219],pp33[221],pp32[223],pp31[225],pp30[227],pp29[229],pp28[231],pp27[233],pp26[235],pp25[237],pp24[239],pp23[241],pp22[243],pp22[244],pp22[245],pp22[246],pp22[247],pp22[248],pp22[249],pp22[250],pp22[251],pp22[252],pp22[253],pp22[254],pp22[255],pp178[100],pp178[101],pp178[102],pp178[103],pp178[104],pp178[105],pp178[106],pp178[107],pp178[108],pp178[109],pp178[110],pp178[111],pp178[112],pp178[113],pp178[114],pp178[115],pp178[116],pp178[117],pp178[118],pp178[119],pp178[120],pp178[121],pp178[122],pp178[123],pp178[124],pp178[125],pp178[126],pp178[127],pp178[128],pp178[129],pp178[130],pp178[131],pp178[132],pp178[133],pp178[134],pp178[135],pp178[136],pp178[137],pp178[138],pp178[139],pp178[140],pp178[141],pp178[142],pp178[143],pp178[144],pp178[145],pp178[146],pp178[147],pp178[148],pp178[149],pp178[150],pp178[151],pp178[152],pp178[153],pp178[154],pp178[155],pp178[156],pp178[157],pp178[158],pp178[159],pp178[160],pp178[161],pp178[162],pp178[163],pp178[164],pp178[165],pp178[166]};
    assign in40_2 = {pp121[46],pp120[48],pp119[50],pp118[52],pp117[54],pp116[56],pp115[58],pp114[60],pp113[62],pp112[64],pp111[66],pp110[68],pp109[70],pp108[72],pp107[74],pp106[76],pp105[78],pp104[80],pp103[82],pp102[84],pp101[86],pp100[88],pp89[100],pp89[101],pp89[102],pp89[103],pp89[104],pp89[105],pp89[106],pp89[107],pp89[108],pp89[109],pp89[110],pp88[112],pp87[114],pp86[116],pp85[118],pp84[120],pp83[122],pp82[124],pp81[126],pp80[128],pp79[130],pp78[132],pp77[134],pp76[136],pp75[138],pp74[140],pp73[142],pp72[144],pp71[146],pp70[148],pp69[150],pp68[152],pp67[154],pp66[156],pp65[158],pp64[160],pp63[162],pp62[164],pp61[166],pp60[168],pp59[170],pp58[172],pp57[174],pp56[176],pp55[178],pp54[180],pp53[182],pp52[184],pp51[186],pp50[188],pp49[190],pp48[192],pp47[194],pp46[196],pp45[198],pp44[200],pp43[202],pp42[204],pp41[206],pp40[208],pp39[210],pp38[212],pp37[214],pp36[216],pp35[218],pp34[220],pp33[222],pp32[224],pp31[226],pp30[228],pp29[230],pp28[232],pp27[234],pp26[236],pp25[238],pp24[240],pp23[242],pp23[243],pp23[244],pp23[245],pp23[246],pp23[247],pp23[248],pp23[249],pp23[250],pp23[251],pp23[252],pp23[253],pp23[254],pp23[255],pp179[100],pp179[101],pp179[102],pp179[103],pp179[104],pp179[105],pp179[106],pp179[107],pp179[108],pp179[109],pp179[110],pp179[111],pp179[112],pp179[113],pp179[114],pp179[115],pp179[116],pp179[117],pp179[118],pp179[119],pp179[120],pp179[121],pp179[122],pp179[123],pp179[124],pp179[125],pp179[126],pp179[127],pp179[128],pp179[129],pp179[130],pp179[131],pp179[132],pp179[133],pp179[134],pp179[135],pp179[136],pp179[137],pp179[138],pp179[139],pp179[140],pp179[141],pp179[142],pp179[143],pp179[144],pp179[145],pp179[146],pp179[147],pp179[148],pp179[149],pp179[150],pp179[151],pp179[152],pp179[153],pp179[154],pp179[155],pp179[156],pp179[157],pp179[158],pp179[159],pp179[160],pp179[161],pp179[162],pp179[163],pp179[164],pp179[165]};
    CLA_178 KS_40(s40, c40, in40_1, in40_2);
    wire[175:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp121[47],pp120[49],pp119[51],pp118[53],pp117[55],pp116[57],pp115[59],pp114[61],pp113[63],pp112[65],pp111[67],pp110[69],pp109[71],pp108[73],pp107[75],pp106[77],pp105[79],pp104[81],pp103[83],pp102[85],pp101[87],pp100[89],pp90[100],pp90[101],pp90[102],pp90[103],pp90[104],pp90[105],pp90[106],pp90[107],pp90[108],pp90[109],pp89[111],pp88[113],pp87[115],pp86[117],pp85[119],pp84[121],pp83[123],pp82[125],pp81[127],pp80[129],pp79[131],pp78[133],pp77[135],pp76[137],pp75[139],pp74[141],pp73[143],pp72[145],pp71[147],pp70[149],pp69[151],pp68[153],pp67[155],pp66[157],pp65[159],pp64[161],pp63[163],pp62[165],pp61[167],pp60[169],pp59[171],pp58[173],pp57[175],pp56[177],pp55[179],pp54[181],pp53[183],pp52[185],pp51[187],pp50[189],pp49[191],pp48[193],pp47[195],pp46[197],pp45[199],pp44[201],pp43[203],pp42[205],pp41[207],pp40[209],pp39[211],pp38[213],pp37[215],pp36[217],pp35[219],pp34[221],pp33[223],pp32[225],pp31[227],pp30[229],pp29[231],pp28[233],pp27[235],pp26[237],pp25[239],pp24[241],pp24[242],pp24[243],pp24[244],pp24[245],pp24[246],pp24[247],pp24[248],pp24[249],pp24[250],pp24[251],pp24[252],pp24[253],pp24[254],pp24[255],pp180[100],pp180[101],pp180[102],pp180[103],pp180[104],pp180[105],pp180[106],pp180[107],pp180[108],pp180[109],pp180[110],pp180[111],pp180[112],pp180[113],pp180[114],pp180[115],pp180[116],pp180[117],pp180[118],pp180[119],pp180[120],pp180[121],pp180[122],pp180[123],pp180[124],pp180[125],pp180[126],pp180[127],pp180[128],pp180[129],pp180[130],pp180[131],pp180[132],pp180[133],pp180[134],pp180[135],pp180[136],pp180[137],pp180[138],pp180[139],pp180[140],pp180[141],pp180[142],pp180[143],pp180[144],pp180[145],pp180[146],pp180[147],pp180[148],pp180[149],pp180[150],pp180[151],pp180[152],pp180[153],pp180[154],pp180[155],pp180[156],pp180[157],pp180[158],pp180[159],pp180[160],pp180[161],pp180[162],pp180[163]};
    assign in41_2 = {pp122[46],pp121[48],pp120[50],pp119[52],pp118[54],pp117[56],pp116[58],pp115[60],pp114[62],pp113[64],pp112[66],pp111[68],pp110[70],pp109[72],pp108[74],pp107[76],pp106[78],pp105[80],pp104[82],pp103[84],pp102[86],pp101[88],pp100[90],pp91[100],pp91[101],pp91[102],pp91[103],pp91[104],pp91[105],pp91[106],pp91[107],pp91[108],pp90[110],pp89[112],pp88[114],pp87[116],pp86[118],pp85[120],pp84[122],pp83[124],pp82[126],pp81[128],pp80[130],pp79[132],pp78[134],pp77[136],pp76[138],pp75[140],pp74[142],pp73[144],pp72[146],pp71[148],pp70[150],pp69[152],pp68[154],pp67[156],pp66[158],pp65[160],pp64[162],pp63[164],pp62[166],pp61[168],pp60[170],pp59[172],pp58[174],pp57[176],pp56[178],pp55[180],pp54[182],pp53[184],pp52[186],pp51[188],pp50[190],pp49[192],pp48[194],pp47[196],pp46[198],pp45[200],pp44[202],pp43[204],pp42[206],pp41[208],pp40[210],pp39[212],pp38[214],pp37[216],pp36[218],pp35[220],pp34[222],pp33[224],pp32[226],pp31[228],pp30[230],pp29[232],pp28[234],pp27[236],pp26[238],pp25[240],pp25[241],pp25[242],pp25[243],pp25[244],pp25[245],pp25[246],pp25[247],pp25[248],pp25[249],pp25[250],pp25[251],pp25[252],pp25[253],pp25[254],pp25[255],pp181[100],pp181[101],pp181[102],pp181[103],pp181[104],pp181[105],pp181[106],pp181[107],pp181[108],pp181[109],pp181[110],pp181[111],pp181[112],pp181[113],pp181[114],pp181[115],pp181[116],pp181[117],pp181[118],pp181[119],pp181[120],pp181[121],pp181[122],pp181[123],pp181[124],pp181[125],pp181[126],pp181[127],pp181[128],pp181[129],pp181[130],pp181[131],pp181[132],pp181[133],pp181[134],pp181[135],pp181[136],pp181[137],pp181[138],pp181[139],pp181[140],pp181[141],pp181[142],pp181[143],pp181[144],pp181[145],pp181[146],pp181[147],pp181[148],pp181[149],pp181[150],pp181[151],pp181[152],pp181[153],pp181[154],pp181[155],pp181[156],pp181[157],pp181[158],pp181[159],pp181[160],pp181[161],pp181[162]};
    CLA_176 KS_41(s41, c41, in41_1, in41_2);
    wire[173:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp122[47],pp121[49],pp120[51],pp119[53],pp118[55],pp117[57],pp116[59],pp115[61],pp114[63],pp113[65],pp112[67],pp111[69],pp110[71],pp109[73],pp108[75],pp107[77],pp106[79],pp105[81],pp104[83],pp103[85],pp102[87],pp101[89],pp100[91],pp92[100],pp92[101],pp92[102],pp92[103],pp92[104],pp92[105],pp92[106],pp92[107],pp91[109],pp90[111],pp89[113],pp88[115],pp87[117],pp86[119],pp85[121],pp84[123],pp83[125],pp82[127],pp81[129],pp80[131],pp79[133],pp78[135],pp77[137],pp76[139],pp75[141],pp74[143],pp73[145],pp72[147],pp71[149],pp70[151],pp69[153],pp68[155],pp67[157],pp66[159],pp65[161],pp64[163],pp63[165],pp62[167],pp61[169],pp60[171],pp59[173],pp58[175],pp57[177],pp56[179],pp55[181],pp54[183],pp53[185],pp52[187],pp51[189],pp50[191],pp49[193],pp48[195],pp47[197],pp46[199],pp45[201],pp44[203],pp43[205],pp42[207],pp41[209],pp40[211],pp39[213],pp38[215],pp37[217],pp36[219],pp35[221],pp34[223],pp33[225],pp32[227],pp31[229],pp30[231],pp29[233],pp28[235],pp27[237],pp26[239],pp26[240],pp26[241],pp26[242],pp26[243],pp26[244],pp26[245],pp26[246],pp26[247],pp26[248],pp26[249],pp26[250],pp26[251],pp26[252],pp26[253],pp26[254],pp26[255],pp182[100],pp182[101],pp182[102],pp182[103],pp182[104],pp182[105],pp182[106],pp182[107],pp182[108],pp182[109],pp182[110],pp182[111],pp182[112],pp182[113],pp182[114],pp182[115],pp182[116],pp182[117],pp182[118],pp182[119],pp182[120],pp182[121],pp182[122],pp182[123],pp182[124],pp182[125],pp182[126],pp182[127],pp182[128],pp182[129],pp182[130],pp182[131],pp182[132],pp182[133],pp182[134],pp182[135],pp182[136],pp182[137],pp182[138],pp182[139],pp182[140],pp182[141],pp182[142],pp182[143],pp182[144],pp182[145],pp182[146],pp182[147],pp182[148],pp182[149],pp182[150],pp182[151],pp182[152],pp182[153],pp182[154],pp182[155],pp182[156],pp182[157],pp182[158],pp182[159],pp182[160]};
    assign in42_2 = {pp123[46],pp122[48],pp121[50],pp120[52],pp119[54],pp118[56],pp117[58],pp116[60],pp115[62],pp114[64],pp113[66],pp112[68],pp111[70],pp110[72],pp109[74],pp108[76],pp107[78],pp106[80],pp105[82],pp104[84],pp103[86],pp102[88],pp101[90],pp100[92],pp93[100],pp93[101],pp93[102],pp93[103],pp93[104],pp93[105],pp93[106],pp92[108],pp91[110],pp90[112],pp89[114],pp88[116],pp87[118],pp86[120],pp85[122],pp84[124],pp83[126],pp82[128],pp81[130],pp80[132],pp79[134],pp78[136],pp77[138],pp76[140],pp75[142],pp74[144],pp73[146],pp72[148],pp71[150],pp70[152],pp69[154],pp68[156],pp67[158],pp66[160],pp65[162],pp64[164],pp63[166],pp62[168],pp61[170],pp60[172],pp59[174],pp58[176],pp57[178],pp56[180],pp55[182],pp54[184],pp53[186],pp52[188],pp51[190],pp50[192],pp49[194],pp48[196],pp47[198],pp46[200],pp45[202],pp44[204],pp43[206],pp42[208],pp41[210],pp40[212],pp39[214],pp38[216],pp37[218],pp36[220],pp35[222],pp34[224],pp33[226],pp32[228],pp31[230],pp30[232],pp29[234],pp28[236],pp27[238],pp27[239],pp27[240],pp27[241],pp27[242],pp27[243],pp27[244],pp27[245],pp27[246],pp27[247],pp27[248],pp27[249],pp27[250],pp27[251],pp27[252],pp27[253],pp27[254],pp27[255],pp183[100],pp183[101],pp183[102],pp183[103],pp183[104],pp183[105],pp183[106],pp183[107],pp183[108],pp183[109],pp183[110],pp183[111],pp183[112],pp183[113],pp183[114],pp183[115],pp183[116],pp183[117],pp183[118],pp183[119],pp183[120],pp183[121],pp183[122],pp183[123],pp183[124],pp183[125],pp183[126],pp183[127],pp183[128],pp183[129],pp183[130],pp183[131],pp183[132],pp183[133],pp183[134],pp183[135],pp183[136],pp183[137],pp183[138],pp183[139],pp183[140],pp183[141],pp183[142],pp183[143],pp183[144],pp183[145],pp183[146],pp183[147],pp183[148],pp183[149],pp183[150],pp183[151],pp183[152],pp183[153],pp183[154],pp183[155],pp183[156],pp183[157],pp183[158],pp183[159]};
    CLA_174 KS_42(s42, c42, in42_1, in42_2);
    wire[171:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp123[47],pp122[49],pp121[51],pp120[53],pp119[55],pp118[57],pp117[59],pp116[61],pp115[63],pp114[65],pp113[67],pp112[69],pp111[71],pp110[73],pp109[75],pp108[77],pp107[79],pp106[81],pp105[83],pp104[85],pp103[87],pp102[89],pp101[91],pp100[93],pp94[100],pp94[101],pp94[102],pp94[103],pp94[104],pp94[105],pp93[107],pp92[109],pp91[111],pp90[113],pp89[115],pp88[117],pp87[119],pp86[121],pp85[123],pp84[125],pp83[127],pp82[129],pp81[131],pp80[133],pp79[135],pp78[137],pp77[139],pp76[141],pp75[143],pp74[145],pp73[147],pp72[149],pp71[151],pp70[153],pp69[155],pp68[157],pp67[159],pp66[161],pp65[163],pp64[165],pp63[167],pp62[169],pp61[171],pp60[173],pp59[175],pp58[177],pp57[179],pp56[181],pp55[183],pp54[185],pp53[187],pp52[189],pp51[191],pp50[193],pp49[195],pp48[197],pp47[199],pp46[201],pp45[203],pp44[205],pp43[207],pp42[209],pp41[211],pp40[213],pp39[215],pp38[217],pp37[219],pp36[221],pp35[223],pp34[225],pp33[227],pp32[229],pp31[231],pp30[233],pp29[235],pp28[237],pp28[238],pp28[239],pp28[240],pp28[241],pp28[242],pp28[243],pp28[244],pp28[245],pp28[246],pp28[247],pp28[248],pp28[249],pp28[250],pp28[251],pp28[252],pp28[253],pp28[254],pp28[255],pp184[100],pp184[101],pp184[102],pp184[103],pp184[104],pp184[105],pp184[106],pp184[107],pp184[108],pp184[109],pp184[110],pp184[111],pp184[112],pp184[113],pp184[114],pp184[115],pp184[116],pp184[117],pp184[118],pp184[119],pp184[120],pp184[121],pp184[122],pp184[123],pp184[124],pp184[125],pp184[126],pp184[127],pp184[128],pp184[129],pp184[130],pp184[131],pp184[132],pp184[133],pp184[134],pp184[135],pp184[136],pp184[137],pp184[138],pp184[139],pp184[140],pp184[141],pp184[142],pp184[143],pp184[144],pp184[145],pp184[146],pp184[147],pp184[148],pp184[149],pp184[150],pp184[151],pp184[152],pp184[153],pp184[154],pp184[155],pp184[156],pp184[157]};
    assign in43_2 = {pp124[46],pp123[48],pp122[50],pp121[52],pp120[54],pp119[56],pp118[58],pp117[60],pp116[62],pp115[64],pp114[66],pp113[68],pp112[70],pp111[72],pp110[74],pp109[76],pp108[78],pp107[80],pp106[82],pp105[84],pp104[86],pp103[88],pp102[90],pp101[92],pp100[94],pp95[100],pp95[101],pp95[102],pp95[103],pp95[104],pp94[106],pp93[108],pp92[110],pp91[112],pp90[114],pp89[116],pp88[118],pp87[120],pp86[122],pp85[124],pp84[126],pp83[128],pp82[130],pp81[132],pp80[134],pp79[136],pp78[138],pp77[140],pp76[142],pp75[144],pp74[146],pp73[148],pp72[150],pp71[152],pp70[154],pp69[156],pp68[158],pp67[160],pp66[162],pp65[164],pp64[166],pp63[168],pp62[170],pp61[172],pp60[174],pp59[176],pp58[178],pp57[180],pp56[182],pp55[184],pp54[186],pp53[188],pp52[190],pp51[192],pp50[194],pp49[196],pp48[198],pp47[200],pp46[202],pp45[204],pp44[206],pp43[208],pp42[210],pp41[212],pp40[214],pp39[216],pp38[218],pp37[220],pp36[222],pp35[224],pp34[226],pp33[228],pp32[230],pp31[232],pp30[234],pp29[236],pp29[237],pp29[238],pp29[239],pp29[240],pp29[241],pp29[242],pp29[243],pp29[244],pp29[245],pp29[246],pp29[247],pp29[248],pp29[249],pp29[250],pp29[251],pp29[252],pp29[253],pp29[254],pp29[255],pp185[100],pp185[101],pp185[102],pp185[103],pp185[104],pp185[105],pp185[106],pp185[107],pp185[108],pp185[109],pp185[110],pp185[111],pp185[112],pp185[113],pp185[114],pp185[115],pp185[116],pp185[117],pp185[118],pp185[119],pp185[120],pp185[121],pp185[122],pp185[123],pp185[124],pp185[125],pp185[126],pp185[127],pp185[128],pp185[129],pp185[130],pp185[131],pp185[132],pp185[133],pp185[134],pp185[135],pp185[136],pp185[137],pp185[138],pp185[139],pp185[140],pp185[141],pp185[142],pp185[143],pp185[144],pp185[145],pp185[146],pp185[147],pp185[148],pp185[149],pp185[150],pp185[151],pp185[152],pp185[153],pp185[154],pp185[155],pp185[156]};
    CLA_172 KS_43(s43, c43, in43_1, in43_2);
    wire[169:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp124[47],pp123[49],pp122[51],pp121[53],pp120[55],pp119[57],pp118[59],pp117[61],pp116[63],pp115[65],pp114[67],pp113[69],pp112[71],pp111[73],pp110[75],pp109[77],pp108[79],pp107[81],pp106[83],pp105[85],pp104[87],pp103[89],pp102[91],pp101[93],pp100[95],pp96[100],pp96[101],pp96[102],pp96[103],pp95[105],pp94[107],pp93[109],pp92[111],pp91[113],pp90[115],pp89[117],pp88[119],pp87[121],pp86[123],pp85[125],pp84[127],pp83[129],pp82[131],pp81[133],pp80[135],pp79[137],pp78[139],pp77[141],pp76[143],pp75[145],pp74[147],pp73[149],pp72[151],pp71[153],pp70[155],pp69[157],pp68[159],pp67[161],pp66[163],pp65[165],pp64[167],pp63[169],pp62[171],pp61[173],pp60[175],pp59[177],pp58[179],pp57[181],pp56[183],pp55[185],pp54[187],pp53[189],pp52[191],pp51[193],pp50[195],pp49[197],pp48[199],pp47[201],pp46[203],pp45[205],pp44[207],pp43[209],pp42[211],pp41[213],pp40[215],pp39[217],pp38[219],pp37[221],pp36[223],pp35[225],pp34[227],pp33[229],pp32[231],pp31[233],pp30[235],pp30[236],pp30[237],pp30[238],pp30[239],pp30[240],pp30[241],pp30[242],pp30[243],pp30[244],pp30[245],pp30[246],pp30[247],pp30[248],pp30[249],pp30[250],pp30[251],pp30[252],pp30[253],pp30[254],pp30[255],pp186[100],pp186[101],pp186[102],pp186[103],pp186[104],pp186[105],pp186[106],pp186[107],pp186[108],pp186[109],pp186[110],pp186[111],pp186[112],pp186[113],pp186[114],pp186[115],pp186[116],pp186[117],pp186[118],pp186[119],pp186[120],pp186[121],pp186[122],pp186[123],pp186[124],pp186[125],pp186[126],pp186[127],pp186[128],pp186[129],pp186[130],pp186[131],pp186[132],pp186[133],pp186[134],pp186[135],pp186[136],pp186[137],pp186[138],pp186[139],pp186[140],pp186[141],pp186[142],pp186[143],pp186[144],pp186[145],pp186[146],pp186[147],pp186[148],pp186[149],pp186[150],pp186[151],pp186[152],pp186[153],pp186[154]};
    assign in44_2 = {pp125[46],pp124[48],pp123[50],pp122[52],pp121[54],pp120[56],pp119[58],pp118[60],pp117[62],pp116[64],pp115[66],pp114[68],pp113[70],pp112[72],pp111[74],pp110[76],pp109[78],pp108[80],pp107[82],pp106[84],pp105[86],pp104[88],pp103[90],pp102[92],pp101[94],pp100[96],pp97[100],pp97[101],pp97[102],pp96[104],pp95[106],pp94[108],pp93[110],pp92[112],pp91[114],pp90[116],pp89[118],pp88[120],pp87[122],pp86[124],pp85[126],pp84[128],pp83[130],pp82[132],pp81[134],pp80[136],pp79[138],pp78[140],pp77[142],pp76[144],pp75[146],pp74[148],pp73[150],pp72[152],pp71[154],pp70[156],pp69[158],pp68[160],pp67[162],pp66[164],pp65[166],pp64[168],pp63[170],pp62[172],pp61[174],pp60[176],pp59[178],pp58[180],pp57[182],pp56[184],pp55[186],pp54[188],pp53[190],pp52[192],pp51[194],pp50[196],pp49[198],pp48[200],pp47[202],pp46[204],pp45[206],pp44[208],pp43[210],pp42[212],pp41[214],pp40[216],pp39[218],pp38[220],pp37[222],pp36[224],pp35[226],pp34[228],pp33[230],pp32[232],pp31[234],pp31[235],pp31[236],pp31[237],pp31[238],pp31[239],pp31[240],pp31[241],pp31[242],pp31[243],pp31[244],pp31[245],pp31[246],pp31[247],pp31[248],pp31[249],pp31[250],pp31[251],pp31[252],pp31[253],pp31[254],pp31[255],pp187[100],pp187[101],pp187[102],pp187[103],pp187[104],pp187[105],pp187[106],pp187[107],pp187[108],pp187[109],pp187[110],pp187[111],pp187[112],pp187[113],pp187[114],pp187[115],pp187[116],pp187[117],pp187[118],pp187[119],pp187[120],pp187[121],pp187[122],pp187[123],pp187[124],pp187[125],pp187[126],pp187[127],pp187[128],pp187[129],pp187[130],pp187[131],pp187[132],pp187[133],pp187[134],pp187[135],pp187[136],pp187[137],pp187[138],pp187[139],pp187[140],pp187[141],pp187[142],pp187[143],pp187[144],pp187[145],pp187[146],pp187[147],pp187[148],pp187[149],pp187[150],pp187[151],pp187[152],pp187[153]};
    CLA_170 KS_44(s44, c44, in44_1, in44_2);
    wire[167:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp125[47],pp124[49],pp123[51],pp122[53],pp121[55],pp120[57],pp119[59],pp118[61],pp117[63],pp116[65],pp115[67],pp114[69],pp113[71],pp112[73],pp111[75],pp110[77],pp109[79],pp108[81],pp107[83],pp106[85],pp105[87],pp104[89],pp103[91],pp102[93],pp101[95],pp100[97],pp98[100],pp98[101],pp97[103],pp96[105],pp95[107],pp94[109],pp93[111],pp92[113],pp91[115],pp90[117],pp89[119],pp88[121],pp87[123],pp86[125],pp85[127],pp84[129],pp83[131],pp82[133],pp81[135],pp80[137],pp79[139],pp78[141],pp77[143],pp76[145],pp75[147],pp74[149],pp73[151],pp72[153],pp71[155],pp70[157],pp69[159],pp68[161],pp67[163],pp66[165],pp65[167],pp64[169],pp63[171],pp62[173],pp61[175],pp60[177],pp59[179],pp58[181],pp57[183],pp56[185],pp55[187],pp54[189],pp53[191],pp52[193],pp51[195],pp50[197],pp49[199],pp48[201],pp47[203],pp46[205],pp45[207],pp44[209],pp43[211],pp42[213],pp41[215],pp40[217],pp39[219],pp38[221],pp37[223],pp36[225],pp35[227],pp34[229],pp33[231],pp32[233],pp32[234],pp32[235],pp32[236],pp32[237],pp32[238],pp32[239],pp32[240],pp32[241],pp32[242],pp32[243],pp32[244],pp32[245],pp32[246],pp32[247],pp32[248],pp32[249],pp32[250],pp32[251],pp32[252],pp32[253],pp32[254],pp32[255],pp188[100],pp188[101],pp188[102],pp188[103],pp188[104],pp188[105],pp188[106],pp188[107],pp188[108],pp188[109],pp188[110],pp188[111],pp188[112],pp188[113],pp188[114],pp188[115],pp188[116],pp188[117],pp188[118],pp188[119],pp188[120],pp188[121],pp188[122],pp188[123],pp188[124],pp188[125],pp188[126],pp188[127],pp188[128],pp188[129],pp188[130],pp188[131],pp188[132],pp188[133],pp188[134],pp188[135],pp188[136],pp188[137],pp188[138],pp188[139],pp188[140],pp188[141],pp188[142],pp188[143],pp188[144],pp188[145],pp188[146],pp188[147],pp188[148],pp188[149],pp188[150],pp188[151]};
    assign in45_2 = {pp126[46],pp125[48],pp124[50],pp123[52],pp122[54],pp121[56],pp120[58],pp119[60],pp118[62],pp117[64],pp116[66],pp115[68],pp114[70],pp113[72],pp112[74],pp111[76],pp110[78],pp109[80],pp108[82],pp107[84],pp106[86],pp105[88],pp104[90],pp103[92],pp102[94],pp101[96],pp100[98],pp99[100],pp98[102],pp97[104],pp96[106],pp95[108],pp94[110],pp93[112],pp92[114],pp91[116],pp90[118],pp89[120],pp88[122],pp87[124],pp86[126],pp85[128],pp84[130],pp83[132],pp82[134],pp81[136],pp80[138],pp79[140],pp78[142],pp77[144],pp76[146],pp75[148],pp74[150],pp73[152],pp72[154],pp71[156],pp70[158],pp69[160],pp68[162],pp67[164],pp66[166],pp65[168],pp64[170],pp63[172],pp62[174],pp61[176],pp60[178],pp59[180],pp58[182],pp57[184],pp56[186],pp55[188],pp54[190],pp53[192],pp52[194],pp51[196],pp50[198],pp49[200],pp48[202],pp47[204],pp46[206],pp45[208],pp44[210],pp43[212],pp42[214],pp41[216],pp40[218],pp39[220],pp38[222],pp37[224],pp36[226],pp35[228],pp34[230],pp33[232],pp33[233],pp33[234],pp33[235],pp33[236],pp33[237],pp33[238],pp33[239],pp33[240],pp33[241],pp33[242],pp33[243],pp33[244],pp33[245],pp33[246],pp33[247],pp33[248],pp33[249],pp33[250],pp33[251],pp33[252],pp33[253],pp33[254],pp33[255],pp189[100],pp189[101],pp189[102],pp189[103],pp189[104],pp189[105],pp189[106],pp189[107],pp189[108],pp189[109],pp189[110],pp189[111],pp189[112],pp189[113],pp189[114],pp189[115],pp189[116],pp189[117],pp189[118],pp189[119],pp189[120],pp189[121],pp189[122],pp189[123],pp189[124],pp189[125],pp189[126],pp189[127],pp189[128],pp189[129],pp189[130],pp189[131],pp189[132],pp189[133],pp189[134],pp189[135],pp189[136],pp189[137],pp189[138],pp189[139],pp189[140],pp189[141],pp189[142],pp189[143],pp189[144],pp189[145],pp189[146],pp189[147],pp189[148],pp189[149],pp189[150]};
    CLA_168 KS_45(s45, c45, in45_1, in45_2);
    wire[165:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp126[47],pp125[49],pp124[51],pp123[53],pp122[55],pp121[57],pp120[59],pp119[61],pp118[63],pp117[65],pp116[67],pp115[69],pp114[71],pp113[73],pp112[75],pp111[77],pp110[79],pp109[81],pp108[83],pp107[85],pp106[87],pp105[89],pp104[91],pp103[93],pp102[95],pp101[97],pp100[99],pp99[101],pp98[103],pp97[105],pp96[107],pp95[109],pp94[111],pp93[113],pp92[115],pp91[117],pp90[119],pp89[121],pp88[123],pp87[125],pp86[127],pp85[129],pp84[131],pp83[133],pp82[135],pp81[137],pp80[139],pp79[141],pp78[143],pp77[145],pp76[147],pp75[149],pp74[151],pp73[153],pp72[155],pp71[157],pp70[159],pp69[161],pp68[163],pp67[165],pp66[167],pp65[169],pp64[171],pp63[173],pp62[175],pp61[177],pp60[179],pp59[181],pp58[183],pp57[185],pp56[187],pp55[189],pp54[191],pp53[193],pp52[195],pp51[197],pp50[199],pp49[201],pp48[203],pp47[205],pp46[207],pp45[209],pp44[211],pp43[213],pp42[215],pp41[217],pp40[219],pp39[221],pp38[223],pp37[225],pp36[227],pp35[229],pp34[231],pp34[232],pp34[233],pp34[234],pp34[235],pp34[236],pp34[237],pp34[238],pp34[239],pp34[240],pp34[241],pp34[242],pp34[243],pp34[244],pp34[245],pp34[246],pp34[247],pp34[248],pp34[249],pp34[250],pp34[251],pp34[252],pp34[253],pp34[254],pp34[255],pp190[100],pp190[101],pp190[102],pp190[103],pp190[104],pp190[105],pp190[106],pp190[107],pp190[108],pp190[109],pp190[110],pp190[111],pp190[112],pp190[113],pp190[114],pp190[115],pp190[116],pp190[117],pp190[118],pp190[119],pp190[120],pp190[121],pp190[122],pp190[123],pp190[124],pp190[125],pp190[126],pp190[127],pp190[128],pp190[129],pp190[130],pp190[131],pp190[132],pp190[133],pp190[134],pp190[135],pp190[136],pp190[137],pp190[138],pp190[139],pp190[140],pp190[141],pp190[142],pp190[143],pp190[144],pp190[145],pp190[146],pp190[147],pp190[148]};
    assign in46_2 = {pp127[46],pp126[48],pp125[50],pp124[52],pp123[54],pp122[56],pp121[58],pp120[60],pp119[62],pp118[64],pp117[66],pp116[68],pp115[70],pp114[72],pp113[74],pp112[76],pp111[78],pp110[80],pp109[82],pp108[84],pp107[86],pp106[88],pp105[90],pp104[92],pp103[94],pp102[96],pp101[98],pp101[99],pp99[102],pp98[104],pp97[106],pp96[108],pp95[110],pp94[112],pp93[114],pp92[116],pp91[118],pp90[120],pp89[122],pp88[124],pp87[126],pp86[128],pp85[130],pp84[132],pp83[134],pp82[136],pp81[138],pp80[140],pp79[142],pp78[144],pp77[146],pp76[148],pp75[150],pp74[152],pp73[154],pp72[156],pp71[158],pp70[160],pp69[162],pp68[164],pp67[166],pp66[168],pp65[170],pp64[172],pp63[174],pp62[176],pp61[178],pp60[180],pp59[182],pp58[184],pp57[186],pp56[188],pp55[190],pp54[192],pp53[194],pp52[196],pp51[198],pp50[200],pp49[202],pp48[204],pp47[206],pp46[208],pp45[210],pp44[212],pp43[214],pp42[216],pp41[218],pp40[220],pp39[222],pp38[224],pp37[226],pp36[228],pp35[230],pp35[231],pp35[232],pp35[233],pp35[234],pp35[235],pp35[236],pp35[237],pp35[238],pp35[239],pp35[240],pp35[241],pp35[242],pp35[243],pp35[244],pp35[245],pp35[246],pp35[247],pp35[248],pp35[249],pp35[250],pp35[251],pp35[252],pp35[253],pp35[254],pp35[255],pp191[100],pp191[101],pp191[102],pp191[103],pp191[104],pp191[105],pp191[106],pp191[107],pp191[108],pp191[109],pp191[110],pp191[111],pp191[112],pp191[113],pp191[114],pp191[115],pp191[116],pp191[117],pp191[118],pp191[119],pp191[120],pp191[121],pp191[122],pp191[123],pp191[124],pp191[125],pp191[126],pp191[127],pp191[128],pp191[129],pp191[130],pp191[131],pp191[132],pp191[133],pp191[134],pp191[135],pp191[136],pp191[137],pp191[138],pp191[139],pp191[140],pp191[141],pp191[142],pp191[143],pp191[144],pp191[145],pp191[146],pp191[147]};
    CLA_166 KS_46(s46, c46, in46_1, in46_2);
    wire[163:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp127[47],pp126[49],pp125[51],pp124[53],pp123[55],pp122[57],pp121[59],pp120[61],pp119[63],pp118[65],pp117[67],pp116[69],pp115[71],pp114[73],pp113[75],pp112[77],pp111[79],pp110[81],pp109[83],pp108[85],pp107[87],pp106[89],pp105[91],pp104[93],pp103[95],pp102[97],pp102[98],pp102[99],pp99[103],pp98[105],pp97[107],pp96[109],pp95[111],pp94[113],pp93[115],pp92[117],pp91[119],pp90[121],pp89[123],pp88[125],pp87[127],pp86[129],pp85[131],pp84[133],pp83[135],pp82[137],pp81[139],pp80[141],pp79[143],pp78[145],pp77[147],pp76[149],pp75[151],pp74[153],pp73[155],pp72[157],pp71[159],pp70[161],pp69[163],pp68[165],pp67[167],pp66[169],pp65[171],pp64[173],pp63[175],pp62[177],pp61[179],pp60[181],pp59[183],pp58[185],pp57[187],pp56[189],pp55[191],pp54[193],pp53[195],pp52[197],pp51[199],pp50[201],pp49[203],pp48[205],pp47[207],pp46[209],pp45[211],pp44[213],pp43[215],pp42[217],pp41[219],pp40[221],pp39[223],pp38[225],pp37[227],pp36[229],pp36[230],pp36[231],pp36[232],pp36[233],pp36[234],pp36[235],pp36[236],pp36[237],pp36[238],pp36[239],pp36[240],pp36[241],pp36[242],pp36[243],pp36[244],pp36[245],pp36[246],pp36[247],pp36[248],pp36[249],pp36[250],pp36[251],pp36[252],pp36[253],pp36[254],pp36[255],pp192[100],pp192[101],pp192[102],pp192[103],pp192[104],pp192[105],pp192[106],pp192[107],pp192[108],pp192[109],pp192[110],pp192[111],pp192[112],pp192[113],pp192[114],pp192[115],pp192[116],pp192[117],pp192[118],pp192[119],pp192[120],pp192[121],pp192[122],pp192[123],pp192[124],pp192[125],pp192[126],pp192[127],pp192[128],pp192[129],pp192[130],pp192[131],pp192[132],pp192[133],pp192[134],pp192[135],pp192[136],pp192[137],pp192[138],pp192[139],pp192[140],pp192[141],pp192[142],pp192[143],pp192[144],pp192[145]};
    assign in47_2 = {pp128[46],pp127[48],pp126[50],pp125[52],pp124[54],pp123[56],pp122[58],pp121[60],pp120[62],pp119[64],pp118[66],pp117[68],pp116[70],pp115[72],pp114[74],pp113[76],pp112[78],pp111[80],pp110[82],pp109[84],pp108[86],pp107[88],pp106[90],pp105[92],pp104[94],pp103[96],pp103[97],pp103[98],pp103[99],pp99[104],pp98[106],pp97[108],pp96[110],pp95[112],pp94[114],pp93[116],pp92[118],pp91[120],pp90[122],pp89[124],pp88[126],pp87[128],pp86[130],pp85[132],pp84[134],pp83[136],pp82[138],pp81[140],pp80[142],pp79[144],pp78[146],pp77[148],pp76[150],pp75[152],pp74[154],pp73[156],pp72[158],pp71[160],pp70[162],pp69[164],pp68[166],pp67[168],pp66[170],pp65[172],pp64[174],pp63[176],pp62[178],pp61[180],pp60[182],pp59[184],pp58[186],pp57[188],pp56[190],pp55[192],pp54[194],pp53[196],pp52[198],pp51[200],pp50[202],pp49[204],pp48[206],pp47[208],pp46[210],pp45[212],pp44[214],pp43[216],pp42[218],pp41[220],pp40[222],pp39[224],pp38[226],pp37[228],pp37[229],pp37[230],pp37[231],pp37[232],pp37[233],pp37[234],pp37[235],pp37[236],pp37[237],pp37[238],pp37[239],pp37[240],pp37[241],pp37[242],pp37[243],pp37[244],pp37[245],pp37[246],pp37[247],pp37[248],pp37[249],pp37[250],pp37[251],pp37[252],pp37[253],pp37[254],pp37[255],pp193[100],pp193[101],pp193[102],pp193[103],pp193[104],pp193[105],pp193[106],pp193[107],pp193[108],pp193[109],pp193[110],pp193[111],pp193[112],pp193[113],pp193[114],pp193[115],pp193[116],pp193[117],pp193[118],pp193[119],pp193[120],pp193[121],pp193[122],pp193[123],pp193[124],pp193[125],pp193[126],pp193[127],pp193[128],pp193[129],pp193[130],pp193[131],pp193[132],pp193[133],pp193[134],pp193[135],pp193[136],pp193[137],pp193[138],pp193[139],pp193[140],pp193[141],pp193[142],pp193[143],pp193[144]};
    CLA_164 KS_47(s47, c47, in47_1, in47_2);
    wire[161:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp128[47],pp127[49],pp126[51],pp125[53],pp124[55],pp123[57],pp122[59],pp121[61],pp120[63],pp119[65],pp118[67],pp117[69],pp116[71],pp115[73],pp114[75],pp113[77],pp112[79],pp111[81],pp110[83],pp109[85],pp108[87],pp107[89],pp106[91],pp105[93],pp104[95],pp104[96],pp104[97],pp104[98],pp104[99],pp99[105],pp98[107],pp97[109],pp96[111],pp95[113],pp94[115],pp93[117],pp92[119],pp91[121],pp90[123],pp89[125],pp88[127],pp87[129],pp86[131],pp85[133],pp84[135],pp83[137],pp82[139],pp81[141],pp80[143],pp79[145],pp78[147],pp77[149],pp76[151],pp75[153],pp74[155],pp73[157],pp72[159],pp71[161],pp70[163],pp69[165],pp68[167],pp67[169],pp66[171],pp65[173],pp64[175],pp63[177],pp62[179],pp61[181],pp60[183],pp59[185],pp58[187],pp57[189],pp56[191],pp55[193],pp54[195],pp53[197],pp52[199],pp51[201],pp50[203],pp49[205],pp48[207],pp47[209],pp46[211],pp45[213],pp44[215],pp43[217],pp42[219],pp41[221],pp40[223],pp39[225],pp38[227],pp38[228],pp38[229],pp38[230],pp38[231],pp38[232],pp38[233],pp38[234],pp38[235],pp38[236],pp38[237],pp38[238],pp38[239],pp38[240],pp38[241],pp38[242],pp38[243],pp38[244],pp38[245],pp38[246],pp38[247],pp38[248],pp38[249],pp38[250],pp38[251],pp38[252],pp38[253],pp38[254],pp38[255],pp194[100],pp194[101],pp194[102],pp194[103],pp194[104],pp194[105],pp194[106],pp194[107],pp194[108],pp194[109],pp194[110],pp194[111],pp194[112],pp194[113],pp194[114],pp194[115],pp194[116],pp194[117],pp194[118],pp194[119],pp194[120],pp194[121],pp194[122],pp194[123],pp194[124],pp194[125],pp194[126],pp194[127],pp194[128],pp194[129],pp194[130],pp194[131],pp194[132],pp194[133],pp194[134],pp194[135],pp194[136],pp194[137],pp194[138],pp194[139],pp194[140],pp194[141],pp194[142]};
    assign in48_2 = {pp129[46],pp128[48],pp127[50],pp126[52],pp125[54],pp124[56],pp123[58],pp122[60],pp121[62],pp120[64],pp119[66],pp118[68],pp117[70],pp116[72],pp115[74],pp114[76],pp113[78],pp112[80],pp111[82],pp110[84],pp109[86],pp108[88],pp107[90],pp106[92],pp105[94],pp105[95],pp105[96],pp105[97],pp105[98],pp105[99],pp99[106],pp98[108],pp97[110],pp96[112],pp95[114],pp94[116],pp93[118],pp92[120],pp91[122],pp90[124],pp89[126],pp88[128],pp87[130],pp86[132],pp85[134],pp84[136],pp83[138],pp82[140],pp81[142],pp80[144],pp79[146],pp78[148],pp77[150],pp76[152],pp75[154],pp74[156],pp73[158],pp72[160],pp71[162],pp70[164],pp69[166],pp68[168],pp67[170],pp66[172],pp65[174],pp64[176],pp63[178],pp62[180],pp61[182],pp60[184],pp59[186],pp58[188],pp57[190],pp56[192],pp55[194],pp54[196],pp53[198],pp52[200],pp51[202],pp50[204],pp49[206],pp48[208],pp47[210],pp46[212],pp45[214],pp44[216],pp43[218],pp42[220],pp41[222],pp40[224],pp39[226],pp39[227],pp39[228],pp39[229],pp39[230],pp39[231],pp39[232],pp39[233],pp39[234],pp39[235],pp39[236],pp39[237],pp39[238],pp39[239],pp39[240],pp39[241],pp39[242],pp39[243],pp39[244],pp39[245],pp39[246],pp39[247],pp39[248],pp39[249],pp39[250],pp39[251],pp39[252],pp39[253],pp39[254],pp39[255],pp195[100],pp195[101],pp195[102],pp195[103],pp195[104],pp195[105],pp195[106],pp195[107],pp195[108],pp195[109],pp195[110],pp195[111],pp195[112],pp195[113],pp195[114],pp195[115],pp195[116],pp195[117],pp195[118],pp195[119],pp195[120],pp195[121],pp195[122],pp195[123],pp195[124],pp195[125],pp195[126],pp195[127],pp195[128],pp195[129],pp195[130],pp195[131],pp195[132],pp195[133],pp195[134],pp195[135],pp195[136],pp195[137],pp195[138],pp195[139],pp195[140],pp195[141]};
    CLA_162 KS_48(s48, c48, in48_1, in48_2);
    wire[159:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp129[47],pp128[49],pp127[51],pp126[53],pp125[55],pp124[57],pp123[59],pp122[61],pp121[63],pp120[65],pp119[67],pp118[69],pp117[71],pp116[73],pp115[75],pp114[77],pp113[79],pp112[81],pp111[83],pp110[85],pp109[87],pp108[89],pp107[91],pp106[93],pp106[94],pp106[95],pp106[96],pp106[97],pp106[98],pp106[99],pp99[107],pp98[109],pp97[111],pp96[113],pp95[115],pp94[117],pp93[119],pp92[121],pp91[123],pp90[125],pp89[127],pp88[129],pp87[131],pp86[133],pp85[135],pp84[137],pp83[139],pp82[141],pp81[143],pp80[145],pp79[147],pp78[149],pp77[151],pp76[153],pp75[155],pp74[157],pp73[159],pp72[161],pp71[163],pp70[165],pp69[167],pp68[169],pp67[171],pp66[173],pp65[175],pp64[177],pp63[179],pp62[181],pp61[183],pp60[185],pp59[187],pp58[189],pp57[191],pp56[193],pp55[195],pp54[197],pp53[199],pp52[201],pp51[203],pp50[205],pp49[207],pp48[209],pp47[211],pp46[213],pp45[215],pp44[217],pp43[219],pp42[221],pp41[223],pp40[225],pp40[226],pp40[227],pp40[228],pp40[229],pp40[230],pp40[231],pp40[232],pp40[233],pp40[234],pp40[235],pp40[236],pp40[237],pp40[238],pp40[239],pp40[240],pp40[241],pp40[242],pp40[243],pp40[244],pp40[245],pp40[246],pp40[247],pp40[248],pp40[249],pp40[250],pp40[251],pp40[252],pp40[253],pp40[254],pp40[255],pp196[100],pp196[101],pp196[102],pp196[103],pp196[104],pp196[105],pp196[106],pp196[107],pp196[108],pp196[109],pp196[110],pp196[111],pp196[112],pp196[113],pp196[114],pp196[115],pp196[116],pp196[117],pp196[118],pp196[119],pp196[120],pp196[121],pp196[122],pp196[123],pp196[124],pp196[125],pp196[126],pp196[127],pp196[128],pp196[129],pp196[130],pp196[131],pp196[132],pp196[133],pp196[134],pp196[135],pp196[136],pp196[137],pp196[138],pp196[139]};
    assign in49_2 = {pp130[46],pp129[48],pp128[50],pp127[52],pp126[54],pp125[56],pp124[58],pp123[60],pp122[62],pp121[64],pp120[66],pp119[68],pp118[70],pp117[72],pp116[74],pp115[76],pp114[78],pp113[80],pp112[82],pp111[84],pp110[86],pp109[88],pp108[90],pp107[92],pp107[93],pp107[94],pp107[95],pp107[96],pp107[97],pp107[98],pp107[99],pp99[108],pp98[110],pp97[112],pp96[114],pp95[116],pp94[118],pp93[120],pp92[122],pp91[124],pp90[126],pp89[128],pp88[130],pp87[132],pp86[134],pp85[136],pp84[138],pp83[140],pp82[142],pp81[144],pp80[146],pp79[148],pp78[150],pp77[152],pp76[154],pp75[156],pp74[158],pp73[160],pp72[162],pp71[164],pp70[166],pp69[168],pp68[170],pp67[172],pp66[174],pp65[176],pp64[178],pp63[180],pp62[182],pp61[184],pp60[186],pp59[188],pp58[190],pp57[192],pp56[194],pp55[196],pp54[198],pp53[200],pp52[202],pp51[204],pp50[206],pp49[208],pp48[210],pp47[212],pp46[214],pp45[216],pp44[218],pp43[220],pp42[222],pp41[224],pp41[225],pp41[226],pp41[227],pp41[228],pp41[229],pp41[230],pp41[231],pp41[232],pp41[233],pp41[234],pp41[235],pp41[236],pp41[237],pp41[238],pp41[239],pp41[240],pp41[241],pp41[242],pp41[243],pp41[244],pp41[245],pp41[246],pp41[247],pp41[248],pp41[249],pp41[250],pp41[251],pp41[252],pp41[253],pp41[254],pp41[255],pp197[100],pp197[101],pp197[102],pp197[103],pp197[104],pp197[105],pp197[106],pp197[107],pp197[108],pp197[109],pp197[110],pp197[111],pp197[112],pp197[113],pp197[114],pp197[115],pp197[116],pp197[117],pp197[118],pp197[119],pp197[120],pp197[121],pp197[122],pp197[123],pp197[124],pp197[125],pp197[126],pp197[127],pp197[128],pp197[129],pp197[130],pp197[131],pp197[132],pp197[133],pp197[134],pp197[135],pp197[136],pp197[137],pp197[138]};
    CLA_160 KS_49(s49, c49, in49_1, in49_2);
    wire[157:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp130[47],pp129[49],pp128[51],pp127[53],pp126[55],pp125[57],pp124[59],pp123[61],pp122[63],pp121[65],pp120[67],pp119[69],pp118[71],pp117[73],pp116[75],pp115[77],pp114[79],pp113[81],pp112[83],pp111[85],pp110[87],pp109[89],pp108[91],pp108[92],pp108[93],pp108[94],pp108[95],pp108[96],pp108[97],pp108[98],pp108[99],pp99[109],pp98[111],pp97[113],pp96[115],pp95[117],pp94[119],pp93[121],pp92[123],pp91[125],pp90[127],pp89[129],pp88[131],pp87[133],pp86[135],pp85[137],pp84[139],pp83[141],pp82[143],pp81[145],pp80[147],pp79[149],pp78[151],pp77[153],pp76[155],pp75[157],pp74[159],pp73[161],pp72[163],pp71[165],pp70[167],pp69[169],pp68[171],pp67[173],pp66[175],pp65[177],pp64[179],pp63[181],pp62[183],pp61[185],pp60[187],pp59[189],pp58[191],pp57[193],pp56[195],pp55[197],pp54[199],pp53[201],pp52[203],pp51[205],pp50[207],pp49[209],pp48[211],pp47[213],pp46[215],pp45[217],pp44[219],pp43[221],pp42[223],pp42[224],pp42[225],pp42[226],pp42[227],pp42[228],pp42[229],pp42[230],pp42[231],pp42[232],pp42[233],pp42[234],pp42[235],pp42[236],pp42[237],pp42[238],pp42[239],pp42[240],pp42[241],pp42[242],pp42[243],pp42[244],pp42[245],pp42[246],pp42[247],pp42[248],pp42[249],pp42[250],pp42[251],pp42[252],pp42[253],pp42[254],pp42[255],pp198[100],pp198[101],pp198[102],pp198[103],pp198[104],pp198[105],pp198[106],pp198[107],pp198[108],pp198[109],pp198[110],pp198[111],pp198[112],pp198[113],pp198[114],pp198[115],pp198[116],pp198[117],pp198[118],pp198[119],pp198[120],pp198[121],pp198[122],pp198[123],pp198[124],pp198[125],pp198[126],pp198[127],pp198[128],pp198[129],pp198[130],pp198[131],pp198[132],pp198[133],pp198[134],pp198[135],pp198[136]};
    assign in50_2 = {pp131[46],pp130[48],pp129[50],pp128[52],pp127[54],pp126[56],pp125[58],pp124[60],pp123[62],pp122[64],pp121[66],pp120[68],pp119[70],pp118[72],pp117[74],pp116[76],pp115[78],pp114[80],pp113[82],pp112[84],pp111[86],pp110[88],pp109[90],pp109[91],pp109[92],pp109[93],pp109[94],pp109[95],pp109[96],pp109[97],pp109[98],pp109[99],pp99[110],pp98[112],pp97[114],pp96[116],pp95[118],pp94[120],pp93[122],pp92[124],pp91[126],pp90[128],pp89[130],pp88[132],pp87[134],pp86[136],pp85[138],pp84[140],pp83[142],pp82[144],pp81[146],pp80[148],pp79[150],pp78[152],pp77[154],pp76[156],pp75[158],pp74[160],pp73[162],pp72[164],pp71[166],pp70[168],pp69[170],pp68[172],pp67[174],pp66[176],pp65[178],pp64[180],pp63[182],pp62[184],pp61[186],pp60[188],pp59[190],pp58[192],pp57[194],pp56[196],pp55[198],pp54[200],pp53[202],pp52[204],pp51[206],pp50[208],pp49[210],pp48[212],pp47[214],pp46[216],pp45[218],pp44[220],pp43[222],pp43[223],pp43[224],pp43[225],pp43[226],pp43[227],pp43[228],pp43[229],pp43[230],pp43[231],pp43[232],pp43[233],pp43[234],pp43[235],pp43[236],pp43[237],pp43[238],pp43[239],pp43[240],pp43[241],pp43[242],pp43[243],pp43[244],pp43[245],pp43[246],pp43[247],pp43[248],pp43[249],pp43[250],pp43[251],pp43[252],pp43[253],pp43[254],pp43[255],pp199[100],pp199[101],pp199[102],pp199[103],pp199[104],pp199[105],pp199[106],pp199[107],pp199[108],pp199[109],pp199[110],pp199[111],pp199[112],pp199[113],pp199[114],pp199[115],pp199[116],pp199[117],pp199[118],pp199[119],pp199[120],pp199[121],pp199[122],pp199[123],pp199[124],pp199[125],pp199[126],pp199[127],pp199[128],pp199[129],pp199[130],pp199[131],pp199[132],pp199[133],pp199[134],pp199[135]};
    CLA_158 KS_50(s50, c50, in50_1, in50_2);
    wire[155:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp131[47],pp130[49],pp129[51],pp128[53],pp127[55],pp126[57],pp125[59],pp124[61],pp123[63],pp122[65],pp121[67],pp120[69],pp119[71],pp118[73],pp117[75],pp116[77],pp115[79],pp114[81],pp113[83],pp112[85],pp111[87],pp110[89],pp110[90],pp110[91],pp110[92],pp110[93],pp110[94],pp110[95],pp110[96],pp110[97],pp110[98],pp110[99],pp99[111],pp98[113],pp97[115],pp96[117],pp95[119],pp94[121],pp93[123],pp92[125],pp91[127],pp90[129],pp89[131],pp88[133],pp87[135],pp86[137],pp85[139],pp84[141],pp83[143],pp82[145],pp81[147],pp80[149],pp79[151],pp78[153],pp77[155],pp76[157],pp75[159],pp74[161],pp73[163],pp72[165],pp71[167],pp70[169],pp69[171],pp68[173],pp67[175],pp66[177],pp65[179],pp64[181],pp63[183],pp62[185],pp61[187],pp60[189],pp59[191],pp58[193],pp57[195],pp56[197],pp55[199],pp54[201],pp53[203],pp52[205],pp51[207],pp50[209],pp49[211],pp48[213],pp47[215],pp46[217],pp45[219],pp44[221],pp44[222],pp44[223],pp44[224],pp44[225],pp44[226],pp44[227],pp44[228],pp44[229],pp44[230],pp44[231],pp44[232],pp44[233],pp44[234],pp44[235],pp44[236],pp44[237],pp44[238],pp44[239],pp44[240],pp44[241],pp44[242],pp44[243],pp44[244],pp44[245],pp44[246],pp44[247],pp44[248],pp44[249],pp44[250],pp44[251],pp44[252],pp44[253],pp44[254],pp44[255],pp200[100],pp200[101],pp200[102],pp200[103],pp200[104],pp200[105],pp200[106],pp200[107],pp200[108],pp200[109],pp200[110],pp200[111],pp200[112],pp200[113],pp200[114],pp200[115],pp200[116],pp200[117],pp200[118],pp200[119],pp200[120],pp200[121],pp200[122],pp200[123],pp200[124],pp200[125],pp200[126],pp200[127],pp200[128],pp200[129],pp200[130],pp200[131],pp200[132],pp200[133]};
    assign in51_2 = {pp132[46],pp131[48],pp130[50],pp129[52],pp128[54],pp127[56],pp126[58],pp125[60],pp124[62],pp123[64],pp122[66],pp121[68],pp120[70],pp119[72],pp118[74],pp117[76],pp116[78],pp115[80],pp114[82],pp113[84],pp112[86],pp111[88],pp111[89],pp111[90],pp111[91],pp111[92],pp111[93],pp111[94],pp111[95],pp111[96],pp111[97],pp111[98],pp111[99],pp99[112],pp98[114],pp97[116],pp96[118],pp95[120],pp94[122],pp93[124],pp92[126],pp91[128],pp90[130],pp89[132],pp88[134],pp87[136],pp86[138],pp85[140],pp84[142],pp83[144],pp82[146],pp81[148],pp80[150],pp79[152],pp78[154],pp77[156],pp76[158],pp75[160],pp74[162],pp73[164],pp72[166],pp71[168],pp70[170],pp69[172],pp68[174],pp67[176],pp66[178],pp65[180],pp64[182],pp63[184],pp62[186],pp61[188],pp60[190],pp59[192],pp58[194],pp57[196],pp56[198],pp55[200],pp54[202],pp53[204],pp52[206],pp51[208],pp50[210],pp49[212],pp48[214],pp47[216],pp46[218],pp45[220],pp45[221],pp45[222],pp45[223],pp45[224],pp45[225],pp45[226],pp45[227],pp45[228],pp45[229],pp45[230],pp45[231],pp45[232],pp45[233],pp45[234],pp45[235],pp45[236],pp45[237],pp45[238],pp45[239],pp45[240],pp45[241],pp45[242],pp45[243],pp45[244],pp45[245],pp45[246],pp45[247],pp45[248],pp45[249],pp45[250],pp45[251],pp45[252],pp45[253],pp45[254],pp45[255],pp201[100],pp201[101],pp201[102],pp201[103],pp201[104],pp201[105],pp201[106],pp201[107],pp201[108],pp201[109],pp201[110],pp201[111],pp201[112],pp201[113],pp201[114],pp201[115],pp201[116],pp201[117],pp201[118],pp201[119],pp201[120],pp201[121],pp201[122],pp201[123],pp201[124],pp201[125],pp201[126],pp201[127],pp201[128],pp201[129],pp201[130],pp201[131],pp201[132]};
    CLA_156 KS_51(s51, c51, in51_1, in51_2);
    wire[153:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp132[47],pp131[49],pp130[51],pp129[53],pp128[55],pp127[57],pp126[59],pp125[61],pp124[63],pp123[65],pp122[67],pp121[69],pp120[71],pp119[73],pp118[75],pp117[77],pp116[79],pp115[81],pp114[83],pp113[85],pp112[87],pp112[88],pp112[89],pp112[90],pp112[91],pp112[92],pp112[93],pp112[94],pp112[95],pp112[96],pp112[97],pp112[98],pp112[99],pp99[113],pp98[115],pp97[117],pp96[119],pp95[121],pp94[123],pp93[125],pp92[127],pp91[129],pp90[131],pp89[133],pp88[135],pp87[137],pp86[139],pp85[141],pp84[143],pp83[145],pp82[147],pp81[149],pp80[151],pp79[153],pp78[155],pp77[157],pp76[159],pp75[161],pp74[163],pp73[165],pp72[167],pp71[169],pp70[171],pp69[173],pp68[175],pp67[177],pp66[179],pp65[181],pp64[183],pp63[185],pp62[187],pp61[189],pp60[191],pp59[193],pp58[195],pp57[197],pp56[199],pp55[201],pp54[203],pp53[205],pp52[207],pp51[209],pp50[211],pp49[213],pp48[215],pp47[217],pp46[219],pp46[220],pp46[221],pp46[222],pp46[223],pp46[224],pp46[225],pp46[226],pp46[227],pp46[228],pp46[229],pp46[230],pp46[231],pp46[232],pp46[233],pp46[234],pp46[235],pp46[236],pp46[237],pp46[238],pp46[239],pp46[240],pp46[241],pp46[242],pp46[243],pp46[244],pp46[245],pp46[246],pp46[247],pp46[248],pp46[249],pp46[250],pp46[251],pp46[252],pp46[253],pp46[254],pp46[255],pp202[100],pp202[101],pp202[102],pp202[103],pp202[104],pp202[105],pp202[106],pp202[107],pp202[108],pp202[109],pp202[110],pp202[111],pp202[112],pp202[113],pp202[114],pp202[115],pp202[116],pp202[117],pp202[118],pp202[119],pp202[120],pp202[121],pp202[122],pp202[123],pp202[124],pp202[125],pp202[126],pp202[127],pp202[128],pp202[129],pp202[130]};
    assign in52_2 = {pp133[46],pp132[48],pp131[50],pp130[52],pp129[54],pp128[56],pp127[58],pp126[60],pp125[62],pp124[64],pp123[66],pp122[68],pp121[70],pp120[72],pp119[74],pp118[76],pp117[78],pp116[80],pp115[82],pp114[84],pp113[86],pp113[87],pp113[88],pp113[89],pp113[90],pp113[91],pp113[92],pp113[93],pp113[94],pp113[95],pp113[96],pp113[97],pp113[98],pp113[99],pp99[114],pp98[116],pp97[118],pp96[120],pp95[122],pp94[124],pp93[126],pp92[128],pp91[130],pp90[132],pp89[134],pp88[136],pp87[138],pp86[140],pp85[142],pp84[144],pp83[146],pp82[148],pp81[150],pp80[152],pp79[154],pp78[156],pp77[158],pp76[160],pp75[162],pp74[164],pp73[166],pp72[168],pp71[170],pp70[172],pp69[174],pp68[176],pp67[178],pp66[180],pp65[182],pp64[184],pp63[186],pp62[188],pp61[190],pp60[192],pp59[194],pp58[196],pp57[198],pp56[200],pp55[202],pp54[204],pp53[206],pp52[208],pp51[210],pp50[212],pp49[214],pp48[216],pp47[218],pp47[219],pp47[220],pp47[221],pp47[222],pp47[223],pp47[224],pp47[225],pp47[226],pp47[227],pp47[228],pp47[229],pp47[230],pp47[231],pp47[232],pp47[233],pp47[234],pp47[235],pp47[236],pp47[237],pp47[238],pp47[239],pp47[240],pp47[241],pp47[242],pp47[243],pp47[244],pp47[245],pp47[246],pp47[247],pp47[248],pp47[249],pp47[250],pp47[251],pp47[252],pp47[253],pp47[254],pp47[255],pp203[100],pp203[101],pp203[102],pp203[103],pp203[104],pp203[105],pp203[106],pp203[107],pp203[108],pp203[109],pp203[110],pp203[111],pp203[112],pp203[113],pp203[114],pp203[115],pp203[116],pp203[117],pp203[118],pp203[119],pp203[120],pp203[121],pp203[122],pp203[123],pp203[124],pp203[125],pp203[126],pp203[127],pp203[128],pp203[129]};
    CLA_154 KS_52(s52, c52, in52_1, in52_2);
    wire[151:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp133[47],pp132[49],pp131[51],pp130[53],pp129[55],pp128[57],pp127[59],pp126[61],pp125[63],pp124[65],pp123[67],pp122[69],pp121[71],pp120[73],pp119[75],pp118[77],pp117[79],pp116[81],pp115[83],pp114[85],pp114[86],pp114[87],pp114[88],pp114[89],pp114[90],pp114[91],pp114[92],pp114[93],pp114[94],pp114[95],pp114[96],pp114[97],pp114[98],pp114[99],pp99[115],pp98[117],pp97[119],pp96[121],pp95[123],pp94[125],pp93[127],pp92[129],pp91[131],pp90[133],pp89[135],pp88[137],pp87[139],pp86[141],pp85[143],pp84[145],pp83[147],pp82[149],pp81[151],pp80[153],pp79[155],pp78[157],pp77[159],pp76[161],pp75[163],pp74[165],pp73[167],pp72[169],pp71[171],pp70[173],pp69[175],pp68[177],pp67[179],pp66[181],pp65[183],pp64[185],pp63[187],pp62[189],pp61[191],pp60[193],pp59[195],pp58[197],pp57[199],pp56[201],pp55[203],pp54[205],pp53[207],pp52[209],pp51[211],pp50[213],pp49[215],pp48[217],pp48[218],pp48[219],pp48[220],pp48[221],pp48[222],pp48[223],pp48[224],pp48[225],pp48[226],pp48[227],pp48[228],pp48[229],pp48[230],pp48[231],pp48[232],pp48[233],pp48[234],pp48[235],pp48[236],pp48[237],pp48[238],pp48[239],pp48[240],pp48[241],pp48[242],pp48[243],pp48[244],pp48[245],pp48[246],pp48[247],pp48[248],pp48[249],pp48[250],pp48[251],pp48[252],pp48[253],pp48[254],pp48[255],pp204[100],pp204[101],pp204[102],pp204[103],pp204[104],pp204[105],pp204[106],pp204[107],pp204[108],pp204[109],pp204[110],pp204[111],pp204[112],pp204[113],pp204[114],pp204[115],pp204[116],pp204[117],pp204[118],pp204[119],pp204[120],pp204[121],pp204[122],pp204[123],pp204[124],pp204[125],pp204[126],pp204[127]};
    assign in53_2 = {pp134[46],pp133[48],pp132[50],pp131[52],pp130[54],pp129[56],pp128[58],pp127[60],pp126[62],pp125[64],pp124[66],pp123[68],pp122[70],pp121[72],pp120[74],pp119[76],pp118[78],pp117[80],pp116[82],pp115[84],pp115[85],pp115[86],pp115[87],pp115[88],pp115[89],pp115[90],pp115[91],pp115[92],pp115[93],pp115[94],pp115[95],pp115[96],pp115[97],pp115[98],pp115[99],pp99[116],pp98[118],pp97[120],pp96[122],pp95[124],pp94[126],pp93[128],pp92[130],pp91[132],pp90[134],pp89[136],pp88[138],pp87[140],pp86[142],pp85[144],pp84[146],pp83[148],pp82[150],pp81[152],pp80[154],pp79[156],pp78[158],pp77[160],pp76[162],pp75[164],pp74[166],pp73[168],pp72[170],pp71[172],pp70[174],pp69[176],pp68[178],pp67[180],pp66[182],pp65[184],pp64[186],pp63[188],pp62[190],pp61[192],pp60[194],pp59[196],pp58[198],pp57[200],pp56[202],pp55[204],pp54[206],pp53[208],pp52[210],pp51[212],pp50[214],pp49[216],pp49[217],pp49[218],pp49[219],pp49[220],pp49[221],pp49[222],pp49[223],pp49[224],pp49[225],pp49[226],pp49[227],pp49[228],pp49[229],pp49[230],pp49[231],pp49[232],pp49[233],pp49[234],pp49[235],pp49[236],pp49[237],pp49[238],pp49[239],pp49[240],pp49[241],pp49[242],pp49[243],pp49[244],pp49[245],pp49[246],pp49[247],pp49[248],pp49[249],pp49[250],pp49[251],pp49[252],pp49[253],pp49[254],pp49[255],pp205[100],pp205[101],pp205[102],pp205[103],pp205[104],pp205[105],pp205[106],pp205[107],pp205[108],pp205[109],pp205[110],pp205[111],pp205[112],pp205[113],pp205[114],pp205[115],pp205[116],pp205[117],pp205[118],pp205[119],pp205[120],pp205[121],pp205[122],pp205[123],pp205[124],pp205[125],pp205[126]};
    CLA_152 KS_53(s53, c53, in53_1, in53_2);
    wire[149:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp134[47],pp133[49],pp132[51],pp131[53],pp130[55],pp129[57],pp128[59],pp127[61],pp126[63],pp125[65],pp124[67],pp123[69],pp122[71],pp121[73],pp120[75],pp119[77],pp118[79],pp117[81],pp116[83],pp116[84],pp116[85],pp116[86],pp116[87],pp116[88],pp116[89],pp116[90],pp116[91],pp116[92],pp116[93],pp116[94],pp116[95],pp116[96],pp116[97],pp116[98],pp116[99],pp99[117],pp98[119],pp97[121],pp96[123],pp95[125],pp94[127],pp93[129],pp92[131],pp91[133],pp90[135],pp89[137],pp88[139],pp87[141],pp86[143],pp85[145],pp84[147],pp83[149],pp82[151],pp81[153],pp80[155],pp79[157],pp78[159],pp77[161],pp76[163],pp75[165],pp74[167],pp73[169],pp72[171],pp71[173],pp70[175],pp69[177],pp68[179],pp67[181],pp66[183],pp65[185],pp64[187],pp63[189],pp62[191],pp61[193],pp60[195],pp59[197],pp58[199],pp57[201],pp56[203],pp55[205],pp54[207],pp53[209],pp52[211],pp51[213],pp50[215],pp50[216],pp50[217],pp50[218],pp50[219],pp50[220],pp50[221],pp50[222],pp50[223],pp50[224],pp50[225],pp50[226],pp50[227],pp50[228],pp50[229],pp50[230],pp50[231],pp50[232],pp50[233],pp50[234],pp50[235],pp50[236],pp50[237],pp50[238],pp50[239],pp50[240],pp50[241],pp50[242],pp50[243],pp50[244],pp50[245],pp50[246],pp50[247],pp50[248],pp50[249],pp50[250],pp50[251],pp50[252],pp50[253],pp50[254],pp50[255],pp206[100],pp206[101],pp206[102],pp206[103],pp206[104],pp206[105],pp206[106],pp206[107],pp206[108],pp206[109],pp206[110],pp206[111],pp206[112],pp206[113],pp206[114],pp206[115],pp206[116],pp206[117],pp206[118],pp206[119],pp206[120],pp206[121],pp206[122],pp206[123],pp206[124]};
    assign in54_2 = {pp135[46],pp134[48],pp133[50],pp132[52],pp131[54],pp130[56],pp129[58],pp128[60],pp127[62],pp126[64],pp125[66],pp124[68],pp123[70],pp122[72],pp121[74],pp120[76],pp119[78],pp118[80],pp117[82],pp117[83],pp117[84],pp117[85],pp117[86],pp117[87],pp117[88],pp117[89],pp117[90],pp117[91],pp117[92],pp117[93],pp117[94],pp117[95],pp117[96],pp117[97],pp117[98],pp117[99],pp99[118],pp98[120],pp97[122],pp96[124],pp95[126],pp94[128],pp93[130],pp92[132],pp91[134],pp90[136],pp89[138],pp88[140],pp87[142],pp86[144],pp85[146],pp84[148],pp83[150],pp82[152],pp81[154],pp80[156],pp79[158],pp78[160],pp77[162],pp76[164],pp75[166],pp74[168],pp73[170],pp72[172],pp71[174],pp70[176],pp69[178],pp68[180],pp67[182],pp66[184],pp65[186],pp64[188],pp63[190],pp62[192],pp61[194],pp60[196],pp59[198],pp58[200],pp57[202],pp56[204],pp55[206],pp54[208],pp53[210],pp52[212],pp51[214],pp51[215],pp51[216],pp51[217],pp51[218],pp51[219],pp51[220],pp51[221],pp51[222],pp51[223],pp51[224],pp51[225],pp51[226],pp51[227],pp51[228],pp51[229],pp51[230],pp51[231],pp51[232],pp51[233],pp51[234],pp51[235],pp51[236],pp51[237],pp51[238],pp51[239],pp51[240],pp51[241],pp51[242],pp51[243],pp51[244],pp51[245],pp51[246],pp51[247],pp51[248],pp51[249],pp51[250],pp51[251],pp51[252],pp51[253],pp51[254],pp51[255],pp207[100],pp207[101],pp207[102],pp207[103],pp207[104],pp207[105],pp207[106],pp207[107],pp207[108],pp207[109],pp207[110],pp207[111],pp207[112],pp207[113],pp207[114],pp207[115],pp207[116],pp207[117],pp207[118],pp207[119],pp207[120],pp207[121],pp207[122],pp207[123]};
    CLA_150 KS_54(s54, c54, in54_1, in54_2);
    wire[147:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp135[47],pp134[49],pp133[51],pp132[53],pp131[55],pp130[57],pp129[59],pp128[61],pp127[63],pp126[65],pp125[67],pp124[69],pp123[71],pp122[73],pp121[75],pp120[77],pp119[79],pp118[81],pp118[82],pp118[83],pp118[84],pp118[85],pp118[86],pp118[87],pp118[88],pp118[89],pp118[90],pp118[91],pp118[92],pp118[93],pp118[94],pp118[95],pp118[96],pp118[97],pp118[98],pp118[99],pp99[119],pp98[121],pp97[123],pp96[125],pp95[127],pp94[129],pp93[131],pp92[133],pp91[135],pp90[137],pp89[139],pp88[141],pp87[143],pp86[145],pp85[147],pp84[149],pp83[151],pp82[153],pp81[155],pp80[157],pp79[159],pp78[161],pp77[163],pp76[165],pp75[167],pp74[169],pp73[171],pp72[173],pp71[175],pp70[177],pp69[179],pp68[181],pp67[183],pp66[185],pp65[187],pp64[189],pp63[191],pp62[193],pp61[195],pp60[197],pp59[199],pp58[201],pp57[203],pp56[205],pp55[207],pp54[209],pp53[211],pp52[213],pp52[214],pp52[215],pp52[216],pp52[217],pp52[218],pp52[219],pp52[220],pp52[221],pp52[222],pp52[223],pp52[224],pp52[225],pp52[226],pp52[227],pp52[228],pp52[229],pp52[230],pp52[231],pp52[232],pp52[233],pp52[234],pp52[235],pp52[236],pp52[237],pp52[238],pp52[239],pp52[240],pp52[241],pp52[242],pp52[243],pp52[244],pp52[245],pp52[246],pp52[247],pp52[248],pp52[249],pp52[250],pp52[251],pp52[252],pp52[253],pp52[254],pp52[255],pp208[100],pp208[101],pp208[102],pp208[103],pp208[104],pp208[105],pp208[106],pp208[107],pp208[108],pp208[109],pp208[110],pp208[111],pp208[112],pp208[113],pp208[114],pp208[115],pp208[116],pp208[117],pp208[118],pp208[119],pp208[120],pp208[121]};
    assign in55_2 = {pp136[46],pp135[48],pp134[50],pp133[52],pp132[54],pp131[56],pp130[58],pp129[60],pp128[62],pp127[64],pp126[66],pp125[68],pp124[70],pp123[72],pp122[74],pp121[76],pp120[78],pp119[80],pp119[81],pp119[82],pp119[83],pp119[84],pp119[85],pp119[86],pp119[87],pp119[88],pp119[89],pp119[90],pp119[91],pp119[92],pp119[93],pp119[94],pp119[95],pp119[96],pp119[97],pp119[98],pp119[99],pp99[120],pp98[122],pp97[124],pp96[126],pp95[128],pp94[130],pp93[132],pp92[134],pp91[136],pp90[138],pp89[140],pp88[142],pp87[144],pp86[146],pp85[148],pp84[150],pp83[152],pp82[154],pp81[156],pp80[158],pp79[160],pp78[162],pp77[164],pp76[166],pp75[168],pp74[170],pp73[172],pp72[174],pp71[176],pp70[178],pp69[180],pp68[182],pp67[184],pp66[186],pp65[188],pp64[190],pp63[192],pp62[194],pp61[196],pp60[198],pp59[200],pp58[202],pp57[204],pp56[206],pp55[208],pp54[210],pp53[212],pp53[213],pp53[214],pp53[215],pp53[216],pp53[217],pp53[218],pp53[219],pp53[220],pp53[221],pp53[222],pp53[223],pp53[224],pp53[225],pp53[226],pp53[227],pp53[228],pp53[229],pp53[230],pp53[231],pp53[232],pp53[233],pp53[234],pp53[235],pp53[236],pp53[237],pp53[238],pp53[239],pp53[240],pp53[241],pp53[242],pp53[243],pp53[244],pp53[245],pp53[246],pp53[247],pp53[248],pp53[249],pp53[250],pp53[251],pp53[252],pp53[253],pp53[254],pp53[255],pp209[100],pp209[101],pp209[102],pp209[103],pp209[104],pp209[105],pp209[106],pp209[107],pp209[108],pp209[109],pp209[110],pp209[111],pp209[112],pp209[113],pp209[114],pp209[115],pp209[116],pp209[117],pp209[118],pp209[119],pp209[120]};
    CLA_148 KS_55(s55, c55, in55_1, in55_2);
    wire[145:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp136[47],pp135[49],pp134[51],pp133[53],pp132[55],pp131[57],pp130[59],pp129[61],pp128[63],pp127[65],pp126[67],pp125[69],pp124[71],pp123[73],pp122[75],pp121[77],pp120[79],pp120[80],pp120[81],pp120[82],pp120[83],pp120[84],pp120[85],pp120[86],pp120[87],pp120[88],pp120[89],pp120[90],pp120[91],pp120[92],pp120[93],pp120[94],pp120[95],pp120[96],pp120[97],pp120[98],pp120[99],pp99[121],pp98[123],pp97[125],pp96[127],pp95[129],pp94[131],pp93[133],pp92[135],pp91[137],pp90[139],pp89[141],pp88[143],pp87[145],pp86[147],pp85[149],pp84[151],pp83[153],pp82[155],pp81[157],pp80[159],pp79[161],pp78[163],pp77[165],pp76[167],pp75[169],pp74[171],pp73[173],pp72[175],pp71[177],pp70[179],pp69[181],pp68[183],pp67[185],pp66[187],pp65[189],pp64[191],pp63[193],pp62[195],pp61[197],pp60[199],pp59[201],pp58[203],pp57[205],pp56[207],pp55[209],pp54[211],pp54[212],pp54[213],pp54[214],pp54[215],pp54[216],pp54[217],pp54[218],pp54[219],pp54[220],pp54[221],pp54[222],pp54[223],pp54[224],pp54[225],pp54[226],pp54[227],pp54[228],pp54[229],pp54[230],pp54[231],pp54[232],pp54[233],pp54[234],pp54[235],pp54[236],pp54[237],pp54[238],pp54[239],pp54[240],pp54[241],pp54[242],pp54[243],pp54[244],pp54[245],pp54[246],pp54[247],pp54[248],pp54[249],pp54[250],pp54[251],pp54[252],pp54[253],pp54[254],pp54[255],pp210[100],pp210[101],pp210[102],pp210[103],pp210[104],pp210[105],pp210[106],pp210[107],pp210[108],pp210[109],pp210[110],pp210[111],pp210[112],pp210[113],pp210[114],pp210[115],pp210[116],pp210[117],pp210[118]};
    assign in56_2 = {pp137[46],pp136[48],pp135[50],pp134[52],pp133[54],pp132[56],pp131[58],pp130[60],pp129[62],pp128[64],pp127[66],pp126[68],pp125[70],pp124[72],pp123[74],pp122[76],pp121[78],pp121[79],pp121[80],pp121[81],pp121[82],pp121[83],pp121[84],pp121[85],pp121[86],pp121[87],pp121[88],pp121[89],pp121[90],pp121[91],pp121[92],pp121[93],pp121[94],pp121[95],pp121[96],pp121[97],pp121[98],pp121[99],pp99[122],pp98[124],pp97[126],pp96[128],pp95[130],pp94[132],pp93[134],pp92[136],pp91[138],pp90[140],pp89[142],pp88[144],pp87[146],pp86[148],pp85[150],pp84[152],pp83[154],pp82[156],pp81[158],pp80[160],pp79[162],pp78[164],pp77[166],pp76[168],pp75[170],pp74[172],pp73[174],pp72[176],pp71[178],pp70[180],pp69[182],pp68[184],pp67[186],pp66[188],pp65[190],pp64[192],pp63[194],pp62[196],pp61[198],pp60[200],pp59[202],pp58[204],pp57[206],pp56[208],pp55[210],pp55[211],pp55[212],pp55[213],pp55[214],pp55[215],pp55[216],pp55[217],pp55[218],pp55[219],pp55[220],pp55[221],pp55[222],pp55[223],pp55[224],pp55[225],pp55[226],pp55[227],pp55[228],pp55[229],pp55[230],pp55[231],pp55[232],pp55[233],pp55[234],pp55[235],pp55[236],pp55[237],pp55[238],pp55[239],pp55[240],pp55[241],pp55[242],pp55[243],pp55[244],pp55[245],pp55[246],pp55[247],pp55[248],pp55[249],pp55[250],pp55[251],pp55[252],pp55[253],pp55[254],pp55[255],pp211[100],pp211[101],pp211[102],pp211[103],pp211[104],pp211[105],pp211[106],pp211[107],pp211[108],pp211[109],pp211[110],pp211[111],pp211[112],pp211[113],pp211[114],pp211[115],pp211[116],pp211[117]};
    CLA_146 KS_56(s56, c56, in56_1, in56_2);
    wire[143:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp137[47],pp136[49],pp135[51],pp134[53],pp133[55],pp132[57],pp131[59],pp130[61],pp129[63],pp128[65],pp127[67],pp126[69],pp125[71],pp124[73],pp123[75],pp122[77],pp122[78],pp122[79],pp122[80],pp122[81],pp122[82],pp122[83],pp122[84],pp122[85],pp122[86],pp122[87],pp122[88],pp122[89],pp122[90],pp122[91],pp122[92],pp122[93],pp122[94],pp122[95],pp122[96],pp122[97],pp122[98],pp122[99],pp99[123],pp98[125],pp97[127],pp96[129],pp95[131],pp94[133],pp93[135],pp92[137],pp91[139],pp90[141],pp89[143],pp88[145],pp87[147],pp86[149],pp85[151],pp84[153],pp83[155],pp82[157],pp81[159],pp80[161],pp79[163],pp78[165],pp77[167],pp76[169],pp75[171],pp74[173],pp73[175],pp72[177],pp71[179],pp70[181],pp69[183],pp68[185],pp67[187],pp66[189],pp65[191],pp64[193],pp63[195],pp62[197],pp61[199],pp60[201],pp59[203],pp58[205],pp57[207],pp56[209],pp56[210],pp56[211],pp56[212],pp56[213],pp56[214],pp56[215],pp56[216],pp56[217],pp56[218],pp56[219],pp56[220],pp56[221],pp56[222],pp56[223],pp56[224],pp56[225],pp56[226],pp56[227],pp56[228],pp56[229],pp56[230],pp56[231],pp56[232],pp56[233],pp56[234],pp56[235],pp56[236],pp56[237],pp56[238],pp56[239],pp56[240],pp56[241],pp56[242],pp56[243],pp56[244],pp56[245],pp56[246],pp56[247],pp56[248],pp56[249],pp56[250],pp56[251],pp56[252],pp56[253],pp56[254],pp56[255],pp212[100],pp212[101],pp212[102],pp212[103],pp212[104],pp212[105],pp212[106],pp212[107],pp212[108],pp212[109],pp212[110],pp212[111],pp212[112],pp212[113],pp212[114],pp212[115]};
    assign in57_2 = {pp138[46],pp137[48],pp136[50],pp135[52],pp134[54],pp133[56],pp132[58],pp131[60],pp130[62],pp129[64],pp128[66],pp127[68],pp126[70],pp125[72],pp124[74],pp123[76],pp123[77],pp123[78],pp123[79],pp123[80],pp123[81],pp123[82],pp123[83],pp123[84],pp123[85],pp123[86],pp123[87],pp123[88],pp123[89],pp123[90],pp123[91],pp123[92],pp123[93],pp123[94],pp123[95],pp123[96],pp123[97],pp123[98],pp123[99],pp99[124],pp98[126],pp97[128],pp96[130],pp95[132],pp94[134],pp93[136],pp92[138],pp91[140],pp90[142],pp89[144],pp88[146],pp87[148],pp86[150],pp85[152],pp84[154],pp83[156],pp82[158],pp81[160],pp80[162],pp79[164],pp78[166],pp77[168],pp76[170],pp75[172],pp74[174],pp73[176],pp72[178],pp71[180],pp70[182],pp69[184],pp68[186],pp67[188],pp66[190],pp65[192],pp64[194],pp63[196],pp62[198],pp61[200],pp60[202],pp59[204],pp58[206],pp57[208],pp57[209],pp57[210],pp57[211],pp57[212],pp57[213],pp57[214],pp57[215],pp57[216],pp57[217],pp57[218],pp57[219],pp57[220],pp57[221],pp57[222],pp57[223],pp57[224],pp57[225],pp57[226],pp57[227],pp57[228],pp57[229],pp57[230],pp57[231],pp57[232],pp57[233],pp57[234],pp57[235],pp57[236],pp57[237],pp57[238],pp57[239],pp57[240],pp57[241],pp57[242],pp57[243],pp57[244],pp57[245],pp57[246],pp57[247],pp57[248],pp57[249],pp57[250],pp57[251],pp57[252],pp57[253],pp57[254],pp57[255],pp213[100],pp213[101],pp213[102],pp213[103],pp213[104],pp213[105],pp213[106],pp213[107],pp213[108],pp213[109],pp213[110],pp213[111],pp213[112],pp213[113],pp213[114]};
    CLA_144 KS_57(s57, c57, in57_1, in57_2);
    wire[141:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp138[47],pp137[49],pp136[51],pp135[53],pp134[55],pp133[57],pp132[59],pp131[61],pp130[63],pp129[65],pp128[67],pp127[69],pp126[71],pp125[73],pp124[75],pp124[76],pp124[77],pp124[78],pp124[79],pp124[80],pp124[81],pp124[82],pp124[83],pp124[84],pp124[85],pp124[86],pp124[87],pp124[88],pp124[89],pp124[90],pp124[91],pp124[92],pp124[93],pp124[94],pp124[95],pp124[96],pp124[97],pp124[98],pp124[99],pp99[125],pp98[127],pp97[129],pp96[131],pp95[133],pp94[135],pp93[137],pp92[139],pp91[141],pp90[143],pp89[145],pp88[147],pp87[149],pp86[151],pp85[153],pp84[155],pp83[157],pp82[159],pp81[161],pp80[163],pp79[165],pp78[167],pp77[169],pp76[171],pp75[173],pp74[175],pp73[177],pp72[179],pp71[181],pp70[183],pp69[185],pp68[187],pp67[189],pp66[191],pp65[193],pp64[195],pp63[197],pp62[199],pp61[201],pp60[203],pp59[205],pp58[207],pp58[208],pp58[209],pp58[210],pp58[211],pp58[212],pp58[213],pp58[214],pp58[215],pp58[216],pp58[217],pp58[218],pp58[219],pp58[220],pp58[221],pp58[222],pp58[223],pp58[224],pp58[225],pp58[226],pp58[227],pp58[228],pp58[229],pp58[230],pp58[231],pp58[232],pp58[233],pp58[234],pp58[235],pp58[236],pp58[237],pp58[238],pp58[239],pp58[240],pp58[241],pp58[242],pp58[243],pp58[244],pp58[245],pp58[246],pp58[247],pp58[248],pp58[249],pp58[250],pp58[251],pp58[252],pp58[253],pp58[254],pp58[255],pp214[100],pp214[101],pp214[102],pp214[103],pp214[104],pp214[105],pp214[106],pp214[107],pp214[108],pp214[109],pp214[110],pp214[111],pp214[112]};
    assign in58_2 = {pp139[46],pp138[48],pp137[50],pp136[52],pp135[54],pp134[56],pp133[58],pp132[60],pp131[62],pp130[64],pp129[66],pp128[68],pp127[70],pp126[72],pp125[74],pp125[75],pp125[76],pp125[77],pp125[78],pp125[79],pp125[80],pp125[81],pp125[82],pp125[83],pp125[84],pp125[85],pp125[86],pp125[87],pp125[88],pp125[89],pp125[90],pp125[91],pp125[92],pp125[93],pp125[94],pp125[95],pp125[96],pp125[97],pp125[98],pp125[99],pp99[126],pp98[128],pp97[130],pp96[132],pp95[134],pp94[136],pp93[138],pp92[140],pp91[142],pp90[144],pp89[146],pp88[148],pp87[150],pp86[152],pp85[154],pp84[156],pp83[158],pp82[160],pp81[162],pp80[164],pp79[166],pp78[168],pp77[170],pp76[172],pp75[174],pp74[176],pp73[178],pp72[180],pp71[182],pp70[184],pp69[186],pp68[188],pp67[190],pp66[192],pp65[194],pp64[196],pp63[198],pp62[200],pp61[202],pp60[204],pp59[206],pp59[207],pp59[208],pp59[209],pp59[210],pp59[211],pp59[212],pp59[213],pp59[214],pp59[215],pp59[216],pp59[217],pp59[218],pp59[219],pp59[220],pp59[221],pp59[222],pp59[223],pp59[224],pp59[225],pp59[226],pp59[227],pp59[228],pp59[229],pp59[230],pp59[231],pp59[232],pp59[233],pp59[234],pp59[235],pp59[236],pp59[237],pp59[238],pp59[239],pp59[240],pp59[241],pp59[242],pp59[243],pp59[244],pp59[245],pp59[246],pp59[247],pp59[248],pp59[249],pp59[250],pp59[251],pp59[252],pp59[253],pp59[254],pp59[255],pp215[100],pp215[101],pp215[102],pp215[103],pp215[104],pp215[105],pp215[106],pp215[107],pp215[108],pp215[109],pp215[110],pp215[111]};
    CLA_142 KS_58(s58, c58, in58_1, in58_2);
    wire[139:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp139[47],pp138[49],pp137[51],pp136[53],pp135[55],pp134[57],pp133[59],pp132[61],pp131[63],pp130[65],pp129[67],pp128[69],pp127[71],pp126[73],pp126[74],pp126[75],pp126[76],pp126[77],pp126[78],pp126[79],pp126[80],pp126[81],pp126[82],pp126[83],pp126[84],pp126[85],pp126[86],pp126[87],pp126[88],pp126[89],pp126[90],pp126[91],pp126[92],pp126[93],pp126[94],pp126[95],pp126[96],pp126[97],pp126[98],pp126[99],pp99[127],pp98[129],pp97[131],pp96[133],pp95[135],pp94[137],pp93[139],pp92[141],pp91[143],pp90[145],pp89[147],pp88[149],pp87[151],pp86[153],pp85[155],pp84[157],pp83[159],pp82[161],pp81[163],pp80[165],pp79[167],pp78[169],pp77[171],pp76[173],pp75[175],pp74[177],pp73[179],pp72[181],pp71[183],pp70[185],pp69[187],pp68[189],pp67[191],pp66[193],pp65[195],pp64[197],pp63[199],pp62[201],pp61[203],pp60[205],pp60[206],pp60[207],pp60[208],pp60[209],pp60[210],pp60[211],pp60[212],pp60[213],pp60[214],pp60[215],pp60[216],pp60[217],pp60[218],pp60[219],pp60[220],pp60[221],pp60[222],pp60[223],pp60[224],pp60[225],pp60[226],pp60[227],pp60[228],pp60[229],pp60[230],pp60[231],pp60[232],pp60[233],pp60[234],pp60[235],pp60[236],pp60[237],pp60[238],pp60[239],pp60[240],pp60[241],pp60[242],pp60[243],pp60[244],pp60[245],pp60[246],pp60[247],pp60[248],pp60[249],pp60[250],pp60[251],pp60[252],pp60[253],pp60[254],pp60[255],pp216[100],pp216[101],pp216[102],pp216[103],pp216[104],pp216[105],pp216[106],pp216[107],pp216[108],pp216[109]};
    assign in59_2 = {pp140[46],pp139[48],pp138[50],pp137[52],pp136[54],pp135[56],pp134[58],pp133[60],pp132[62],pp131[64],pp130[66],pp129[68],pp128[70],pp127[72],pp127[73],pp127[74],pp127[75],pp127[76],pp127[77],pp127[78],pp127[79],pp127[80],pp127[81],pp127[82],pp127[83],pp127[84],pp127[85],pp127[86],pp127[87],pp127[88],pp127[89],pp127[90],pp127[91],pp127[92],pp127[93],pp127[94],pp127[95],pp127[96],pp127[97],pp127[98],pp127[99],pp99[128],pp98[130],pp97[132],pp96[134],pp95[136],pp94[138],pp93[140],pp92[142],pp91[144],pp90[146],pp89[148],pp88[150],pp87[152],pp86[154],pp85[156],pp84[158],pp83[160],pp82[162],pp81[164],pp80[166],pp79[168],pp78[170],pp77[172],pp76[174],pp75[176],pp74[178],pp73[180],pp72[182],pp71[184],pp70[186],pp69[188],pp68[190],pp67[192],pp66[194],pp65[196],pp64[198],pp63[200],pp62[202],pp61[204],pp61[205],pp61[206],pp61[207],pp61[208],pp61[209],pp61[210],pp61[211],pp61[212],pp61[213],pp61[214],pp61[215],pp61[216],pp61[217],pp61[218],pp61[219],pp61[220],pp61[221],pp61[222],pp61[223],pp61[224],pp61[225],pp61[226],pp61[227],pp61[228],pp61[229],pp61[230],pp61[231],pp61[232],pp61[233],pp61[234],pp61[235],pp61[236],pp61[237],pp61[238],pp61[239],pp61[240],pp61[241],pp61[242],pp61[243],pp61[244],pp61[245],pp61[246],pp61[247],pp61[248],pp61[249],pp61[250],pp61[251],pp61[252],pp61[253],pp61[254],pp61[255],pp217[100],pp217[101],pp217[102],pp217[103],pp217[104],pp217[105],pp217[106],pp217[107],pp217[108]};
    CLA_140 KS_59(s59, c59, in59_1, in59_2);
    wire[137:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp140[47],pp139[49],pp138[51],pp137[53],pp136[55],pp135[57],pp134[59],pp133[61],pp132[63],pp131[65],pp130[67],pp129[69],pp128[71],pp128[72],pp128[73],pp128[74],pp128[75],pp128[76],pp128[77],pp128[78],pp128[79],pp128[80],pp128[81],pp128[82],pp128[83],pp128[84],pp128[85],pp128[86],pp128[87],pp128[88],pp128[89],pp128[90],pp128[91],pp128[92],pp128[93],pp128[94],pp128[95],pp128[96],pp128[97],pp128[98],pp128[99],pp99[129],pp98[131],pp97[133],pp96[135],pp95[137],pp94[139],pp93[141],pp92[143],pp91[145],pp90[147],pp89[149],pp88[151],pp87[153],pp86[155],pp85[157],pp84[159],pp83[161],pp82[163],pp81[165],pp80[167],pp79[169],pp78[171],pp77[173],pp76[175],pp75[177],pp74[179],pp73[181],pp72[183],pp71[185],pp70[187],pp69[189],pp68[191],pp67[193],pp66[195],pp65[197],pp64[199],pp63[201],pp62[203],pp62[204],pp62[205],pp62[206],pp62[207],pp62[208],pp62[209],pp62[210],pp62[211],pp62[212],pp62[213],pp62[214],pp62[215],pp62[216],pp62[217],pp62[218],pp62[219],pp62[220],pp62[221],pp62[222],pp62[223],pp62[224],pp62[225],pp62[226],pp62[227],pp62[228],pp62[229],pp62[230],pp62[231],pp62[232],pp62[233],pp62[234],pp62[235],pp62[236],pp62[237],pp62[238],pp62[239],pp62[240],pp62[241],pp62[242],pp62[243],pp62[244],pp62[245],pp62[246],pp62[247],pp62[248],pp62[249],pp62[250],pp62[251],pp62[252],pp62[253],pp62[254],pp62[255],pp218[100],pp218[101],pp218[102],pp218[103],pp218[104],pp218[105],pp218[106]};
    assign in60_2 = {pp141[46],pp140[48],pp139[50],pp138[52],pp137[54],pp136[56],pp135[58],pp134[60],pp133[62],pp132[64],pp131[66],pp130[68],pp129[70],pp129[71],pp129[72],pp129[73],pp129[74],pp129[75],pp129[76],pp129[77],pp129[78],pp129[79],pp129[80],pp129[81],pp129[82],pp129[83],pp129[84],pp129[85],pp129[86],pp129[87],pp129[88],pp129[89],pp129[90],pp129[91],pp129[92],pp129[93],pp129[94],pp129[95],pp129[96],pp129[97],pp129[98],pp129[99],pp99[130],pp98[132],pp97[134],pp96[136],pp95[138],pp94[140],pp93[142],pp92[144],pp91[146],pp90[148],pp89[150],pp88[152],pp87[154],pp86[156],pp85[158],pp84[160],pp83[162],pp82[164],pp81[166],pp80[168],pp79[170],pp78[172],pp77[174],pp76[176],pp75[178],pp74[180],pp73[182],pp72[184],pp71[186],pp70[188],pp69[190],pp68[192],pp67[194],pp66[196],pp65[198],pp64[200],pp63[202],pp63[203],pp63[204],pp63[205],pp63[206],pp63[207],pp63[208],pp63[209],pp63[210],pp63[211],pp63[212],pp63[213],pp63[214],pp63[215],pp63[216],pp63[217],pp63[218],pp63[219],pp63[220],pp63[221],pp63[222],pp63[223],pp63[224],pp63[225],pp63[226],pp63[227],pp63[228],pp63[229],pp63[230],pp63[231],pp63[232],pp63[233],pp63[234],pp63[235],pp63[236],pp63[237],pp63[238],pp63[239],pp63[240],pp63[241],pp63[242],pp63[243],pp63[244],pp63[245],pp63[246],pp63[247],pp63[248],pp63[249],pp63[250],pp63[251],pp63[252],pp63[253],pp63[254],pp63[255],pp219[100],pp219[101],pp219[102],pp219[103],pp219[104],pp219[105]};
    CLA_138 KS_60(s60, c60, in60_1, in60_2);
    wire[135:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp141[47],pp140[49],pp139[51],pp138[53],pp137[55],pp136[57],pp135[59],pp134[61],pp133[63],pp132[65],pp131[67],pp130[69],pp130[70],pp130[71],pp130[72],pp130[73],pp130[74],pp130[75],pp130[76],pp130[77],pp130[78],pp130[79],pp130[80],pp130[81],pp130[82],pp130[83],pp130[84],pp130[85],pp130[86],pp130[87],pp130[88],pp130[89],pp130[90],pp130[91],pp130[92],pp130[93],pp130[94],pp130[95],pp130[96],pp130[97],pp130[98],pp130[99],pp99[131],pp98[133],pp97[135],pp96[137],pp95[139],pp94[141],pp93[143],pp92[145],pp91[147],pp90[149],pp89[151],pp88[153],pp87[155],pp86[157],pp85[159],pp84[161],pp83[163],pp82[165],pp81[167],pp80[169],pp79[171],pp78[173],pp77[175],pp76[177],pp75[179],pp74[181],pp73[183],pp72[185],pp71[187],pp70[189],pp69[191],pp68[193],pp67[195],pp66[197],pp65[199],pp64[201],pp64[202],pp64[203],pp64[204],pp64[205],pp64[206],pp64[207],pp64[208],pp64[209],pp64[210],pp64[211],pp64[212],pp64[213],pp64[214],pp64[215],pp64[216],pp64[217],pp64[218],pp64[219],pp64[220],pp64[221],pp64[222],pp64[223],pp64[224],pp64[225],pp64[226],pp64[227],pp64[228],pp64[229],pp64[230],pp64[231],pp64[232],pp64[233],pp64[234],pp64[235],pp64[236],pp64[237],pp64[238],pp64[239],pp64[240],pp64[241],pp64[242],pp64[243],pp64[244],pp64[245],pp64[246],pp64[247],pp64[248],pp64[249],pp64[250],pp64[251],pp64[252],pp64[253],pp64[254],pp64[255],pp220[100],pp220[101],pp220[102],pp220[103]};
    assign in61_2 = {pp142[46],pp141[48],pp140[50],pp139[52],pp138[54],pp137[56],pp136[58],pp135[60],pp134[62],pp133[64],pp132[66],pp131[68],pp131[69],pp131[70],pp131[71],pp131[72],pp131[73],pp131[74],pp131[75],pp131[76],pp131[77],pp131[78],pp131[79],pp131[80],pp131[81],pp131[82],pp131[83],pp131[84],pp131[85],pp131[86],pp131[87],pp131[88],pp131[89],pp131[90],pp131[91],pp131[92],pp131[93],pp131[94],pp131[95],pp131[96],pp131[97],pp131[98],pp131[99],pp99[132],pp98[134],pp97[136],pp96[138],pp95[140],pp94[142],pp93[144],pp92[146],pp91[148],pp90[150],pp89[152],pp88[154],pp87[156],pp86[158],pp85[160],pp84[162],pp83[164],pp82[166],pp81[168],pp80[170],pp79[172],pp78[174],pp77[176],pp76[178],pp75[180],pp74[182],pp73[184],pp72[186],pp71[188],pp70[190],pp69[192],pp68[194],pp67[196],pp66[198],pp65[200],pp65[201],pp65[202],pp65[203],pp65[204],pp65[205],pp65[206],pp65[207],pp65[208],pp65[209],pp65[210],pp65[211],pp65[212],pp65[213],pp65[214],pp65[215],pp65[216],pp65[217],pp65[218],pp65[219],pp65[220],pp65[221],pp65[222],pp65[223],pp65[224],pp65[225],pp65[226],pp65[227],pp65[228],pp65[229],pp65[230],pp65[231],pp65[232],pp65[233],pp65[234],pp65[235],pp65[236],pp65[237],pp65[238],pp65[239],pp65[240],pp65[241],pp65[242],pp65[243],pp65[244],pp65[245],pp65[246],pp65[247],pp65[248],pp65[249],pp65[250],pp65[251],pp65[252],pp65[253],pp65[254],pp65[255],pp221[100],pp221[101],pp221[102]};
    CLA_136 KS_61(s61, c61, in61_1, in61_2);
    wire[133:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp142[47],pp141[49],pp140[51],pp139[53],pp138[55],pp137[57],pp136[59],pp135[61],pp134[63],pp133[65],pp132[67],pp132[68],pp132[69],pp132[70],pp132[71],pp132[72],pp132[73],pp132[74],pp132[75],pp132[76],pp132[77],pp132[78],pp132[79],pp132[80],pp132[81],pp132[82],pp132[83],pp132[84],pp132[85],pp132[86],pp132[87],pp132[88],pp132[89],pp132[90],pp132[91],pp132[92],pp132[93],pp132[94],pp132[95],pp132[96],pp132[97],pp132[98],pp132[99],pp99[133],pp98[135],pp97[137],pp96[139],pp95[141],pp94[143],pp93[145],pp92[147],pp91[149],pp90[151],pp89[153],pp88[155],pp87[157],pp86[159],pp85[161],pp84[163],pp83[165],pp82[167],pp81[169],pp80[171],pp79[173],pp78[175],pp77[177],pp76[179],pp75[181],pp74[183],pp73[185],pp72[187],pp71[189],pp70[191],pp69[193],pp68[195],pp67[197],pp66[199],pp66[200],pp66[201],pp66[202],pp66[203],pp66[204],pp66[205],pp66[206],pp66[207],pp66[208],pp66[209],pp66[210],pp66[211],pp66[212],pp66[213],pp66[214],pp66[215],pp66[216],pp66[217],pp66[218],pp66[219],pp66[220],pp66[221],pp66[222],pp66[223],pp66[224],pp66[225],pp66[226],pp66[227],pp66[228],pp66[229],pp66[230],pp66[231],pp66[232],pp66[233],pp66[234],pp66[235],pp66[236],pp66[237],pp66[238],pp66[239],pp66[240],pp66[241],pp66[242],pp66[243],pp66[244],pp66[245],pp66[246],pp66[247],pp66[248],pp66[249],pp66[250],pp66[251],pp66[252],pp66[253],pp66[254],pp66[255],pp222[100]};
    assign in62_2 = {pp143[46],pp142[48],pp141[50],pp140[52],pp139[54],pp138[56],pp137[58],pp136[60],pp135[62],pp134[64],pp133[66],pp133[67],pp133[68],pp133[69],pp133[70],pp133[71],pp133[72],pp133[73],pp133[74],pp133[75],pp133[76],pp133[77],pp133[78],pp133[79],pp133[80],pp133[81],pp133[82],pp133[83],pp133[84],pp133[85],pp133[86],pp133[87],pp133[88],pp133[89],pp133[90],pp133[91],pp133[92],pp133[93],pp133[94],pp133[95],pp133[96],pp133[97],pp133[98],pp133[99],pp99[134],pp98[136],pp97[138],pp96[140],pp95[142],pp94[144],pp93[146],pp92[148],pp91[150],pp90[152],pp89[154],pp88[156],pp87[158],pp86[160],pp85[162],pp84[164],pp83[166],pp82[168],pp81[170],pp80[172],pp79[174],pp78[176],pp77[178],pp76[180],pp75[182],pp74[184],pp73[186],pp72[188],pp71[190],pp70[192],pp69[194],pp68[196],pp67[198],pp67[199],pp67[200],pp67[201],pp67[202],pp67[203],pp67[204],pp67[205],pp67[206],pp67[207],pp67[208],pp67[209],pp67[210],pp67[211],pp67[212],pp67[213],pp67[214],pp67[215],pp67[216],pp67[217],pp67[218],pp67[219],pp67[220],pp67[221],pp67[222],pp67[223],pp67[224],pp67[225],pp67[226],pp67[227],pp67[228],pp67[229],pp67[230],pp67[231],pp67[232],pp67[233],pp67[234],pp67[235],pp67[236],pp67[237],pp67[238],pp67[239],pp67[240],pp67[241],pp67[242],pp67[243],pp67[244],pp67[245],pp67[246],pp67[247],pp67[248],pp67[249],pp67[250],pp67[251],pp67[252],pp67[253],pp67[254],pp67[255]};
    CLA_134 KS_62(s62, c62, in62_1, in62_2);
    wire[131:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp143[47],pp142[49],pp141[51],pp140[53],pp139[55],pp138[57],pp137[59],pp136[61],pp135[63],pp134[65],pp134[66],pp134[67],pp134[68],pp134[69],pp134[70],pp134[71],pp134[72],pp134[73],pp134[74],pp134[75],pp134[76],pp134[77],pp134[78],pp134[79],pp134[80],pp134[81],pp134[82],pp134[83],pp134[84],pp134[85],pp134[86],pp134[87],pp134[88],pp134[89],pp134[90],pp134[91],pp134[92],pp134[93],pp134[94],pp134[95],pp134[96],pp134[97],pp134[98],pp134[99],pp99[135],pp98[137],pp97[139],pp96[141],pp95[143],pp94[145],pp93[147],pp92[149],pp91[151],pp90[153],pp89[155],pp88[157],pp87[159],pp86[161],pp85[163],pp84[165],pp83[167],pp82[169],pp81[171],pp80[173],pp79[175],pp78[177],pp77[179],pp76[181],pp75[183],pp74[185],pp73[187],pp72[189],pp71[191],pp70[193],pp69[195],pp68[197],pp68[198],pp68[199],pp68[200],pp68[201],pp68[202],pp68[203],pp68[204],pp68[205],pp68[206],pp68[207],pp68[208],pp68[209],pp68[210],pp68[211],pp68[212],pp68[213],pp68[214],pp68[215],pp68[216],pp68[217],pp68[218],pp68[219],pp68[220],pp68[221],pp68[222],pp68[223],pp68[224],pp68[225],pp68[226],pp68[227],pp68[228],pp68[229],pp68[230],pp68[231],pp68[232],pp68[233],pp68[234],pp68[235],pp68[236],pp68[237],pp68[238],pp68[239],pp68[240],pp68[241],pp68[242],pp68[243],pp68[244],pp68[245],pp68[246],pp68[247],pp68[248],pp68[249],pp68[250],pp68[251],pp68[252],pp68[253]};
    assign in63_2 = {pp144[46],pp143[48],pp142[50],pp141[52],pp140[54],pp139[56],pp138[58],pp137[60],pp136[62],pp135[64],pp135[65],pp135[66],pp135[67],pp135[68],pp135[69],pp135[70],pp135[71],pp135[72],pp135[73],pp135[74],pp135[75],pp135[76],pp135[77],pp135[78],pp135[79],pp135[80],pp135[81],pp135[82],pp135[83],pp135[84],pp135[85],pp135[86],pp135[87],pp135[88],pp135[89],pp135[90],pp135[91],pp135[92],pp135[93],pp135[94],pp135[95],pp135[96],pp135[97],pp135[98],pp135[99],pp99[136],pp98[138],pp97[140],pp96[142],pp95[144],pp94[146],pp93[148],pp92[150],pp91[152],pp90[154],pp89[156],pp88[158],pp87[160],pp86[162],pp85[164],pp84[166],pp83[168],pp82[170],pp81[172],pp80[174],pp79[176],pp78[178],pp77[180],pp76[182],pp75[184],pp74[186],pp73[188],pp72[190],pp71[192],pp70[194],pp69[196],pp69[197],pp69[198],pp69[199],pp69[200],pp69[201],pp69[202],pp69[203],pp69[204],pp69[205],pp69[206],pp69[207],pp69[208],pp69[209],pp69[210],pp69[211],pp69[212],pp69[213],pp69[214],pp69[215],pp69[216],pp69[217],pp69[218],pp69[219],pp69[220],pp69[221],pp69[222],pp69[223],pp69[224],pp69[225],pp69[226],pp69[227],pp69[228],pp69[229],pp69[230],pp69[231],pp69[232],pp69[233],pp69[234],pp69[235],pp69[236],pp69[237],pp69[238],pp69[239],pp69[240],pp69[241],pp69[242],pp69[243],pp69[244],pp69[245],pp69[246],pp69[247],pp69[248],pp69[249],pp69[250],pp69[251],pp69[252]};
    CLA_132 KS_63(s63, c63, in63_1, in63_2);
    wire[129:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp144[47],pp143[49],pp142[51],pp141[53],pp140[55],pp139[57],pp138[59],pp137[61],pp136[63],pp136[64],pp136[65],pp136[66],pp136[67],pp136[68],pp136[69],pp136[70],pp136[71],pp136[72],pp136[73],pp136[74],pp136[75],pp136[76],pp136[77],pp136[78],pp136[79],pp136[80],pp136[81],pp136[82],pp136[83],pp136[84],pp136[85],pp136[86],pp136[87],pp136[88],pp136[89],pp136[90],pp136[91],pp136[92],pp136[93],pp136[94],pp136[95],pp136[96],pp136[97],pp136[98],pp136[99],pp99[137],pp98[139],pp97[141],pp96[143],pp95[145],pp94[147],pp93[149],pp92[151],pp91[153],pp90[155],pp89[157],pp88[159],pp87[161],pp86[163],pp85[165],pp84[167],pp83[169],pp82[171],pp81[173],pp80[175],pp79[177],pp78[179],pp77[181],pp76[183],pp75[185],pp74[187],pp73[189],pp72[191],pp71[193],pp70[195],pp70[196],pp70[197],pp70[198],pp70[199],pp70[200],pp70[201],pp70[202],pp70[203],pp70[204],pp70[205],pp70[206],pp70[207],pp70[208],pp70[209],pp70[210],pp70[211],pp70[212],pp70[213],pp70[214],pp70[215],pp70[216],pp70[217],pp70[218],pp70[219],pp70[220],pp70[221],pp70[222],pp70[223],pp70[224],pp70[225],pp70[226],pp70[227],pp70[228],pp70[229],pp70[230],pp70[231],pp70[232],pp70[233],pp70[234],pp70[235],pp70[236],pp70[237],pp70[238],pp70[239],pp70[240],pp70[241],pp70[242],pp70[243],pp70[244],pp70[245],pp70[246],pp70[247],pp70[248],pp70[249],pp70[250]};
    assign in64_2 = {pp145[46],pp144[48],pp143[50],pp142[52],pp141[54],pp140[56],pp139[58],pp138[60],pp137[62],pp137[63],pp137[64],pp137[65],pp137[66],pp137[67],pp137[68],pp137[69],pp137[70],pp137[71],pp137[72],pp137[73],pp137[74],pp137[75],pp137[76],pp137[77],pp137[78],pp137[79],pp137[80],pp137[81],pp137[82],pp137[83],pp137[84],pp137[85],pp137[86],pp137[87],pp137[88],pp137[89],pp137[90],pp137[91],pp137[92],pp137[93],pp137[94],pp137[95],pp137[96],pp137[97],pp137[98],pp137[99],pp99[138],pp98[140],pp97[142],pp96[144],pp95[146],pp94[148],pp93[150],pp92[152],pp91[154],pp90[156],pp89[158],pp88[160],pp87[162],pp86[164],pp85[166],pp84[168],pp83[170],pp82[172],pp81[174],pp80[176],pp79[178],pp78[180],pp77[182],pp76[184],pp75[186],pp74[188],pp73[190],pp72[192],pp71[194],pp71[195],pp71[196],pp71[197],pp71[198],pp71[199],pp71[200],pp71[201],pp71[202],pp71[203],pp71[204],pp71[205],pp71[206],pp71[207],pp71[208],pp71[209],pp71[210],pp71[211],pp71[212],pp71[213],pp71[214],pp71[215],pp71[216],pp71[217],pp71[218],pp71[219],pp71[220],pp71[221],pp71[222],pp71[223],pp71[224],pp71[225],pp71[226],pp71[227],pp71[228],pp71[229],pp71[230],pp71[231],pp71[232],pp71[233],pp71[234],pp71[235],pp71[236],pp71[237],pp71[238],pp71[239],pp71[240],pp71[241],pp71[242],pp71[243],pp71[244],pp71[245],pp71[246],pp71[247],pp71[248],pp71[249]};
    CLA_130 KS_64(s64, c64, in64_1, in64_2);
    wire[127:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp145[47],pp144[49],pp143[51],pp142[53],pp141[55],pp140[57],pp139[59],pp138[61],pp138[62],pp138[63],pp138[64],pp138[65],pp138[66],pp138[67],pp138[68],pp138[69],pp138[70],pp138[71],pp138[72],pp138[73],pp138[74],pp138[75],pp138[76],pp138[77],pp138[78],pp138[79],pp138[80],pp138[81],pp138[82],pp138[83],pp138[84],pp138[85],pp138[86],pp138[87],pp138[88],pp138[89],pp138[90],pp138[91],pp138[92],pp138[93],pp138[94],pp138[95],pp138[96],pp138[97],pp138[98],pp138[99],pp99[139],pp98[141],pp97[143],pp96[145],pp95[147],pp94[149],pp93[151],pp92[153],pp91[155],pp90[157],pp89[159],pp88[161],pp87[163],pp86[165],pp85[167],pp84[169],pp83[171],pp82[173],pp81[175],pp80[177],pp79[179],pp78[181],pp77[183],pp76[185],pp75[187],pp74[189],pp73[191],pp72[193],pp72[194],pp72[195],pp72[196],pp72[197],pp72[198],pp72[199],pp72[200],pp72[201],pp72[202],pp72[203],pp72[204],pp72[205],pp72[206],pp72[207],pp72[208],pp72[209],pp72[210],pp72[211],pp72[212],pp72[213],pp72[214],pp72[215],pp72[216],pp72[217],pp72[218],pp72[219],pp72[220],pp72[221],pp72[222],pp72[223],pp72[224],pp72[225],pp72[226],pp72[227],pp72[228],pp72[229],pp72[230],pp72[231],pp72[232],pp72[233],pp72[234],pp72[235],pp72[236],pp72[237],pp72[238],pp72[239],pp72[240],pp72[241],pp72[242],pp72[243],pp72[244],pp72[245],pp72[246],pp72[247]};
    assign in65_2 = {pp146[46],pp145[48],pp144[50],pp143[52],pp142[54],pp141[56],pp140[58],pp139[60],pp139[61],pp139[62],pp139[63],pp139[64],pp139[65],pp139[66],pp139[67],pp139[68],pp139[69],pp139[70],pp139[71],pp139[72],pp139[73],pp139[74],pp139[75],pp139[76],pp139[77],pp139[78],pp139[79],pp139[80],pp139[81],pp139[82],pp139[83],pp139[84],pp139[85],pp139[86],pp139[87],pp139[88],pp139[89],pp139[90],pp139[91],pp139[92],pp139[93],pp139[94],pp139[95],pp139[96],pp139[97],pp139[98],pp139[99],pp99[140],pp98[142],pp97[144],pp96[146],pp95[148],pp94[150],pp93[152],pp92[154],pp91[156],pp90[158],pp89[160],pp88[162],pp87[164],pp86[166],pp85[168],pp84[170],pp83[172],pp82[174],pp81[176],pp80[178],pp79[180],pp78[182],pp77[184],pp76[186],pp75[188],pp74[190],pp73[192],pp73[193],pp73[194],pp73[195],pp73[196],pp73[197],pp73[198],pp73[199],pp73[200],pp73[201],pp73[202],pp73[203],pp73[204],pp73[205],pp73[206],pp73[207],pp73[208],pp73[209],pp73[210],pp73[211],pp73[212],pp73[213],pp73[214],pp73[215],pp73[216],pp73[217],pp73[218],pp73[219],pp73[220],pp73[221],pp73[222],pp73[223],pp73[224],pp73[225],pp73[226],pp73[227],pp73[228],pp73[229],pp73[230],pp73[231],pp73[232],pp73[233],pp73[234],pp73[235],pp73[236],pp73[237],pp73[238],pp73[239],pp73[240],pp73[241],pp73[242],pp73[243],pp73[244],pp73[245],pp73[246]};
    CLA_128 KS_65(s65, c65, in65_1, in65_2);
    wire[125:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp146[47],pp145[49],pp144[51],pp143[53],pp142[55],pp141[57],pp140[59],pp140[60],pp140[61],pp140[62],pp140[63],pp140[64],pp140[65],pp140[66],pp140[67],pp140[68],pp140[69],pp140[70],pp140[71],pp140[72],pp140[73],pp140[74],pp140[75],pp140[76],pp140[77],pp140[78],pp140[79],pp140[80],pp140[81],pp140[82],pp140[83],pp140[84],pp140[85],pp140[86],pp140[87],pp140[88],pp140[89],pp140[90],pp140[91],pp140[92],pp140[93],pp140[94],pp140[95],pp140[96],pp140[97],pp140[98],pp140[99],pp99[141],pp98[143],pp97[145],pp96[147],pp95[149],pp94[151],pp93[153],pp92[155],pp91[157],pp90[159],pp89[161],pp88[163],pp87[165],pp86[167],pp85[169],pp84[171],pp83[173],pp82[175],pp81[177],pp80[179],pp79[181],pp78[183],pp77[185],pp76[187],pp75[189],pp74[191],pp74[192],pp74[193],pp74[194],pp74[195],pp74[196],pp74[197],pp74[198],pp74[199],pp74[200],pp74[201],pp74[202],pp74[203],pp74[204],pp74[205],pp74[206],pp74[207],pp74[208],pp74[209],pp74[210],pp74[211],pp74[212],pp74[213],pp74[214],pp74[215],pp74[216],pp74[217],pp74[218],pp74[219],pp74[220],pp74[221],pp74[222],pp74[223],pp74[224],pp74[225],pp74[226],pp74[227],pp74[228],pp74[229],pp74[230],pp74[231],pp74[232],pp74[233],pp74[234],pp74[235],pp74[236],pp74[237],pp74[238],pp74[239],pp74[240],pp74[241],pp74[242],pp74[243],pp74[244]};
    assign in66_2 = {pp147[46],pp146[48],pp145[50],pp144[52],pp143[54],pp142[56],pp141[58],pp141[59],pp141[60],pp141[61],pp141[62],pp141[63],pp141[64],pp141[65],pp141[66],pp141[67],pp141[68],pp141[69],pp141[70],pp141[71],pp141[72],pp141[73],pp141[74],pp141[75],pp141[76],pp141[77],pp141[78],pp141[79],pp141[80],pp141[81],pp141[82],pp141[83],pp141[84],pp141[85],pp141[86],pp141[87],pp141[88],pp141[89],pp141[90],pp141[91],pp141[92],pp141[93],pp141[94],pp141[95],pp141[96],pp141[97],pp141[98],pp141[99],pp99[142],pp98[144],pp97[146],pp96[148],pp95[150],pp94[152],pp93[154],pp92[156],pp91[158],pp90[160],pp89[162],pp88[164],pp87[166],pp86[168],pp85[170],pp84[172],pp83[174],pp82[176],pp81[178],pp80[180],pp79[182],pp78[184],pp77[186],pp76[188],pp75[190],pp75[191],pp75[192],pp75[193],pp75[194],pp75[195],pp75[196],pp75[197],pp75[198],pp75[199],pp75[200],pp75[201],pp75[202],pp75[203],pp75[204],pp75[205],pp75[206],pp75[207],pp75[208],pp75[209],pp75[210],pp75[211],pp75[212],pp75[213],pp75[214],pp75[215],pp75[216],pp75[217],pp75[218],pp75[219],pp75[220],pp75[221],pp75[222],pp75[223],pp75[224],pp75[225],pp75[226],pp75[227],pp75[228],pp75[229],pp75[230],pp75[231],pp75[232],pp75[233],pp75[234],pp75[235],pp75[236],pp75[237],pp75[238],pp75[239],pp75[240],pp75[241],pp75[242],pp75[243]};
    CLA_126 KS_66(s66, c66, in66_1, in66_2);
    wire[123:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp147[47],pp146[49],pp145[51],pp144[53],pp143[55],pp142[57],pp142[58],pp142[59],pp142[60],pp142[61],pp142[62],pp142[63],pp142[64],pp142[65],pp142[66],pp142[67],pp142[68],pp142[69],pp142[70],pp142[71],pp142[72],pp142[73],pp142[74],pp142[75],pp142[76],pp142[77],pp142[78],pp142[79],pp142[80],pp142[81],pp142[82],pp142[83],pp142[84],pp142[85],pp142[86],pp142[87],pp142[88],pp142[89],pp142[90],pp142[91],pp142[92],pp142[93],pp142[94],pp142[95],pp142[96],pp142[97],pp142[98],pp142[99],pp99[143],pp98[145],pp97[147],pp96[149],pp95[151],pp94[153],pp93[155],pp92[157],pp91[159],pp90[161],pp89[163],pp88[165],pp87[167],pp86[169],pp85[171],pp84[173],pp83[175],pp82[177],pp81[179],pp80[181],pp79[183],pp78[185],pp77[187],pp76[189],pp76[190],pp76[191],pp76[192],pp76[193],pp76[194],pp76[195],pp76[196],pp76[197],pp76[198],pp76[199],pp76[200],pp76[201],pp76[202],pp76[203],pp76[204],pp76[205],pp76[206],pp76[207],pp76[208],pp76[209],pp76[210],pp76[211],pp76[212],pp76[213],pp76[214],pp76[215],pp76[216],pp76[217],pp76[218],pp76[219],pp76[220],pp76[221],pp76[222],pp76[223],pp76[224],pp76[225],pp76[226],pp76[227],pp76[228],pp76[229],pp76[230],pp76[231],pp76[232],pp76[233],pp76[234],pp76[235],pp76[236],pp76[237],pp76[238],pp76[239],pp76[240],pp76[241]};
    assign in67_2 = {pp148[46],pp147[48],pp146[50],pp145[52],pp144[54],pp143[56],pp143[57],pp143[58],pp143[59],pp143[60],pp143[61],pp143[62],pp143[63],pp143[64],pp143[65],pp143[66],pp143[67],pp143[68],pp143[69],pp143[70],pp143[71],pp143[72],pp143[73],pp143[74],pp143[75],pp143[76],pp143[77],pp143[78],pp143[79],pp143[80],pp143[81],pp143[82],pp143[83],pp143[84],pp143[85],pp143[86],pp143[87],pp143[88],pp143[89],pp143[90],pp143[91],pp143[92],pp143[93],pp143[94],pp143[95],pp143[96],pp143[97],pp143[98],pp143[99],pp99[144],pp98[146],pp97[148],pp96[150],pp95[152],pp94[154],pp93[156],pp92[158],pp91[160],pp90[162],pp89[164],pp88[166],pp87[168],pp86[170],pp85[172],pp84[174],pp83[176],pp82[178],pp81[180],pp80[182],pp79[184],pp78[186],pp77[188],pp77[189],pp77[190],pp77[191],pp77[192],pp77[193],pp77[194],pp77[195],pp77[196],pp77[197],pp77[198],pp77[199],pp77[200],pp77[201],pp77[202],pp77[203],pp77[204],pp77[205],pp77[206],pp77[207],pp77[208],pp77[209],pp77[210],pp77[211],pp77[212],pp77[213],pp77[214],pp77[215],pp77[216],pp77[217],pp77[218],pp77[219],pp77[220],pp77[221],pp77[222],pp77[223],pp77[224],pp77[225],pp77[226],pp77[227],pp77[228],pp77[229],pp77[230],pp77[231],pp77[232],pp77[233],pp77[234],pp77[235],pp77[236],pp77[237],pp77[238],pp77[239],pp77[240]};
    CLA_124 KS_67(s67, c67, in67_1, in67_2);
    wire[121:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp148[47],pp147[49],pp146[51],pp145[53],pp144[55],pp144[56],pp144[57],pp144[58],pp144[59],pp144[60],pp144[61],pp144[62],pp144[63],pp144[64],pp144[65],pp144[66],pp144[67],pp144[68],pp144[69],pp144[70],pp144[71],pp144[72],pp144[73],pp144[74],pp144[75],pp144[76],pp144[77],pp144[78],pp144[79],pp144[80],pp144[81],pp144[82],pp144[83],pp144[84],pp144[85],pp144[86],pp144[87],pp144[88],pp144[89],pp144[90],pp144[91],pp144[92],pp144[93],pp144[94],pp144[95],pp144[96],pp144[97],pp144[98],pp144[99],pp99[145],pp98[147],pp97[149],pp96[151],pp95[153],pp94[155],pp93[157],pp92[159],pp91[161],pp90[163],pp89[165],pp88[167],pp87[169],pp86[171],pp85[173],pp84[175],pp83[177],pp82[179],pp81[181],pp80[183],pp79[185],pp78[187],pp78[188],pp78[189],pp78[190],pp78[191],pp78[192],pp78[193],pp78[194],pp78[195],pp78[196],pp78[197],pp78[198],pp78[199],pp78[200],pp78[201],pp78[202],pp78[203],pp78[204],pp78[205],pp78[206],pp78[207],pp78[208],pp78[209],pp78[210],pp78[211],pp78[212],pp78[213],pp78[214],pp78[215],pp78[216],pp78[217],pp78[218],pp78[219],pp78[220],pp78[221],pp78[222],pp78[223],pp78[224],pp78[225],pp78[226],pp78[227],pp78[228],pp78[229],pp78[230],pp78[231],pp78[232],pp78[233],pp78[234],pp78[235],pp78[236],pp78[237],pp78[238]};
    assign in68_2 = {pp149[46],pp148[48],pp147[50],pp146[52],pp145[54],pp145[55],pp145[56],pp145[57],pp145[58],pp145[59],pp145[60],pp145[61],pp145[62],pp145[63],pp145[64],pp145[65],pp145[66],pp145[67],pp145[68],pp145[69],pp145[70],pp145[71],pp145[72],pp145[73],pp145[74],pp145[75],pp145[76],pp145[77],pp145[78],pp145[79],pp145[80],pp145[81],pp145[82],pp145[83],pp145[84],pp145[85],pp145[86],pp145[87],pp145[88],pp145[89],pp145[90],pp145[91],pp145[92],pp145[93],pp145[94],pp145[95],pp145[96],pp145[97],pp145[98],pp145[99],pp99[146],pp98[148],pp97[150],pp96[152],pp95[154],pp94[156],pp93[158],pp92[160],pp91[162],pp90[164],pp89[166],pp88[168],pp87[170],pp86[172],pp85[174],pp84[176],pp83[178],pp82[180],pp81[182],pp80[184],pp79[186],pp79[187],pp79[188],pp79[189],pp79[190],pp79[191],pp79[192],pp79[193],pp79[194],pp79[195],pp79[196],pp79[197],pp79[198],pp79[199],pp79[200],pp79[201],pp79[202],pp79[203],pp79[204],pp79[205],pp79[206],pp79[207],pp79[208],pp79[209],pp79[210],pp79[211],pp79[212],pp79[213],pp79[214],pp79[215],pp79[216],pp79[217],pp79[218],pp79[219],pp79[220],pp79[221],pp79[222],pp79[223],pp79[224],pp79[225],pp79[226],pp79[227],pp79[228],pp79[229],pp79[230],pp79[231],pp79[232],pp79[233],pp79[234],pp79[235],pp79[236],pp79[237]};
    CLA_122 KS_68(s68, c68, in68_1, in68_2);
    wire[119:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp149[47],pp148[49],pp147[51],pp146[53],pp146[54],pp146[55],pp146[56],pp146[57],pp146[58],pp146[59],pp146[60],pp146[61],pp146[62],pp146[63],pp146[64],pp146[65],pp146[66],pp146[67],pp146[68],pp146[69],pp146[70],pp146[71],pp146[72],pp146[73],pp146[74],pp146[75],pp146[76],pp146[77],pp146[78],pp146[79],pp146[80],pp146[81],pp146[82],pp146[83],pp146[84],pp146[85],pp146[86],pp146[87],pp146[88],pp146[89],pp146[90],pp146[91],pp146[92],pp146[93],pp146[94],pp146[95],pp146[96],pp146[97],pp146[98],pp146[99],pp99[147],pp98[149],pp97[151],pp96[153],pp95[155],pp94[157],pp93[159],pp92[161],pp91[163],pp90[165],pp89[167],pp88[169],pp87[171],pp86[173],pp85[175],pp84[177],pp83[179],pp82[181],pp81[183],pp80[185],pp80[186],pp80[187],pp80[188],pp80[189],pp80[190],pp80[191],pp80[192],pp80[193],pp80[194],pp80[195],pp80[196],pp80[197],pp80[198],pp80[199],pp80[200],pp80[201],pp80[202],pp80[203],pp80[204],pp80[205],pp80[206],pp80[207],pp80[208],pp80[209],pp80[210],pp80[211],pp80[212],pp80[213],pp80[214],pp80[215],pp80[216],pp80[217],pp80[218],pp80[219],pp80[220],pp80[221],pp80[222],pp80[223],pp80[224],pp80[225],pp80[226],pp80[227],pp80[228],pp80[229],pp80[230],pp80[231],pp80[232],pp80[233],pp80[234],pp80[235]};
    assign in69_2 = {pp150[46],pp149[48],pp148[50],pp147[52],pp147[53],pp147[54],pp147[55],pp147[56],pp147[57],pp147[58],pp147[59],pp147[60],pp147[61],pp147[62],pp147[63],pp147[64],pp147[65],pp147[66],pp147[67],pp147[68],pp147[69],pp147[70],pp147[71],pp147[72],pp147[73],pp147[74],pp147[75],pp147[76],pp147[77],pp147[78],pp147[79],pp147[80],pp147[81],pp147[82],pp147[83],pp147[84],pp147[85],pp147[86],pp147[87],pp147[88],pp147[89],pp147[90],pp147[91],pp147[92],pp147[93],pp147[94],pp147[95],pp147[96],pp147[97],pp147[98],pp147[99],pp99[148],pp98[150],pp97[152],pp96[154],pp95[156],pp94[158],pp93[160],pp92[162],pp91[164],pp90[166],pp89[168],pp88[170],pp87[172],pp86[174],pp85[176],pp84[178],pp83[180],pp82[182],pp81[184],pp81[185],pp81[186],pp81[187],pp81[188],pp81[189],pp81[190],pp81[191],pp81[192],pp81[193],pp81[194],pp81[195],pp81[196],pp81[197],pp81[198],pp81[199],pp81[200],pp81[201],pp81[202],pp81[203],pp81[204],pp81[205],pp81[206],pp81[207],pp81[208],pp81[209],pp81[210],pp81[211],pp81[212],pp81[213],pp81[214],pp81[215],pp81[216],pp81[217],pp81[218],pp81[219],pp81[220],pp81[221],pp81[222],pp81[223],pp81[224],pp81[225],pp81[226],pp81[227],pp81[228],pp81[229],pp81[230],pp81[231],pp81[232],pp81[233],pp81[234]};
    CLA_120 KS_69(s69, c69, in69_1, in69_2);
    wire[117:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp150[47],pp149[49],pp148[51],pp148[52],pp148[53],pp148[54],pp148[55],pp148[56],pp148[57],pp148[58],pp148[59],pp148[60],pp148[61],pp148[62],pp148[63],pp148[64],pp148[65],pp148[66],pp148[67],pp148[68],pp148[69],pp148[70],pp148[71],pp148[72],pp148[73],pp148[74],pp148[75],pp148[76],pp148[77],pp148[78],pp148[79],pp148[80],pp148[81],pp148[82],pp148[83],pp148[84],pp148[85],pp148[86],pp148[87],pp148[88],pp148[89],pp148[90],pp148[91],pp148[92],pp148[93],pp148[94],pp148[95],pp148[96],pp148[97],pp148[98],pp148[99],pp99[149],pp98[151],pp97[153],pp96[155],pp95[157],pp94[159],pp93[161],pp92[163],pp91[165],pp90[167],pp89[169],pp88[171],pp87[173],pp86[175],pp85[177],pp84[179],pp83[181],pp82[183],pp82[184],pp82[185],pp82[186],pp82[187],pp82[188],pp82[189],pp82[190],pp82[191],pp82[192],pp82[193],pp82[194],pp82[195],pp82[196],pp82[197],pp82[198],pp82[199],pp82[200],pp82[201],pp82[202],pp82[203],pp82[204],pp82[205],pp82[206],pp82[207],pp82[208],pp82[209],pp82[210],pp82[211],pp82[212],pp82[213],pp82[214],pp82[215],pp82[216],pp82[217],pp82[218],pp82[219],pp82[220],pp82[221],pp82[222],pp82[223],pp82[224],pp82[225],pp82[226],pp82[227],pp82[228],pp82[229],pp82[230],pp82[231],pp82[232]};
    assign in70_2 = {pp151[46],pp150[48],pp149[50],pp149[51],pp149[52],pp149[53],pp149[54],pp149[55],pp149[56],pp149[57],pp149[58],pp149[59],pp149[60],pp149[61],pp149[62],pp149[63],pp149[64],pp149[65],pp149[66],pp149[67],pp149[68],pp149[69],pp149[70],pp149[71],pp149[72],pp149[73],pp149[74],pp149[75],pp149[76],pp149[77],pp149[78],pp149[79],pp149[80],pp149[81],pp149[82],pp149[83],pp149[84],pp149[85],pp149[86],pp149[87],pp149[88],pp149[89],pp149[90],pp149[91],pp149[92],pp149[93],pp149[94],pp149[95],pp149[96],pp149[97],pp149[98],pp149[99],pp99[150],pp98[152],pp97[154],pp96[156],pp95[158],pp94[160],pp93[162],pp92[164],pp91[166],pp90[168],pp89[170],pp88[172],pp87[174],pp86[176],pp85[178],pp84[180],pp83[182],pp83[183],pp83[184],pp83[185],pp83[186],pp83[187],pp83[188],pp83[189],pp83[190],pp83[191],pp83[192],pp83[193],pp83[194],pp83[195],pp83[196],pp83[197],pp83[198],pp83[199],pp83[200],pp83[201],pp83[202],pp83[203],pp83[204],pp83[205],pp83[206],pp83[207],pp83[208],pp83[209],pp83[210],pp83[211],pp83[212],pp83[213],pp83[214],pp83[215],pp83[216],pp83[217],pp83[218],pp83[219],pp83[220],pp83[221],pp83[222],pp83[223],pp83[224],pp83[225],pp83[226],pp83[227],pp83[228],pp83[229],pp83[230],pp83[231]};
    CLA_118 KS_70(s70, c70, in70_1, in70_2);
    wire[115:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp151[47],pp150[49],pp150[50],pp150[51],pp150[52],pp150[53],pp150[54],pp150[55],pp150[56],pp150[57],pp150[58],pp150[59],pp150[60],pp150[61],pp150[62],pp150[63],pp150[64],pp150[65],pp150[66],pp150[67],pp150[68],pp150[69],pp150[70],pp150[71],pp150[72],pp150[73],pp150[74],pp150[75],pp150[76],pp150[77],pp150[78],pp150[79],pp150[80],pp150[81],pp150[82],pp150[83],pp150[84],pp150[85],pp150[86],pp150[87],pp150[88],pp150[89],pp150[90],pp150[91],pp150[92],pp150[93],pp150[94],pp150[95],pp150[96],pp150[97],pp150[98],pp150[99],pp99[151],pp98[153],pp97[155],pp96[157],pp95[159],pp94[161],pp93[163],pp92[165],pp91[167],pp90[169],pp89[171],pp88[173],pp87[175],pp86[177],pp85[179],pp84[181],pp84[182],pp84[183],pp84[184],pp84[185],pp84[186],pp84[187],pp84[188],pp84[189],pp84[190],pp84[191],pp84[192],pp84[193],pp84[194],pp84[195],pp84[196],pp84[197],pp84[198],pp84[199],pp84[200],pp84[201],pp84[202],pp84[203],pp84[204],pp84[205],pp84[206],pp84[207],pp84[208],pp84[209],pp84[210],pp84[211],pp84[212],pp84[213],pp84[214],pp84[215],pp84[216],pp84[217],pp84[218],pp84[219],pp84[220],pp84[221],pp84[222],pp84[223],pp84[224],pp84[225],pp84[226],pp84[227],pp84[228],pp84[229]};
    assign in71_2 = {pp152[46],pp151[48],pp151[49],pp151[50],pp151[51],pp151[52],pp151[53],pp151[54],pp151[55],pp151[56],pp151[57],pp151[58],pp151[59],pp151[60],pp151[61],pp151[62],pp151[63],pp151[64],pp151[65],pp151[66],pp151[67],pp151[68],pp151[69],pp151[70],pp151[71],pp151[72],pp151[73],pp151[74],pp151[75],pp151[76],pp151[77],pp151[78],pp151[79],pp151[80],pp151[81],pp151[82],pp151[83],pp151[84],pp151[85],pp151[86],pp151[87],pp151[88],pp151[89],pp151[90],pp151[91],pp151[92],pp151[93],pp151[94],pp151[95],pp151[96],pp151[97],pp151[98],pp151[99],pp99[152],pp98[154],pp97[156],pp96[158],pp95[160],pp94[162],pp93[164],pp92[166],pp91[168],pp90[170],pp89[172],pp88[174],pp87[176],pp86[178],pp85[180],pp85[181],pp85[182],pp85[183],pp85[184],pp85[185],pp85[186],pp85[187],pp85[188],pp85[189],pp85[190],pp85[191],pp85[192],pp85[193],pp85[194],pp85[195],pp85[196],pp85[197],pp85[198],pp85[199],pp85[200],pp85[201],pp85[202],pp85[203],pp85[204],pp85[205],pp85[206],pp85[207],pp85[208],pp85[209],pp85[210],pp85[211],pp85[212],pp85[213],pp85[214],pp85[215],pp85[216],pp85[217],pp85[218],pp85[219],pp85[220],pp85[221],pp85[222],pp85[223],pp85[224],pp85[225],pp85[226],pp85[227],pp85[228]};
    CLA_116 KS_71(s71, c71, in71_1, in71_2);
    wire[113:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp152[47],pp152[48],pp152[49],pp152[50],pp152[51],pp152[52],pp152[53],pp152[54],pp152[55],pp152[56],pp152[57],pp152[58],pp152[59],pp152[60],pp152[61],pp152[62],pp152[63],pp152[64],pp152[65],pp152[66],pp152[67],pp152[68],pp152[69],pp152[70],pp152[71],pp152[72],pp152[73],pp152[74],pp152[75],pp152[76],pp152[77],pp152[78],pp152[79],pp152[80],pp152[81],pp152[82],pp152[83],pp152[84],pp152[85],pp152[86],pp152[87],pp152[88],pp152[89],pp152[90],pp152[91],pp152[92],pp152[93],pp152[94],pp152[95],pp152[96],pp152[97],pp152[98],pp152[99],pp99[153],pp98[155],pp97[157],pp96[159],pp95[161],pp94[163],pp93[165],pp92[167],pp91[169],pp90[171],pp89[173],pp88[175],pp87[177],pp86[179],pp86[180],pp86[181],pp86[182],pp86[183],pp86[184],pp86[185],pp86[186],pp86[187],pp86[188],pp86[189],pp86[190],pp86[191],pp86[192],pp86[193],pp86[194],pp86[195],pp86[196],pp86[197],pp86[198],pp86[199],pp86[200],pp86[201],pp86[202],pp86[203],pp86[204],pp86[205],pp86[206],pp86[207],pp86[208],pp86[209],pp86[210],pp86[211],pp86[212],pp86[213],pp86[214],pp86[215],pp86[216],pp86[217],pp86[218],pp86[219],pp86[220],pp86[221],pp86[222],pp86[223],pp86[224],pp86[225],pp86[226]};
    assign in72_2 = {pp153[46],pp153[47],pp153[48],pp153[49],pp153[50],pp153[51],pp153[52],pp153[53],pp153[54],pp153[55],pp153[56],pp153[57],pp153[58],pp153[59],pp153[60],pp153[61],pp153[62],pp153[63],pp153[64],pp153[65],pp153[66],pp153[67],pp153[68],pp153[69],pp153[70],pp153[71],pp153[72],pp153[73],pp153[74],pp153[75],pp153[76],pp153[77],pp153[78],pp153[79],pp153[80],pp153[81],pp153[82],pp153[83],pp153[84],pp153[85],pp153[86],pp153[87],pp153[88],pp153[89],pp153[90],pp153[91],pp153[92],pp153[93],pp153[94],pp153[95],pp153[96],pp153[97],pp153[98],pp153[99],pp99[154],pp98[156],pp97[158],pp96[160],pp95[162],pp94[164],pp93[166],pp92[168],pp91[170],pp90[172],pp89[174],pp88[176],pp87[178],pp87[179],pp87[180],pp87[181],pp87[182],pp87[183],pp87[184],pp87[185],pp87[186],pp87[187],pp87[188],pp87[189],pp87[190],pp87[191],pp87[192],pp87[193],pp87[194],pp87[195],pp87[196],pp87[197],pp87[198],pp87[199],pp87[200],pp87[201],pp87[202],pp87[203],pp87[204],pp87[205],pp87[206],pp87[207],pp87[208],pp87[209],pp87[210],pp87[211],pp87[212],pp87[213],pp87[214],pp87[215],pp87[216],pp87[217],pp87[218],pp87[219],pp87[220],pp87[221],pp87[222],pp87[223],pp87[224],pp87[225]};
    CLA_114 KS_72(s72, c72, in72_1, in72_2);
    wire[111:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp154[46],pp154[47],pp154[48],pp154[49],pp154[50],pp154[51],pp154[52],pp154[53],pp154[54],pp154[55],pp154[56],pp154[57],pp154[58],pp154[59],pp154[60],pp154[61],pp154[62],pp154[63],pp154[64],pp154[65],pp154[66],pp154[67],pp154[68],pp154[69],pp154[70],pp154[71],pp154[72],pp154[73],pp154[74],pp154[75],pp154[76],pp154[77],pp154[78],pp154[79],pp154[80],pp154[81],pp154[82],pp154[83],pp154[84],pp154[85],pp154[86],pp154[87],pp154[88],pp154[89],pp154[90],pp154[91],pp154[92],pp154[93],pp154[94],pp154[95],pp154[96],pp154[97],pp154[98],pp154[99],pp99[155],pp98[157],pp97[159],pp96[161],pp95[163],pp94[165],pp93[167],pp92[169],pp91[171],pp90[173],pp89[175],pp88[177],pp88[178],pp88[179],pp88[180],pp88[181],pp88[182],pp88[183],pp88[184],pp88[185],pp88[186],pp88[187],pp88[188],pp88[189],pp88[190],pp88[191],pp88[192],pp88[193],pp88[194],pp88[195],pp88[196],pp88[197],pp88[198],pp88[199],pp88[200],pp88[201],pp88[202],pp88[203],pp88[204],pp88[205],pp88[206],pp88[207],pp88[208],pp88[209],pp88[210],pp88[211],pp88[212],pp88[213],pp88[214],pp88[215],pp88[216],pp88[217],pp88[218],pp88[219],pp88[220],pp88[221],pp88[222],pp88[223]};
    assign in73_2 = {pp155[45],pp155[46],pp155[47],pp155[48],pp155[49],pp155[50],pp155[51],pp155[52],pp155[53],pp155[54],pp155[55],pp155[56],pp155[57],pp155[58],pp155[59],pp155[60],pp155[61],pp155[62],pp155[63],pp155[64],pp155[65],pp155[66],pp155[67],pp155[68],pp155[69],pp155[70],pp155[71],pp155[72],pp155[73],pp155[74],pp155[75],pp155[76],pp155[77],pp155[78],pp155[79],pp155[80],pp155[81],pp155[82],pp155[83],pp155[84],pp155[85],pp155[86],pp155[87],pp155[88],pp155[89],pp155[90],pp155[91],pp155[92],pp155[93],pp155[94],pp155[95],pp155[96],pp155[97],pp155[98],pp155[99],pp99[156],pp98[158],pp97[160],pp96[162],pp95[164],pp94[166],pp93[168],pp92[170],pp91[172],pp90[174],pp89[176],pp89[177],pp89[178],pp89[179],pp89[180],pp89[181],pp89[182],pp89[183],pp89[184],pp89[185],pp89[186],pp89[187],pp89[188],pp89[189],pp89[190],pp89[191],pp89[192],pp89[193],pp89[194],pp89[195],pp89[196],pp89[197],pp89[198],pp89[199],pp89[200],pp89[201],pp89[202],pp89[203],pp89[204],pp89[205],pp89[206],pp89[207],pp89[208],pp89[209],pp89[210],pp89[211],pp89[212],pp89[213],pp89[214],pp89[215],pp89[216],pp89[217],pp89[218],pp89[219],pp89[220],pp89[221],pp89[222]};
    CLA_112 KS_73(s73, c73, in73_1, in73_2);
    wire[109:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp156[45],pp156[46],pp156[47],pp156[48],pp156[49],pp156[50],pp156[51],pp156[52],pp156[53],pp156[54],pp156[55],pp156[56],pp156[57],pp156[58],pp156[59],pp156[60],pp156[61],pp156[62],pp156[63],pp156[64],pp156[65],pp156[66],pp156[67],pp156[68],pp156[69],pp156[70],pp156[71],pp156[72],pp156[73],pp156[74],pp156[75],pp156[76],pp156[77],pp156[78],pp156[79],pp156[80],pp156[81],pp156[82],pp156[83],pp156[84],pp156[85],pp156[86],pp156[87],pp156[88],pp156[89],pp156[90],pp156[91],pp156[92],pp156[93],pp156[94],pp156[95],pp156[96],pp156[97],pp156[98],pp156[99],pp99[157],pp98[159],pp97[161],pp96[163],pp95[165],pp94[167],pp93[169],pp92[171],pp91[173],pp90[175],pp90[176],pp90[177],pp90[178],pp90[179],pp90[180],pp90[181],pp90[182],pp90[183],pp90[184],pp90[185],pp90[186],pp90[187],pp90[188],pp90[189],pp90[190],pp90[191],pp90[192],pp90[193],pp90[194],pp90[195],pp90[196],pp90[197],pp90[198],pp90[199],pp90[200],pp90[201],pp90[202],pp90[203],pp90[204],pp90[205],pp90[206],pp90[207],pp90[208],pp90[209],pp90[210],pp90[211],pp90[212],pp90[213],pp90[214],pp90[215],pp90[216],pp90[217],pp90[218],pp90[219],pp90[220]};
    assign in74_2 = {pp157[44],pp157[45],pp157[46],pp157[47],pp157[48],pp157[49],pp157[50],pp157[51],pp157[52],pp157[53],pp157[54],pp157[55],pp157[56],pp157[57],pp157[58],pp157[59],pp157[60],pp157[61],pp157[62],pp157[63],pp157[64],pp157[65],pp157[66],pp157[67],pp157[68],pp157[69],pp157[70],pp157[71],pp157[72],pp157[73],pp157[74],pp157[75],pp157[76],pp157[77],pp157[78],pp157[79],pp157[80],pp157[81],pp157[82],pp157[83],pp157[84],pp157[85],pp157[86],pp157[87],pp157[88],pp157[89],pp157[90],pp157[91],pp157[92],pp157[93],pp157[94],pp157[95],pp157[96],pp157[97],pp157[98],pp157[99],pp99[158],pp98[160],pp97[162],pp96[164],pp95[166],pp94[168],pp93[170],pp92[172],pp91[174],pp91[175],pp91[176],pp91[177],pp91[178],pp91[179],pp91[180],pp91[181],pp91[182],pp91[183],pp91[184],pp91[185],pp91[186],pp91[187],pp91[188],pp91[189],pp91[190],pp91[191],pp91[192],pp91[193],pp91[194],pp91[195],pp91[196],pp91[197],pp91[198],pp91[199],pp91[200],pp91[201],pp91[202],pp91[203],pp91[204],pp91[205],pp91[206],pp91[207],pp91[208],pp91[209],pp91[210],pp91[211],pp91[212],pp91[213],pp91[214],pp91[215],pp91[216],pp91[217],pp91[218],pp91[219]};
    CLA_110 KS_74(s74, c74, in74_1, in74_2);
    wire[107:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp158[44],pp158[45],pp158[46],pp158[47],pp158[48],pp158[49],pp158[50],pp158[51],pp158[52],pp158[53],pp158[54],pp158[55],pp158[56],pp158[57],pp158[58],pp158[59],pp158[60],pp158[61],pp158[62],pp158[63],pp158[64],pp158[65],pp158[66],pp158[67],pp158[68],pp158[69],pp158[70],pp158[71],pp158[72],pp158[73],pp158[74],pp158[75],pp158[76],pp158[77],pp158[78],pp158[79],pp158[80],pp158[81],pp158[82],pp158[83],pp158[84],pp158[85],pp158[86],pp158[87],pp158[88],pp158[89],pp158[90],pp158[91],pp158[92],pp158[93],pp158[94],pp158[95],pp158[96],pp158[97],pp158[98],pp158[99],pp99[159],pp98[161],pp97[163],pp96[165],pp95[167],pp94[169],pp93[171],pp92[173],pp92[174],pp92[175],pp92[176],pp92[177],pp92[178],pp92[179],pp92[180],pp92[181],pp92[182],pp92[183],pp92[184],pp92[185],pp92[186],pp92[187],pp92[188],pp92[189],pp92[190],pp92[191],pp92[192],pp92[193],pp92[194],pp92[195],pp92[196],pp92[197],pp92[198],pp92[199],pp92[200],pp92[201],pp92[202],pp92[203],pp92[204],pp92[205],pp92[206],pp92[207],pp92[208],pp92[209],pp92[210],pp92[211],pp92[212],pp92[213],pp92[214],pp92[215],pp92[216],pp92[217]};
    assign in75_2 = {pp159[43],pp159[44],pp159[45],pp159[46],pp159[47],pp159[48],pp159[49],pp159[50],pp159[51],pp159[52],pp159[53],pp159[54],pp159[55],pp159[56],pp159[57],pp159[58],pp159[59],pp159[60],pp159[61],pp159[62],pp159[63],pp159[64],pp159[65],pp159[66],pp159[67],pp159[68],pp159[69],pp159[70],pp159[71],pp159[72],pp159[73],pp159[74],pp159[75],pp159[76],pp159[77],pp159[78],pp159[79],pp159[80],pp159[81],pp159[82],pp159[83],pp159[84],pp159[85],pp159[86],pp159[87],pp159[88],pp159[89],pp159[90],pp159[91],pp159[92],pp159[93],pp159[94],pp159[95],pp159[96],pp159[97],pp159[98],pp159[99],pp99[160],pp98[162],pp97[164],pp96[166],pp95[168],pp94[170],pp93[172],pp93[173],pp93[174],pp93[175],pp93[176],pp93[177],pp93[178],pp93[179],pp93[180],pp93[181],pp93[182],pp93[183],pp93[184],pp93[185],pp93[186],pp93[187],pp93[188],pp93[189],pp93[190],pp93[191],pp93[192],pp93[193],pp93[194],pp93[195],pp93[196],pp93[197],pp93[198],pp93[199],pp93[200],pp93[201],pp93[202],pp93[203],pp93[204],pp93[205],pp93[206],pp93[207],pp93[208],pp93[209],pp93[210],pp93[211],pp93[212],pp93[213],pp93[214],pp93[215],pp93[216]};
    CLA_108 KS_75(s75, c75, in75_1, in75_2);
    wire[105:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp160[43],pp160[44],pp160[45],pp160[46],pp160[47],pp160[48],pp160[49],pp160[50],pp160[51],pp160[52],pp160[53],pp160[54],pp160[55],pp160[56],pp160[57],pp160[58],pp160[59],pp160[60],pp160[61],pp160[62],pp160[63],pp160[64],pp160[65],pp160[66],pp160[67],pp160[68],pp160[69],pp160[70],pp160[71],pp160[72],pp160[73],pp160[74],pp160[75],pp160[76],pp160[77],pp160[78],pp160[79],pp160[80],pp160[81],pp160[82],pp160[83],pp160[84],pp160[85],pp160[86],pp160[87],pp160[88],pp160[89],pp160[90],pp160[91],pp160[92],pp160[93],pp160[94],pp160[95],pp160[96],pp160[97],pp160[98],pp160[99],pp99[161],pp98[163],pp97[165],pp96[167],pp95[169],pp94[171],pp94[172],pp94[173],pp94[174],pp94[175],pp94[176],pp94[177],pp94[178],pp94[179],pp94[180],pp94[181],pp94[182],pp94[183],pp94[184],pp94[185],pp94[186],pp94[187],pp94[188],pp94[189],pp94[190],pp94[191],pp94[192],pp94[193],pp94[194],pp94[195],pp94[196],pp94[197],pp94[198],pp94[199],pp94[200],pp94[201],pp94[202],pp94[203],pp94[204],pp94[205],pp94[206],pp94[207],pp94[208],pp94[209],pp94[210],pp94[211],pp94[212],pp94[213],pp94[214]};
    assign in76_2 = {pp161[42],pp161[43],pp161[44],pp161[45],pp161[46],pp161[47],pp161[48],pp161[49],pp161[50],pp161[51],pp161[52],pp161[53],pp161[54],pp161[55],pp161[56],pp161[57],pp161[58],pp161[59],pp161[60],pp161[61],pp161[62],pp161[63],pp161[64],pp161[65],pp161[66],pp161[67],pp161[68],pp161[69],pp161[70],pp161[71],pp161[72],pp161[73],pp161[74],pp161[75],pp161[76],pp161[77],pp161[78],pp161[79],pp161[80],pp161[81],pp161[82],pp161[83],pp161[84],pp161[85],pp161[86],pp161[87],pp161[88],pp161[89],pp161[90],pp161[91],pp161[92],pp161[93],pp161[94],pp161[95],pp161[96],pp161[97],pp161[98],pp161[99],pp99[162],pp98[164],pp97[166],pp96[168],pp95[170],pp95[171],pp95[172],pp95[173],pp95[174],pp95[175],pp95[176],pp95[177],pp95[178],pp95[179],pp95[180],pp95[181],pp95[182],pp95[183],pp95[184],pp95[185],pp95[186],pp95[187],pp95[188],pp95[189],pp95[190],pp95[191],pp95[192],pp95[193],pp95[194],pp95[195],pp95[196],pp95[197],pp95[198],pp95[199],pp95[200],pp95[201],pp95[202],pp95[203],pp95[204],pp95[205],pp95[206],pp95[207],pp95[208],pp95[209],pp95[210],pp95[211],pp95[212],pp95[213]};
    CLA_106 KS_76(s76, c76, in76_1, in76_2);
    wire[103:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp162[42],pp162[43],pp162[44],pp162[45],pp162[46],pp162[47],pp162[48],pp162[49],pp162[50],pp162[51],pp162[52],pp162[53],pp162[54],pp162[55],pp162[56],pp162[57],pp162[58],pp162[59],pp162[60],pp162[61],pp162[62],pp162[63],pp162[64],pp162[65],pp162[66],pp162[67],pp162[68],pp162[69],pp162[70],pp162[71],pp162[72],pp162[73],pp162[74],pp162[75],pp162[76],pp162[77],pp162[78],pp162[79],pp162[80],pp162[81],pp162[82],pp162[83],pp162[84],pp162[85],pp162[86],pp162[87],pp162[88],pp162[89],pp162[90],pp162[91],pp162[92],pp162[93],pp162[94],pp162[95],pp162[96],pp162[97],pp162[98],pp162[99],pp99[163],pp98[165],pp97[167],pp96[169],pp96[170],pp96[171],pp96[172],pp96[173],pp96[174],pp96[175],pp96[176],pp96[177],pp96[178],pp96[179],pp96[180],pp96[181],pp96[182],pp96[183],pp96[184],pp96[185],pp96[186],pp96[187],pp96[188],pp96[189],pp96[190],pp96[191],pp96[192],pp96[193],pp96[194],pp96[195],pp96[196],pp96[197],pp96[198],pp96[199],pp96[200],pp96[201],pp96[202],pp96[203],pp96[204],pp96[205],pp96[206],pp96[207],pp96[208],pp96[209],pp96[210],pp96[211]};
    assign in77_2 = {pp163[41],pp163[42],pp163[43],pp163[44],pp163[45],pp163[46],pp163[47],pp163[48],pp163[49],pp163[50],pp163[51],pp163[52],pp163[53],pp163[54],pp163[55],pp163[56],pp163[57],pp163[58],pp163[59],pp163[60],pp163[61],pp163[62],pp163[63],pp163[64],pp163[65],pp163[66],pp163[67],pp163[68],pp163[69],pp163[70],pp163[71],pp163[72],pp163[73],pp163[74],pp163[75],pp163[76],pp163[77],pp163[78],pp163[79],pp163[80],pp163[81],pp163[82],pp163[83],pp163[84],pp163[85],pp163[86],pp163[87],pp163[88],pp163[89],pp163[90],pp163[91],pp163[92],pp163[93],pp163[94],pp163[95],pp163[96],pp163[97],pp163[98],pp163[99],pp99[164],pp98[166],pp97[168],pp97[169],pp97[170],pp97[171],pp97[172],pp97[173],pp97[174],pp97[175],pp97[176],pp97[177],pp97[178],pp97[179],pp97[180],pp97[181],pp97[182],pp97[183],pp97[184],pp97[185],pp97[186],pp97[187],pp97[188],pp97[189],pp97[190],pp97[191],pp97[192],pp97[193],pp97[194],pp97[195],pp97[196],pp97[197],pp97[198],pp97[199],pp97[200],pp97[201],pp97[202],pp97[203],pp97[204],pp97[205],pp97[206],pp97[207],pp97[208],pp97[209],pp97[210]};
    CLA_104 KS_77(s77, c77, in77_1, in77_2);
    wire[101:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp164[41],pp164[42],pp164[43],pp164[44],pp164[45],pp164[46],pp164[47],pp164[48],pp164[49],pp164[50],pp164[51],pp164[52],pp164[53],pp164[54],pp164[55],pp164[56],pp164[57],pp164[58],pp164[59],pp164[60],pp164[61],pp164[62],pp164[63],pp164[64],pp164[65],pp164[66],pp164[67],pp164[68],pp164[69],pp164[70],pp164[71],pp164[72],pp164[73],pp164[74],pp164[75],pp164[76],pp164[77],pp164[78],pp164[79],pp164[80],pp164[81],pp164[82],pp164[83],pp164[84],pp164[85],pp164[86],pp164[87],pp164[88],pp164[89],pp164[90],pp164[91],pp164[92],pp164[93],pp164[94],pp164[95],pp164[96],pp164[97],pp164[98],pp164[99],pp99[165],pp98[167],pp98[168],pp98[169],pp98[170],pp98[171],pp98[172],pp98[173],pp98[174],pp98[175],pp98[176],pp98[177],pp98[178],pp98[179],pp98[180],pp98[181],pp98[182],pp98[183],pp98[184],pp98[185],pp98[186],pp98[187],pp98[188],pp98[189],pp98[190],pp98[191],pp98[192],pp98[193],pp98[194],pp98[195],pp98[196],pp98[197],pp98[198],pp98[199],pp98[200],pp98[201],pp98[202],pp98[203],pp98[204],pp98[205],pp98[206],pp98[207],pp98[208]};
    assign in78_2 = {pp165[40],pp165[41],pp165[42],pp165[43],pp165[44],pp165[45],pp165[46],pp165[47],pp165[48],pp165[49],pp165[50],pp165[51],pp165[52],pp165[53],pp165[54],pp165[55],pp165[56],pp165[57],pp165[58],pp165[59],pp165[60],pp165[61],pp165[62],pp165[63],pp165[64],pp165[65],pp165[66],pp165[67],pp165[68],pp165[69],pp165[70],pp165[71],pp165[72],pp165[73],pp165[74],pp165[75],pp165[76],pp165[77],pp165[78],pp165[79],pp165[80],pp165[81],pp165[82],pp165[83],pp165[84],pp165[85],pp165[86],pp165[87],pp165[88],pp165[89],pp165[90],pp165[91],pp165[92],pp165[93],pp165[94],pp165[95],pp165[96],pp165[97],pp165[98],pp165[99],pp99[166],pp99[167],pp99[168],pp99[169],pp99[170],pp99[171],pp99[172],pp99[173],pp99[174],pp99[175],pp99[176],pp99[177],pp99[178],pp99[179],pp99[180],pp99[181],pp99[182],pp99[183],pp99[184],pp99[185],pp99[186],pp99[187],pp99[188],pp99[189],pp99[190],pp99[191],pp99[192],pp99[193],pp99[194],pp99[195],pp99[196],pp99[197],pp99[198],pp99[199],pp99[200],pp99[201],pp99[202],pp99[203],pp99[204],pp99[205],pp99[206],pp99[207]};
    CLA_102 KS_78(s78, c78, in78_1, in78_2);
    wire[99:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp166[40],pp166[41],pp166[42],pp166[43],pp166[44],pp166[45],pp166[46],pp166[47],pp166[48],pp166[49],pp166[50],pp166[51],pp166[52],pp166[53],pp166[54],pp166[55],pp166[56],pp166[57],pp166[58],pp166[59],pp166[60],pp166[61],pp166[62],pp166[63],pp166[64],pp166[65],pp166[66],pp166[67],pp166[68],pp166[69],pp166[70],pp166[71],pp166[72],pp166[73],pp166[74],pp166[75],pp166[76],pp166[77],pp166[78],pp166[79],pp166[80],pp166[81],pp166[82],pp166[83],pp166[84],pp166[85],pp166[86],pp166[87],pp166[88],pp166[89],pp166[90],pp166[91],pp166[92],pp166[93],pp166[94],pp166[95],pp166[96],pp166[97],pp166[98],pp166[99],pp167[99],pp168[99],pp169[99],pp170[99],pp171[99],pp172[99],pp173[99],pp174[99],pp175[99],pp176[99],pp177[99],pp178[99],pp179[99],pp180[99],pp181[99],pp182[99],pp183[99],pp184[99],pp185[99],pp186[99],pp187[99],pp188[99],pp189[99],pp190[99],pp191[99],pp192[99],pp193[99],pp194[99],pp195[99],pp196[99],pp197[99],pp198[99],pp199[99],pp200[99],pp201[99],pp202[99],pp203[99],pp204[99],pp205[99],pp206[99]};
    assign in79_2 = {pp167[39],pp167[40],pp167[41],pp167[42],pp167[43],pp167[44],pp167[45],pp167[46],pp167[47],pp167[48],pp167[49],pp167[50],pp167[51],pp167[52],pp167[53],pp167[54],pp167[55],pp167[56],pp167[57],pp167[58],pp167[59],pp167[60],pp167[61],pp167[62],pp167[63],pp167[64],pp167[65],pp167[66],pp167[67],pp167[68],pp167[69],pp167[70],pp167[71],pp167[72],pp167[73],pp167[74],pp167[75],pp167[76],pp167[77],pp167[78],pp167[79],pp167[80],pp167[81],pp167[82],pp167[83],pp167[84],pp167[85],pp167[86],pp167[87],pp167[88],pp167[89],pp167[90],pp167[91],pp167[92],pp167[93],pp167[94],pp167[95],pp167[96],pp167[97],pp167[98],pp168[98],pp169[98],pp170[98],pp171[98],pp172[98],pp173[98],pp174[98],pp175[98],pp176[98],pp177[98],pp178[98],pp179[98],pp180[98],pp181[98],pp182[98],pp183[98],pp184[98],pp185[98],pp186[98],pp187[98],pp188[98],pp189[98],pp190[98],pp191[98],pp192[98],pp193[98],pp194[98],pp195[98],pp196[98],pp197[98],pp198[98],pp199[98],pp200[98],pp201[98],pp202[98],pp203[98],pp204[98],pp205[98],pp206[98],pp207[98]};
    CLA_100 KS_79(s79, c79, in79_1, in79_2);
    wire[97:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp168[39],pp168[40],pp168[41],pp168[42],pp168[43],pp168[44],pp168[45],pp168[46],pp168[47],pp168[48],pp168[49],pp168[50],pp168[51],pp168[52],pp168[53],pp168[54],pp168[55],pp168[56],pp168[57],pp168[58],pp168[59],pp168[60],pp168[61],pp168[62],pp168[63],pp168[64],pp168[65],pp168[66],pp168[67],pp168[68],pp168[69],pp168[70],pp168[71],pp168[72],pp168[73],pp168[74],pp168[75],pp168[76],pp168[77],pp168[78],pp168[79],pp168[80],pp168[81],pp168[82],pp168[83],pp168[84],pp168[85],pp168[86],pp168[87],pp168[88],pp168[89],pp168[90],pp168[91],pp168[92],pp168[93],pp168[94],pp168[95],pp168[96],pp168[97],pp169[97],pp170[97],pp171[97],pp172[97],pp173[97],pp174[97],pp175[97],pp176[97],pp177[97],pp178[97],pp179[97],pp180[97],pp181[97],pp182[97],pp183[97],pp184[97],pp185[97],pp186[97],pp187[97],pp188[97],pp189[97],pp190[97],pp191[97],pp192[97],pp193[97],pp194[97],pp195[97],pp196[97],pp197[97],pp198[97],pp199[97],pp200[97],pp201[97],pp202[97],pp203[97],pp204[97],pp205[97],pp206[97],pp207[97]};
    assign in80_2 = {pp169[38],pp169[39],pp169[40],pp169[41],pp169[42],pp169[43],pp169[44],pp169[45],pp169[46],pp169[47],pp169[48],pp169[49],pp169[50],pp169[51],pp169[52],pp169[53],pp169[54],pp169[55],pp169[56],pp169[57],pp169[58],pp169[59],pp169[60],pp169[61],pp169[62],pp169[63],pp169[64],pp169[65],pp169[66],pp169[67],pp169[68],pp169[69],pp169[70],pp169[71],pp169[72],pp169[73],pp169[74],pp169[75],pp169[76],pp169[77],pp169[78],pp169[79],pp169[80],pp169[81],pp169[82],pp169[83],pp169[84],pp169[85],pp169[86],pp169[87],pp169[88],pp169[89],pp169[90],pp169[91],pp169[92],pp169[93],pp169[94],pp169[95],pp169[96],pp170[96],pp171[96],pp172[96],pp173[96],pp174[96],pp175[96],pp176[96],pp177[96],pp178[96],pp179[96],pp180[96],pp181[96],pp182[96],pp183[96],pp184[96],pp185[96],pp186[96],pp187[96],pp188[96],pp189[96],pp190[96],pp191[96],pp192[96],pp193[96],pp194[96],pp195[96],pp196[96],pp197[96],pp198[96],pp199[96],pp200[96],pp201[96],pp202[96],pp203[96],pp204[96],pp205[96],pp206[96],pp207[96],pp208[96]};
    CLA_98 KS_80(s80, c80, in80_1, in80_2);
    wire[95:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp170[38],pp170[39],pp170[40],pp170[41],pp170[42],pp170[43],pp170[44],pp170[45],pp170[46],pp170[47],pp170[48],pp170[49],pp170[50],pp170[51],pp170[52],pp170[53],pp170[54],pp170[55],pp170[56],pp170[57],pp170[58],pp170[59],pp170[60],pp170[61],pp170[62],pp170[63],pp170[64],pp170[65],pp170[66],pp170[67],pp170[68],pp170[69],pp170[70],pp170[71],pp170[72],pp170[73],pp170[74],pp170[75],pp170[76],pp170[77],pp170[78],pp170[79],pp170[80],pp170[81],pp170[82],pp170[83],pp170[84],pp170[85],pp170[86],pp170[87],pp170[88],pp170[89],pp170[90],pp170[91],pp170[92],pp170[93],pp170[94],pp170[95],pp171[95],pp172[95],pp173[95],pp174[95],pp175[95],pp176[95],pp177[95],pp178[95],pp179[95],pp180[95],pp181[95],pp182[95],pp183[95],pp184[95],pp185[95],pp186[95],pp187[95],pp188[95],pp189[95],pp190[95],pp191[95],pp192[95],pp193[95],pp194[95],pp195[95],pp196[95],pp197[95],pp198[95],pp199[95],pp200[95],pp201[95],pp202[95],pp203[95],pp204[95],pp205[95],pp206[95],pp207[95],pp208[95]};
    assign in81_2 = {pp171[37],pp171[38],pp171[39],pp171[40],pp171[41],pp171[42],pp171[43],pp171[44],pp171[45],pp171[46],pp171[47],pp171[48],pp171[49],pp171[50],pp171[51],pp171[52],pp171[53],pp171[54],pp171[55],pp171[56],pp171[57],pp171[58],pp171[59],pp171[60],pp171[61],pp171[62],pp171[63],pp171[64],pp171[65],pp171[66],pp171[67],pp171[68],pp171[69],pp171[70],pp171[71],pp171[72],pp171[73],pp171[74],pp171[75],pp171[76],pp171[77],pp171[78],pp171[79],pp171[80],pp171[81],pp171[82],pp171[83],pp171[84],pp171[85],pp171[86],pp171[87],pp171[88],pp171[89],pp171[90],pp171[91],pp171[92],pp171[93],pp171[94],pp172[94],pp173[94],pp174[94],pp175[94],pp176[94],pp177[94],pp178[94],pp179[94],pp180[94],pp181[94],pp182[94],pp183[94],pp184[94],pp185[94],pp186[94],pp187[94],pp188[94],pp189[94],pp190[94],pp191[94],pp192[94],pp193[94],pp194[94],pp195[94],pp196[94],pp197[94],pp198[94],pp199[94],pp200[94],pp201[94],pp202[94],pp203[94],pp204[94],pp205[94],pp206[94],pp207[94],pp208[94],pp209[94]};
    CLA_96 KS_81(s81, c81, in81_1, in81_2);
    wire[93:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp172[37],pp172[38],pp172[39],pp172[40],pp172[41],pp172[42],pp172[43],pp172[44],pp172[45],pp172[46],pp172[47],pp172[48],pp172[49],pp172[50],pp172[51],pp172[52],pp172[53],pp172[54],pp172[55],pp172[56],pp172[57],pp172[58],pp172[59],pp172[60],pp172[61],pp172[62],pp172[63],pp172[64],pp172[65],pp172[66],pp172[67],pp172[68],pp172[69],pp172[70],pp172[71],pp172[72],pp172[73],pp172[74],pp172[75],pp172[76],pp172[77],pp172[78],pp172[79],pp172[80],pp172[81],pp172[82],pp172[83],pp172[84],pp172[85],pp172[86],pp172[87],pp172[88],pp172[89],pp172[90],pp172[91],pp172[92],pp172[93],pp173[93],pp174[93],pp175[93],pp176[93],pp177[93],pp178[93],pp179[93],pp180[93],pp181[93],pp182[93],pp183[93],pp184[93],pp185[93],pp186[93],pp187[93],pp188[93],pp189[93],pp190[93],pp191[93],pp192[93],pp193[93],pp194[93],pp195[93],pp196[93],pp197[93],pp198[93],pp199[93],pp200[93],pp201[93],pp202[93],pp203[93],pp204[93],pp205[93],pp206[93],pp207[93],pp208[93],pp209[93]};
    assign in82_2 = {pp173[36],pp173[37],pp173[38],pp173[39],pp173[40],pp173[41],pp173[42],pp173[43],pp173[44],pp173[45],pp173[46],pp173[47],pp173[48],pp173[49],pp173[50],pp173[51],pp173[52],pp173[53],pp173[54],pp173[55],pp173[56],pp173[57],pp173[58],pp173[59],pp173[60],pp173[61],pp173[62],pp173[63],pp173[64],pp173[65],pp173[66],pp173[67],pp173[68],pp173[69],pp173[70],pp173[71],pp173[72],pp173[73],pp173[74],pp173[75],pp173[76],pp173[77],pp173[78],pp173[79],pp173[80],pp173[81],pp173[82],pp173[83],pp173[84],pp173[85],pp173[86],pp173[87],pp173[88],pp173[89],pp173[90],pp173[91],pp173[92],pp174[92],pp175[92],pp176[92],pp177[92],pp178[92],pp179[92],pp180[92],pp181[92],pp182[92],pp183[92],pp184[92],pp185[92],pp186[92],pp187[92],pp188[92],pp189[92],pp190[92],pp191[92],pp192[92],pp193[92],pp194[92],pp195[92],pp196[92],pp197[92],pp198[92],pp199[92],pp200[92],pp201[92],pp202[92],pp203[92],pp204[92],pp205[92],pp206[92],pp207[92],pp208[92],pp209[92],pp210[92]};
    CLA_94 KS_82(s82, c82, in82_1, in82_2);
    wire[91:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp174[36],pp174[37],pp174[38],pp174[39],pp174[40],pp174[41],pp174[42],pp174[43],pp174[44],pp174[45],pp174[46],pp174[47],pp174[48],pp174[49],pp174[50],pp174[51],pp174[52],pp174[53],pp174[54],pp174[55],pp174[56],pp174[57],pp174[58],pp174[59],pp174[60],pp174[61],pp174[62],pp174[63],pp174[64],pp174[65],pp174[66],pp174[67],pp174[68],pp174[69],pp174[70],pp174[71],pp174[72],pp174[73],pp174[74],pp174[75],pp174[76],pp174[77],pp174[78],pp174[79],pp174[80],pp174[81],pp174[82],pp174[83],pp174[84],pp174[85],pp174[86],pp174[87],pp174[88],pp174[89],pp174[90],pp174[91],pp175[91],pp176[91],pp177[91],pp178[91],pp179[91],pp180[91],pp181[91],pp182[91],pp183[91],pp184[91],pp185[91],pp186[91],pp187[91],pp188[91],pp189[91],pp190[91],pp191[91],pp192[91],pp193[91],pp194[91],pp195[91],pp196[91],pp197[91],pp198[91],pp199[91],pp200[91],pp201[91],pp202[91],pp203[91],pp204[91],pp205[91],pp206[91],pp207[91],pp208[91],pp209[91],pp210[91]};
    assign in83_2 = {pp175[35],pp175[36],pp175[37],pp175[38],pp175[39],pp175[40],pp175[41],pp175[42],pp175[43],pp175[44],pp175[45],pp175[46],pp175[47],pp175[48],pp175[49],pp175[50],pp175[51],pp175[52],pp175[53],pp175[54],pp175[55],pp175[56],pp175[57],pp175[58],pp175[59],pp175[60],pp175[61],pp175[62],pp175[63],pp175[64],pp175[65],pp175[66],pp175[67],pp175[68],pp175[69],pp175[70],pp175[71],pp175[72],pp175[73],pp175[74],pp175[75],pp175[76],pp175[77],pp175[78],pp175[79],pp175[80],pp175[81],pp175[82],pp175[83],pp175[84],pp175[85],pp175[86],pp175[87],pp175[88],pp175[89],pp175[90],pp176[90],pp177[90],pp178[90],pp179[90],pp180[90],pp181[90],pp182[90],pp183[90],pp184[90],pp185[90],pp186[90],pp187[90],pp188[90],pp189[90],pp190[90],pp191[90],pp192[90],pp193[90],pp194[90],pp195[90],pp196[90],pp197[90],pp198[90],pp199[90],pp200[90],pp201[90],pp202[90],pp203[90],pp204[90],pp205[90],pp206[90],pp207[90],pp208[90],pp209[90],pp210[90],pp211[90]};
    CLA_92 KS_83(s83, c83, in83_1, in83_2);
    wire[89:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp176[35],pp176[36],pp176[37],pp176[38],pp176[39],pp176[40],pp176[41],pp176[42],pp176[43],pp176[44],pp176[45],pp176[46],pp176[47],pp176[48],pp176[49],pp176[50],pp176[51],pp176[52],pp176[53],pp176[54],pp176[55],pp176[56],pp176[57],pp176[58],pp176[59],pp176[60],pp176[61],pp176[62],pp176[63],pp176[64],pp176[65],pp176[66],pp176[67],pp176[68],pp176[69],pp176[70],pp176[71],pp176[72],pp176[73],pp176[74],pp176[75],pp176[76],pp176[77],pp176[78],pp176[79],pp176[80],pp176[81],pp176[82],pp176[83],pp176[84],pp176[85],pp176[86],pp176[87],pp176[88],pp176[89],pp177[89],pp178[89],pp179[89],pp180[89],pp181[89],pp182[89],pp183[89],pp184[89],pp185[89],pp186[89],pp187[89],pp188[89],pp189[89],pp190[89],pp191[89],pp192[89],pp193[89],pp194[89],pp195[89],pp196[89],pp197[89],pp198[89],pp199[89],pp200[89],pp201[89],pp202[89],pp203[89],pp204[89],pp205[89],pp206[89],pp207[89],pp208[89],pp209[89],pp210[89],pp211[89]};
    assign in84_2 = {pp177[34],pp177[35],pp177[36],pp177[37],pp177[38],pp177[39],pp177[40],pp177[41],pp177[42],pp177[43],pp177[44],pp177[45],pp177[46],pp177[47],pp177[48],pp177[49],pp177[50],pp177[51],pp177[52],pp177[53],pp177[54],pp177[55],pp177[56],pp177[57],pp177[58],pp177[59],pp177[60],pp177[61],pp177[62],pp177[63],pp177[64],pp177[65],pp177[66],pp177[67],pp177[68],pp177[69],pp177[70],pp177[71],pp177[72],pp177[73],pp177[74],pp177[75],pp177[76],pp177[77],pp177[78],pp177[79],pp177[80],pp177[81],pp177[82],pp177[83],pp177[84],pp177[85],pp177[86],pp177[87],pp177[88],pp178[88],pp179[88],pp180[88],pp181[88],pp182[88],pp183[88],pp184[88],pp185[88],pp186[88],pp187[88],pp188[88],pp189[88],pp190[88],pp191[88],pp192[88],pp193[88],pp194[88],pp195[88],pp196[88],pp197[88],pp198[88],pp199[88],pp200[88],pp201[88],pp202[88],pp203[88],pp204[88],pp205[88],pp206[88],pp207[88],pp208[88],pp209[88],pp210[88],pp211[88],pp212[88]};
    CLA_90 KS_84(s84, c84, in84_1, in84_2);
    wire[87:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp178[34],pp178[35],pp178[36],pp178[37],pp178[38],pp178[39],pp178[40],pp178[41],pp178[42],pp178[43],pp178[44],pp178[45],pp178[46],pp178[47],pp178[48],pp178[49],pp178[50],pp178[51],pp178[52],pp178[53],pp178[54],pp178[55],pp178[56],pp178[57],pp178[58],pp178[59],pp178[60],pp178[61],pp178[62],pp178[63],pp178[64],pp178[65],pp178[66],pp178[67],pp178[68],pp178[69],pp178[70],pp178[71],pp178[72],pp178[73],pp178[74],pp178[75],pp178[76],pp178[77],pp178[78],pp178[79],pp178[80],pp178[81],pp178[82],pp178[83],pp178[84],pp178[85],pp178[86],pp178[87],pp179[87],pp180[87],pp181[87],pp182[87],pp183[87],pp184[87],pp185[87],pp186[87],pp187[87],pp188[87],pp189[87],pp190[87],pp191[87],pp192[87],pp193[87],pp194[87],pp195[87],pp196[87],pp197[87],pp198[87],pp199[87],pp200[87],pp201[87],pp202[87],pp203[87],pp204[87],pp205[87],pp206[87],pp207[87],pp208[87],pp209[87],pp210[87],pp211[87],pp212[87]};
    assign in85_2 = {pp179[33],pp179[34],pp179[35],pp179[36],pp179[37],pp179[38],pp179[39],pp179[40],pp179[41],pp179[42],pp179[43],pp179[44],pp179[45],pp179[46],pp179[47],pp179[48],pp179[49],pp179[50],pp179[51],pp179[52],pp179[53],pp179[54],pp179[55],pp179[56],pp179[57],pp179[58],pp179[59],pp179[60],pp179[61],pp179[62],pp179[63],pp179[64],pp179[65],pp179[66],pp179[67],pp179[68],pp179[69],pp179[70],pp179[71],pp179[72],pp179[73],pp179[74],pp179[75],pp179[76],pp179[77],pp179[78],pp179[79],pp179[80],pp179[81],pp179[82],pp179[83],pp179[84],pp179[85],pp179[86],pp180[86],pp181[86],pp182[86],pp183[86],pp184[86],pp185[86],pp186[86],pp187[86],pp188[86],pp189[86],pp190[86],pp191[86],pp192[86],pp193[86],pp194[86],pp195[86],pp196[86],pp197[86],pp198[86],pp199[86],pp200[86],pp201[86],pp202[86],pp203[86],pp204[86],pp205[86],pp206[86],pp207[86],pp208[86],pp209[86],pp210[86],pp211[86],pp212[86],pp213[86]};
    CLA_88 KS_85(s85, c85, in85_1, in85_2);
    wire[85:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp180[33],pp180[34],pp180[35],pp180[36],pp180[37],pp180[38],pp180[39],pp180[40],pp180[41],pp180[42],pp180[43],pp180[44],pp180[45],pp180[46],pp180[47],pp180[48],pp180[49],pp180[50],pp180[51],pp180[52],pp180[53],pp180[54],pp180[55],pp180[56],pp180[57],pp180[58],pp180[59],pp180[60],pp180[61],pp180[62],pp180[63],pp180[64],pp180[65],pp180[66],pp180[67],pp180[68],pp180[69],pp180[70],pp180[71],pp180[72],pp180[73],pp180[74],pp180[75],pp180[76],pp180[77],pp180[78],pp180[79],pp180[80],pp180[81],pp180[82],pp180[83],pp180[84],pp180[85],pp181[85],pp182[85],pp183[85],pp184[85],pp185[85],pp186[85],pp187[85],pp188[85],pp189[85],pp190[85],pp191[85],pp192[85],pp193[85],pp194[85],pp195[85],pp196[85],pp197[85],pp198[85],pp199[85],pp200[85],pp201[85],pp202[85],pp203[85],pp204[85],pp205[85],pp206[85],pp207[85],pp208[85],pp209[85],pp210[85],pp211[85],pp212[85],pp213[85]};
    assign in86_2 = {pp181[32],pp181[33],pp181[34],pp181[35],pp181[36],pp181[37],pp181[38],pp181[39],pp181[40],pp181[41],pp181[42],pp181[43],pp181[44],pp181[45],pp181[46],pp181[47],pp181[48],pp181[49],pp181[50],pp181[51],pp181[52],pp181[53],pp181[54],pp181[55],pp181[56],pp181[57],pp181[58],pp181[59],pp181[60],pp181[61],pp181[62],pp181[63],pp181[64],pp181[65],pp181[66],pp181[67],pp181[68],pp181[69],pp181[70],pp181[71],pp181[72],pp181[73],pp181[74],pp181[75],pp181[76],pp181[77],pp181[78],pp181[79],pp181[80],pp181[81],pp181[82],pp181[83],pp181[84],pp182[84],pp183[84],pp184[84],pp185[84],pp186[84],pp187[84],pp188[84],pp189[84],pp190[84],pp191[84],pp192[84],pp193[84],pp194[84],pp195[84],pp196[84],pp197[84],pp198[84],pp199[84],pp200[84],pp201[84],pp202[84],pp203[84],pp204[84],pp205[84],pp206[84],pp207[84],pp208[84],pp209[84],pp210[84],pp211[84],pp212[84],pp213[84],pp214[84]};
    CLA_86 KS_86(s86, c86, in86_1, in86_2);
    wire[83:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp182[32],pp182[33],pp182[34],pp182[35],pp182[36],pp182[37],pp182[38],pp182[39],pp182[40],pp182[41],pp182[42],pp182[43],pp182[44],pp182[45],pp182[46],pp182[47],pp182[48],pp182[49],pp182[50],pp182[51],pp182[52],pp182[53],pp182[54],pp182[55],pp182[56],pp182[57],pp182[58],pp182[59],pp182[60],pp182[61],pp182[62],pp182[63],pp182[64],pp182[65],pp182[66],pp182[67],pp182[68],pp182[69],pp182[70],pp182[71],pp182[72],pp182[73],pp182[74],pp182[75],pp182[76],pp182[77],pp182[78],pp182[79],pp182[80],pp182[81],pp182[82],pp182[83],pp183[83],pp184[83],pp185[83],pp186[83],pp187[83],pp188[83],pp189[83],pp190[83],pp191[83],pp192[83],pp193[83],pp194[83],pp195[83],pp196[83],pp197[83],pp198[83],pp199[83],pp200[83],pp201[83],pp202[83],pp203[83],pp204[83],pp205[83],pp206[83],pp207[83],pp208[83],pp209[83],pp210[83],pp211[83],pp212[83],pp213[83],pp214[83]};
    assign in87_2 = {pp183[31],pp183[32],pp183[33],pp183[34],pp183[35],pp183[36],pp183[37],pp183[38],pp183[39],pp183[40],pp183[41],pp183[42],pp183[43],pp183[44],pp183[45],pp183[46],pp183[47],pp183[48],pp183[49],pp183[50],pp183[51],pp183[52],pp183[53],pp183[54],pp183[55],pp183[56],pp183[57],pp183[58],pp183[59],pp183[60],pp183[61],pp183[62],pp183[63],pp183[64],pp183[65],pp183[66],pp183[67],pp183[68],pp183[69],pp183[70],pp183[71],pp183[72],pp183[73],pp183[74],pp183[75],pp183[76],pp183[77],pp183[78],pp183[79],pp183[80],pp183[81],pp183[82],pp184[82],pp185[82],pp186[82],pp187[82],pp188[82],pp189[82],pp190[82],pp191[82],pp192[82],pp193[82],pp194[82],pp195[82],pp196[82],pp197[82],pp198[82],pp199[82],pp200[82],pp201[82],pp202[82],pp203[82],pp204[82],pp205[82],pp206[82],pp207[82],pp208[82],pp209[82],pp210[82],pp211[82],pp212[82],pp213[82],pp214[82],pp215[82]};
    CLA_84 KS_87(s87, c87, in87_1, in87_2);
    wire[81:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp184[31],pp184[32],pp184[33],pp184[34],pp184[35],pp184[36],pp184[37],pp184[38],pp184[39],pp184[40],pp184[41],pp184[42],pp184[43],pp184[44],pp184[45],pp184[46],pp184[47],pp184[48],pp184[49],pp184[50],pp184[51],pp184[52],pp184[53],pp184[54],pp184[55],pp184[56],pp184[57],pp184[58],pp184[59],pp184[60],pp184[61],pp184[62],pp184[63],pp184[64],pp184[65],pp184[66],pp184[67],pp184[68],pp184[69],pp184[70],pp184[71],pp184[72],pp184[73],pp184[74],pp184[75],pp184[76],pp184[77],pp184[78],pp184[79],pp184[80],pp184[81],pp185[81],pp186[81],pp187[81],pp188[81],pp189[81],pp190[81],pp191[81],pp192[81],pp193[81],pp194[81],pp195[81],pp196[81],pp197[81],pp198[81],pp199[81],pp200[81],pp201[81],pp202[81],pp203[81],pp204[81],pp205[81],pp206[81],pp207[81],pp208[81],pp209[81],pp210[81],pp211[81],pp212[81],pp213[81],pp214[81],pp215[81]};
    assign in88_2 = {pp185[30],pp185[31],pp185[32],pp185[33],pp185[34],pp185[35],pp185[36],pp185[37],pp185[38],pp185[39],pp185[40],pp185[41],pp185[42],pp185[43],pp185[44],pp185[45],pp185[46],pp185[47],pp185[48],pp185[49],pp185[50],pp185[51],pp185[52],pp185[53],pp185[54],pp185[55],pp185[56],pp185[57],pp185[58],pp185[59],pp185[60],pp185[61],pp185[62],pp185[63],pp185[64],pp185[65],pp185[66],pp185[67],pp185[68],pp185[69],pp185[70],pp185[71],pp185[72],pp185[73],pp185[74],pp185[75],pp185[76],pp185[77],pp185[78],pp185[79],pp185[80],pp186[80],pp187[80],pp188[80],pp189[80],pp190[80],pp191[80],pp192[80],pp193[80],pp194[80],pp195[80],pp196[80],pp197[80],pp198[80],pp199[80],pp200[80],pp201[80],pp202[80],pp203[80],pp204[80],pp205[80],pp206[80],pp207[80],pp208[80],pp209[80],pp210[80],pp211[80],pp212[80],pp213[80],pp214[80],pp215[80],pp216[80]};
    CLA_82 KS_88(s88, c88, in88_1, in88_2);
    wire[79:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp186[30],pp186[31],pp186[32],pp186[33],pp186[34],pp186[35],pp186[36],pp186[37],pp186[38],pp186[39],pp186[40],pp186[41],pp186[42],pp186[43],pp186[44],pp186[45],pp186[46],pp186[47],pp186[48],pp186[49],pp186[50],pp186[51],pp186[52],pp186[53],pp186[54],pp186[55],pp186[56],pp186[57],pp186[58],pp186[59],pp186[60],pp186[61],pp186[62],pp186[63],pp186[64],pp186[65],pp186[66],pp186[67],pp186[68],pp186[69],pp186[70],pp186[71],pp186[72],pp186[73],pp186[74],pp186[75],pp186[76],pp186[77],pp186[78],pp186[79],pp187[79],pp188[79],pp189[79],pp190[79],pp191[79],pp192[79],pp193[79],pp194[79],pp195[79],pp196[79],pp197[79],pp198[79],pp199[79],pp200[79],pp201[79],pp202[79],pp203[79],pp204[79],pp205[79],pp206[79],pp207[79],pp208[79],pp209[79],pp210[79],pp211[79],pp212[79],pp213[79],pp214[79],pp215[79],pp216[79]};
    assign in89_2 = {pp187[29],pp187[30],pp187[31],pp187[32],pp187[33],pp187[34],pp187[35],pp187[36],pp187[37],pp187[38],pp187[39],pp187[40],pp187[41],pp187[42],pp187[43],pp187[44],pp187[45],pp187[46],pp187[47],pp187[48],pp187[49],pp187[50],pp187[51],pp187[52],pp187[53],pp187[54],pp187[55],pp187[56],pp187[57],pp187[58],pp187[59],pp187[60],pp187[61],pp187[62],pp187[63],pp187[64],pp187[65],pp187[66],pp187[67],pp187[68],pp187[69],pp187[70],pp187[71],pp187[72],pp187[73],pp187[74],pp187[75],pp187[76],pp187[77],pp187[78],pp188[78],pp189[78],pp190[78],pp191[78],pp192[78],pp193[78],pp194[78],pp195[78],pp196[78],pp197[78],pp198[78],pp199[78],pp200[78],pp201[78],pp202[78],pp203[78],pp204[78],pp205[78],pp206[78],pp207[78],pp208[78],pp209[78],pp210[78],pp211[78],pp212[78],pp213[78],pp214[78],pp215[78],pp216[78],pp217[78]};
    CLA_80 KS_89(s89, c89, in89_1, in89_2);
    wire[77:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp188[29],pp188[30],pp188[31],pp188[32],pp188[33],pp188[34],pp188[35],pp188[36],pp188[37],pp188[38],pp188[39],pp188[40],pp188[41],pp188[42],pp188[43],pp188[44],pp188[45],pp188[46],pp188[47],pp188[48],pp188[49],pp188[50],pp188[51],pp188[52],pp188[53],pp188[54],pp188[55],pp188[56],pp188[57],pp188[58],pp188[59],pp188[60],pp188[61],pp188[62],pp188[63],pp188[64],pp188[65],pp188[66],pp188[67],pp188[68],pp188[69],pp188[70],pp188[71],pp188[72],pp188[73],pp188[74],pp188[75],pp188[76],pp188[77],pp189[77],pp190[77],pp191[77],pp192[77],pp193[77],pp194[77],pp195[77],pp196[77],pp197[77],pp198[77],pp199[77],pp200[77],pp201[77],pp202[77],pp203[77],pp204[77],pp205[77],pp206[77],pp207[77],pp208[77],pp209[77],pp210[77],pp211[77],pp212[77],pp213[77],pp214[77],pp215[77],pp216[77],pp217[77]};
    assign in90_2 = {pp189[28],pp189[29],pp189[30],pp189[31],pp189[32],pp189[33],pp189[34],pp189[35],pp189[36],pp189[37],pp189[38],pp189[39],pp189[40],pp189[41],pp189[42],pp189[43],pp189[44],pp189[45],pp189[46],pp189[47],pp189[48],pp189[49],pp189[50],pp189[51],pp189[52],pp189[53],pp189[54],pp189[55],pp189[56],pp189[57],pp189[58],pp189[59],pp189[60],pp189[61],pp189[62],pp189[63],pp189[64],pp189[65],pp189[66],pp189[67],pp189[68],pp189[69],pp189[70],pp189[71],pp189[72],pp189[73],pp189[74],pp189[75],pp189[76],pp190[76],pp191[76],pp192[76],pp193[76],pp194[76],pp195[76],pp196[76],pp197[76],pp198[76],pp199[76],pp200[76],pp201[76],pp202[76],pp203[76],pp204[76],pp205[76],pp206[76],pp207[76],pp208[76],pp209[76],pp210[76],pp211[76],pp212[76],pp213[76],pp214[76],pp215[76],pp216[76],pp217[76],pp218[76]};
    CLA_78 KS_90(s90, c90, in90_1, in90_2);
    wire[75:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp190[28],pp190[29],pp190[30],pp190[31],pp190[32],pp190[33],pp190[34],pp190[35],pp190[36],pp190[37],pp190[38],pp190[39],pp190[40],pp190[41],pp190[42],pp190[43],pp190[44],pp190[45],pp190[46],pp190[47],pp190[48],pp190[49],pp190[50],pp190[51],pp190[52],pp190[53],pp190[54],pp190[55],pp190[56],pp190[57],pp190[58],pp190[59],pp190[60],pp190[61],pp190[62],pp190[63],pp190[64],pp190[65],pp190[66],pp190[67],pp190[68],pp190[69],pp190[70],pp190[71],pp190[72],pp190[73],pp190[74],pp190[75],pp191[75],pp192[75],pp193[75],pp194[75],pp195[75],pp196[75],pp197[75],pp198[75],pp199[75],pp200[75],pp201[75],pp202[75],pp203[75],pp204[75],pp205[75],pp206[75],pp207[75],pp208[75],pp209[75],pp210[75],pp211[75],pp212[75],pp213[75],pp214[75],pp215[75],pp216[75],pp217[75],pp218[75]};
    assign in91_2 = {pp191[27],pp191[28],pp191[29],pp191[30],pp191[31],pp191[32],pp191[33],pp191[34],pp191[35],pp191[36],pp191[37],pp191[38],pp191[39],pp191[40],pp191[41],pp191[42],pp191[43],pp191[44],pp191[45],pp191[46],pp191[47],pp191[48],pp191[49],pp191[50],pp191[51],pp191[52],pp191[53],pp191[54],pp191[55],pp191[56],pp191[57],pp191[58],pp191[59],pp191[60],pp191[61],pp191[62],pp191[63],pp191[64],pp191[65],pp191[66],pp191[67],pp191[68],pp191[69],pp191[70],pp191[71],pp191[72],pp191[73],pp191[74],pp192[74],pp193[74],pp194[74],pp195[74],pp196[74],pp197[74],pp198[74],pp199[74],pp200[74],pp201[74],pp202[74],pp203[74],pp204[74],pp205[74],pp206[74],pp207[74],pp208[74],pp209[74],pp210[74],pp211[74],pp212[74],pp213[74],pp214[74],pp215[74],pp216[74],pp217[74],pp218[74],pp219[74]};
    CLA_76 KS_91(s91, c91, in91_1, in91_2);
    wire[73:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp192[27],pp192[28],pp192[29],pp192[30],pp192[31],pp192[32],pp192[33],pp192[34],pp192[35],pp192[36],pp192[37],pp192[38],pp192[39],pp192[40],pp192[41],pp192[42],pp192[43],pp192[44],pp192[45],pp192[46],pp192[47],pp192[48],pp192[49],pp192[50],pp192[51],pp192[52],pp192[53],pp192[54],pp192[55],pp192[56],pp192[57],pp192[58],pp192[59],pp192[60],pp192[61],pp192[62],pp192[63],pp192[64],pp192[65],pp192[66],pp192[67],pp192[68],pp192[69],pp192[70],pp192[71],pp192[72],pp192[73],pp193[73],pp194[73],pp195[73],pp196[73],pp197[73],pp198[73],pp199[73],pp200[73],pp201[73],pp202[73],pp203[73],pp204[73],pp205[73],pp206[73],pp207[73],pp208[73],pp209[73],pp210[73],pp211[73],pp212[73],pp213[73],pp214[73],pp215[73],pp216[73],pp217[73],pp218[73],pp219[73]};
    assign in92_2 = {pp193[26],pp193[27],pp193[28],pp193[29],pp193[30],pp193[31],pp193[32],pp193[33],pp193[34],pp193[35],pp193[36],pp193[37],pp193[38],pp193[39],pp193[40],pp193[41],pp193[42],pp193[43],pp193[44],pp193[45],pp193[46],pp193[47],pp193[48],pp193[49],pp193[50],pp193[51],pp193[52],pp193[53],pp193[54],pp193[55],pp193[56],pp193[57],pp193[58],pp193[59],pp193[60],pp193[61],pp193[62],pp193[63],pp193[64],pp193[65],pp193[66],pp193[67],pp193[68],pp193[69],pp193[70],pp193[71],pp193[72],pp194[72],pp195[72],pp196[72],pp197[72],pp198[72],pp199[72],pp200[72],pp201[72],pp202[72],pp203[72],pp204[72],pp205[72],pp206[72],pp207[72],pp208[72],pp209[72],pp210[72],pp211[72],pp212[72],pp213[72],pp214[72],pp215[72],pp216[72],pp217[72],pp218[72],pp219[72],pp220[72]};
    CLA_74 KS_92(s92, c92, in92_1, in92_2);
    wire[71:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp194[26],pp194[27],pp194[28],pp194[29],pp194[30],pp194[31],pp194[32],pp194[33],pp194[34],pp194[35],pp194[36],pp194[37],pp194[38],pp194[39],pp194[40],pp194[41],pp194[42],pp194[43],pp194[44],pp194[45],pp194[46],pp194[47],pp194[48],pp194[49],pp194[50],pp194[51],pp194[52],pp194[53],pp194[54],pp194[55],pp194[56],pp194[57],pp194[58],pp194[59],pp194[60],pp194[61],pp194[62],pp194[63],pp194[64],pp194[65],pp194[66],pp194[67],pp194[68],pp194[69],pp194[70],pp194[71],pp195[71],pp196[71],pp197[71],pp198[71],pp199[71],pp200[71],pp201[71],pp202[71],pp203[71],pp204[71],pp205[71],pp206[71],pp207[71],pp208[71],pp209[71],pp210[71],pp211[71],pp212[71],pp213[71],pp214[71],pp215[71],pp216[71],pp217[71],pp218[71],pp219[71],pp220[71]};
    assign in93_2 = {pp195[25],pp195[26],pp195[27],pp195[28],pp195[29],pp195[30],pp195[31],pp195[32],pp195[33],pp195[34],pp195[35],pp195[36],pp195[37],pp195[38],pp195[39],pp195[40],pp195[41],pp195[42],pp195[43],pp195[44],pp195[45],pp195[46],pp195[47],pp195[48],pp195[49],pp195[50],pp195[51],pp195[52],pp195[53],pp195[54],pp195[55],pp195[56],pp195[57],pp195[58],pp195[59],pp195[60],pp195[61],pp195[62],pp195[63],pp195[64],pp195[65],pp195[66],pp195[67],pp195[68],pp195[69],pp195[70],pp196[70],pp197[70],pp198[70],pp199[70],pp200[70],pp201[70],pp202[70],pp203[70],pp204[70],pp205[70],pp206[70],pp207[70],pp208[70],pp209[70],pp210[70],pp211[70],pp212[70],pp213[70],pp214[70],pp215[70],pp216[70],pp217[70],pp218[70],pp219[70],pp220[70],pp221[70]};
    CLA_72 KS_93(s93, c93, in93_1, in93_2);
    wire[69:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp196[25],pp196[26],pp196[27],pp196[28],pp196[29],pp196[30],pp196[31],pp196[32],pp196[33],pp196[34],pp196[35],pp196[36],pp196[37],pp196[38],pp196[39],pp196[40],pp196[41],pp196[42],pp196[43],pp196[44],pp196[45],pp196[46],pp196[47],pp196[48],pp196[49],pp196[50],pp196[51],pp196[52],pp196[53],pp196[54],pp196[55],pp196[56],pp196[57],pp196[58],pp196[59],pp196[60],pp196[61],pp196[62],pp196[63],pp196[64],pp196[65],pp196[66],pp196[67],pp196[68],pp196[69],pp197[69],pp198[69],pp199[69],pp200[69],pp201[69],pp202[69],pp203[69],pp204[69],pp205[69],pp206[69],pp207[69],pp208[69],pp209[69],pp210[69],pp211[69],pp212[69],pp213[69],pp214[69],pp215[69],pp216[69],pp217[69],pp218[69],pp219[69],pp220[69],pp221[69]};
    assign in94_2 = {pp197[24],pp197[25],pp197[26],pp197[27],pp197[28],pp197[29],pp197[30],pp197[31],pp197[32],pp197[33],pp197[34],pp197[35],pp197[36],pp197[37],pp197[38],pp197[39],pp197[40],pp197[41],pp197[42],pp197[43],pp197[44],pp197[45],pp197[46],pp197[47],pp197[48],pp197[49],pp197[50],pp197[51],pp197[52],pp197[53],pp197[54],pp197[55],pp197[56],pp197[57],pp197[58],pp197[59],pp197[60],pp197[61],pp197[62],pp197[63],pp197[64],pp197[65],pp197[66],pp197[67],pp197[68],pp198[68],pp199[68],pp200[68],pp201[68],pp202[68],pp203[68],pp204[68],pp205[68],pp206[68],pp207[68],pp208[68],pp209[68],pp210[68],pp211[68],pp212[68],pp213[68],pp214[68],pp215[68],pp216[68],pp217[68],pp218[68],pp219[68],pp220[68],pp221[68],pp222[68]};
    CLA_70 KS_94(s94, c94, in94_1, in94_2);
    wire[67:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp198[24],pp198[25],pp198[26],pp198[27],pp198[28],pp198[29],pp198[30],pp198[31],pp198[32],pp198[33],pp198[34],pp198[35],pp198[36],pp198[37],pp198[38],pp198[39],pp198[40],pp198[41],pp198[42],pp198[43],pp198[44],pp198[45],pp198[46],pp198[47],pp198[48],pp198[49],pp198[50],pp198[51],pp198[52],pp198[53],pp198[54],pp198[55],pp198[56],pp198[57],pp198[58],pp198[59],pp198[60],pp198[61],pp198[62],pp198[63],pp198[64],pp198[65],pp198[66],pp198[67],pp199[67],pp200[67],pp201[67],pp202[67],pp203[67],pp204[67],pp205[67],pp206[67],pp207[67],pp208[67],pp209[67],pp210[67],pp211[67],pp212[67],pp213[67],pp214[67],pp215[67],pp216[67],pp217[67],pp218[67],pp219[67],pp220[67],pp221[67],pp222[67]};
    assign in95_2 = {pp199[23],pp199[24],pp199[25],pp199[26],pp199[27],pp199[28],pp199[29],pp199[30],pp199[31],pp199[32],pp199[33],pp199[34],pp199[35],pp199[36],pp199[37],pp199[38],pp199[39],pp199[40],pp199[41],pp199[42],pp199[43],pp199[44],pp199[45],pp199[46],pp199[47],pp199[48],pp199[49],pp199[50],pp199[51],pp199[52],pp199[53],pp199[54],pp199[55],pp199[56],pp199[57],pp199[58],pp199[59],pp199[60],pp199[61],pp199[62],pp199[63],pp199[64],pp199[65],pp199[66],pp200[66],pp201[66],pp202[66],pp203[66],pp204[66],pp205[66],pp206[66],pp207[66],pp208[66],pp209[66],pp210[66],pp211[66],pp212[66],pp213[66],pp214[66],pp215[66],pp216[66],pp217[66],pp218[66],pp219[66],pp220[66],pp221[66],pp222[66],pp223[66]};
    CLA_68 KS_95(s95, c95, in95_1, in95_2);
    wire[65:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp200[23],pp200[24],pp200[25],pp200[26],pp200[27],pp200[28],pp200[29],pp200[30],pp200[31],pp200[32],pp200[33],pp200[34],pp200[35],pp200[36],pp200[37],pp200[38],pp200[39],pp200[40],pp200[41],pp200[42],pp200[43],pp200[44],pp200[45],pp200[46],pp200[47],pp200[48],pp200[49],pp200[50],pp200[51],pp200[52],pp200[53],pp200[54],pp200[55],pp200[56],pp200[57],pp200[58],pp200[59],pp200[60],pp200[61],pp200[62],pp200[63],pp200[64],pp200[65],pp201[65],pp202[65],pp203[65],pp204[65],pp205[65],pp206[65],pp207[65],pp208[65],pp209[65],pp210[65],pp211[65],pp212[65],pp213[65],pp214[65],pp215[65],pp216[65],pp217[65],pp218[65],pp219[65],pp220[65],pp221[65],pp222[65],pp223[65]};
    assign in96_2 = {pp201[22],pp201[23],pp201[24],pp201[25],pp201[26],pp201[27],pp201[28],pp201[29],pp201[30],pp201[31],pp201[32],pp201[33],pp201[34],pp201[35],pp201[36],pp201[37],pp201[38],pp201[39],pp201[40],pp201[41],pp201[42],pp201[43],pp201[44],pp201[45],pp201[46],pp201[47],pp201[48],pp201[49],pp201[50],pp201[51],pp201[52],pp201[53],pp201[54],pp201[55],pp201[56],pp201[57],pp201[58],pp201[59],pp201[60],pp201[61],pp201[62],pp201[63],pp201[64],pp202[64],pp203[64],pp204[64],pp205[64],pp206[64],pp207[64],pp208[64],pp209[64],pp210[64],pp211[64],pp212[64],pp213[64],pp214[64],pp215[64],pp216[64],pp217[64],pp218[64],pp219[64],pp220[64],pp221[64],pp222[64],pp223[64],pp224[64]};
    CLA_66 KS_96(s96, c96, in96_1, in96_2);
    wire[63:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp202[22],pp202[23],pp202[24],pp202[25],pp202[26],pp202[27],pp202[28],pp202[29],pp202[30],pp202[31],pp202[32],pp202[33],pp202[34],pp202[35],pp202[36],pp202[37],pp202[38],pp202[39],pp202[40],pp202[41],pp202[42],pp202[43],pp202[44],pp202[45],pp202[46],pp202[47],pp202[48],pp202[49],pp202[50],pp202[51],pp202[52],pp202[53],pp202[54],pp202[55],pp202[56],pp202[57],pp202[58],pp202[59],pp202[60],pp202[61],pp202[62],pp202[63],pp203[63],pp204[63],pp205[63],pp206[63],pp207[63],pp208[63],pp209[63],pp210[63],pp211[63],pp212[63],pp213[63],pp214[63],pp215[63],pp216[63],pp217[63],pp218[63],pp219[63],pp220[63],pp221[63],pp222[63],pp223[63],pp224[63]};
    assign in97_2 = {pp203[21],pp203[22],pp203[23],pp203[24],pp203[25],pp203[26],pp203[27],pp203[28],pp203[29],pp203[30],pp203[31],pp203[32],pp203[33],pp203[34],pp203[35],pp203[36],pp203[37],pp203[38],pp203[39],pp203[40],pp203[41],pp203[42],pp203[43],pp203[44],pp203[45],pp203[46],pp203[47],pp203[48],pp203[49],pp203[50],pp203[51],pp203[52],pp203[53],pp203[54],pp203[55],pp203[56],pp203[57],pp203[58],pp203[59],pp203[60],pp203[61],pp203[62],pp204[62],pp205[62],pp206[62],pp207[62],pp208[62],pp209[62],pp210[62],pp211[62],pp212[62],pp213[62],pp214[62],pp215[62],pp216[62],pp217[62],pp218[62],pp219[62],pp220[62],pp221[62],pp222[62],pp223[62],pp224[62],pp225[62]};
    CLA_64 KS_97(s97, c97, in97_1, in97_2);
    wire[61:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp204[21],pp204[22],pp204[23],pp204[24],pp204[25],pp204[26],pp204[27],pp204[28],pp204[29],pp204[30],pp204[31],pp204[32],pp204[33],pp204[34],pp204[35],pp204[36],pp204[37],pp204[38],pp204[39],pp204[40],pp204[41],pp204[42],pp204[43],pp204[44],pp204[45],pp204[46],pp204[47],pp204[48],pp204[49],pp204[50],pp204[51],pp204[52],pp204[53],pp204[54],pp204[55],pp204[56],pp204[57],pp204[58],pp204[59],pp204[60],pp204[61],pp205[61],pp206[61],pp207[61],pp208[61],pp209[61],pp210[61],pp211[61],pp212[61],pp213[61],pp214[61],pp215[61],pp216[61],pp217[61],pp218[61],pp219[61],pp220[61],pp221[61],pp222[61],pp223[61],pp224[61],pp225[61]};
    assign in98_2 = {pp205[20],pp205[21],pp205[22],pp205[23],pp205[24],pp205[25],pp205[26],pp205[27],pp205[28],pp205[29],pp205[30],pp205[31],pp205[32],pp205[33],pp205[34],pp205[35],pp205[36],pp205[37],pp205[38],pp205[39],pp205[40],pp205[41],pp205[42],pp205[43],pp205[44],pp205[45],pp205[46],pp205[47],pp205[48],pp205[49],pp205[50],pp205[51],pp205[52],pp205[53],pp205[54],pp205[55],pp205[56],pp205[57],pp205[58],pp205[59],pp205[60],pp206[60],pp207[60],pp208[60],pp209[60],pp210[60],pp211[60],pp212[60],pp213[60],pp214[60],pp215[60],pp216[60],pp217[60],pp218[60],pp219[60],pp220[60],pp221[60],pp222[60],pp223[60],pp224[60],pp225[60],pp226[60]};
    CLA_62 KS_98(s98, c98, in98_1, in98_2);
    wire[59:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp206[20],pp206[21],pp206[22],pp206[23],pp206[24],pp206[25],pp206[26],pp206[27],pp206[28],pp206[29],pp206[30],pp206[31],pp206[32],pp206[33],pp206[34],pp206[35],pp206[36],pp206[37],pp206[38],pp206[39],pp206[40],pp206[41],pp206[42],pp206[43],pp206[44],pp206[45],pp206[46],pp206[47],pp206[48],pp206[49],pp206[50],pp206[51],pp206[52],pp206[53],pp206[54],pp206[55],pp206[56],pp206[57],pp206[58],pp206[59],pp207[59],pp208[59],pp209[59],pp210[59],pp211[59],pp212[59],pp213[59],pp214[59],pp215[59],pp216[59],pp217[59],pp218[59],pp219[59],pp220[59],pp221[59],pp222[59],pp223[59],pp224[59],pp225[59],pp226[59]};
    assign in99_2 = {pp207[19],pp207[20],pp207[21],pp207[22],pp207[23],pp207[24],pp207[25],pp207[26],pp207[27],pp207[28],pp207[29],pp207[30],pp207[31],pp207[32],pp207[33],pp207[34],pp207[35],pp207[36],pp207[37],pp207[38],pp207[39],pp207[40],pp207[41],pp207[42],pp207[43],pp207[44],pp207[45],pp207[46],pp207[47],pp207[48],pp207[49],pp207[50],pp207[51],pp207[52],pp207[53],pp207[54],pp207[55],pp207[56],pp207[57],pp207[58],pp208[58],pp209[58],pp210[58],pp211[58],pp212[58],pp213[58],pp214[58],pp215[58],pp216[58],pp217[58],pp218[58],pp219[58],pp220[58],pp221[58],pp222[58],pp223[58],pp224[58],pp225[58],pp226[58],pp227[58]};
    CLA_60 KS_99(s99, c99, in99_1, in99_2);
    wire[57:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp208[19],pp208[20],pp208[21],pp208[22],pp208[23],pp208[24],pp208[25],pp208[26],pp208[27],pp208[28],pp208[29],pp208[30],pp208[31],pp208[32],pp208[33],pp208[34],pp208[35],pp208[36],pp208[37],pp208[38],pp208[39],pp208[40],pp208[41],pp208[42],pp208[43],pp208[44],pp208[45],pp208[46],pp208[47],pp208[48],pp208[49],pp208[50],pp208[51],pp208[52],pp208[53],pp208[54],pp208[55],pp208[56],pp208[57],pp209[57],pp210[57],pp211[57],pp212[57],pp213[57],pp214[57],pp215[57],pp216[57],pp217[57],pp218[57],pp219[57],pp220[57],pp221[57],pp222[57],pp223[57],pp224[57],pp225[57],pp226[57],pp227[57]};
    assign in100_2 = {pp209[18],pp209[19],pp209[20],pp209[21],pp209[22],pp209[23],pp209[24],pp209[25],pp209[26],pp209[27],pp209[28],pp209[29],pp209[30],pp209[31],pp209[32],pp209[33],pp209[34],pp209[35],pp209[36],pp209[37],pp209[38],pp209[39],pp209[40],pp209[41],pp209[42],pp209[43],pp209[44],pp209[45],pp209[46],pp209[47],pp209[48],pp209[49],pp209[50],pp209[51],pp209[52],pp209[53],pp209[54],pp209[55],pp209[56],pp210[56],pp211[56],pp212[56],pp213[56],pp214[56],pp215[56],pp216[56],pp217[56],pp218[56],pp219[56],pp220[56],pp221[56],pp222[56],pp223[56],pp224[56],pp225[56],pp226[56],pp227[56],pp228[56]};
    CLA_58 KS_100(s100, c100, in100_1, in100_2);
    wire[55:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp210[18],pp210[19],pp210[20],pp210[21],pp210[22],pp210[23],pp210[24],pp210[25],pp210[26],pp210[27],pp210[28],pp210[29],pp210[30],pp210[31],pp210[32],pp210[33],pp210[34],pp210[35],pp210[36],pp210[37],pp210[38],pp210[39],pp210[40],pp210[41],pp210[42],pp210[43],pp210[44],pp210[45],pp210[46],pp210[47],pp210[48],pp210[49],pp210[50],pp210[51],pp210[52],pp210[53],pp210[54],pp210[55],pp211[55],pp212[55],pp213[55],pp214[55],pp215[55],pp216[55],pp217[55],pp218[55],pp219[55],pp220[55],pp221[55],pp222[55],pp223[55],pp224[55],pp225[55],pp226[55],pp227[55],pp228[55]};
    assign in101_2 = {pp211[17],pp211[18],pp211[19],pp211[20],pp211[21],pp211[22],pp211[23],pp211[24],pp211[25],pp211[26],pp211[27],pp211[28],pp211[29],pp211[30],pp211[31],pp211[32],pp211[33],pp211[34],pp211[35],pp211[36],pp211[37],pp211[38],pp211[39],pp211[40],pp211[41],pp211[42],pp211[43],pp211[44],pp211[45],pp211[46],pp211[47],pp211[48],pp211[49],pp211[50],pp211[51],pp211[52],pp211[53],pp211[54],pp212[54],pp213[54],pp214[54],pp215[54],pp216[54],pp217[54],pp218[54],pp219[54],pp220[54],pp221[54],pp222[54],pp223[54],pp224[54],pp225[54],pp226[54],pp227[54],pp228[54],pp229[54]};
    CLA_56 KS_101(s101, c101, in101_1, in101_2);
    wire[53:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp212[17],pp212[18],pp212[19],pp212[20],pp212[21],pp212[22],pp212[23],pp212[24],pp212[25],pp212[26],pp212[27],pp212[28],pp212[29],pp212[30],pp212[31],pp212[32],pp212[33],pp212[34],pp212[35],pp212[36],pp212[37],pp212[38],pp212[39],pp212[40],pp212[41],pp212[42],pp212[43],pp212[44],pp212[45],pp212[46],pp212[47],pp212[48],pp212[49],pp212[50],pp212[51],pp212[52],pp212[53],pp213[53],pp214[53],pp215[53],pp216[53],pp217[53],pp218[53],pp219[53],pp220[53],pp221[53],pp222[53],pp223[53],pp224[53],pp225[53],pp226[53],pp227[53],pp228[53],pp229[53]};
    assign in102_2 = {pp213[16],pp213[17],pp213[18],pp213[19],pp213[20],pp213[21],pp213[22],pp213[23],pp213[24],pp213[25],pp213[26],pp213[27],pp213[28],pp213[29],pp213[30],pp213[31],pp213[32],pp213[33],pp213[34],pp213[35],pp213[36],pp213[37],pp213[38],pp213[39],pp213[40],pp213[41],pp213[42],pp213[43],pp213[44],pp213[45],pp213[46],pp213[47],pp213[48],pp213[49],pp213[50],pp213[51],pp213[52],pp214[52],pp215[52],pp216[52],pp217[52],pp218[52],pp219[52],pp220[52],pp221[52],pp222[52],pp223[52],pp224[52],pp225[52],pp226[52],pp227[52],pp228[52],pp229[52],pp230[52]};
    CLA_54 KS_102(s102, c102, in102_1, in102_2);
    wire[51:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp214[16],pp214[17],pp214[18],pp214[19],pp214[20],pp214[21],pp214[22],pp214[23],pp214[24],pp214[25],pp214[26],pp214[27],pp214[28],pp214[29],pp214[30],pp214[31],pp214[32],pp214[33],pp214[34],pp214[35],pp214[36],pp214[37],pp214[38],pp214[39],pp214[40],pp214[41],pp214[42],pp214[43],pp214[44],pp214[45],pp214[46],pp214[47],pp214[48],pp214[49],pp214[50],pp214[51],pp215[51],pp216[51],pp217[51],pp218[51],pp219[51],pp220[51],pp221[51],pp222[51],pp223[51],pp224[51],pp225[51],pp226[51],pp227[51],pp228[51],pp229[51],pp230[51]};
    assign in103_2 = {pp215[15],pp215[16],pp215[17],pp215[18],pp215[19],pp215[20],pp215[21],pp215[22],pp215[23],pp215[24],pp215[25],pp215[26],pp215[27],pp215[28],pp215[29],pp215[30],pp215[31],pp215[32],pp215[33],pp215[34],pp215[35],pp215[36],pp215[37],pp215[38],pp215[39],pp215[40],pp215[41],pp215[42],pp215[43],pp215[44],pp215[45],pp215[46],pp215[47],pp215[48],pp215[49],pp215[50],pp216[50],pp217[50],pp218[50],pp219[50],pp220[50],pp221[50],pp222[50],pp223[50],pp224[50],pp225[50],pp226[50],pp227[50],pp228[50],pp229[50],pp230[50],pp231[50]};
    CLA_52 KS_103(s103, c103, in103_1, in103_2);
    wire[49:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp216[15],pp216[16],pp216[17],pp216[18],pp216[19],pp216[20],pp216[21],pp216[22],pp216[23],pp216[24],pp216[25],pp216[26],pp216[27],pp216[28],pp216[29],pp216[30],pp216[31],pp216[32],pp216[33],pp216[34],pp216[35],pp216[36],pp216[37],pp216[38],pp216[39],pp216[40],pp216[41],pp216[42],pp216[43],pp216[44],pp216[45],pp216[46],pp216[47],pp216[48],pp216[49],pp217[49],pp218[49],pp219[49],pp220[49],pp221[49],pp222[49],pp223[49],pp224[49],pp225[49],pp226[49],pp227[49],pp228[49],pp229[49],pp230[49],pp231[49]};
    assign in104_2 = {pp217[14],pp217[15],pp217[16],pp217[17],pp217[18],pp217[19],pp217[20],pp217[21],pp217[22],pp217[23],pp217[24],pp217[25],pp217[26],pp217[27],pp217[28],pp217[29],pp217[30],pp217[31],pp217[32],pp217[33],pp217[34],pp217[35],pp217[36],pp217[37],pp217[38],pp217[39],pp217[40],pp217[41],pp217[42],pp217[43],pp217[44],pp217[45],pp217[46],pp217[47],pp217[48],pp218[48],pp219[48],pp220[48],pp221[48],pp222[48],pp223[48],pp224[48],pp225[48],pp226[48],pp227[48],pp228[48],pp229[48],pp230[48],pp231[48],pp232[48]};
    CLA_50 KS_104(s104, c104, in104_1, in104_2);
    wire[47:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp218[14],pp218[15],pp218[16],pp218[17],pp218[18],pp218[19],pp218[20],pp218[21],pp218[22],pp218[23],pp218[24],pp218[25],pp218[26],pp218[27],pp218[28],pp218[29],pp218[30],pp218[31],pp218[32],pp218[33],pp218[34],pp218[35],pp218[36],pp218[37],pp218[38],pp218[39],pp218[40],pp218[41],pp218[42],pp218[43],pp218[44],pp218[45],pp218[46],pp218[47],pp219[47],pp220[47],pp221[47],pp222[47],pp223[47],pp224[47],pp225[47],pp226[47],pp227[47],pp228[47],pp229[47],pp230[47],pp231[47],pp232[47]};
    assign in105_2 = {pp219[13],pp219[14],pp219[15],pp219[16],pp219[17],pp219[18],pp219[19],pp219[20],pp219[21],pp219[22],pp219[23],pp219[24],pp219[25],pp219[26],pp219[27],pp219[28],pp219[29],pp219[30],pp219[31],pp219[32],pp219[33],pp219[34],pp219[35],pp219[36],pp219[37],pp219[38],pp219[39],pp219[40],pp219[41],pp219[42],pp219[43],pp219[44],pp219[45],pp219[46],pp220[46],pp221[46],pp222[46],pp223[46],pp224[46],pp225[46],pp226[46],pp227[46],pp228[46],pp229[46],pp230[46],pp231[46],pp232[46],pp233[46]};
    CLA_48 KS_105(s105, c105, in105_1, in105_2);
    wire[45:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp220[13],pp220[14],pp220[15],pp220[16],pp220[17],pp220[18],pp220[19],pp220[20],pp220[21],pp220[22],pp220[23],pp220[24],pp220[25],pp220[26],pp220[27],pp220[28],pp220[29],pp220[30],pp220[31],pp220[32],pp220[33],pp220[34],pp220[35],pp220[36],pp220[37],pp220[38],pp220[39],pp220[40],pp220[41],pp220[42],pp220[43],pp220[44],pp220[45],pp221[45],pp222[45],pp223[45],pp224[45],pp225[45],pp226[45],pp227[45],pp228[45],pp229[45],pp230[45],pp231[45],pp232[45],pp233[45]};
    assign in106_2 = {pp221[12],pp221[13],pp221[14],pp221[15],pp221[16],pp221[17],pp221[18],pp221[19],pp221[20],pp221[21],pp221[22],pp221[23],pp221[24],pp221[25],pp221[26],pp221[27],pp221[28],pp221[29],pp221[30],pp221[31],pp221[32],pp221[33],pp221[34],pp221[35],pp221[36],pp221[37],pp221[38],pp221[39],pp221[40],pp221[41],pp221[42],pp221[43],pp221[44],pp222[44],pp223[44],pp224[44],pp225[44],pp226[44],pp227[44],pp228[44],pp229[44],pp230[44],pp231[44],pp232[44],pp233[44],pp234[44]};
    CLA_46 KS_106(s106, c106, in106_1, in106_2);
    wire[43:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp222[12],pp222[13],pp222[14],pp222[15],pp222[16],pp222[17],pp222[18],pp222[19],pp222[20],pp222[21],pp222[22],pp222[23],pp222[24],pp222[25],pp222[26],pp222[27],pp222[28],pp222[29],pp222[30],pp222[31],pp222[32],pp222[33],pp222[34],pp222[35],pp222[36],pp222[37],pp222[38],pp222[39],pp222[40],pp222[41],pp222[42],pp222[43],pp223[43],pp224[43],pp225[43],pp226[43],pp227[43],pp228[43],pp229[43],pp230[43],pp231[43],pp232[43],pp233[43],pp234[43]};
    assign in107_2 = {pp223[11],pp223[12],pp223[13],pp223[14],pp223[15],pp223[16],pp223[17],pp223[18],pp223[19],pp223[20],pp223[21],pp223[22],pp223[23],pp223[24],pp223[25],pp223[26],pp223[27],pp223[28],pp223[29],pp223[30],pp223[31],pp223[32],pp223[33],pp223[34],pp223[35],pp223[36],pp223[37],pp223[38],pp223[39],pp223[40],pp223[41],pp223[42],pp224[42],pp225[42],pp226[42],pp227[42],pp228[42],pp229[42],pp230[42],pp231[42],pp232[42],pp233[42],pp234[42],pp235[42]};
    CLA_44 KS_107(s107, c107, in107_1, in107_2);
    wire[41:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp224[11],pp224[12],pp224[13],pp224[14],pp224[15],pp224[16],pp224[17],pp224[18],pp224[19],pp224[20],pp224[21],pp224[22],pp224[23],pp224[24],pp224[25],pp224[26],pp224[27],pp224[28],pp224[29],pp224[30],pp224[31],pp224[32],pp224[33],pp224[34],pp224[35],pp224[36],pp224[37],pp224[38],pp224[39],pp224[40],pp224[41],pp225[41],pp226[41],pp227[41],pp228[41],pp229[41],pp230[41],pp231[41],pp232[41],pp233[41],pp234[41],pp235[41]};
    assign in108_2 = {pp225[10],pp225[11],pp225[12],pp225[13],pp225[14],pp225[15],pp225[16],pp225[17],pp225[18],pp225[19],pp225[20],pp225[21],pp225[22],pp225[23],pp225[24],pp225[25],pp225[26],pp225[27],pp225[28],pp225[29],pp225[30],pp225[31],pp225[32],pp225[33],pp225[34],pp225[35],pp225[36],pp225[37],pp225[38],pp225[39],pp225[40],pp226[40],pp227[40],pp228[40],pp229[40],pp230[40],pp231[40],pp232[40],pp233[40],pp234[40],pp235[40],pp236[40]};
    CLA_42 KS_108(s108, c108, in108_1, in108_2);
    wire[39:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp226[10],pp226[11],pp226[12],pp226[13],pp226[14],pp226[15],pp226[16],pp226[17],pp226[18],pp226[19],pp226[20],pp226[21],pp226[22],pp226[23],pp226[24],pp226[25],pp226[26],pp226[27],pp226[28],pp226[29],pp226[30],pp226[31],pp226[32],pp226[33],pp226[34],pp226[35],pp226[36],pp226[37],pp226[38],pp226[39],pp227[39],pp228[39],pp229[39],pp230[39],pp231[39],pp232[39],pp233[39],pp234[39],pp235[39],pp236[39]};
    assign in109_2 = {pp0[236],pp227[10],pp227[11],pp227[12],pp227[13],pp227[14],pp227[15],pp227[16],pp227[17],pp227[18],pp227[19],pp227[20],pp227[21],pp227[22],pp227[23],pp227[24],pp227[25],pp227[26],pp227[27],pp227[28],pp227[29],pp227[30],pp227[31],pp227[32],pp227[33],pp227[34],pp227[35],pp227[36],pp227[37],pp227[38],pp228[38],pp229[38],pp230[38],pp231[38],pp232[38],pp233[38],pp234[38],pp235[38],pp236[38],pp237[38]};
    CLA_40 KS_109(s109, c109, in109_1, in109_2);
    wire[37:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp0[237],pp228[10],pp228[11],pp228[12],pp228[13],pp228[14],pp228[15],pp228[16],pp228[17],pp228[18],pp228[19],pp228[20],pp228[21],pp228[22],pp228[23],pp228[24],pp228[25],pp228[26],pp228[27],pp228[28],pp228[29],pp228[30],pp228[31],pp228[32],pp228[33],pp228[34],pp228[35],pp228[36],pp228[37],pp229[37],pp230[37],pp231[37],pp232[37],pp233[37],pp234[37],pp235[37],pp236[37],pp237[37]};
    assign in110_2 = {pp1[236],pp0[238],pp229[10],pp229[11],pp229[12],pp229[13],pp229[14],pp229[15],pp229[16],pp229[17],pp229[18],pp229[19],pp229[20],pp229[21],pp229[22],pp229[23],pp229[24],pp229[25],pp229[26],pp229[27],pp229[28],pp229[29],pp229[30],pp229[31],pp229[32],pp229[33],pp229[34],pp229[35],pp229[36],pp230[36],pp231[36],pp232[36],pp233[36],pp234[36],pp235[36],pp236[36],pp237[36],pp238[36]};
    CLA_38 KS_110(s110, c110, in110_1, in110_2);
    wire[35:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp1[237],pp0[239],pp230[10],pp230[11],pp230[12],pp230[13],pp230[14],pp230[15],pp230[16],pp230[17],pp230[18],pp230[19],pp230[20],pp230[21],pp230[22],pp230[23],pp230[24],pp230[25],pp230[26],pp230[27],pp230[28],pp230[29],pp230[30],pp230[31],pp230[32],pp230[33],pp230[34],pp230[35],pp231[35],pp232[35],pp233[35],pp234[35],pp235[35],pp236[35],pp237[35],pp238[35]};
    assign in111_2 = {pp2[236],pp1[238],pp0[240],pp231[10],pp231[11],pp231[12],pp231[13],pp231[14],pp231[15],pp231[16],pp231[17],pp231[18],pp231[19],pp231[20],pp231[21],pp231[22],pp231[23],pp231[24],pp231[25],pp231[26],pp231[27],pp231[28],pp231[29],pp231[30],pp231[31],pp231[32],pp231[33],pp231[34],pp232[34],pp233[34],pp234[34],pp235[34],pp236[34],pp237[34],pp238[34],pp239[34]};
    CLA_36 KS_111(s111, c111, in111_1, in111_2);
    wire[33:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp2[237],pp1[239],pp0[241],pp232[10],pp232[11],pp232[12],pp232[13],pp232[14],pp232[15],pp232[16],pp232[17],pp232[18],pp232[19],pp232[20],pp232[21],pp232[22],pp232[23],pp232[24],pp232[25],pp232[26],pp232[27],pp232[28],pp232[29],pp232[30],pp232[31],pp232[32],pp232[33],pp233[33],pp234[33],pp235[33],pp236[33],pp237[33],pp238[33],pp239[33]};
    assign in112_2 = {pp3[236],pp2[238],pp1[240],pp0[242],pp233[10],pp233[11],pp233[12],pp233[13],pp233[14],pp233[15],pp233[16],pp233[17],pp233[18],pp233[19],pp233[20],pp233[21],pp233[22],pp233[23],pp233[24],pp233[25],pp233[26],pp233[27],pp233[28],pp233[29],pp233[30],pp233[31],pp233[32],pp234[32],pp235[32],pp236[32],pp237[32],pp238[32],pp239[32],pp240[32]};
    CLA_34 KS_112(s112, c112, in112_1, in112_2);
    wire[31:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp3[237],pp2[239],pp1[241],pp0[243],pp234[10],pp234[11],pp234[12],pp234[13],pp234[14],pp234[15],pp234[16],pp234[17],pp234[18],pp234[19],pp234[20],pp234[21],pp234[22],pp234[23],pp234[24],pp234[25],pp234[26],pp234[27],pp234[28],pp234[29],pp234[30],pp234[31],pp235[31],pp236[31],pp237[31],pp238[31],pp239[31],pp240[31]};
    assign in113_2 = {pp4[236],pp3[238],pp2[240],pp1[242],pp0[244],pp235[10],pp235[11],pp235[12],pp235[13],pp235[14],pp235[15],pp235[16],pp235[17],pp235[18],pp235[19],pp235[20],pp235[21],pp235[22],pp235[23],pp235[24],pp235[25],pp235[26],pp235[27],pp235[28],pp235[29],pp235[30],pp236[30],pp237[30],pp238[30],pp239[30],pp240[30],pp241[30]};
    CLA_32 KS_113(s113, c113, in113_1, in113_2);
    wire[29:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp4[237],pp3[239],pp2[241],pp1[243],pp0[245],pp236[10],pp236[11],pp236[12],pp236[13],pp236[14],pp236[15],pp236[16],pp236[17],pp236[18],pp236[19],pp236[20],pp236[21],pp236[22],pp236[23],pp236[24],pp236[25],pp236[26],pp236[27],pp236[28],pp236[29],pp237[29],pp238[29],pp239[29],pp240[29],pp241[29]};
    assign in114_2 = {pp5[236],pp4[238],pp3[240],pp2[242],pp1[244],pp0[246],pp237[10],pp237[11],pp237[12],pp237[13],pp237[14],pp237[15],pp237[16],pp237[17],pp237[18],pp237[19],pp237[20],pp237[21],pp237[22],pp237[23],pp237[24],pp237[25],pp237[26],pp237[27],pp237[28],pp238[28],pp239[28],pp240[28],pp241[28],pp242[28]};
    CLA_30 KS_114(s114, c114, in114_1, in114_2);
    wire[27:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp5[237],pp4[239],pp3[241],pp2[243],pp1[245],pp0[247],pp238[10],pp238[11],pp238[12],pp238[13],pp238[14],pp238[15],pp238[16],pp238[17],pp238[18],pp238[19],pp238[20],pp238[21],pp238[22],pp238[23],pp238[24],pp238[25],pp238[26],pp238[27],pp239[27],pp240[27],pp241[27],pp242[27]};
    assign in115_2 = {pp6[236],pp5[238],pp4[240],pp3[242],pp2[244],pp1[246],pp0[248],pp239[10],pp239[11],pp239[12],pp239[13],pp239[14],pp239[15],pp239[16],pp239[17],pp239[18],pp239[19],pp239[20],pp239[21],pp239[22],pp239[23],pp239[24],pp239[25],pp239[26],pp240[26],pp241[26],pp242[26],pp243[26]};
    CLA_28 KS_115(s115, c115, in115_1, in115_2);
    wire[25:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp6[237],pp5[239],pp4[241],pp3[243],pp2[245],pp1[247],pp0[249],pp240[10],pp240[11],pp240[12],pp240[13],pp240[14],pp240[15],pp240[16],pp240[17],pp240[18],pp240[19],pp240[20],pp240[21],pp240[22],pp240[23],pp240[24],pp240[25],pp241[25],pp242[25],pp243[25]};
    assign in116_2 = {pp7[236],pp6[238],pp5[240],pp4[242],pp3[244],pp2[246],pp1[248],pp0[250],pp241[10],pp241[11],pp241[12],pp241[13],pp241[14],pp241[15],pp241[16],pp241[17],pp241[18],pp241[19],pp241[20],pp241[21],pp241[22],pp241[23],pp241[24],pp242[24],pp243[24],pp244[24]};
    CLA_26 KS_116(s116, c116, in116_1, in116_2);
    wire[23:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp7[237],pp6[239],pp5[241],pp4[243],pp3[245],pp2[247],pp1[249],pp0[251],pp242[10],pp242[11],pp242[12],pp242[13],pp242[14],pp242[15],pp242[16],pp242[17],pp242[18],pp242[19],pp242[20],pp242[21],pp242[22],pp242[23],pp243[23],pp244[23]};
    assign in117_2 = {pp8[236],pp7[238],pp6[240],pp5[242],pp4[244],pp3[246],pp2[248],pp1[250],pp0[252],pp243[10],pp243[11],pp243[12],pp243[13],pp243[14],pp243[15],pp243[16],pp243[17],pp243[18],pp243[19],pp243[20],pp243[21],pp243[22],pp244[22],pp245[22]};
    CLA_24 KS_117(s117, c117, in117_1, in117_2);
    wire[21:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp8[237],pp7[239],pp6[241],pp5[243],pp4[245],pp3[247],pp2[249],pp1[251],pp0[253],pp244[10],pp244[11],pp244[12],pp244[13],pp244[14],pp244[15],pp244[16],pp244[17],pp244[18],pp244[19],pp244[20],pp244[21],pp245[21]};
    assign in118_2 = {pp9[236],pp8[238],pp7[240],pp6[242],pp5[244],pp4[246],pp3[248],pp2[250],pp1[252],pp0[254],pp245[10],pp245[11],pp245[12],pp245[13],pp245[14],pp245[15],pp245[16],pp245[17],pp245[18],pp245[19],pp245[20],pp246[20]};
    CLA_22 KS_118(s118, c118, in118_1, in118_2);
    wire[19:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp9[237],pp8[239],pp7[241],pp6[243],pp5[245],pp4[247],pp3[249],pp2[251],pp1[253],pp0[255],pp246[10],pp246[11],pp246[12],pp246[13],pp246[14],pp246[15],pp246[16],pp246[17],pp246[18],pp246[19]};
    assign in119_2 = {pp237[9],pp9[238],pp8[240],pp7[242],pp6[244],pp5[246],pp4[248],pp3[250],pp2[252],pp1[254],pp1[255],pp247[10],pp247[11],pp247[12],pp247[13],pp247[14],pp247[15],pp247[16],pp247[17],pp247[18]};
    CLA_20 KS_119(s119, c119, in119_1, in119_2);
    wire[17:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {pp238[9],pp9[239],pp8[241],pp7[243],pp6[245],pp5[247],pp4[249],pp3[251],pp2[253],pp2[254],pp2[255],pp248[10],pp248[11],pp248[12],pp248[13],pp248[14],pp248[15],pp248[16]};
    assign in120_2 = {pp239[8],pp239[9],pp9[240],pp8[242],pp7[244],pp6[246],pp5[248],pp4[250],pp3[252],pp3[253],pp3[254],pp3[255],pp249[10],pp249[11],pp249[12],pp249[13],pp249[14],pp249[15]};
    CLA_18 KS_120(s120, c120, in120_1, in120_2);
    wire[15:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp240[8],pp240[9],pp9[241],pp8[243],pp7[245],pp6[247],pp5[249],pp4[251],pp4[252],pp4[253],pp4[254],pp4[255],pp250[10],pp250[11],pp250[12],pp250[13]};
    assign in121_2 = {pp241[7],pp241[8],pp241[9],pp9[242],pp8[244],pp7[246],pp6[248],pp5[250],pp5[251],pp5[252],pp5[253],pp5[254],pp5[255],pp251[10],pp251[11],pp251[12]};
    CLA_16 KS_121(s121, c121, in121_1, in121_2);
    wire[13:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp242[7],pp242[8],pp242[9],pp9[243],pp8[245],pp7[247],pp6[249],pp6[250],pp6[251],pp6[252],pp6[253],pp6[254],pp6[255],pp252[10]};
    assign in122_2 = {pp243[6],pp243[7],pp243[8],pp243[9],pp9[244],pp8[246],pp7[248],pp7[249],pp7[250],pp7[251],pp7[252],pp7[253],pp7[254],pp7[255]};
    CLA_14 KS_122(s122, c122, in122_1, in122_2);
    wire[11:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp244[6],pp244[7],pp244[8],pp244[9],pp9[245],pp8[247],pp8[248],pp8[249],pp8[250],pp8[251],pp8[252],pp8[253]};
    assign in123_2 = {pp245[5],pp245[6],pp245[7],pp245[8],pp245[9],pp9[246],pp9[247],pp9[248],pp9[249],pp9[250],pp9[251],pp9[252]};
    CLA_12 KS_123(s123, c123, in123_1, in123_2);
    wire[9:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp246[5],pp246[6],pp246[7],pp246[8],pp246[9],pp247[9],pp248[9],pp249[9],pp250[9],pp251[9]};
    assign in124_2 = {pp247[4],pp247[5],pp247[6],pp247[7],pp247[8],pp248[8],pp249[8],pp250[8],pp251[8],pp252[8]};
    CLA_10 KS_124(s124, c124, in124_1, in124_2);
    wire[7:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp248[4],pp248[5],pp248[6],pp248[7],pp249[7],pp250[7],pp251[7],pp252[7]};
    assign in125_2 = {pp249[3],pp249[4],pp249[5],pp249[6],pp250[6],pp251[6],pp252[6],pp253[6]};
    CLA_8 KS_125(s125, c125, in125_1, in125_2);
    wire[5:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp250[3],pp250[4],pp250[5],pp251[5],pp252[5],pp253[5]};
    assign in126_2 = {pp251[2],pp251[3],pp251[4],pp252[4],pp253[4],pp254[4]};
    CLA_6 KS_126(s126, c126, in126_1, in126_2);
    wire[3:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {pp252[2],pp252[3],pp253[3],pp254[3]};
    assign in127_2 = {pp253[1],pp253[2],pp254[2],pp255[2]};
    CLA_4 KS_127(s127, c127, in127_1, in127_2);
    wire[1:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {pp254[1],pp255[1]};
    assign in128_2 = {pp255[0],s10[119]};
    CLA_2 KS_128(s128, c128, in128_1, in128_2);

    /*Stage 2*/
    wire[383:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp10[54],pp10[55],pp10[56],pp10[57],pp10[58],pp10[59],pp10[60],pp10[61],pp10[62],pp10[63],pp10[64],pp10[65],pp10[66],pp10[67],pp10[68],pp10[69],pp10[70],pp10[71],pp10[72],pp10[73],pp10[74],pp10[75],pp10[76],pp10[77],pp10[78],pp10[79],pp10[80],pp10[81],pp10[82],pp10[83],pp10[84],pp10[85],pp10[86],pp10[87],pp10[88],pp10[89],pp0[100],pp0[101],pp0[102],pp0[103],pp0[104],pp0[105],pp0[106],pp0[107],pp0[108],pp0[109],pp10[100],pp10[101],pp10[102],pp10[103],pp10[104],pp10[105],pp10[106],pp10[107],pp10[108],pp10[109],pp10[110],pp10[111],pp10[112],pp10[113],pp10[114],pp10[115],pp10[116],pp10[117],pp12[116],pp14[115],pp16[114],pp18[113],pp20[112],pp22[111],pp24[110],pp26[109],pp28[108],pp30[107],pp32[106],pp34[105],pp36[104],pp38[103],pp40[102],pp42[101],pp44[100],pp100[45],pp101[45],pp102[45],pp103[45],pp104[45],pp105[45],pp106[45],pp107[45],pp108[45],pp109[45],pp110[45],pp111[45],pp112[45],pp113[45],pp114[45],pp115[45],pp116[45],pp117[45],pp118[45],pp119[45],pp120[45],pp121[45],pp122[45],pp123[45],pp124[45],pp125[45],pp126[45],pp127[45],pp128[45],pp129[45],pp130[45],pp131[45],pp132[45],pp133[45],pp134[45],pp135[45],pp136[45],pp137[45],pp138[45],pp139[45],pp140[45],pp141[45],pp142[45],pp143[45],pp144[45],pp145[45],pp146[45],pp147[45],pp148[45],pp149[45],pp150[45],pp151[45],pp152[45],pp153[45],pp154[45],pp156[44],pp158[43],pp160[42],pp162[41],pp164[40],pp166[39],pp168[38],pp170[37],pp172[36],pp174[35],pp176[34],pp178[33],pp180[32],pp182[31],pp184[30],pp186[29],pp188[28],pp190[27],pp192[26],pp194[25],pp196[24],pp198[23],pp200[22],pp202[21],pp204[20],pp206[19],pp208[18],pp210[17],pp212[16],pp214[15],pp216[14],pp218[13],pp220[12],pp222[11],pp224[10],pp0[235],pp1[235],pp2[235],pp3[235],pp4[235],pp5[235],pp6[235],pp7[235],pp8[235],pp9[235],pp236[9],pp238[8],pp240[7],pp242[6],pp244[5],pp246[4],pp248[3],pp250[2],pp252[1],pp254[0],s10[118],s11[118],s10[120],pp255[3],pp254[5],pp253[7],pp252[9],pp8[254],pp252[11],pp250[14],pp248[17],pp247[19],pp246[21],pp245[23],pp244[25],pp243[27],pp242[29],pp241[31],pp240[33],pp239[35],pp238[37],pp237[39],pp236[41],pp235[43],pp234[45],pp233[47],pp232[49],pp231[51],pp230[53],pp229[55],pp228[57],pp227[59],pp226[61],pp225[63],pp224[65],pp223[67],pp222[69],pp221[71],pp220[73],pp219[75],pp218[77],pp217[79],pp216[81],pp215[83],pp214[85],pp213[87],pp212[89],pp211[91],pp210[93],pp209[95],pp208[97],pp207[99],pp98[209],pp96[212],pp94[215],pp92[218],pp90[221],pp88[224],pp86[227],pp84[230],pp82[233],pp80[236],pp78[239],pp76[242],pp74[245],pp72[248],pp70[251],pp68[254],pp222[101],pp220[104],pp218[107],pp216[110],pp214[113],pp212[116],pp210[119],pp208[122],pp206[125],pp204[128],pp202[131],pp200[134],pp198[137],pp196[140],pp194[143],pp192[146],pp190[149],pp188[152],pp186[155],pp184[158],pp182[161],pp180[164],pp178[167],pp176[170],pp174[173],pp172[176],pp170[179],pp168[182],pp166[185],pp164[188],pp162[191],pp160[194],pp158[197],pp157[199],pp156[201],pp155[203],pp154[205],pp153[207],pp152[209],pp151[211],pp150[213],pp149[215],pp148[217],pp147[219],pp146[221],pp145[223],pp144[225],pp143[227],pp142[229],pp141[231],pp140[233],pp139[235],pp138[237],pp137[239],pp136[241],pp135[243],pp134[245],pp133[247],pp132[249],pp131[251],pp130[253],pp129[255],pp130[255],pp131[255],pp132[255],pp133[255],pp134[255],pp135[255],pp136[255],pp137[255],pp138[255],pp139[255],pp140[255],pp141[255],pp142[255],pp143[255],pp144[255],pp145[255],pp146[255],pp147[255],pp148[255],pp149[255],pp150[255],pp151[255],pp152[255],pp153[255],pp154[255],pp155[255],pp156[255],pp157[255],pp158[255],pp159[255],pp160[255],pp161[255],pp162[255],pp163[255],pp164[255],pp165[255],pp166[255],pp167[255],pp168[255],pp169[255],pp170[255],pp171[255],pp172[255],pp173[255],pp174[255],pp175[255],pp176[255],pp177[255],pp178[255],pp179[255],pp180[255],pp181[255],pp182[255],pp183[255],pp184[255],pp185[255],pp186[255],pp187[255],pp188[255],pp189[255],pp190[255],pp191[255],pp192[255]};
    assign in129_2 = {pp11[53],pp11[54],pp11[55],pp11[56],pp11[57],pp11[58],pp11[59],pp11[60],pp11[61],pp11[62],pp11[63],pp11[64],pp11[65],pp11[66],pp11[67],pp11[68],pp11[69],pp11[70],pp11[71],pp11[72],pp11[73],pp11[74],pp11[75],pp11[76],pp11[77],pp11[78],pp11[79],pp11[80],pp11[81],pp11[82],pp11[83],pp11[84],pp11[85],pp11[86],pp11[87],pp11[88],pp10[90],pp1[100],pp1[101],pp1[102],pp1[103],pp1[104],pp1[105],pp1[106],pp1[107],pp1[108],pp100[10],pp11[100],pp11[101],pp11[102],pp11[103],pp11[104],pp11[105],pp11[106],pp11[107],pp11[108],pp11[109],pp11[110],pp11[111],pp11[112],pp11[113],pp11[114],pp11[115],pp11[116],pp13[115],pp15[114],pp17[113],pp19[112],pp21[111],pp23[110],pp25[109],pp27[108],pp29[107],pp31[106],pp33[105],pp35[104],pp37[103],pp39[102],pp41[101],pp43[100],pp100[44],pp101[44],pp102[44],pp103[44],pp104[44],pp105[44],pp106[44],pp107[44],pp108[44],pp109[44],pp110[44],pp111[44],pp112[44],pp113[44],pp114[44],pp115[44],pp116[44],pp117[44],pp118[44],pp119[44],pp120[44],pp121[44],pp122[44],pp123[44],pp124[44],pp125[44],pp126[44],pp127[44],pp128[44],pp129[44],pp130[44],pp131[44],pp132[44],pp133[44],pp134[44],pp135[44],pp136[44],pp137[44],pp138[44],pp139[44],pp140[44],pp141[44],pp142[44],pp143[44],pp144[44],pp145[44],pp146[44],pp147[44],pp148[44],pp149[44],pp150[44],pp151[44],pp152[44],pp153[44],pp154[44],pp155[44],pp157[43],pp159[42],pp161[41],pp163[40],pp165[39],pp167[38],pp169[37],pp171[36],pp173[35],pp175[34],pp177[33],pp179[32],pp181[31],pp183[30],pp185[29],pp187[28],pp189[27],pp191[26],pp193[25],pp195[24],pp197[23],pp199[22],pp201[21],pp203[20],pp205[19],pp207[18],pp209[17],pp211[16],pp213[15],pp215[14],pp217[13],pp219[12],pp221[11],pp223[10],pp0[234],pp1[234],pp2[234],pp3[234],pp4[234],pp5[234],pp6[234],pp7[234],pp8[234],pp9[234],pp235[9],pp237[8],pp239[7],pp241[6],pp243[5],pp245[4],pp247[3],pp249[2],pp251[1],pp253[0],s10[117],s11[117],s12[117],s11[119],s10[121],pp255[4],pp254[6],pp253[8],pp9[253],pp253[10],pp251[13],pp249[16],pp248[18],pp247[20],pp246[22],pp245[24],pp244[26],pp243[28],pp242[30],pp241[32],pp240[34],pp239[36],pp238[38],pp237[40],pp236[42],pp235[44],pp234[46],pp233[48],pp232[50],pp231[52],pp230[54],pp229[56],pp228[58],pp227[60],pp226[62],pp225[64],pp224[66],pp223[68],pp222[70],pp221[72],pp220[74],pp219[76],pp218[78],pp217[80],pp216[82],pp215[84],pp214[86],pp213[88],pp212[90],pp211[92],pp210[94],pp209[96],pp208[98],pp99[208],pp97[211],pp95[214],pp93[217],pp91[220],pp89[223],pp87[226],pp85[229],pp83[232],pp81[235],pp79[238],pp77[241],pp75[244],pp73[247],pp71[250],pp69[253],pp223[100],pp221[103],pp219[106],pp217[109],pp215[112],pp213[115],pp211[118],pp209[121],pp207[124],pp205[127],pp203[130],pp201[133],pp199[136],pp197[139],pp195[142],pp193[145],pp191[148],pp189[151],pp187[154],pp185[157],pp183[160],pp181[163],pp179[166],pp177[169],pp175[172],pp173[175],pp171[178],pp169[181],pp167[184],pp165[187],pp163[190],pp161[193],pp159[196],pp158[198],pp157[200],pp156[202],pp155[204],pp154[206],pp153[208],pp152[210],pp151[212],pp150[214],pp149[216],pp148[218],pp147[220],pp146[222],pp145[224],pp144[226],pp143[228],pp142[230],pp141[232],pp140[234],pp139[236],pp138[238],pp137[240],pp136[242],pp135[244],pp134[246],pp133[248],pp132[250],pp131[252],pp130[254],pp131[254],pp132[254],pp133[254],pp134[254],pp135[254],pp136[254],pp137[254],pp138[254],pp139[254],pp140[254],pp141[254],pp142[254],pp143[254],pp144[254],pp145[254],pp146[254],pp147[254],pp148[254],pp149[254],pp150[254],pp151[254],pp152[254],pp153[254],pp154[254],pp155[254],pp156[254],pp157[254],pp158[254],pp159[254],pp160[254],pp161[254],pp162[254],pp163[254],pp164[254],pp165[254],pp166[254],pp167[254],pp168[254],pp169[254],pp170[254],pp171[254],pp172[254],pp173[254],pp174[254],pp175[254],pp176[254],pp177[254],pp178[254],pp179[254],pp180[254],pp181[254],pp182[254],pp183[254],pp184[254],pp185[254],pp186[254],pp187[254],pp188[254],pp189[254],pp190[254],pp191[254],pp192[254],pp193[254]};
    CLA_384 KS_129(s129, c129, in129_1, in129_2);
    wire[381:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp12[53],pp12[54],pp12[55],pp12[56],pp12[57],pp12[58],pp12[59],pp12[60],pp12[61],pp12[62],pp12[63],pp12[64],pp12[65],pp12[66],pp12[67],pp12[68],pp12[69],pp12[70],pp12[71],pp12[72],pp12[73],pp12[74],pp12[75],pp12[76],pp12[77],pp12[78],pp12[79],pp12[80],pp12[81],pp12[82],pp12[83],pp12[84],pp12[85],pp12[86],pp12[87],pp11[89],pp10[91],pp2[100],pp2[101],pp2[102],pp2[103],pp2[104],pp2[105],pp2[106],pp2[107],pp0[110],pp100[11],pp12[100],pp12[101],pp12[102],pp12[103],pp12[104],pp12[105],pp12[106],pp12[107],pp12[108],pp12[109],pp12[110],pp12[111],pp12[112],pp12[113],pp12[114],pp12[115],pp14[114],pp16[113],pp18[112],pp20[111],pp22[110],pp24[109],pp26[108],pp28[107],pp30[106],pp32[105],pp34[104],pp36[103],pp38[102],pp40[101],pp42[100],pp100[43],pp101[43],pp102[43],pp103[43],pp104[43],pp105[43],pp106[43],pp107[43],pp108[43],pp109[43],pp110[43],pp111[43],pp112[43],pp113[43],pp114[43],pp115[43],pp116[43],pp117[43],pp118[43],pp119[43],pp120[43],pp121[43],pp122[43],pp123[43],pp124[43],pp125[43],pp126[43],pp127[43],pp128[43],pp129[43],pp130[43],pp131[43],pp132[43],pp133[43],pp134[43],pp135[43],pp136[43],pp137[43],pp138[43],pp139[43],pp140[43],pp141[43],pp142[43],pp143[43],pp144[43],pp145[43],pp146[43],pp147[43],pp148[43],pp149[43],pp150[43],pp151[43],pp152[43],pp153[43],pp154[43],pp155[43],pp156[43],pp158[42],pp160[41],pp162[40],pp164[39],pp166[38],pp168[37],pp170[36],pp172[35],pp174[34],pp176[33],pp178[32],pp180[31],pp182[30],pp184[29],pp186[28],pp188[27],pp190[26],pp192[25],pp194[24],pp196[23],pp198[22],pp200[21],pp202[20],pp204[19],pp206[18],pp208[17],pp210[16],pp212[15],pp214[14],pp216[13],pp218[12],pp220[11],pp222[10],s129[169],s129[170],s129[171],s129[172],s129[173],s129[174],s129[175],s129[176],s129[177],s129[178],s129[179],s129[180],s129[181],s129[182],s129[183],s129[184],s129[185],s129[186],s129[187],s129[188],s129[189],s129[190],s129[191],s129[192],s129[193],s129[194],s129[195],s129[196],s129[197],s129[198],s129[199],pp252[12],pp250[15],pp249[17],pp248[19],pp247[21],pp246[23],pp245[25],pp244[27],pp243[29],pp242[31],pp241[33],pp240[35],pp239[37],pp238[39],pp237[41],pp236[43],pp235[45],pp234[47],pp233[49],pp232[51],pp231[53],pp230[55],pp229[57],pp228[59],pp227[61],pp226[63],pp225[65],pp224[67],pp223[69],pp222[71],pp221[73],pp220[75],pp219[77],pp218[79],pp217[81],pp216[83],pp215[85],pp214[87],pp213[89],pp212[91],pp211[93],pp210[95],pp209[97],pp208[99],pp98[210],pp96[213],pp94[216],pp92[219],pp90[222],pp88[225],pp86[228],pp84[231],pp82[234],pp80[237],pp78[240],pp76[243],pp74[246],pp72[249],pp70[252],pp68[255],pp222[102],pp220[105],pp218[108],pp216[111],pp214[114],pp212[117],pp210[120],pp208[123],pp206[126],pp204[129],pp202[132],pp200[135],pp198[138],pp196[141],pp194[144],pp192[147],pp190[150],pp188[153],pp186[156],pp184[159],pp182[162],pp180[165],pp178[168],pp176[171],pp174[174],pp172[177],pp170[180],pp168[183],pp166[186],pp164[189],pp162[192],pp160[195],pp159[197],pp158[199],pp157[201],pp156[203],pp155[205],pp154[207],pp153[209],pp152[211],pp151[213],pp150[215],pp149[217],pp148[219],pp147[221],pp146[223],pp145[225],pp144[227],pp143[229],pp142[231],pp141[233],pp140[235],pp139[237],pp138[239],pp137[241],pp136[243],pp135[245],pp134[247],pp133[249],pp132[251],pp131[253],pp132[253],pp133[253],pp134[253],pp135[253],pp136[253],pp137[253],pp138[253],pp139[253],pp140[253],pp141[253],pp142[253],pp143[253],pp144[253],pp145[253],pp146[253],pp147[253],pp148[253],pp149[253],pp150[253],pp151[253],pp152[253],pp153[253],pp154[253],pp155[253],pp156[253],pp157[253],pp158[253],pp159[253],pp160[253],pp161[253],pp162[253],pp163[253],pp164[253],pp165[253],pp166[253],pp167[253],pp168[253],pp169[253],pp170[253],pp171[253],pp172[253],pp173[253],pp174[253],pp175[253],pp176[253],pp177[253],pp178[253],pp179[253],pp180[253],pp181[253],pp182[253],pp183[253],pp184[253],pp185[253],pp186[253],pp187[253],pp188[253],pp189[253],pp190[253],pp191[253],pp192[253],pp193[253]};
    assign in130_2 = {pp13[52],pp13[53],pp13[54],pp13[55],pp13[56],pp13[57],pp13[58],pp13[59],pp13[60],pp13[61],pp13[62],pp13[63],pp13[64],pp13[65],pp13[66],pp13[67],pp13[68],pp13[69],pp13[70],pp13[71],pp13[72],pp13[73],pp13[74],pp13[75],pp13[76],pp13[77],pp13[78],pp13[79],pp13[80],pp13[81],pp13[82],pp13[83],pp13[84],pp13[85],pp13[86],pp12[88],pp11[90],pp10[92],pp3[100],pp3[101],pp3[102],pp3[103],pp3[104],pp3[105],pp3[106],pp1[109],pp101[10],pp100[12],pp13[100],pp13[101],pp13[102],pp13[103],pp13[104],pp13[105],pp13[106],pp13[107],pp13[108],pp13[109],pp13[110],pp13[111],pp13[112],pp13[113],pp13[114],pp15[113],pp17[112],pp19[111],pp21[110],pp23[109],pp25[108],pp27[107],pp29[106],pp31[105],pp33[104],pp35[103],pp37[102],pp39[101],pp41[100],pp100[42],pp101[42],pp102[42],pp103[42],pp104[42],pp105[42],pp106[42],pp107[42],pp108[42],pp109[42],pp110[42],pp111[42],pp112[42],pp113[42],pp114[42],pp115[42],pp116[42],pp117[42],pp118[42],pp119[42],pp120[42],pp121[42],pp122[42],pp123[42],pp124[42],pp125[42],pp126[42],pp127[42],pp128[42],pp129[42],pp130[42],pp131[42],pp132[42],pp133[42],pp134[42],pp135[42],pp136[42],pp137[42],pp138[42],pp139[42],pp140[42],pp141[42],pp142[42],pp143[42],pp144[42],pp145[42],pp146[42],pp147[42],pp148[42],pp149[42],pp150[42],pp151[42],pp152[42],pp153[42],pp154[42],pp155[42],pp156[42],pp157[42],pp159[41],pp161[40],pp163[39],pp165[38],pp167[37],pp169[36],pp171[35],pp173[34],pp175[33],pp177[32],pp179[31],pp181[30],pp183[29],pp185[28],pp187[27],pp189[26],pp191[25],pp193[24],pp195[23],pp197[22],pp199[21],pp201[20],pp203[19],pp205[18],pp207[17],pp209[16],pp211[15],pp213[14],pp215[13],pp217[12],pp219[11],pp221[10],s129[168],pp0[233],pp1[233],pp2[233],pp3[233],pp4[233],pp5[233],pp6[233],pp7[233],pp8[233],pp9[233],pp234[9],pp236[8],pp238[7],pp240[6],pp242[5],pp244[4],pp246[3],pp248[2],pp250[1],pp252[0],s10[116],s11[116],s12[116],s13[116],s12[118],s11[120],s10[122],pp255[5],pp254[7],pp253[9],pp8[255],pp253[11],pp251[14],pp250[16],pp249[18],pp248[20],pp247[22],pp246[24],pp245[26],pp244[28],pp243[30],pp242[32],pp241[34],pp240[36],pp239[38],pp238[40],pp237[42],pp236[44],pp235[46],pp234[48],pp233[50],pp232[52],pp231[54],pp230[56],pp229[58],pp228[60],pp227[62],pp226[64],pp225[66],pp224[68],pp223[70],pp222[72],pp221[74],pp220[76],pp219[78],pp218[80],pp217[82],pp216[84],pp215[86],pp214[88],pp213[90],pp212[92],pp211[94],pp210[96],pp209[98],pp99[209],pp97[212],pp95[215],pp93[218],pp91[221],pp89[224],pp87[227],pp85[230],pp83[233],pp81[236],pp79[239],pp77[242],pp75[245],pp73[248],pp71[251],pp69[254],pp223[101],pp221[104],pp219[107],pp217[110],pp215[113],pp213[116],pp211[119],pp209[122],pp207[125],pp205[128],pp203[131],pp201[134],pp199[137],pp197[140],pp195[143],pp193[146],pp191[149],pp189[152],pp187[155],pp185[158],pp183[161],pp181[164],pp179[167],pp177[170],pp175[173],pp173[176],pp171[179],pp169[182],pp167[185],pp165[188],pp163[191],pp161[194],pp160[196],pp159[198],pp158[200],pp157[202],pp156[204],pp155[206],pp154[208],pp153[210],pp152[212],pp151[214],pp150[216],pp149[218],pp148[220],pp147[222],pp146[224],pp145[226],pp144[228],pp143[230],pp142[232],pp141[234],pp140[236],pp139[238],pp138[240],pp137[242],pp136[244],pp135[246],pp134[248],pp133[250],pp132[252],pp133[252],pp134[252],pp135[252],pp136[252],pp137[252],pp138[252],pp139[252],pp140[252],pp141[252],pp142[252],pp143[252],pp144[252],pp145[252],pp146[252],pp147[252],pp148[252],pp149[252],pp150[252],pp151[252],pp152[252],pp153[252],pp154[252],pp155[252],pp156[252],pp157[252],pp158[252],pp159[252],pp160[252],pp161[252],pp162[252],pp163[252],pp164[252],pp165[252],pp166[252],pp167[252],pp168[252],pp169[252],pp170[252],pp171[252],pp172[252],pp173[252],pp174[252],pp175[252],pp176[252],pp177[252],pp178[252],pp179[252],pp180[252],pp181[252],pp182[252],pp183[252],pp184[252],pp185[252],pp186[252],pp187[252],pp188[252],pp189[252],pp190[252],pp191[252],pp192[252],pp193[252],pp194[252]};
    CLA_382 KS_130(s130, c130, in130_1, in130_2);
    wire[379:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp14[52],pp14[53],pp14[54],pp14[55],pp14[56],pp14[57],pp14[58],pp14[59],pp14[60],pp14[61],pp14[62],pp14[63],pp14[64],pp14[65],pp14[66],pp14[67],pp14[68],pp14[69],pp14[70],pp14[71],pp14[72],pp14[73],pp14[74],pp14[75],pp14[76],pp14[77],pp14[78],pp14[79],pp14[80],pp14[81],pp14[82],pp14[83],pp14[84],pp14[85],pp13[87],pp12[89],pp11[91],pp10[93],pp4[100],pp4[101],pp4[102],pp4[103],pp4[104],pp4[105],pp2[108],pp0[111],pp101[11],pp100[13],pp14[100],pp14[101],pp14[102],pp14[103],pp14[104],pp14[105],pp14[106],pp14[107],pp14[108],pp14[109],pp14[110],pp14[111],pp14[112],pp14[113],pp16[112],pp18[111],pp20[110],pp22[109],pp24[108],pp26[107],pp28[106],pp30[105],pp32[104],pp34[103],pp36[102],pp38[101],pp40[100],pp100[41],pp101[41],pp102[41],pp103[41],pp104[41],pp105[41],pp106[41],pp107[41],pp108[41],pp109[41],pp110[41],pp111[41],pp112[41],pp113[41],pp114[41],pp115[41],pp116[41],pp117[41],pp118[41],pp119[41],pp120[41],pp121[41],pp122[41],pp123[41],pp124[41],pp125[41],pp126[41],pp127[41],pp128[41],pp129[41],pp130[41],pp131[41],pp132[41],pp133[41],pp134[41],pp135[41],pp136[41],pp137[41],pp138[41],pp139[41],pp140[41],pp141[41],pp142[41],pp143[41],pp144[41],pp145[41],pp146[41],pp147[41],pp148[41],pp149[41],pp150[41],pp151[41],pp152[41],pp153[41],pp154[41],pp155[41],pp156[41],pp157[41],pp158[41],pp160[40],pp162[39],pp164[38],pp166[37],pp168[36],pp170[35],pp172[34],pp174[33],pp176[32],pp178[31],pp180[30],pp182[29],pp184[28],pp186[27],pp188[26],pp190[25],pp192[24],pp194[23],pp196[22],pp198[21],pp200[20],pp202[19],pp204[18],pp206[17],pp208[16],pp210[15],pp212[14],pp214[13],pp216[12],pp218[11],pp220[10],s129[167],s130[167],s130[168],s130[169],s130[170],s130[171],s130[172],s130[173],s130[174],s130[175],s130[176],s130[177],s130[178],s130[179],s130[180],s130[181],s130[182],s130[183],s130[184],s130[185],s130[186],s130[187],s130[188],s130[189],s130[190],s130[191],s130[192],s130[193],s130[194],s130[195],s130[196],s130[197],s130[198],pp254[10],pp252[13],pp251[15],pp250[17],pp249[19],pp248[21],pp247[23],pp246[25],pp245[27],pp244[29],pp243[31],pp242[33],pp241[35],pp240[37],pp239[39],pp238[41],pp237[43],pp236[45],pp235[47],pp234[49],pp233[51],pp232[53],pp231[55],pp230[57],pp229[59],pp228[61],pp227[63],pp226[65],pp225[67],pp224[69],pp223[71],pp222[73],pp221[75],pp220[77],pp219[79],pp218[81],pp217[83],pp216[85],pp215[87],pp214[89],pp213[91],pp212[93],pp211[95],pp210[97],pp209[99],pp98[211],pp96[214],pp94[217],pp92[220],pp90[223],pp88[226],pp86[229],pp84[232],pp82[235],pp80[238],pp78[241],pp76[244],pp74[247],pp72[250],pp70[253],pp224[100],pp222[103],pp220[106],pp218[109],pp216[112],pp214[115],pp212[118],pp210[121],pp208[124],pp206[127],pp204[130],pp202[133],pp200[136],pp198[139],pp196[142],pp194[145],pp192[148],pp190[151],pp188[154],pp186[157],pp184[160],pp182[163],pp180[166],pp178[169],pp176[172],pp174[175],pp172[178],pp170[181],pp168[184],pp166[187],pp164[190],pp162[193],pp161[195],pp160[197],pp159[199],pp158[201],pp157[203],pp156[205],pp155[207],pp154[209],pp153[211],pp152[213],pp151[215],pp150[217],pp149[219],pp148[221],pp147[223],pp146[225],pp145[227],pp144[229],pp143[231],pp142[233],pp141[235],pp140[237],pp139[239],pp138[241],pp137[243],pp136[245],pp135[247],pp134[249],pp133[251],pp134[251],pp135[251],pp136[251],pp137[251],pp138[251],pp139[251],pp140[251],pp141[251],pp142[251],pp143[251],pp144[251],pp145[251],pp146[251],pp147[251],pp148[251],pp149[251],pp150[251],pp151[251],pp152[251],pp153[251],pp154[251],pp155[251],pp156[251],pp157[251],pp158[251],pp159[251],pp160[251],pp161[251],pp162[251],pp163[251],pp164[251],pp165[251],pp166[251],pp167[251],pp168[251],pp169[251],pp170[251],pp171[251],pp172[251],pp173[251],pp174[251],pp175[251],pp176[251],pp177[251],pp178[251],pp179[251],pp180[251],pp181[251],pp182[251],pp183[251],pp184[251],pp185[251],pp186[251],pp187[251],pp188[251],pp189[251],pp190[251],pp191[251],pp192[251],pp193[251],pp194[251]};
    assign in131_2 = {pp15[51],pp15[52],pp15[53],pp15[54],pp15[55],pp15[56],pp15[57],pp15[58],pp15[59],pp15[60],pp15[61],pp15[62],pp15[63],pp15[64],pp15[65],pp15[66],pp15[67],pp15[68],pp15[69],pp15[70],pp15[71],pp15[72],pp15[73],pp15[74],pp15[75],pp15[76],pp15[77],pp15[78],pp15[79],pp15[80],pp15[81],pp15[82],pp15[83],pp15[84],pp14[86],pp13[88],pp12[90],pp11[92],pp10[94],pp5[100],pp5[101],pp5[102],pp5[103],pp5[104],pp3[107],pp1[110],pp102[10],pp101[12],pp100[14],pp15[100],pp15[101],pp15[102],pp15[103],pp15[104],pp15[105],pp15[106],pp15[107],pp15[108],pp15[109],pp15[110],pp15[111],pp15[112],pp17[111],pp19[110],pp21[109],pp23[108],pp25[107],pp27[106],pp29[105],pp31[104],pp33[103],pp35[102],pp37[101],pp39[100],pp100[40],pp101[40],pp102[40],pp103[40],pp104[40],pp105[40],pp106[40],pp107[40],pp108[40],pp109[40],pp110[40],pp111[40],pp112[40],pp113[40],pp114[40],pp115[40],pp116[40],pp117[40],pp118[40],pp119[40],pp120[40],pp121[40],pp122[40],pp123[40],pp124[40],pp125[40],pp126[40],pp127[40],pp128[40],pp129[40],pp130[40],pp131[40],pp132[40],pp133[40],pp134[40],pp135[40],pp136[40],pp137[40],pp138[40],pp139[40],pp140[40],pp141[40],pp142[40],pp143[40],pp144[40],pp145[40],pp146[40],pp147[40],pp148[40],pp149[40],pp150[40],pp151[40],pp152[40],pp153[40],pp154[40],pp155[40],pp156[40],pp157[40],pp158[40],pp159[40],pp161[39],pp163[38],pp165[37],pp167[36],pp169[35],pp171[34],pp173[33],pp175[32],pp177[31],pp179[30],pp181[29],pp183[28],pp185[27],pp187[26],pp189[25],pp191[24],pp193[23],pp195[22],pp197[21],pp199[20],pp201[19],pp203[18],pp205[17],pp207[16],pp209[15],pp211[14],pp213[13],pp215[12],pp217[11],pp219[10],s129[166],s130[166],pp0[232],pp1[232],pp2[232],pp3[232],pp4[232],pp5[232],pp6[232],pp7[232],pp8[232],pp9[232],pp233[9],pp235[8],pp237[7],pp239[6],pp241[5],pp243[4],pp245[3],pp247[2],pp249[1],pp251[0],s10[115],s11[115],s12[115],s13[115],s14[115],s13[117],s12[119],s11[121],s10[123],pp255[6],pp254[8],pp9[254],s129[200],pp253[12],pp252[14],pp251[16],pp250[18],pp249[20],pp248[22],pp247[24],pp246[26],pp245[28],pp244[30],pp243[32],pp242[34],pp241[36],pp240[38],pp239[40],pp238[42],pp237[44],pp236[46],pp235[48],pp234[50],pp233[52],pp232[54],pp231[56],pp230[58],pp229[60],pp228[62],pp227[64],pp226[66],pp225[68],pp224[70],pp223[72],pp222[74],pp221[76],pp220[78],pp219[80],pp218[82],pp217[84],pp216[86],pp215[88],pp214[90],pp213[92],pp212[94],pp211[96],pp210[98],pp99[210],pp97[213],pp95[216],pp93[219],pp91[222],pp89[225],pp87[228],pp85[231],pp83[234],pp81[237],pp79[240],pp77[243],pp75[246],pp73[249],pp71[252],pp69[255],pp223[102],pp221[105],pp219[108],pp217[111],pp215[114],pp213[117],pp211[120],pp209[123],pp207[126],pp205[129],pp203[132],pp201[135],pp199[138],pp197[141],pp195[144],pp193[147],pp191[150],pp189[153],pp187[156],pp185[159],pp183[162],pp181[165],pp179[168],pp177[171],pp175[174],pp173[177],pp171[180],pp169[183],pp167[186],pp165[189],pp163[192],pp162[194],pp161[196],pp160[198],pp159[200],pp158[202],pp157[204],pp156[206],pp155[208],pp154[210],pp153[212],pp152[214],pp151[216],pp150[218],pp149[220],pp148[222],pp147[224],pp146[226],pp145[228],pp144[230],pp143[232],pp142[234],pp141[236],pp140[238],pp139[240],pp138[242],pp137[244],pp136[246],pp135[248],pp134[250],pp135[250],pp136[250],pp137[250],pp138[250],pp139[250],pp140[250],pp141[250],pp142[250],pp143[250],pp144[250],pp145[250],pp146[250],pp147[250],pp148[250],pp149[250],pp150[250],pp151[250],pp152[250],pp153[250],pp154[250],pp155[250],pp156[250],pp157[250],pp158[250],pp159[250],pp160[250],pp161[250],pp162[250],pp163[250],pp164[250],pp165[250],pp166[250],pp167[250],pp168[250],pp169[250],pp170[250],pp171[250],pp172[250],pp173[250],pp174[250],pp175[250],pp176[250],pp177[250],pp178[250],pp179[250],pp180[250],pp181[250],pp182[250],pp183[250],pp184[250],pp185[250],pp186[250],pp187[250],pp188[250],pp189[250],pp190[250],pp191[250],pp192[250],pp193[250],pp194[250],pp195[250]};
    CLA_380 KS_131(s131, c131, in131_1, in131_2);
    wire[377:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp16[51],pp16[52],pp16[53],pp16[54],pp16[55],pp16[56],pp16[57],pp16[58],pp16[59],pp16[60],pp16[61],pp16[62],pp16[63],pp16[64],pp16[65],pp16[66],pp16[67],pp16[68],pp16[69],pp16[70],pp16[71],pp16[72],pp16[73],pp16[74],pp16[75],pp16[76],pp16[77],pp16[78],pp16[79],pp16[80],pp16[81],pp16[82],pp16[83],pp15[85],pp14[87],pp13[89],pp12[91],pp11[93],pp10[95],pp6[100],pp6[101],pp6[102],pp6[103],pp4[106],pp2[109],pp0[112],pp102[11],pp101[13],pp100[15],pp16[100],pp16[101],pp16[102],pp16[103],pp16[104],pp16[105],pp16[106],pp16[107],pp16[108],pp16[109],pp16[110],pp16[111],pp18[110],pp20[109],pp22[108],pp24[107],pp26[106],pp28[105],pp30[104],pp32[103],pp34[102],pp36[101],pp38[100],pp100[39],pp101[39],pp102[39],pp103[39],pp104[39],pp105[39],pp106[39],pp107[39],pp108[39],pp109[39],pp110[39],pp111[39],pp112[39],pp113[39],pp114[39],pp115[39],pp116[39],pp117[39],pp118[39],pp119[39],pp120[39],pp121[39],pp122[39],pp123[39],pp124[39],pp125[39],pp126[39],pp127[39],pp128[39],pp129[39],pp130[39],pp131[39],pp132[39],pp133[39],pp134[39],pp135[39],pp136[39],pp137[39],pp138[39],pp139[39],pp140[39],pp141[39],pp142[39],pp143[39],pp144[39],pp145[39],pp146[39],pp147[39],pp148[39],pp149[39],pp150[39],pp151[39],pp152[39],pp153[39],pp154[39],pp155[39],pp156[39],pp157[39],pp158[39],pp159[39],pp160[39],pp162[38],pp164[37],pp166[36],pp168[35],pp170[34],pp172[33],pp174[32],pp176[31],pp178[30],pp180[29],pp182[28],pp184[27],pp186[26],pp188[25],pp190[24],pp192[23],pp194[22],pp196[21],pp198[20],pp200[19],pp202[18],pp204[17],pp206[16],pp208[15],pp210[14],pp212[13],pp214[12],pp216[11],pp218[10],s129[165],s130[165],s131[165],s131[166],s131[167],s131[168],s131[169],s131[170],s131[171],s131[172],s131[173],s131[174],s131[175],s131[176],s131[177],s131[178],s131[179],s131[180],s131[181],s131[182],s131[183],s131[184],s131[185],s131[186],s131[187],s131[188],s131[189],s131[190],s131[191],s131[192],s131[193],s131[194],s131[195],s131[196],s131[197],s130[199],pp254[11],pp253[13],pp252[15],pp251[17],pp250[19],pp249[21],pp248[23],pp247[25],pp246[27],pp245[29],pp244[31],pp243[33],pp242[35],pp241[37],pp240[39],pp239[41],pp238[43],pp237[45],pp236[47],pp235[49],pp234[51],pp233[53],pp232[55],pp231[57],pp230[59],pp229[61],pp228[63],pp227[65],pp226[67],pp225[69],pp224[71],pp223[73],pp222[75],pp221[77],pp220[79],pp219[81],pp218[83],pp217[85],pp216[87],pp215[89],pp214[91],pp213[93],pp212[95],pp211[97],pp210[99],pp98[212],pp96[215],pp94[218],pp92[221],pp90[224],pp88[227],pp86[230],pp84[233],pp82[236],pp80[239],pp78[242],pp76[245],pp74[248],pp72[251],pp70[254],pp224[101],pp222[104],pp220[107],pp218[110],pp216[113],pp214[116],pp212[119],pp210[122],pp208[125],pp206[128],pp204[131],pp202[134],pp200[137],pp198[140],pp196[143],pp194[146],pp192[149],pp190[152],pp188[155],pp186[158],pp184[161],pp182[164],pp180[167],pp178[170],pp176[173],pp174[176],pp172[179],pp170[182],pp168[185],pp166[188],pp164[191],pp163[193],pp162[195],pp161[197],pp160[199],pp159[201],pp158[203],pp157[205],pp156[207],pp155[209],pp154[211],pp153[213],pp152[215],pp151[217],pp150[219],pp149[221],pp148[223],pp147[225],pp146[227],pp145[229],pp144[231],pp143[233],pp142[235],pp141[237],pp140[239],pp139[241],pp138[243],pp137[245],pp136[247],pp135[249],pp136[249],pp137[249],pp138[249],pp139[249],pp140[249],pp141[249],pp142[249],pp143[249],pp144[249],pp145[249],pp146[249],pp147[249],pp148[249],pp149[249],pp150[249],pp151[249],pp152[249],pp153[249],pp154[249],pp155[249],pp156[249],pp157[249],pp158[249],pp159[249],pp160[249],pp161[249],pp162[249],pp163[249],pp164[249],pp165[249],pp166[249],pp167[249],pp168[249],pp169[249],pp170[249],pp171[249],pp172[249],pp173[249],pp174[249],pp175[249],pp176[249],pp177[249],pp178[249],pp179[249],pp180[249],pp181[249],pp182[249],pp183[249],pp184[249],pp185[249],pp186[249],pp187[249],pp188[249],pp189[249],pp190[249],pp191[249],pp192[249],pp193[249],pp194[249],pp195[249]};
    assign in132_2 = {pp17[50],pp17[51],pp17[52],pp17[53],pp17[54],pp17[55],pp17[56],pp17[57],pp17[58],pp17[59],pp17[60],pp17[61],pp17[62],pp17[63],pp17[64],pp17[65],pp17[66],pp17[67],pp17[68],pp17[69],pp17[70],pp17[71],pp17[72],pp17[73],pp17[74],pp17[75],pp17[76],pp17[77],pp17[78],pp17[79],pp17[80],pp17[81],pp17[82],pp16[84],pp15[86],pp14[88],pp13[90],pp12[92],pp11[94],pp10[96],pp7[100],pp7[101],pp7[102],pp5[105],pp3[108],pp1[111],pp103[10],pp102[12],pp101[14],pp100[16],pp17[100],pp17[101],pp17[102],pp17[103],pp17[104],pp17[105],pp17[106],pp17[107],pp17[108],pp17[109],pp17[110],pp19[109],pp21[108],pp23[107],pp25[106],pp27[105],pp29[104],pp31[103],pp33[102],pp35[101],pp37[100],pp100[38],pp101[38],pp102[38],pp103[38],pp104[38],pp105[38],pp106[38],pp107[38],pp108[38],pp109[38],pp110[38],pp111[38],pp112[38],pp113[38],pp114[38],pp115[38],pp116[38],pp117[38],pp118[38],pp119[38],pp120[38],pp121[38],pp122[38],pp123[38],pp124[38],pp125[38],pp126[38],pp127[38],pp128[38],pp129[38],pp130[38],pp131[38],pp132[38],pp133[38],pp134[38],pp135[38],pp136[38],pp137[38],pp138[38],pp139[38],pp140[38],pp141[38],pp142[38],pp143[38],pp144[38],pp145[38],pp146[38],pp147[38],pp148[38],pp149[38],pp150[38],pp151[38],pp152[38],pp153[38],pp154[38],pp155[38],pp156[38],pp157[38],pp158[38],pp159[38],pp160[38],pp161[38],pp163[37],pp165[36],pp167[35],pp169[34],pp171[33],pp173[32],pp175[31],pp177[30],pp179[29],pp181[28],pp183[27],pp185[26],pp187[25],pp189[24],pp191[23],pp193[22],pp195[21],pp197[20],pp199[19],pp201[18],pp203[17],pp205[16],pp207[15],pp209[14],pp211[13],pp213[12],pp215[11],pp217[10],s129[164],s130[164],s131[164],pp0[231],pp1[231],pp2[231],pp3[231],pp4[231],pp5[231],pp6[231],pp7[231],pp8[231],pp9[231],pp232[9],pp234[8],pp236[7],pp238[6],pp240[5],pp242[4],pp244[3],pp246[2],pp248[1],pp250[0],s10[114],s11[114],s12[114],s13[114],s14[114],s15[114],s14[116],s13[118],s12[120],s11[122],s10[124],pp255[7],pp254[9],s131[198],pp255[10],pp254[12],pp253[14],pp252[16],pp251[18],pp250[20],pp249[22],pp248[24],pp247[26],pp246[28],pp245[30],pp244[32],pp243[34],pp242[36],pp241[38],pp240[40],pp239[42],pp238[44],pp237[46],pp236[48],pp235[50],pp234[52],pp233[54],pp232[56],pp231[58],pp230[60],pp229[62],pp228[64],pp227[66],pp226[68],pp225[70],pp224[72],pp223[74],pp222[76],pp221[78],pp220[80],pp219[82],pp218[84],pp217[86],pp216[88],pp215[90],pp214[92],pp213[94],pp212[96],pp211[98],pp99[211],pp97[214],pp95[217],pp93[220],pp91[223],pp89[226],pp87[229],pp85[232],pp83[235],pp81[238],pp79[241],pp77[244],pp75[247],pp73[250],pp71[253],pp225[100],pp223[103],pp221[106],pp219[109],pp217[112],pp215[115],pp213[118],pp211[121],pp209[124],pp207[127],pp205[130],pp203[133],pp201[136],pp199[139],pp197[142],pp195[145],pp193[148],pp191[151],pp189[154],pp187[157],pp185[160],pp183[163],pp181[166],pp179[169],pp177[172],pp175[175],pp173[178],pp171[181],pp169[184],pp167[187],pp165[190],pp164[192],pp163[194],pp162[196],pp161[198],pp160[200],pp159[202],pp158[204],pp157[206],pp156[208],pp155[210],pp154[212],pp153[214],pp152[216],pp151[218],pp150[220],pp149[222],pp148[224],pp147[226],pp146[228],pp145[230],pp144[232],pp143[234],pp142[236],pp141[238],pp140[240],pp139[242],pp138[244],pp137[246],pp136[248],pp137[248],pp138[248],pp139[248],pp140[248],pp141[248],pp142[248],pp143[248],pp144[248],pp145[248],pp146[248],pp147[248],pp148[248],pp149[248],pp150[248],pp151[248],pp152[248],pp153[248],pp154[248],pp155[248],pp156[248],pp157[248],pp158[248],pp159[248],pp160[248],pp161[248],pp162[248],pp163[248],pp164[248],pp165[248],pp166[248],pp167[248],pp168[248],pp169[248],pp170[248],pp171[248],pp172[248],pp173[248],pp174[248],pp175[248],pp176[248],pp177[248],pp178[248],pp179[248],pp180[248],pp181[248],pp182[248],pp183[248],pp184[248],pp185[248],pp186[248],pp187[248],pp188[248],pp189[248],pp190[248],pp191[248],pp192[248],pp193[248],pp194[248],pp195[248],pp196[248]};
    CLA_378 KS_132(s132, c132, in132_1, in132_2);
    wire[375:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp18[50],pp18[51],pp18[52],pp18[53],pp18[54],pp18[55],pp18[56],pp18[57],pp18[58],pp18[59],pp18[60],pp18[61],pp18[62],pp18[63],pp18[64],pp18[65],pp18[66],pp18[67],pp18[68],pp18[69],pp18[70],pp18[71],pp18[72],pp18[73],pp18[74],pp18[75],pp18[76],pp18[77],pp18[78],pp18[79],pp18[80],pp18[81],pp17[83],pp16[85],pp15[87],pp14[89],pp13[91],pp12[93],pp11[95],pp10[97],pp8[100],pp8[101],pp6[104],pp4[107],pp2[110],pp0[113],pp103[11],pp102[13],pp101[15],pp100[17],pp18[100],pp18[101],pp18[102],pp18[103],pp18[104],pp18[105],pp18[106],pp18[107],pp18[108],pp18[109],pp20[108],pp22[107],pp24[106],pp26[105],pp28[104],pp30[103],pp32[102],pp34[101],pp36[100],pp100[37],pp101[37],pp102[37],pp103[37],pp104[37],pp105[37],pp106[37],pp107[37],pp108[37],pp109[37],pp110[37],pp111[37],pp112[37],pp113[37],pp114[37],pp115[37],pp116[37],pp117[37],pp118[37],pp119[37],pp120[37],pp121[37],pp122[37],pp123[37],pp124[37],pp125[37],pp126[37],pp127[37],pp128[37],pp129[37],pp130[37],pp131[37],pp132[37],pp133[37],pp134[37],pp135[37],pp136[37],pp137[37],pp138[37],pp139[37],pp140[37],pp141[37],pp142[37],pp143[37],pp144[37],pp145[37],pp146[37],pp147[37],pp148[37],pp149[37],pp150[37],pp151[37],pp152[37],pp153[37],pp154[37],pp155[37],pp156[37],pp157[37],pp158[37],pp159[37],pp160[37],pp161[37],pp162[37],pp164[36],pp166[35],pp168[34],pp170[33],pp172[32],pp174[31],pp176[30],pp178[29],pp180[28],pp182[27],pp184[26],pp186[25],pp188[24],pp190[23],pp192[22],pp194[21],pp196[20],pp198[19],pp200[18],pp202[17],pp204[16],pp206[15],pp208[14],pp210[13],pp212[12],pp214[11],pp216[10],s129[163],s130[163],s131[163],s132[163],s132[164],s132[165],s132[166],s132[167],s132[168],s132[169],s132[170],s132[171],s132[172],s132[173],s132[174],s132[175],s132[176],s132[177],s132[178],s132[179],s132[180],s132[181],s132[182],s132[183],s132[184],s132[185],s132[186],s132[187],s132[188],s132[189],s132[190],s132[191],s132[192],s132[193],s132[194],s132[195],s132[196],s132[197],s129[201],pp255[11],pp254[13],pp253[15],pp252[17],pp251[19],pp250[21],pp249[23],pp248[25],pp247[27],pp246[29],pp245[31],pp244[33],pp243[35],pp242[37],pp241[39],pp240[41],pp239[43],pp238[45],pp237[47],pp236[49],pp235[51],pp234[53],pp233[55],pp232[57],pp231[59],pp230[61],pp229[63],pp228[65],pp227[67],pp226[69],pp225[71],pp224[73],pp223[75],pp222[77],pp221[79],pp220[81],pp219[83],pp218[85],pp217[87],pp216[89],pp215[91],pp214[93],pp213[95],pp212[97],pp211[99],pp98[213],pp96[216],pp94[219],pp92[222],pp90[225],pp88[228],pp86[231],pp84[234],pp82[237],pp80[240],pp78[243],pp76[246],pp74[249],pp72[252],pp70[255],pp224[102],pp222[105],pp220[108],pp218[111],pp216[114],pp214[117],pp212[120],pp210[123],pp208[126],pp206[129],pp204[132],pp202[135],pp200[138],pp198[141],pp196[144],pp194[147],pp192[150],pp190[153],pp188[156],pp186[159],pp184[162],pp182[165],pp180[168],pp178[171],pp176[174],pp174[177],pp172[180],pp170[183],pp168[186],pp166[189],pp165[191],pp164[193],pp163[195],pp162[197],pp161[199],pp160[201],pp159[203],pp158[205],pp157[207],pp156[209],pp155[211],pp154[213],pp153[215],pp152[217],pp151[219],pp150[221],pp149[223],pp148[225],pp147[227],pp146[229],pp145[231],pp144[233],pp143[235],pp142[237],pp141[239],pp140[241],pp139[243],pp138[245],pp137[247],pp138[247],pp139[247],pp140[247],pp141[247],pp142[247],pp143[247],pp144[247],pp145[247],pp146[247],pp147[247],pp148[247],pp149[247],pp150[247],pp151[247],pp152[247],pp153[247],pp154[247],pp155[247],pp156[247],pp157[247],pp158[247],pp159[247],pp160[247],pp161[247],pp162[247],pp163[247],pp164[247],pp165[247],pp166[247],pp167[247],pp168[247],pp169[247],pp170[247],pp171[247],pp172[247],pp173[247],pp174[247],pp175[247],pp176[247],pp177[247],pp178[247],pp179[247],pp180[247],pp181[247],pp182[247],pp183[247],pp184[247],pp185[247],pp186[247],pp187[247],pp188[247],pp189[247],pp190[247],pp191[247],pp192[247],pp193[247],pp194[247],pp195[247],pp196[247]};
    assign in133_2 = {pp19[49],pp19[50],pp19[51],pp19[52],pp19[53],pp19[54],pp19[55],pp19[56],pp19[57],pp19[58],pp19[59],pp19[60],pp19[61],pp19[62],pp19[63],pp19[64],pp19[65],pp19[66],pp19[67],pp19[68],pp19[69],pp19[70],pp19[71],pp19[72],pp19[73],pp19[74],pp19[75],pp19[76],pp19[77],pp19[78],pp19[79],pp19[80],pp18[82],pp17[84],pp16[86],pp15[88],pp14[90],pp13[92],pp12[94],pp11[96],pp10[98],pp9[100],pp7[103],pp5[106],pp3[109],pp1[112],pp104[10],pp103[12],pp102[14],pp101[16],pp100[18],pp19[100],pp19[101],pp19[102],pp19[103],pp19[104],pp19[105],pp19[106],pp19[107],pp19[108],pp21[107],pp23[106],pp25[105],pp27[104],pp29[103],pp31[102],pp33[101],pp35[100],pp100[36],pp101[36],pp102[36],pp103[36],pp104[36],pp105[36],pp106[36],pp107[36],pp108[36],pp109[36],pp110[36],pp111[36],pp112[36],pp113[36],pp114[36],pp115[36],pp116[36],pp117[36],pp118[36],pp119[36],pp120[36],pp121[36],pp122[36],pp123[36],pp124[36],pp125[36],pp126[36],pp127[36],pp128[36],pp129[36],pp130[36],pp131[36],pp132[36],pp133[36],pp134[36],pp135[36],pp136[36],pp137[36],pp138[36],pp139[36],pp140[36],pp141[36],pp142[36],pp143[36],pp144[36],pp145[36],pp146[36],pp147[36],pp148[36],pp149[36],pp150[36],pp151[36],pp152[36],pp153[36],pp154[36],pp155[36],pp156[36],pp157[36],pp158[36],pp159[36],pp160[36],pp161[36],pp162[36],pp163[36],pp165[35],pp167[34],pp169[33],pp171[32],pp173[31],pp175[30],pp177[29],pp179[28],pp181[27],pp183[26],pp185[25],pp187[24],pp189[23],pp191[22],pp193[21],pp195[20],pp197[19],pp199[18],pp201[17],pp203[16],pp205[15],pp207[14],pp209[13],pp211[12],pp213[11],pp215[10],s129[162],s130[162],s131[162],s132[162],pp0[230],pp1[230],pp2[230],pp3[230],pp4[230],pp5[230],pp6[230],pp7[230],pp8[230],pp9[230],pp231[9],pp233[8],pp235[7],pp237[6],pp239[5],pp241[4],pp243[3],pp245[2],pp247[1],pp249[0],s10[113],s11[113],s12[113],s13[113],s14[113],s15[113],s16[113],s15[115],s14[117],s13[119],s12[121],s11[123],s10[125],pp255[8],pp9[255],s130[200],s129[202],pp255[12],pp254[14],pp253[16],pp252[18],pp251[20],pp250[22],pp249[24],pp248[26],pp247[28],pp246[30],pp245[32],pp244[34],pp243[36],pp242[38],pp241[40],pp240[42],pp239[44],pp238[46],pp237[48],pp236[50],pp235[52],pp234[54],pp233[56],pp232[58],pp231[60],pp230[62],pp229[64],pp228[66],pp227[68],pp226[70],pp225[72],pp224[74],pp223[76],pp222[78],pp221[80],pp220[82],pp219[84],pp218[86],pp217[88],pp216[90],pp215[92],pp214[94],pp213[96],pp212[98],pp99[212],pp97[215],pp95[218],pp93[221],pp91[224],pp89[227],pp87[230],pp85[233],pp83[236],pp81[239],pp79[242],pp77[245],pp75[248],pp73[251],pp71[254],pp225[101],pp223[104],pp221[107],pp219[110],pp217[113],pp215[116],pp213[119],pp211[122],pp209[125],pp207[128],pp205[131],pp203[134],pp201[137],pp199[140],pp197[143],pp195[146],pp193[149],pp191[152],pp189[155],pp187[158],pp185[161],pp183[164],pp181[167],pp179[170],pp177[173],pp175[176],pp173[179],pp171[182],pp169[185],pp167[188],pp166[190],pp165[192],pp164[194],pp163[196],pp162[198],pp161[200],pp160[202],pp159[204],pp158[206],pp157[208],pp156[210],pp155[212],pp154[214],pp153[216],pp152[218],pp151[220],pp150[222],pp149[224],pp148[226],pp147[228],pp146[230],pp145[232],pp144[234],pp143[236],pp142[238],pp141[240],pp140[242],pp139[244],pp138[246],pp139[246],pp140[246],pp141[246],pp142[246],pp143[246],pp144[246],pp145[246],pp146[246],pp147[246],pp148[246],pp149[246],pp150[246],pp151[246],pp152[246],pp153[246],pp154[246],pp155[246],pp156[246],pp157[246],pp158[246],pp159[246],pp160[246],pp161[246],pp162[246],pp163[246],pp164[246],pp165[246],pp166[246],pp167[246],pp168[246],pp169[246],pp170[246],pp171[246],pp172[246],pp173[246],pp174[246],pp175[246],pp176[246],pp177[246],pp178[246],pp179[246],pp180[246],pp181[246],pp182[246],pp183[246],pp184[246],pp185[246],pp186[246],pp187[246],pp188[246],pp189[246],pp190[246],pp191[246],pp192[246],pp193[246],pp194[246],pp195[246],pp196[246],pp197[246]};
    CLA_376 KS_133(s133, c133, in133_1, in133_2);
    wire[373:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp20[49],pp20[50],pp20[51],pp20[52],pp20[53],pp20[54],pp20[55],pp20[56],pp20[57],pp20[58],pp20[59],pp20[60],pp20[61],pp20[62],pp20[63],pp20[64],pp20[65],pp20[66],pp20[67],pp20[68],pp20[69],pp20[70],pp20[71],pp20[72],pp20[73],pp20[74],pp20[75],pp20[76],pp20[77],pp20[78],pp20[79],pp19[81],pp18[83],pp17[85],pp16[87],pp15[89],pp14[91],pp13[93],pp12[95],pp11[97],pp10[99],pp8[102],pp6[105],pp4[108],pp2[111],pp0[114],pp104[11],pp103[13],pp102[15],pp101[17],pp100[19],pp20[100],pp20[101],pp20[102],pp20[103],pp20[104],pp20[105],pp20[106],pp20[107],pp22[106],pp24[105],pp26[104],pp28[103],pp30[102],pp32[101],pp34[100],pp100[35],pp101[35],pp102[35],pp103[35],pp104[35],pp105[35],pp106[35],pp107[35],pp108[35],pp109[35],pp110[35],pp111[35],pp112[35],pp113[35],pp114[35],pp115[35],pp116[35],pp117[35],pp118[35],pp119[35],pp120[35],pp121[35],pp122[35],pp123[35],pp124[35],pp125[35],pp126[35],pp127[35],pp128[35],pp129[35],pp130[35],pp131[35],pp132[35],pp133[35],pp134[35],pp135[35],pp136[35],pp137[35],pp138[35],pp139[35],pp140[35],pp141[35],pp142[35],pp143[35],pp144[35],pp145[35],pp146[35],pp147[35],pp148[35],pp149[35],pp150[35],pp151[35],pp152[35],pp153[35],pp154[35],pp155[35],pp156[35],pp157[35],pp158[35],pp159[35],pp160[35],pp161[35],pp162[35],pp163[35],pp164[35],pp166[34],pp168[33],pp170[32],pp172[31],pp174[30],pp176[29],pp178[28],pp180[27],pp182[26],pp184[25],pp186[24],pp188[23],pp190[22],pp192[21],pp194[20],pp196[19],pp198[18],pp200[17],pp202[16],pp204[15],pp206[14],pp208[13],pp210[12],pp212[11],pp214[10],s129[161],s130[161],s131[161],s132[161],s133[161],s133[162],s133[163],s133[164],s133[165],s133[166],s133[167],s133[168],s133[169],s133[170],s133[171],s133[172],s133[173],s133[174],s133[175],s133[176],s133[177],s133[178],s133[179],s133[180],s133[181],s133[182],s133[183],s133[184],s133[185],s133[186],s133[187],s133[188],s133[189],s133[190],s133[191],s133[192],s133[193],s133[194],s133[195],s133[196],s131[199],s130[201],s129[203],pp255[13],pp254[15],pp253[17],pp252[19],pp251[21],pp250[23],pp249[25],pp248[27],pp247[29],pp246[31],pp245[33],pp244[35],pp243[37],pp242[39],pp241[41],pp240[43],pp239[45],pp238[47],pp237[49],pp236[51],pp235[53],pp234[55],pp233[57],pp232[59],pp231[61],pp230[63],pp229[65],pp228[67],pp227[69],pp226[71],pp225[73],pp224[75],pp223[77],pp222[79],pp221[81],pp220[83],pp219[85],pp218[87],pp217[89],pp216[91],pp215[93],pp214[95],pp213[97],pp212[99],pp98[214],pp96[217],pp94[220],pp92[223],pp90[226],pp88[229],pp86[232],pp84[235],pp82[238],pp80[241],pp78[244],pp76[247],pp74[250],pp72[253],pp226[100],pp224[103],pp222[106],pp220[109],pp218[112],pp216[115],pp214[118],pp212[121],pp210[124],pp208[127],pp206[130],pp204[133],pp202[136],pp200[139],pp198[142],pp196[145],pp194[148],pp192[151],pp190[154],pp188[157],pp186[160],pp184[163],pp182[166],pp180[169],pp178[172],pp176[175],pp174[178],pp172[181],pp170[184],pp168[187],pp167[189],pp166[191],pp165[193],pp164[195],pp163[197],pp162[199],pp161[201],pp160[203],pp159[205],pp158[207],pp157[209],pp156[211],pp155[213],pp154[215],pp153[217],pp152[219],pp151[221],pp150[223],pp149[225],pp148[227],pp147[229],pp146[231],pp145[233],pp144[235],pp143[237],pp142[239],pp141[241],pp140[243],pp139[245],pp140[245],pp141[245],pp142[245],pp143[245],pp144[245],pp145[245],pp146[245],pp147[245],pp148[245],pp149[245],pp150[245],pp151[245],pp152[245],pp153[245],pp154[245],pp155[245],pp156[245],pp157[245],pp158[245],pp159[245],pp160[245],pp161[245],pp162[245],pp163[245],pp164[245],pp165[245],pp166[245],pp167[245],pp168[245],pp169[245],pp170[245],pp171[245],pp172[245],pp173[245],pp174[245],pp175[245],pp176[245],pp177[245],pp178[245],pp179[245],pp180[245],pp181[245],pp182[245],pp183[245],pp184[245],pp185[245],pp186[245],pp187[245],pp188[245],pp189[245],pp190[245],pp191[245],pp192[245],pp193[245],pp194[245],pp195[245],pp196[245],pp197[245]};
    assign in134_2 = {pp21[48],pp21[49],pp21[50],pp21[51],pp21[52],pp21[53],pp21[54],pp21[55],pp21[56],pp21[57],pp21[58],pp21[59],pp21[60],pp21[61],pp21[62],pp21[63],pp21[64],pp21[65],pp21[66],pp21[67],pp21[68],pp21[69],pp21[70],pp21[71],pp21[72],pp21[73],pp21[74],pp21[75],pp21[76],pp21[77],pp21[78],pp20[80],pp19[82],pp18[84],pp17[86],pp16[88],pp15[90],pp14[92],pp13[94],pp12[96],pp11[98],pp9[101],pp7[104],pp5[107],pp3[110],pp1[113],pp105[10],pp104[12],pp103[14],pp102[16],pp101[18],pp100[20],pp21[100],pp21[101],pp21[102],pp21[103],pp21[104],pp21[105],pp21[106],pp23[105],pp25[104],pp27[103],pp29[102],pp31[101],pp33[100],pp100[34],pp101[34],pp102[34],pp103[34],pp104[34],pp105[34],pp106[34],pp107[34],pp108[34],pp109[34],pp110[34],pp111[34],pp112[34],pp113[34],pp114[34],pp115[34],pp116[34],pp117[34],pp118[34],pp119[34],pp120[34],pp121[34],pp122[34],pp123[34],pp124[34],pp125[34],pp126[34],pp127[34],pp128[34],pp129[34],pp130[34],pp131[34],pp132[34],pp133[34],pp134[34],pp135[34],pp136[34],pp137[34],pp138[34],pp139[34],pp140[34],pp141[34],pp142[34],pp143[34],pp144[34],pp145[34],pp146[34],pp147[34],pp148[34],pp149[34],pp150[34],pp151[34],pp152[34],pp153[34],pp154[34],pp155[34],pp156[34],pp157[34],pp158[34],pp159[34],pp160[34],pp161[34],pp162[34],pp163[34],pp164[34],pp165[34],pp167[33],pp169[32],pp171[31],pp173[30],pp175[29],pp177[28],pp179[27],pp181[26],pp183[25],pp185[24],pp187[23],pp189[22],pp191[21],pp193[20],pp195[19],pp197[18],pp199[17],pp201[16],pp203[15],pp205[14],pp207[13],pp209[12],pp211[11],pp213[10],s129[160],s130[160],s131[160],s132[160],s133[160],pp0[229],pp1[229],pp2[229],pp3[229],pp4[229],pp5[229],pp6[229],pp7[229],pp8[229],pp9[229],pp230[9],pp232[8],pp234[7],pp236[6],pp238[5],pp240[4],pp242[3],pp244[2],pp246[1],pp248[0],s10[112],s11[112],s12[112],s13[112],s14[112],s15[112],s16[112],s17[112],s16[114],s15[116],s14[118],s13[120],s12[122],s11[124],s10[126],pp255[9],s132[198],s131[200],s130[202],s129[204],pp255[14],pp254[16],pp253[18],pp252[20],pp251[22],pp250[24],pp249[26],pp248[28],pp247[30],pp246[32],pp245[34],pp244[36],pp243[38],pp242[40],pp241[42],pp240[44],pp239[46],pp238[48],pp237[50],pp236[52],pp235[54],pp234[56],pp233[58],pp232[60],pp231[62],pp230[64],pp229[66],pp228[68],pp227[70],pp226[72],pp225[74],pp224[76],pp223[78],pp222[80],pp221[82],pp220[84],pp219[86],pp218[88],pp217[90],pp216[92],pp215[94],pp214[96],pp213[98],pp99[213],pp97[216],pp95[219],pp93[222],pp91[225],pp89[228],pp87[231],pp85[234],pp83[237],pp81[240],pp79[243],pp77[246],pp75[249],pp73[252],pp71[255],pp225[102],pp223[105],pp221[108],pp219[111],pp217[114],pp215[117],pp213[120],pp211[123],pp209[126],pp207[129],pp205[132],pp203[135],pp201[138],pp199[141],pp197[144],pp195[147],pp193[150],pp191[153],pp189[156],pp187[159],pp185[162],pp183[165],pp181[168],pp179[171],pp177[174],pp175[177],pp173[180],pp171[183],pp169[186],pp168[188],pp167[190],pp166[192],pp165[194],pp164[196],pp163[198],pp162[200],pp161[202],pp160[204],pp159[206],pp158[208],pp157[210],pp156[212],pp155[214],pp154[216],pp153[218],pp152[220],pp151[222],pp150[224],pp149[226],pp148[228],pp147[230],pp146[232],pp145[234],pp144[236],pp143[238],pp142[240],pp141[242],pp140[244],pp141[244],pp142[244],pp143[244],pp144[244],pp145[244],pp146[244],pp147[244],pp148[244],pp149[244],pp150[244],pp151[244],pp152[244],pp153[244],pp154[244],pp155[244],pp156[244],pp157[244],pp158[244],pp159[244],pp160[244],pp161[244],pp162[244],pp163[244],pp164[244],pp165[244],pp166[244],pp167[244],pp168[244],pp169[244],pp170[244],pp171[244],pp172[244],pp173[244],pp174[244],pp175[244],pp176[244],pp177[244],pp178[244],pp179[244],pp180[244],pp181[244],pp182[244],pp183[244],pp184[244],pp185[244],pp186[244],pp187[244],pp188[244],pp189[244],pp190[244],pp191[244],pp192[244],pp193[244],pp194[244],pp195[244],pp196[244],pp197[244],pp198[244]};
    CLA_374 KS_134(s134, c134, in134_1, in134_2);
    wire[371:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp22[48],pp22[49],pp22[50],pp22[51],pp22[52],pp22[53],pp22[54],pp22[55],pp22[56],pp22[57],pp22[58],pp22[59],pp22[60],pp22[61],pp22[62],pp22[63],pp22[64],pp22[65],pp22[66],pp22[67],pp22[68],pp22[69],pp22[70],pp22[71],pp22[72],pp22[73],pp22[74],pp22[75],pp22[76],pp22[77],pp21[79],pp20[81],pp19[83],pp18[85],pp17[87],pp16[89],pp15[91],pp14[93],pp13[95],pp12[97],pp11[99],pp8[103],pp6[106],pp4[109],pp2[112],pp0[115],pp105[11],pp104[13],pp103[15],pp102[17],pp101[19],pp100[21],pp22[100],pp22[101],pp22[102],pp22[103],pp22[104],pp22[105],pp24[104],pp26[103],pp28[102],pp30[101],pp32[100],pp100[33],pp101[33],pp102[33],pp103[33],pp104[33],pp105[33],pp106[33],pp107[33],pp108[33],pp109[33],pp110[33],pp111[33],pp112[33],pp113[33],pp114[33],pp115[33],pp116[33],pp117[33],pp118[33],pp119[33],pp120[33],pp121[33],pp122[33],pp123[33],pp124[33],pp125[33],pp126[33],pp127[33],pp128[33],pp129[33],pp130[33],pp131[33],pp132[33],pp133[33],pp134[33],pp135[33],pp136[33],pp137[33],pp138[33],pp139[33],pp140[33],pp141[33],pp142[33],pp143[33],pp144[33],pp145[33],pp146[33],pp147[33],pp148[33],pp149[33],pp150[33],pp151[33],pp152[33],pp153[33],pp154[33],pp155[33],pp156[33],pp157[33],pp158[33],pp159[33],pp160[33],pp161[33],pp162[33],pp163[33],pp164[33],pp165[33],pp166[33],pp168[32],pp170[31],pp172[30],pp174[29],pp176[28],pp178[27],pp180[26],pp182[25],pp184[24],pp186[23],pp188[22],pp190[21],pp192[20],pp194[19],pp196[18],pp198[17],pp200[16],pp202[15],pp204[14],pp206[13],pp208[12],pp210[11],pp212[10],s129[159],s130[159],s131[159],s132[159],s133[159],s134[159],s134[160],s134[161],s134[162],s134[163],s134[164],s134[165],s134[166],s134[167],s134[168],s134[169],s134[170],s134[171],s134[172],s134[173],s134[174],s134[175],s134[176],s134[177],s134[178],s134[179],s134[180],s134[181],s134[182],s134[183],s134[184],s134[185],s134[186],s134[187],s134[188],s134[189],s134[190],s134[191],s134[192],s134[193],s134[194],s134[195],s133[197],s132[199],s131[201],s130[203],s129[205],pp255[15],pp254[17],pp253[19],pp252[21],pp251[23],pp250[25],pp249[27],pp248[29],pp247[31],pp246[33],pp245[35],pp244[37],pp243[39],pp242[41],pp241[43],pp240[45],pp239[47],pp238[49],pp237[51],pp236[53],pp235[55],pp234[57],pp233[59],pp232[61],pp231[63],pp230[65],pp229[67],pp228[69],pp227[71],pp226[73],pp225[75],pp224[77],pp223[79],pp222[81],pp221[83],pp220[85],pp219[87],pp218[89],pp217[91],pp216[93],pp215[95],pp214[97],pp213[99],pp98[215],pp96[218],pp94[221],pp92[224],pp90[227],pp88[230],pp86[233],pp84[236],pp82[239],pp80[242],pp78[245],pp76[248],pp74[251],pp72[254],pp226[101],pp224[104],pp222[107],pp220[110],pp218[113],pp216[116],pp214[119],pp212[122],pp210[125],pp208[128],pp206[131],pp204[134],pp202[137],pp200[140],pp198[143],pp196[146],pp194[149],pp192[152],pp190[155],pp188[158],pp186[161],pp184[164],pp182[167],pp180[170],pp178[173],pp176[176],pp174[179],pp172[182],pp170[185],pp169[187],pp168[189],pp167[191],pp166[193],pp165[195],pp164[197],pp163[199],pp162[201],pp161[203],pp160[205],pp159[207],pp158[209],pp157[211],pp156[213],pp155[215],pp154[217],pp153[219],pp152[221],pp151[223],pp150[225],pp149[227],pp148[229],pp147[231],pp146[233],pp145[235],pp144[237],pp143[239],pp142[241],pp141[243],pp142[243],pp143[243],pp144[243],pp145[243],pp146[243],pp147[243],pp148[243],pp149[243],pp150[243],pp151[243],pp152[243],pp153[243],pp154[243],pp155[243],pp156[243],pp157[243],pp158[243],pp159[243],pp160[243],pp161[243],pp162[243],pp163[243],pp164[243],pp165[243],pp166[243],pp167[243],pp168[243],pp169[243],pp170[243],pp171[243],pp172[243],pp173[243],pp174[243],pp175[243],pp176[243],pp177[243],pp178[243],pp179[243],pp180[243],pp181[243],pp182[243],pp183[243],pp184[243],pp185[243],pp186[243],pp187[243],pp188[243],pp189[243],pp190[243],pp191[243],pp192[243],pp193[243],pp194[243],pp195[243],pp196[243],pp197[243],pp198[243]};
    assign in135_2 = {pp23[47],pp23[48],pp23[49],pp23[50],pp23[51],pp23[52],pp23[53],pp23[54],pp23[55],pp23[56],pp23[57],pp23[58],pp23[59],pp23[60],pp23[61],pp23[62],pp23[63],pp23[64],pp23[65],pp23[66],pp23[67],pp23[68],pp23[69],pp23[70],pp23[71],pp23[72],pp23[73],pp23[74],pp23[75],pp23[76],pp22[78],pp21[80],pp20[82],pp19[84],pp18[86],pp17[88],pp16[90],pp15[92],pp14[94],pp13[96],pp12[98],pp9[102],pp7[105],pp5[108],pp3[111],pp1[114],pp106[10],pp105[12],pp104[14],pp103[16],pp102[18],pp101[20],pp100[22],pp23[100],pp23[101],pp23[102],pp23[103],pp23[104],pp25[103],pp27[102],pp29[101],pp31[100],pp100[32],pp101[32],pp102[32],pp103[32],pp104[32],pp105[32],pp106[32],pp107[32],pp108[32],pp109[32],pp110[32],pp111[32],pp112[32],pp113[32],pp114[32],pp115[32],pp116[32],pp117[32],pp118[32],pp119[32],pp120[32],pp121[32],pp122[32],pp123[32],pp124[32],pp125[32],pp126[32],pp127[32],pp128[32],pp129[32],pp130[32],pp131[32],pp132[32],pp133[32],pp134[32],pp135[32],pp136[32],pp137[32],pp138[32],pp139[32],pp140[32],pp141[32],pp142[32],pp143[32],pp144[32],pp145[32],pp146[32],pp147[32],pp148[32],pp149[32],pp150[32],pp151[32],pp152[32],pp153[32],pp154[32],pp155[32],pp156[32],pp157[32],pp158[32],pp159[32],pp160[32],pp161[32],pp162[32],pp163[32],pp164[32],pp165[32],pp166[32],pp167[32],pp169[31],pp171[30],pp173[29],pp175[28],pp177[27],pp179[26],pp181[25],pp183[24],pp185[23],pp187[22],pp189[21],pp191[20],pp193[19],pp195[18],pp197[17],pp199[16],pp201[15],pp203[14],pp205[13],pp207[12],pp209[11],pp211[10],s129[158],s130[158],s131[158],s132[158],s133[158],s134[158],pp0[228],pp1[228],pp2[228],pp3[228],pp4[228],pp5[228],pp6[228],pp7[228],pp8[228],pp9[228],pp229[9],pp231[8],pp233[7],pp235[6],pp237[5],pp239[4],pp241[3],pp243[2],pp245[1],pp247[0],s10[111],s11[111],s12[111],s13[111],s14[111],s15[111],s16[111],s17[111],s18[111],s17[113],s16[115],s15[117],s14[119],s13[121],s12[123],s11[125],s10[127],s134[196],s133[198],s132[200],s131[202],s130[204],s129[206],pp255[16],pp254[18],pp253[20],pp252[22],pp251[24],pp250[26],pp249[28],pp248[30],pp247[32],pp246[34],pp245[36],pp244[38],pp243[40],pp242[42],pp241[44],pp240[46],pp239[48],pp238[50],pp237[52],pp236[54],pp235[56],pp234[58],pp233[60],pp232[62],pp231[64],pp230[66],pp229[68],pp228[70],pp227[72],pp226[74],pp225[76],pp224[78],pp223[80],pp222[82],pp221[84],pp220[86],pp219[88],pp218[90],pp217[92],pp216[94],pp215[96],pp214[98],pp99[214],pp97[217],pp95[220],pp93[223],pp91[226],pp89[229],pp87[232],pp85[235],pp83[238],pp81[241],pp79[244],pp77[247],pp75[250],pp73[253],pp227[100],pp225[103],pp223[106],pp221[109],pp219[112],pp217[115],pp215[118],pp213[121],pp211[124],pp209[127],pp207[130],pp205[133],pp203[136],pp201[139],pp199[142],pp197[145],pp195[148],pp193[151],pp191[154],pp189[157],pp187[160],pp185[163],pp183[166],pp181[169],pp179[172],pp177[175],pp175[178],pp173[181],pp171[184],pp170[186],pp169[188],pp168[190],pp167[192],pp166[194],pp165[196],pp164[198],pp163[200],pp162[202],pp161[204],pp160[206],pp159[208],pp158[210],pp157[212],pp156[214],pp155[216],pp154[218],pp153[220],pp152[222],pp151[224],pp150[226],pp149[228],pp148[230],pp147[232],pp146[234],pp145[236],pp144[238],pp143[240],pp142[242],pp143[242],pp144[242],pp145[242],pp146[242],pp147[242],pp148[242],pp149[242],pp150[242],pp151[242],pp152[242],pp153[242],pp154[242],pp155[242],pp156[242],pp157[242],pp158[242],pp159[242],pp160[242],pp161[242],pp162[242],pp163[242],pp164[242],pp165[242],pp166[242],pp167[242],pp168[242],pp169[242],pp170[242],pp171[242],pp172[242],pp173[242],pp174[242],pp175[242],pp176[242],pp177[242],pp178[242],pp179[242],pp180[242],pp181[242],pp182[242],pp183[242],pp184[242],pp185[242],pp186[242],pp187[242],pp188[242],pp189[242],pp190[242],pp191[242],pp192[242],pp193[242],pp194[242],pp195[242],pp196[242],pp197[242],pp198[242],pp199[242]};
    CLA_372 KS_135(s135, c135, in135_1, in135_2);
    wire[369:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp24[47],pp24[48],pp24[49],pp24[50],pp24[51],pp24[52],pp24[53],pp24[54],pp24[55],pp24[56],pp24[57],pp24[58],pp24[59],pp24[60],pp24[61],pp24[62],pp24[63],pp24[64],pp24[65],pp24[66],pp24[67],pp24[68],pp24[69],pp24[70],pp24[71],pp24[72],pp24[73],pp24[74],pp24[75],pp23[77],pp22[79],pp21[81],pp20[83],pp19[85],pp18[87],pp17[89],pp16[91],pp15[93],pp14[95],pp13[97],pp12[99],pp8[104],pp6[107],pp4[110],pp2[113],pp0[116],pp106[11],pp105[13],pp104[15],pp103[17],pp102[19],pp101[21],pp100[23],pp24[100],pp24[101],pp24[102],pp24[103],pp26[102],pp28[101],pp30[100],pp100[31],pp101[31],pp102[31],pp103[31],pp104[31],pp105[31],pp106[31],pp107[31],pp108[31],pp109[31],pp110[31],pp111[31],pp112[31],pp113[31],pp114[31],pp115[31],pp116[31],pp117[31],pp118[31],pp119[31],pp120[31],pp121[31],pp122[31],pp123[31],pp124[31],pp125[31],pp126[31],pp127[31],pp128[31],pp129[31],pp130[31],pp131[31],pp132[31],pp133[31],pp134[31],pp135[31],pp136[31],pp137[31],pp138[31],pp139[31],pp140[31],pp141[31],pp142[31],pp143[31],pp144[31],pp145[31],pp146[31],pp147[31],pp148[31],pp149[31],pp150[31],pp151[31],pp152[31],pp153[31],pp154[31],pp155[31],pp156[31],pp157[31],pp158[31],pp159[31],pp160[31],pp161[31],pp162[31],pp163[31],pp164[31],pp165[31],pp166[31],pp167[31],pp168[31],pp170[30],pp172[29],pp174[28],pp176[27],pp178[26],pp180[25],pp182[24],pp184[23],pp186[22],pp188[21],pp190[20],pp192[19],pp194[18],pp196[17],pp198[16],pp200[15],pp202[14],pp204[13],pp206[12],pp208[11],pp210[10],s129[157],s130[157],s131[157],s132[157],s133[157],s134[157],s135[157],s135[158],s135[159],s135[160],s135[161],s135[162],s135[163],s135[164],s135[165],s135[166],s135[167],s135[168],s135[169],s135[170],s135[171],s135[172],s135[173],s135[174],s135[175],s135[176],s135[177],s135[178],s135[179],s135[180],s135[181],s135[182],s135[183],s135[184],s135[185],s135[186],s135[187],s135[188],s135[189],s135[190],s135[191],s135[192],s135[193],s135[194],s135[195],s134[197],s133[199],s132[201],s131[203],s130[205],s129[207],pp255[17],pp254[19],pp253[21],pp252[23],pp251[25],pp250[27],pp249[29],pp248[31],pp247[33],pp246[35],pp245[37],pp244[39],pp243[41],pp242[43],pp241[45],pp240[47],pp239[49],pp238[51],pp237[53],pp236[55],pp235[57],pp234[59],pp233[61],pp232[63],pp231[65],pp230[67],pp229[69],pp228[71],pp227[73],pp226[75],pp225[77],pp224[79],pp223[81],pp222[83],pp221[85],pp220[87],pp219[89],pp218[91],pp217[93],pp216[95],pp215[97],pp214[99],pp98[216],pp96[219],pp94[222],pp92[225],pp90[228],pp88[231],pp86[234],pp84[237],pp82[240],pp80[243],pp78[246],pp76[249],pp74[252],pp72[255],pp226[102],pp224[105],pp222[108],pp220[111],pp218[114],pp216[117],pp214[120],pp212[123],pp210[126],pp208[129],pp206[132],pp204[135],pp202[138],pp200[141],pp198[144],pp196[147],pp194[150],pp192[153],pp190[156],pp188[159],pp186[162],pp184[165],pp182[168],pp180[171],pp178[174],pp176[177],pp174[180],pp172[183],pp171[185],pp170[187],pp169[189],pp168[191],pp167[193],pp166[195],pp165[197],pp164[199],pp163[201],pp162[203],pp161[205],pp160[207],pp159[209],pp158[211],pp157[213],pp156[215],pp155[217],pp154[219],pp153[221],pp152[223],pp151[225],pp150[227],pp149[229],pp148[231],pp147[233],pp146[235],pp145[237],pp144[239],pp143[241],pp144[241],pp145[241],pp146[241],pp147[241],pp148[241],pp149[241],pp150[241],pp151[241],pp152[241],pp153[241],pp154[241],pp155[241],pp156[241],pp157[241],pp158[241],pp159[241],pp160[241],pp161[241],pp162[241],pp163[241],pp164[241],pp165[241],pp166[241],pp167[241],pp168[241],pp169[241],pp170[241],pp171[241],pp172[241],pp173[241],pp174[241],pp175[241],pp176[241],pp177[241],pp178[241],pp179[241],pp180[241],pp181[241],pp182[241],pp183[241],pp184[241],pp185[241],pp186[241],pp187[241],pp188[241],pp189[241],pp190[241],pp191[241],pp192[241],pp193[241],pp194[241],pp195[241],pp196[241],pp197[241],pp198[241],pp199[241]};
    assign in136_2 = {pp25[46],pp25[47],pp25[48],pp25[49],pp25[50],pp25[51],pp25[52],pp25[53],pp25[54],pp25[55],pp25[56],pp25[57],pp25[58],pp25[59],pp25[60],pp25[61],pp25[62],pp25[63],pp25[64],pp25[65],pp25[66],pp25[67],pp25[68],pp25[69],pp25[70],pp25[71],pp25[72],pp25[73],pp25[74],pp24[76],pp23[78],pp22[80],pp21[82],pp20[84],pp19[86],pp18[88],pp17[90],pp16[92],pp15[94],pp14[96],pp13[98],pp9[103],pp7[106],pp5[109],pp3[112],pp1[115],pp107[10],pp106[12],pp105[14],pp104[16],pp103[18],pp102[20],pp101[22],pp100[24],pp25[100],pp25[101],pp25[102],pp27[101],pp29[100],pp100[30],pp101[30],pp102[30],pp103[30],pp104[30],pp105[30],pp106[30],pp107[30],pp108[30],pp109[30],pp110[30],pp111[30],pp112[30],pp113[30],pp114[30],pp115[30],pp116[30],pp117[30],pp118[30],pp119[30],pp120[30],pp121[30],pp122[30],pp123[30],pp124[30],pp125[30],pp126[30],pp127[30],pp128[30],pp129[30],pp130[30],pp131[30],pp132[30],pp133[30],pp134[30],pp135[30],pp136[30],pp137[30],pp138[30],pp139[30],pp140[30],pp141[30],pp142[30],pp143[30],pp144[30],pp145[30],pp146[30],pp147[30],pp148[30],pp149[30],pp150[30],pp151[30],pp152[30],pp153[30],pp154[30],pp155[30],pp156[30],pp157[30],pp158[30],pp159[30],pp160[30],pp161[30],pp162[30],pp163[30],pp164[30],pp165[30],pp166[30],pp167[30],pp168[30],pp169[30],pp171[29],pp173[28],pp175[27],pp177[26],pp179[25],pp181[24],pp183[23],pp185[22],pp187[21],pp189[20],pp191[19],pp193[18],pp195[17],pp197[16],pp199[15],pp201[14],pp203[13],pp205[12],pp207[11],pp209[10],s129[156],s130[156],s131[156],s132[156],s133[156],s134[156],s135[156],pp0[227],pp1[227],pp2[227],pp3[227],pp4[227],pp5[227],pp6[227],pp7[227],pp8[227],pp9[227],pp228[9],pp230[8],pp232[7],pp234[6],pp236[5],pp238[4],pp240[3],pp242[2],pp244[1],pp246[0],s10[110],s11[110],s12[110],s13[110],s14[110],s15[110],s16[110],s17[110],s18[110],s19[110],s18[112],s17[114],s16[116],s15[118],s14[120],s13[122],s12[124],s11[126],s10[128],s135[196],s134[198],s133[200],s132[202],s131[204],s130[206],s129[208],pp255[18],pp254[20],pp253[22],pp252[24],pp251[26],pp250[28],pp249[30],pp248[32],pp247[34],pp246[36],pp245[38],pp244[40],pp243[42],pp242[44],pp241[46],pp240[48],pp239[50],pp238[52],pp237[54],pp236[56],pp235[58],pp234[60],pp233[62],pp232[64],pp231[66],pp230[68],pp229[70],pp228[72],pp227[74],pp226[76],pp225[78],pp224[80],pp223[82],pp222[84],pp221[86],pp220[88],pp219[90],pp218[92],pp217[94],pp216[96],pp215[98],pp99[215],pp97[218],pp95[221],pp93[224],pp91[227],pp89[230],pp87[233],pp85[236],pp83[239],pp81[242],pp79[245],pp77[248],pp75[251],pp73[254],pp227[101],pp225[104],pp223[107],pp221[110],pp219[113],pp217[116],pp215[119],pp213[122],pp211[125],pp209[128],pp207[131],pp205[134],pp203[137],pp201[140],pp199[143],pp197[146],pp195[149],pp193[152],pp191[155],pp189[158],pp187[161],pp185[164],pp183[167],pp181[170],pp179[173],pp177[176],pp175[179],pp173[182],pp172[184],pp171[186],pp170[188],pp169[190],pp168[192],pp167[194],pp166[196],pp165[198],pp164[200],pp163[202],pp162[204],pp161[206],pp160[208],pp159[210],pp158[212],pp157[214],pp156[216],pp155[218],pp154[220],pp153[222],pp152[224],pp151[226],pp150[228],pp149[230],pp148[232],pp147[234],pp146[236],pp145[238],pp144[240],pp145[240],pp146[240],pp147[240],pp148[240],pp149[240],pp150[240],pp151[240],pp152[240],pp153[240],pp154[240],pp155[240],pp156[240],pp157[240],pp158[240],pp159[240],pp160[240],pp161[240],pp162[240],pp163[240],pp164[240],pp165[240],pp166[240],pp167[240],pp168[240],pp169[240],pp170[240],pp171[240],pp172[240],pp173[240],pp174[240],pp175[240],pp176[240],pp177[240],pp178[240],pp179[240],pp180[240],pp181[240],pp182[240],pp183[240],pp184[240],pp185[240],pp186[240],pp187[240],pp188[240],pp189[240],pp190[240],pp191[240],pp192[240],pp193[240],pp194[240],pp195[240],pp196[240],pp197[240],pp198[240],pp199[240],pp200[240]};
    CLA_370 KS_136(s136, c136, in136_1, in136_2);
    wire[367:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp26[46],pp26[47],pp26[48],pp26[49],pp26[50],pp26[51],pp26[52],pp26[53],pp26[54],pp26[55],pp26[56],pp26[57],pp26[58],pp26[59],pp26[60],pp26[61],pp26[62],pp26[63],pp26[64],pp26[65],pp26[66],pp26[67],pp26[68],pp26[69],pp26[70],pp26[71],pp26[72],pp26[73],pp25[75],pp24[77],pp23[79],pp22[81],pp21[83],pp20[85],pp19[87],pp18[89],pp17[91],pp16[93],pp15[95],pp14[97],pp13[99],pp8[105],pp6[108],pp4[111],pp2[114],pp0[117],pp107[11],pp106[13],pp105[15],pp104[17],pp103[19],pp102[21],pp101[23],pp100[25],pp26[100],pp26[101],pp28[100],pp100[29],pp101[29],pp102[29],pp103[29],pp104[29],pp105[29],pp106[29],pp107[29],pp108[29],pp109[29],pp110[29],pp111[29],pp112[29],pp113[29],pp114[29],pp115[29],pp116[29],pp117[29],pp118[29],pp119[29],pp120[29],pp121[29],pp122[29],pp123[29],pp124[29],pp125[29],pp126[29],pp127[29],pp128[29],pp129[29],pp130[29],pp131[29],pp132[29],pp133[29],pp134[29],pp135[29],pp136[29],pp137[29],pp138[29],pp139[29],pp140[29],pp141[29],pp142[29],pp143[29],pp144[29],pp145[29],pp146[29],pp147[29],pp148[29],pp149[29],pp150[29],pp151[29],pp152[29],pp153[29],pp154[29],pp155[29],pp156[29],pp157[29],pp158[29],pp159[29],pp160[29],pp161[29],pp162[29],pp163[29],pp164[29],pp165[29],pp166[29],pp167[29],pp168[29],pp169[29],pp170[29],pp172[28],pp174[27],pp176[26],pp178[25],pp180[24],pp182[23],pp184[22],pp186[21],pp188[20],pp190[19],pp192[18],pp194[17],pp196[16],pp198[15],pp200[14],pp202[13],pp204[12],pp206[11],pp208[10],s129[155],s130[155],s131[155],s132[155],s133[155],s134[155],s135[155],s136[155],s136[156],s136[157],s136[158],s136[159],s136[160],s136[161],s136[162],s136[163],s136[164],s136[165],s136[166],s136[167],s136[168],s136[169],s136[170],s136[171],s136[172],s136[173],s136[174],s136[175],s136[176],s136[177],s136[178],s136[179],s136[180],s136[181],s136[182],s136[183],s136[184],s136[185],s136[186],s136[187],s136[188],s136[189],s136[190],s136[191],s136[192],s136[193],s136[194],s136[195],s135[197],s134[199],s133[201],s132[203],s131[205],s130[207],s129[209],pp255[19],pp254[21],pp253[23],pp252[25],pp251[27],pp250[29],pp249[31],pp248[33],pp247[35],pp246[37],pp245[39],pp244[41],pp243[43],pp242[45],pp241[47],pp240[49],pp239[51],pp238[53],pp237[55],pp236[57],pp235[59],pp234[61],pp233[63],pp232[65],pp231[67],pp230[69],pp229[71],pp228[73],pp227[75],pp226[77],pp225[79],pp224[81],pp223[83],pp222[85],pp221[87],pp220[89],pp219[91],pp218[93],pp217[95],pp216[97],pp215[99],pp98[217],pp96[220],pp94[223],pp92[226],pp90[229],pp88[232],pp86[235],pp84[238],pp82[241],pp80[244],pp78[247],pp76[250],pp74[253],pp228[100],pp226[103],pp224[106],pp222[109],pp220[112],pp218[115],pp216[118],pp214[121],pp212[124],pp210[127],pp208[130],pp206[133],pp204[136],pp202[139],pp200[142],pp198[145],pp196[148],pp194[151],pp192[154],pp190[157],pp188[160],pp186[163],pp184[166],pp182[169],pp180[172],pp178[175],pp176[178],pp174[181],pp173[183],pp172[185],pp171[187],pp170[189],pp169[191],pp168[193],pp167[195],pp166[197],pp165[199],pp164[201],pp163[203],pp162[205],pp161[207],pp160[209],pp159[211],pp158[213],pp157[215],pp156[217],pp155[219],pp154[221],pp153[223],pp152[225],pp151[227],pp150[229],pp149[231],pp148[233],pp147[235],pp146[237],pp145[239],pp146[239],pp147[239],pp148[239],pp149[239],pp150[239],pp151[239],pp152[239],pp153[239],pp154[239],pp155[239],pp156[239],pp157[239],pp158[239],pp159[239],pp160[239],pp161[239],pp162[239],pp163[239],pp164[239],pp165[239],pp166[239],pp167[239],pp168[239],pp169[239],pp170[239],pp171[239],pp172[239],pp173[239],pp174[239],pp175[239],pp176[239],pp177[239],pp178[239],pp179[239],pp180[239],pp181[239],pp182[239],pp183[239],pp184[239],pp185[239],pp186[239],pp187[239],pp188[239],pp189[239],pp190[239],pp191[239],pp192[239],pp193[239],pp194[239],pp195[239],pp196[239],pp197[239],pp198[239],pp199[239],pp200[239]};
    assign in137_2 = {pp27[45],pp27[46],pp27[47],pp27[48],pp27[49],pp27[50],pp27[51],pp27[52],pp27[53],pp27[54],pp27[55],pp27[56],pp27[57],pp27[58],pp27[59],pp27[60],pp27[61],pp27[62],pp27[63],pp27[64],pp27[65],pp27[66],pp27[67],pp27[68],pp27[69],pp27[70],pp27[71],pp27[72],pp26[74],pp25[76],pp24[78],pp23[80],pp22[82],pp21[84],pp20[86],pp19[88],pp18[90],pp17[92],pp16[94],pp15[96],pp14[98],pp9[104],pp7[107],pp5[110],pp3[113],pp1[116],pp108[10],pp107[12],pp106[14],pp105[16],pp104[18],pp103[20],pp102[22],pp101[24],pp100[26],pp27[100],pp100[28],pp101[28],pp102[28],pp103[28],pp104[28],pp105[28],pp106[28],pp107[28],pp108[28],pp109[28],pp110[28],pp111[28],pp112[28],pp113[28],pp114[28],pp115[28],pp116[28],pp117[28],pp118[28],pp119[28],pp120[28],pp121[28],pp122[28],pp123[28],pp124[28],pp125[28],pp126[28],pp127[28],pp128[28],pp129[28],pp130[28],pp131[28],pp132[28],pp133[28],pp134[28],pp135[28],pp136[28],pp137[28],pp138[28],pp139[28],pp140[28],pp141[28],pp142[28],pp143[28],pp144[28],pp145[28],pp146[28],pp147[28],pp148[28],pp149[28],pp150[28],pp151[28],pp152[28],pp153[28],pp154[28],pp155[28],pp156[28],pp157[28],pp158[28],pp159[28],pp160[28],pp161[28],pp162[28],pp163[28],pp164[28],pp165[28],pp166[28],pp167[28],pp168[28],pp169[28],pp170[28],pp171[28],pp173[27],pp175[26],pp177[25],pp179[24],pp181[23],pp183[22],pp185[21],pp187[20],pp189[19],pp191[18],pp193[17],pp195[16],pp197[15],pp199[14],pp201[13],pp203[12],pp205[11],pp207[10],s129[154],s130[154],s131[154],s132[154],s133[154],s134[154],s135[154],s136[154],pp0[226],pp1[226],pp2[226],pp3[226],pp4[226],pp5[226],pp6[226],pp7[226],pp8[226],pp9[226],pp227[9],pp229[8],pp231[7],pp233[6],pp235[5],pp237[4],pp239[3],pp241[2],pp243[1],pp245[0],s10[109],s11[109],s12[109],s13[109],s14[109],s15[109],s16[109],s17[109],s18[109],s19[109],s20[109],s19[111],s18[113],s17[115],s16[117],s15[119],s14[121],s13[123],s12[125],s11[127],s10[129],s136[196],s135[198],s134[200],s133[202],s132[204],s131[206],s130[208],s129[210],pp255[20],pp254[22],pp253[24],pp252[26],pp251[28],pp250[30],pp249[32],pp248[34],pp247[36],pp246[38],pp245[40],pp244[42],pp243[44],pp242[46],pp241[48],pp240[50],pp239[52],pp238[54],pp237[56],pp236[58],pp235[60],pp234[62],pp233[64],pp232[66],pp231[68],pp230[70],pp229[72],pp228[74],pp227[76],pp226[78],pp225[80],pp224[82],pp223[84],pp222[86],pp221[88],pp220[90],pp219[92],pp218[94],pp217[96],pp216[98],pp99[216],pp97[219],pp95[222],pp93[225],pp91[228],pp89[231],pp87[234],pp85[237],pp83[240],pp81[243],pp79[246],pp77[249],pp75[252],pp73[255],pp227[102],pp225[105],pp223[108],pp221[111],pp219[114],pp217[117],pp215[120],pp213[123],pp211[126],pp209[129],pp207[132],pp205[135],pp203[138],pp201[141],pp199[144],pp197[147],pp195[150],pp193[153],pp191[156],pp189[159],pp187[162],pp185[165],pp183[168],pp181[171],pp179[174],pp177[177],pp175[180],pp174[182],pp173[184],pp172[186],pp171[188],pp170[190],pp169[192],pp168[194],pp167[196],pp166[198],pp165[200],pp164[202],pp163[204],pp162[206],pp161[208],pp160[210],pp159[212],pp158[214],pp157[216],pp156[218],pp155[220],pp154[222],pp153[224],pp152[226],pp151[228],pp150[230],pp149[232],pp148[234],pp147[236],pp146[238],pp147[238],pp148[238],pp149[238],pp150[238],pp151[238],pp152[238],pp153[238],pp154[238],pp155[238],pp156[238],pp157[238],pp158[238],pp159[238],pp160[238],pp161[238],pp162[238],pp163[238],pp164[238],pp165[238],pp166[238],pp167[238],pp168[238],pp169[238],pp170[238],pp171[238],pp172[238],pp173[238],pp174[238],pp175[238],pp176[238],pp177[238],pp178[238],pp179[238],pp180[238],pp181[238],pp182[238],pp183[238],pp184[238],pp185[238],pp186[238],pp187[238],pp188[238],pp189[238],pp190[238],pp191[238],pp192[238],pp193[238],pp194[238],pp195[238],pp196[238],pp197[238],pp198[238],pp199[238],pp200[238],pp201[238]};
    CLA_368 KS_137(s137, c137, in137_1, in137_2);
    wire[365:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp28[45],pp28[46],pp28[47],pp28[48],pp28[49],pp28[50],pp28[51],pp28[52],pp28[53],pp28[54],pp28[55],pp28[56],pp28[57],pp28[58],pp28[59],pp28[60],pp28[61],pp28[62],pp28[63],pp28[64],pp28[65],pp28[66],pp28[67],pp28[68],pp28[69],pp28[70],pp28[71],pp27[73],pp26[75],pp25[77],pp24[79],pp23[81],pp22[83],pp21[85],pp20[87],pp19[89],pp18[91],pp17[93],pp16[95],pp15[97],pp14[99],pp8[106],pp6[109],pp4[112],pp2[115],pp0[118],pp108[11],pp107[13],pp106[15],pp105[17],pp104[19],pp103[21],pp102[23],pp101[25],pp100[27],pp101[27],pp102[27],pp103[27],pp104[27],pp105[27],pp106[27],pp107[27],pp108[27],pp109[27],pp110[27],pp111[27],pp112[27],pp113[27],pp114[27],pp115[27],pp116[27],pp117[27],pp118[27],pp119[27],pp120[27],pp121[27],pp122[27],pp123[27],pp124[27],pp125[27],pp126[27],pp127[27],pp128[27],pp129[27],pp130[27],pp131[27],pp132[27],pp133[27],pp134[27],pp135[27],pp136[27],pp137[27],pp138[27],pp139[27],pp140[27],pp141[27],pp142[27],pp143[27],pp144[27],pp145[27],pp146[27],pp147[27],pp148[27],pp149[27],pp150[27],pp151[27],pp152[27],pp153[27],pp154[27],pp155[27],pp156[27],pp157[27],pp158[27],pp159[27],pp160[27],pp161[27],pp162[27],pp163[27],pp164[27],pp165[27],pp166[27],pp167[27],pp168[27],pp169[27],pp170[27],pp171[27],pp172[27],pp174[26],pp176[25],pp178[24],pp180[23],pp182[22],pp184[21],pp186[20],pp188[19],pp190[18],pp192[17],pp194[16],pp196[15],pp198[14],pp200[13],pp202[12],pp204[11],pp206[10],s129[153],s130[153],s131[153],s132[153],s133[153],s134[153],s135[153],s136[153],s137[153],s137[154],s137[155],s137[156],s137[157],s137[158],s137[159],s137[160],s137[161],s137[162],s137[163],s137[164],s137[165],s137[166],s137[167],s137[168],s137[169],s137[170],s137[171],s137[172],s137[173],s137[174],s137[175],s137[176],s137[177],s137[178],s137[179],s137[180],s137[181],s137[182],s137[183],s137[184],s137[185],s137[186],s137[187],s137[188],s137[189],s137[190],s137[191],s137[192],s137[193],s137[194],s137[195],s136[197],s135[199],s134[201],s133[203],s132[205],s131[207],s130[209],s129[211],pp255[21],pp254[23],pp253[25],pp252[27],pp251[29],pp250[31],pp249[33],pp248[35],pp247[37],pp246[39],pp245[41],pp244[43],pp243[45],pp242[47],pp241[49],pp240[51],pp239[53],pp238[55],pp237[57],pp236[59],pp235[61],pp234[63],pp233[65],pp232[67],pp231[69],pp230[71],pp229[73],pp228[75],pp227[77],pp226[79],pp225[81],pp224[83],pp223[85],pp222[87],pp221[89],pp220[91],pp219[93],pp218[95],pp217[97],pp216[99],pp98[218],pp96[221],pp94[224],pp92[227],pp90[230],pp88[233],pp86[236],pp84[239],pp82[242],pp80[245],pp78[248],pp76[251],pp74[254],pp228[101],pp226[104],pp224[107],pp222[110],pp220[113],pp218[116],pp216[119],pp214[122],pp212[125],pp210[128],pp208[131],pp206[134],pp204[137],pp202[140],pp200[143],pp198[146],pp196[149],pp194[152],pp192[155],pp190[158],pp188[161],pp186[164],pp184[167],pp182[170],pp180[173],pp178[176],pp176[179],pp175[181],pp174[183],pp173[185],pp172[187],pp171[189],pp170[191],pp169[193],pp168[195],pp167[197],pp166[199],pp165[201],pp164[203],pp163[205],pp162[207],pp161[209],pp160[211],pp159[213],pp158[215],pp157[217],pp156[219],pp155[221],pp154[223],pp153[225],pp152[227],pp151[229],pp150[231],pp149[233],pp148[235],pp147[237],pp148[237],pp149[237],pp150[237],pp151[237],pp152[237],pp153[237],pp154[237],pp155[237],pp156[237],pp157[237],pp158[237],pp159[237],pp160[237],pp161[237],pp162[237],pp163[237],pp164[237],pp165[237],pp166[237],pp167[237],pp168[237],pp169[237],pp170[237],pp171[237],pp172[237],pp173[237],pp174[237],pp175[237],pp176[237],pp177[237],pp178[237],pp179[237],pp180[237],pp181[237],pp182[237],pp183[237],pp184[237],pp185[237],pp186[237],pp187[237],pp188[237],pp189[237],pp190[237],pp191[237],pp192[237],pp193[237],pp194[237],pp195[237],pp196[237],pp197[237],pp198[237],pp199[237],pp200[237],pp201[237]};
    assign in138_2 = {pp29[44],pp29[45],pp29[46],pp29[47],pp29[48],pp29[49],pp29[50],pp29[51],pp29[52],pp29[53],pp29[54],pp29[55],pp29[56],pp29[57],pp29[58],pp29[59],pp29[60],pp29[61],pp29[62],pp29[63],pp29[64],pp29[65],pp29[66],pp29[67],pp29[68],pp29[69],pp29[70],pp28[72],pp27[74],pp26[76],pp25[78],pp24[80],pp23[82],pp22[84],pp21[86],pp20[88],pp19[90],pp18[92],pp17[94],pp16[96],pp15[98],pp9[105],pp7[108],pp5[111],pp3[114],pp1[117],pp109[10],pp108[12],pp107[14],pp106[16],pp105[18],pp104[20],pp103[22],pp102[24],pp101[26],pp102[26],pp103[26],pp104[26],pp105[26],pp106[26],pp107[26],pp108[26],pp109[26],pp110[26],pp111[26],pp112[26],pp113[26],pp114[26],pp115[26],pp116[26],pp117[26],pp118[26],pp119[26],pp120[26],pp121[26],pp122[26],pp123[26],pp124[26],pp125[26],pp126[26],pp127[26],pp128[26],pp129[26],pp130[26],pp131[26],pp132[26],pp133[26],pp134[26],pp135[26],pp136[26],pp137[26],pp138[26],pp139[26],pp140[26],pp141[26],pp142[26],pp143[26],pp144[26],pp145[26],pp146[26],pp147[26],pp148[26],pp149[26],pp150[26],pp151[26],pp152[26],pp153[26],pp154[26],pp155[26],pp156[26],pp157[26],pp158[26],pp159[26],pp160[26],pp161[26],pp162[26],pp163[26],pp164[26],pp165[26],pp166[26],pp167[26],pp168[26],pp169[26],pp170[26],pp171[26],pp172[26],pp173[26],pp175[25],pp177[24],pp179[23],pp181[22],pp183[21],pp185[20],pp187[19],pp189[18],pp191[17],pp193[16],pp195[15],pp197[14],pp199[13],pp201[12],pp203[11],pp205[10],s129[152],s130[152],s131[152],s132[152],s133[152],s134[152],s135[152],s136[152],s137[152],pp0[225],pp1[225],pp2[225],pp3[225],pp4[225],pp5[225],pp6[225],pp7[225],pp8[225],pp9[225],pp226[9],pp228[8],pp230[7],pp232[6],pp234[5],pp236[4],pp238[3],pp240[2],pp242[1],pp244[0],s10[108],s11[108],s12[108],s13[108],s14[108],s15[108],s16[108],s17[108],s18[108],s19[108],s20[108],s21[108],s20[110],s19[112],s18[114],s17[116],s16[118],s15[120],s14[122],s13[124],s12[126],s11[128],s10[130],s137[196],s136[198],s135[200],s134[202],s133[204],s132[206],s131[208],s130[210],s129[212],pp255[22],pp254[24],pp253[26],pp252[28],pp251[30],pp250[32],pp249[34],pp248[36],pp247[38],pp246[40],pp245[42],pp244[44],pp243[46],pp242[48],pp241[50],pp240[52],pp239[54],pp238[56],pp237[58],pp236[60],pp235[62],pp234[64],pp233[66],pp232[68],pp231[70],pp230[72],pp229[74],pp228[76],pp227[78],pp226[80],pp225[82],pp224[84],pp223[86],pp222[88],pp221[90],pp220[92],pp219[94],pp218[96],pp217[98],pp99[217],pp97[220],pp95[223],pp93[226],pp91[229],pp89[232],pp87[235],pp85[238],pp83[241],pp81[244],pp79[247],pp77[250],pp75[253],pp229[100],pp227[103],pp225[106],pp223[109],pp221[112],pp219[115],pp217[118],pp215[121],pp213[124],pp211[127],pp209[130],pp207[133],pp205[136],pp203[139],pp201[142],pp199[145],pp197[148],pp195[151],pp193[154],pp191[157],pp189[160],pp187[163],pp185[166],pp183[169],pp181[172],pp179[175],pp177[178],pp176[180],pp175[182],pp174[184],pp173[186],pp172[188],pp171[190],pp170[192],pp169[194],pp168[196],pp167[198],pp166[200],pp165[202],pp164[204],pp163[206],pp162[208],pp161[210],pp160[212],pp159[214],pp158[216],pp157[218],pp156[220],pp155[222],pp154[224],pp153[226],pp152[228],pp151[230],pp150[232],pp149[234],pp148[236],pp149[236],pp150[236],pp151[236],pp152[236],pp153[236],pp154[236],pp155[236],pp156[236],pp157[236],pp158[236],pp159[236],pp160[236],pp161[236],pp162[236],pp163[236],pp164[236],pp165[236],pp166[236],pp167[236],pp168[236],pp169[236],pp170[236],pp171[236],pp172[236],pp173[236],pp174[236],pp175[236],pp176[236],pp177[236],pp178[236],pp179[236],pp180[236],pp181[236],pp182[236],pp183[236],pp184[236],pp185[236],pp186[236],pp187[236],pp188[236],pp189[236],pp190[236],pp191[236],pp192[236],pp193[236],pp194[236],pp195[236],pp196[236],pp197[236],pp198[236],pp199[236],pp200[236],pp201[236],pp202[236]};
    CLA_366 KS_138(s138, c138, in138_1, in138_2);
    wire[363:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp30[44],pp30[45],pp30[46],pp30[47],pp30[48],pp30[49],pp30[50],pp30[51],pp30[52],pp30[53],pp30[54],pp30[55],pp30[56],pp30[57],pp30[58],pp30[59],pp30[60],pp30[61],pp30[62],pp30[63],pp30[64],pp30[65],pp30[66],pp30[67],pp30[68],pp30[69],pp29[71],pp28[73],pp27[75],pp26[77],pp25[79],pp24[81],pp23[83],pp22[85],pp21[87],pp20[89],pp19[91],pp18[93],pp17[95],pp16[97],pp15[99],pp8[107],pp6[110],pp4[113],pp2[116],pp0[119],pp109[11],pp108[13],pp107[15],pp106[17],pp105[19],pp104[21],pp103[23],pp102[25],pp103[25],pp104[25],pp105[25],pp106[25],pp107[25],pp108[25],pp109[25],pp110[25],pp111[25],pp112[25],pp113[25],pp114[25],pp115[25],pp116[25],pp117[25],pp118[25],pp119[25],pp120[25],pp121[25],pp122[25],pp123[25],pp124[25],pp125[25],pp126[25],pp127[25],pp128[25],pp129[25],pp130[25],pp131[25],pp132[25],pp133[25],pp134[25],pp135[25],pp136[25],pp137[25],pp138[25],pp139[25],pp140[25],pp141[25],pp142[25],pp143[25],pp144[25],pp145[25],pp146[25],pp147[25],pp148[25],pp149[25],pp150[25],pp151[25],pp152[25],pp153[25],pp154[25],pp155[25],pp156[25],pp157[25],pp158[25],pp159[25],pp160[25],pp161[25],pp162[25],pp163[25],pp164[25],pp165[25],pp166[25],pp167[25],pp168[25],pp169[25],pp170[25],pp171[25],pp172[25],pp173[25],pp174[25],pp176[24],pp178[23],pp180[22],pp182[21],pp184[20],pp186[19],pp188[18],pp190[17],pp192[16],pp194[15],pp196[14],pp198[13],pp200[12],pp202[11],pp204[10],s129[151],s130[151],s131[151],s132[151],s133[151],s134[151],s135[151],s136[151],s137[151],s138[151],s138[152],s138[153],s138[154],s138[155],s138[156],s138[157],s138[158],s138[159],s138[160],s138[161],s138[162],s138[163],s138[164],s138[165],s138[166],s138[167],s138[168],s138[169],s138[170],s138[171],s138[172],s138[173],s138[174],s138[175],s138[176],s138[177],s138[178],s138[179],s138[180],s138[181],s138[182],s138[183],s138[184],s138[185],s138[186],s138[187],s138[188],s138[189],s138[190],s138[191],s138[192],s138[193],s138[194],s138[195],s137[197],s136[199],s135[201],s134[203],s133[205],s132[207],s131[209],s130[211],s129[213],pp255[23],pp254[25],pp253[27],pp252[29],pp251[31],pp250[33],pp249[35],pp248[37],pp247[39],pp246[41],pp245[43],pp244[45],pp243[47],pp242[49],pp241[51],pp240[53],pp239[55],pp238[57],pp237[59],pp236[61],pp235[63],pp234[65],pp233[67],pp232[69],pp231[71],pp230[73],pp229[75],pp228[77],pp227[79],pp226[81],pp225[83],pp224[85],pp223[87],pp222[89],pp221[91],pp220[93],pp219[95],pp218[97],pp217[99],pp98[219],pp96[222],pp94[225],pp92[228],pp90[231],pp88[234],pp86[237],pp84[240],pp82[243],pp80[246],pp78[249],pp76[252],pp74[255],pp228[102],pp226[105],pp224[108],pp222[111],pp220[114],pp218[117],pp216[120],pp214[123],pp212[126],pp210[129],pp208[132],pp206[135],pp204[138],pp202[141],pp200[144],pp198[147],pp196[150],pp194[153],pp192[156],pp190[159],pp188[162],pp186[165],pp184[168],pp182[171],pp180[174],pp178[177],pp177[179],pp176[181],pp175[183],pp174[185],pp173[187],pp172[189],pp171[191],pp170[193],pp169[195],pp168[197],pp167[199],pp166[201],pp165[203],pp164[205],pp163[207],pp162[209],pp161[211],pp160[213],pp159[215],pp158[217],pp157[219],pp156[221],pp155[223],pp154[225],pp153[227],pp152[229],pp151[231],pp150[233],pp149[235],pp150[235],pp151[235],pp152[235],pp153[235],pp154[235],pp155[235],pp156[235],pp157[235],pp158[235],pp159[235],pp160[235],pp161[235],pp162[235],pp163[235],pp164[235],pp165[235],pp166[235],pp167[235],pp168[235],pp169[235],pp170[235],pp171[235],pp172[235],pp173[235],pp174[235],pp175[235],pp176[235],pp177[235],pp178[235],pp179[235],pp180[235],pp181[235],pp182[235],pp183[235],pp184[235],pp185[235],pp186[235],pp187[235],pp188[235],pp189[235],pp190[235],pp191[235],pp192[235],pp193[235],pp194[235],pp195[235],pp196[235],pp197[235],pp198[235],pp199[235],pp200[235],pp201[235],pp202[235]};
    assign in139_2 = {pp31[43],pp31[44],pp31[45],pp31[46],pp31[47],pp31[48],pp31[49],pp31[50],pp31[51],pp31[52],pp31[53],pp31[54],pp31[55],pp31[56],pp31[57],pp31[58],pp31[59],pp31[60],pp31[61],pp31[62],pp31[63],pp31[64],pp31[65],pp31[66],pp31[67],pp31[68],pp30[70],pp29[72],pp28[74],pp27[76],pp26[78],pp25[80],pp24[82],pp23[84],pp22[86],pp21[88],pp20[90],pp19[92],pp18[94],pp17[96],pp16[98],pp9[106],pp7[109],pp5[112],pp3[115],pp1[118],pp110[10],pp109[12],pp108[14],pp107[16],pp106[18],pp105[20],pp104[22],pp103[24],pp104[24],pp105[24],pp106[24],pp107[24],pp108[24],pp109[24],pp110[24],pp111[24],pp112[24],pp113[24],pp114[24],pp115[24],pp116[24],pp117[24],pp118[24],pp119[24],pp120[24],pp121[24],pp122[24],pp123[24],pp124[24],pp125[24],pp126[24],pp127[24],pp128[24],pp129[24],pp130[24],pp131[24],pp132[24],pp133[24],pp134[24],pp135[24],pp136[24],pp137[24],pp138[24],pp139[24],pp140[24],pp141[24],pp142[24],pp143[24],pp144[24],pp145[24],pp146[24],pp147[24],pp148[24],pp149[24],pp150[24],pp151[24],pp152[24],pp153[24],pp154[24],pp155[24],pp156[24],pp157[24],pp158[24],pp159[24],pp160[24],pp161[24],pp162[24],pp163[24],pp164[24],pp165[24],pp166[24],pp167[24],pp168[24],pp169[24],pp170[24],pp171[24],pp172[24],pp173[24],pp174[24],pp175[24],pp177[23],pp179[22],pp181[21],pp183[20],pp185[19],pp187[18],pp189[17],pp191[16],pp193[15],pp195[14],pp197[13],pp199[12],pp201[11],pp203[10],s129[150],s130[150],s131[150],s132[150],s133[150],s134[150],s135[150],s136[150],s137[150],s138[150],pp0[224],pp1[224],pp2[224],pp3[224],pp4[224],pp5[224],pp6[224],pp7[224],pp8[224],pp9[224],pp225[9],pp227[8],pp229[7],pp231[6],pp233[5],pp235[4],pp237[3],pp239[2],pp241[1],pp243[0],s10[107],s11[107],s12[107],s13[107],s14[107],s15[107],s16[107],s17[107],s18[107],s19[107],s20[107],s21[107],s22[107],s21[109],s20[111],s19[113],s18[115],s17[117],s16[119],s15[121],s14[123],s13[125],s12[127],s11[129],s10[131],s138[196],s137[198],s136[200],s135[202],s134[204],s133[206],s132[208],s131[210],s130[212],s129[214],pp255[24],pp254[26],pp253[28],pp252[30],pp251[32],pp250[34],pp249[36],pp248[38],pp247[40],pp246[42],pp245[44],pp244[46],pp243[48],pp242[50],pp241[52],pp240[54],pp239[56],pp238[58],pp237[60],pp236[62],pp235[64],pp234[66],pp233[68],pp232[70],pp231[72],pp230[74],pp229[76],pp228[78],pp227[80],pp226[82],pp225[84],pp224[86],pp223[88],pp222[90],pp221[92],pp220[94],pp219[96],pp218[98],pp99[218],pp97[221],pp95[224],pp93[227],pp91[230],pp89[233],pp87[236],pp85[239],pp83[242],pp81[245],pp79[248],pp77[251],pp75[254],pp229[101],pp227[104],pp225[107],pp223[110],pp221[113],pp219[116],pp217[119],pp215[122],pp213[125],pp211[128],pp209[131],pp207[134],pp205[137],pp203[140],pp201[143],pp199[146],pp197[149],pp195[152],pp193[155],pp191[158],pp189[161],pp187[164],pp185[167],pp183[170],pp181[173],pp179[176],pp178[178],pp177[180],pp176[182],pp175[184],pp174[186],pp173[188],pp172[190],pp171[192],pp170[194],pp169[196],pp168[198],pp167[200],pp166[202],pp165[204],pp164[206],pp163[208],pp162[210],pp161[212],pp160[214],pp159[216],pp158[218],pp157[220],pp156[222],pp155[224],pp154[226],pp153[228],pp152[230],pp151[232],pp150[234],pp151[234],pp152[234],pp153[234],pp154[234],pp155[234],pp156[234],pp157[234],pp158[234],pp159[234],pp160[234],pp161[234],pp162[234],pp163[234],pp164[234],pp165[234],pp166[234],pp167[234],pp168[234],pp169[234],pp170[234],pp171[234],pp172[234],pp173[234],pp174[234],pp175[234],pp176[234],pp177[234],pp178[234],pp179[234],pp180[234],pp181[234],pp182[234],pp183[234],pp184[234],pp185[234],pp186[234],pp187[234],pp188[234],pp189[234],pp190[234],pp191[234],pp192[234],pp193[234],pp194[234],pp195[234],pp196[234],pp197[234],pp198[234],pp199[234],pp200[234],pp201[234],pp202[234],pp203[234]};
    CLA_364 KS_139(s139, c139, in139_1, in139_2);
    wire[361:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp32[43],pp32[44],pp32[45],pp32[46],pp32[47],pp32[48],pp32[49],pp32[50],pp32[51],pp32[52],pp32[53],pp32[54],pp32[55],pp32[56],pp32[57],pp32[58],pp32[59],pp32[60],pp32[61],pp32[62],pp32[63],pp32[64],pp32[65],pp32[66],pp32[67],pp31[69],pp30[71],pp29[73],pp28[75],pp27[77],pp26[79],pp25[81],pp24[83],pp23[85],pp22[87],pp21[89],pp20[91],pp19[93],pp18[95],pp17[97],pp16[99],pp8[108],pp6[111],pp4[114],pp2[117],pp0[120],pp110[11],pp109[13],pp108[15],pp107[17],pp106[19],pp105[21],pp104[23],pp105[23],pp106[23],pp107[23],pp108[23],pp109[23],pp110[23],pp111[23],pp112[23],pp113[23],pp114[23],pp115[23],pp116[23],pp117[23],pp118[23],pp119[23],pp120[23],pp121[23],pp122[23],pp123[23],pp124[23],pp125[23],pp126[23],pp127[23],pp128[23],pp129[23],pp130[23],pp131[23],pp132[23],pp133[23],pp134[23],pp135[23],pp136[23],pp137[23],pp138[23],pp139[23],pp140[23],pp141[23],pp142[23],pp143[23],pp144[23],pp145[23],pp146[23],pp147[23],pp148[23],pp149[23],pp150[23],pp151[23],pp152[23],pp153[23],pp154[23],pp155[23],pp156[23],pp157[23],pp158[23],pp159[23],pp160[23],pp161[23],pp162[23],pp163[23],pp164[23],pp165[23],pp166[23],pp167[23],pp168[23],pp169[23],pp170[23],pp171[23],pp172[23],pp173[23],pp174[23],pp175[23],pp176[23],pp178[22],pp180[21],pp182[20],pp184[19],pp186[18],pp188[17],pp190[16],pp192[15],pp194[14],pp196[13],pp198[12],pp200[11],pp202[10],s129[149],s130[149],s131[149],s132[149],s133[149],s134[149],s135[149],s136[149],s137[149],s138[149],s139[149],s139[150],s139[151],s139[152],s139[153],s139[154],s139[155],s139[156],s139[157],s139[158],s139[159],s139[160],s139[161],s139[162],s139[163],s139[164],s139[165],s139[166],s139[167],s139[168],s139[169],s139[170],s139[171],s139[172],s139[173],s139[174],s139[175],s139[176],s139[177],s139[178],s139[179],s139[180],s139[181],s139[182],s139[183],s139[184],s139[185],s139[186],s139[187],s139[188],s139[189],s139[190],s139[191],s139[192],s139[193],s139[194],s139[195],s138[197],s137[199],s136[201],s135[203],s134[205],s133[207],s132[209],s131[211],s130[213],s129[215],pp255[25],pp254[27],pp253[29],pp252[31],pp251[33],pp250[35],pp249[37],pp248[39],pp247[41],pp246[43],pp245[45],pp244[47],pp243[49],pp242[51],pp241[53],pp240[55],pp239[57],pp238[59],pp237[61],pp236[63],pp235[65],pp234[67],pp233[69],pp232[71],pp231[73],pp230[75],pp229[77],pp228[79],pp227[81],pp226[83],pp225[85],pp224[87],pp223[89],pp222[91],pp221[93],pp220[95],pp219[97],pp218[99],pp98[220],pp96[223],pp94[226],pp92[229],pp90[232],pp88[235],pp86[238],pp84[241],pp82[244],pp80[247],pp78[250],pp76[253],pp230[100],pp228[103],pp226[106],pp224[109],pp222[112],pp220[115],pp218[118],pp216[121],pp214[124],pp212[127],pp210[130],pp208[133],pp206[136],pp204[139],pp202[142],pp200[145],pp198[148],pp196[151],pp194[154],pp192[157],pp190[160],pp188[163],pp186[166],pp184[169],pp182[172],pp180[175],pp179[177],pp178[179],pp177[181],pp176[183],pp175[185],pp174[187],pp173[189],pp172[191],pp171[193],pp170[195],pp169[197],pp168[199],pp167[201],pp166[203],pp165[205],pp164[207],pp163[209],pp162[211],pp161[213],pp160[215],pp159[217],pp158[219],pp157[221],pp156[223],pp155[225],pp154[227],pp153[229],pp152[231],pp151[233],pp152[233],pp153[233],pp154[233],pp155[233],pp156[233],pp157[233],pp158[233],pp159[233],pp160[233],pp161[233],pp162[233],pp163[233],pp164[233],pp165[233],pp166[233],pp167[233],pp168[233],pp169[233],pp170[233],pp171[233],pp172[233],pp173[233],pp174[233],pp175[233],pp176[233],pp177[233],pp178[233],pp179[233],pp180[233],pp181[233],pp182[233],pp183[233],pp184[233],pp185[233],pp186[233],pp187[233],pp188[233],pp189[233],pp190[233],pp191[233],pp192[233],pp193[233],pp194[233],pp195[233],pp196[233],pp197[233],pp198[233],pp199[233],pp200[233],pp201[233],pp202[233],pp203[233]};
    assign in140_2 = {pp33[42],pp33[43],pp33[44],pp33[45],pp33[46],pp33[47],pp33[48],pp33[49],pp33[50],pp33[51],pp33[52],pp33[53],pp33[54],pp33[55],pp33[56],pp33[57],pp33[58],pp33[59],pp33[60],pp33[61],pp33[62],pp33[63],pp33[64],pp33[65],pp33[66],pp32[68],pp31[70],pp30[72],pp29[74],pp28[76],pp27[78],pp26[80],pp25[82],pp24[84],pp23[86],pp22[88],pp21[90],pp20[92],pp19[94],pp18[96],pp17[98],pp9[107],pp7[110],pp5[113],pp3[116],pp1[119],pp111[10],pp110[12],pp109[14],pp108[16],pp107[18],pp106[20],pp105[22],pp106[22],pp107[22],pp108[22],pp109[22],pp110[22],pp111[22],pp112[22],pp113[22],pp114[22],pp115[22],pp116[22],pp117[22],pp118[22],pp119[22],pp120[22],pp121[22],pp122[22],pp123[22],pp124[22],pp125[22],pp126[22],pp127[22],pp128[22],pp129[22],pp130[22],pp131[22],pp132[22],pp133[22],pp134[22],pp135[22],pp136[22],pp137[22],pp138[22],pp139[22],pp140[22],pp141[22],pp142[22],pp143[22],pp144[22],pp145[22],pp146[22],pp147[22],pp148[22],pp149[22],pp150[22],pp151[22],pp152[22],pp153[22],pp154[22],pp155[22],pp156[22],pp157[22],pp158[22],pp159[22],pp160[22],pp161[22],pp162[22],pp163[22],pp164[22],pp165[22],pp166[22],pp167[22],pp168[22],pp169[22],pp170[22],pp171[22],pp172[22],pp173[22],pp174[22],pp175[22],pp176[22],pp177[22],pp179[21],pp181[20],pp183[19],pp185[18],pp187[17],pp189[16],pp191[15],pp193[14],pp195[13],pp197[12],pp199[11],pp201[10],s129[148],s130[148],s131[148],s132[148],s133[148],s134[148],s135[148],s136[148],s137[148],s138[148],s139[148],pp0[223],pp1[223],pp2[223],pp3[223],pp4[223],pp5[223],pp6[223],pp7[223],pp8[223],pp9[223],pp224[9],pp226[8],pp228[7],pp230[6],pp232[5],pp234[4],pp236[3],pp238[2],pp240[1],pp242[0],s10[106],s11[106],s12[106],s13[106],s14[106],s15[106],s16[106],s17[106],s18[106],s19[106],s20[106],s21[106],s22[106],s23[106],s22[108],s21[110],s20[112],s19[114],s18[116],s17[118],s16[120],s15[122],s14[124],s13[126],s12[128],s11[130],s10[132],s139[196],s138[198],s137[200],s136[202],s135[204],s134[206],s133[208],s132[210],s131[212],s130[214],s129[216],pp255[26],pp254[28],pp253[30],pp252[32],pp251[34],pp250[36],pp249[38],pp248[40],pp247[42],pp246[44],pp245[46],pp244[48],pp243[50],pp242[52],pp241[54],pp240[56],pp239[58],pp238[60],pp237[62],pp236[64],pp235[66],pp234[68],pp233[70],pp232[72],pp231[74],pp230[76],pp229[78],pp228[80],pp227[82],pp226[84],pp225[86],pp224[88],pp223[90],pp222[92],pp221[94],pp220[96],pp219[98],pp99[219],pp97[222],pp95[225],pp93[228],pp91[231],pp89[234],pp87[237],pp85[240],pp83[243],pp81[246],pp79[249],pp77[252],pp75[255],pp229[102],pp227[105],pp225[108],pp223[111],pp221[114],pp219[117],pp217[120],pp215[123],pp213[126],pp211[129],pp209[132],pp207[135],pp205[138],pp203[141],pp201[144],pp199[147],pp197[150],pp195[153],pp193[156],pp191[159],pp189[162],pp187[165],pp185[168],pp183[171],pp181[174],pp180[176],pp179[178],pp178[180],pp177[182],pp176[184],pp175[186],pp174[188],pp173[190],pp172[192],pp171[194],pp170[196],pp169[198],pp168[200],pp167[202],pp166[204],pp165[206],pp164[208],pp163[210],pp162[212],pp161[214],pp160[216],pp159[218],pp158[220],pp157[222],pp156[224],pp155[226],pp154[228],pp153[230],pp152[232],pp153[232],pp154[232],pp155[232],pp156[232],pp157[232],pp158[232],pp159[232],pp160[232],pp161[232],pp162[232],pp163[232],pp164[232],pp165[232],pp166[232],pp167[232],pp168[232],pp169[232],pp170[232],pp171[232],pp172[232],pp173[232],pp174[232],pp175[232],pp176[232],pp177[232],pp178[232],pp179[232],pp180[232],pp181[232],pp182[232],pp183[232],pp184[232],pp185[232],pp186[232],pp187[232],pp188[232],pp189[232],pp190[232],pp191[232],pp192[232],pp193[232],pp194[232],pp195[232],pp196[232],pp197[232],pp198[232],pp199[232],pp200[232],pp201[232],pp202[232],pp203[232],pp204[232]};
    CLA_362 KS_140(s140, c140, in140_1, in140_2);
    wire[359:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp34[42],pp34[43],pp34[44],pp34[45],pp34[46],pp34[47],pp34[48],pp34[49],pp34[50],pp34[51],pp34[52],pp34[53],pp34[54],pp34[55],pp34[56],pp34[57],pp34[58],pp34[59],pp34[60],pp34[61],pp34[62],pp34[63],pp34[64],pp34[65],pp33[67],pp32[69],pp31[71],pp30[73],pp29[75],pp28[77],pp27[79],pp26[81],pp25[83],pp24[85],pp23[87],pp22[89],pp21[91],pp20[93],pp19[95],pp18[97],pp17[99],pp8[109],pp6[112],pp4[115],pp2[118],pp0[121],pp111[11],pp110[13],pp109[15],pp108[17],pp107[19],pp106[21],pp107[21],pp108[21],pp109[21],pp110[21],pp111[21],pp112[21],pp113[21],pp114[21],pp115[21],pp116[21],pp117[21],pp118[21],pp119[21],pp120[21],pp121[21],pp122[21],pp123[21],pp124[21],pp125[21],pp126[21],pp127[21],pp128[21],pp129[21],pp130[21],pp131[21],pp132[21],pp133[21],pp134[21],pp135[21],pp136[21],pp137[21],pp138[21],pp139[21],pp140[21],pp141[21],pp142[21],pp143[21],pp144[21],pp145[21],pp146[21],pp147[21],pp148[21],pp149[21],pp150[21],pp151[21],pp152[21],pp153[21],pp154[21],pp155[21],pp156[21],pp157[21],pp158[21],pp159[21],pp160[21],pp161[21],pp162[21],pp163[21],pp164[21],pp165[21],pp166[21],pp167[21],pp168[21],pp169[21],pp170[21],pp171[21],pp172[21],pp173[21],pp174[21],pp175[21],pp176[21],pp177[21],pp178[21],pp180[20],pp182[19],pp184[18],pp186[17],pp188[16],pp190[15],pp192[14],pp194[13],pp196[12],pp198[11],pp200[10],s129[147],s130[147],s131[147],s132[147],s133[147],s134[147],s135[147],s136[147],s137[147],s138[147],s139[147],s140[147],s140[148],s140[149],s140[150],s140[151],s140[152],s140[153],s140[154],s140[155],s140[156],s140[157],s140[158],s140[159],s140[160],s140[161],s140[162],s140[163],s140[164],s140[165],s140[166],s140[167],s140[168],s140[169],s140[170],s140[171],s140[172],s140[173],s140[174],s140[175],s140[176],s140[177],s140[178],s140[179],s140[180],s140[181],s140[182],s140[183],s140[184],s140[185],s140[186],s140[187],s140[188],s140[189],s140[190],s140[191],s140[192],s140[193],s140[194],s140[195],s139[197],s138[199],s137[201],s136[203],s135[205],s134[207],s133[209],s132[211],s131[213],s130[215],s129[217],pp255[27],pp254[29],pp253[31],pp252[33],pp251[35],pp250[37],pp249[39],pp248[41],pp247[43],pp246[45],pp245[47],pp244[49],pp243[51],pp242[53],pp241[55],pp240[57],pp239[59],pp238[61],pp237[63],pp236[65],pp235[67],pp234[69],pp233[71],pp232[73],pp231[75],pp230[77],pp229[79],pp228[81],pp227[83],pp226[85],pp225[87],pp224[89],pp223[91],pp222[93],pp221[95],pp220[97],pp219[99],pp98[221],pp96[224],pp94[227],pp92[230],pp90[233],pp88[236],pp86[239],pp84[242],pp82[245],pp80[248],pp78[251],pp76[254],pp230[101],pp228[104],pp226[107],pp224[110],pp222[113],pp220[116],pp218[119],pp216[122],pp214[125],pp212[128],pp210[131],pp208[134],pp206[137],pp204[140],pp202[143],pp200[146],pp198[149],pp196[152],pp194[155],pp192[158],pp190[161],pp188[164],pp186[167],pp184[170],pp182[173],pp181[175],pp180[177],pp179[179],pp178[181],pp177[183],pp176[185],pp175[187],pp174[189],pp173[191],pp172[193],pp171[195],pp170[197],pp169[199],pp168[201],pp167[203],pp166[205],pp165[207],pp164[209],pp163[211],pp162[213],pp161[215],pp160[217],pp159[219],pp158[221],pp157[223],pp156[225],pp155[227],pp154[229],pp153[231],pp154[231],pp155[231],pp156[231],pp157[231],pp158[231],pp159[231],pp160[231],pp161[231],pp162[231],pp163[231],pp164[231],pp165[231],pp166[231],pp167[231],pp168[231],pp169[231],pp170[231],pp171[231],pp172[231],pp173[231],pp174[231],pp175[231],pp176[231],pp177[231],pp178[231],pp179[231],pp180[231],pp181[231],pp182[231],pp183[231],pp184[231],pp185[231],pp186[231],pp187[231],pp188[231],pp189[231],pp190[231],pp191[231],pp192[231],pp193[231],pp194[231],pp195[231],pp196[231],pp197[231],pp198[231],pp199[231],pp200[231],pp201[231],pp202[231],pp203[231],pp204[231]};
    assign in141_2 = {pp35[41],pp35[42],pp35[43],pp35[44],pp35[45],pp35[46],pp35[47],pp35[48],pp35[49],pp35[50],pp35[51],pp35[52],pp35[53],pp35[54],pp35[55],pp35[56],pp35[57],pp35[58],pp35[59],pp35[60],pp35[61],pp35[62],pp35[63],pp35[64],pp34[66],pp33[68],pp32[70],pp31[72],pp30[74],pp29[76],pp28[78],pp27[80],pp26[82],pp25[84],pp24[86],pp23[88],pp22[90],pp21[92],pp20[94],pp19[96],pp18[98],pp9[108],pp7[111],pp5[114],pp3[117],pp1[120],pp112[10],pp111[12],pp110[14],pp109[16],pp108[18],pp107[20],pp108[20],pp109[20],pp110[20],pp111[20],pp112[20],pp113[20],pp114[20],pp115[20],pp116[20],pp117[20],pp118[20],pp119[20],pp120[20],pp121[20],pp122[20],pp123[20],pp124[20],pp125[20],pp126[20],pp127[20],pp128[20],pp129[20],pp130[20],pp131[20],pp132[20],pp133[20],pp134[20],pp135[20],pp136[20],pp137[20],pp138[20],pp139[20],pp140[20],pp141[20],pp142[20],pp143[20],pp144[20],pp145[20],pp146[20],pp147[20],pp148[20],pp149[20],pp150[20],pp151[20],pp152[20],pp153[20],pp154[20],pp155[20],pp156[20],pp157[20],pp158[20],pp159[20],pp160[20],pp161[20],pp162[20],pp163[20],pp164[20],pp165[20],pp166[20],pp167[20],pp168[20],pp169[20],pp170[20],pp171[20],pp172[20],pp173[20],pp174[20],pp175[20],pp176[20],pp177[20],pp178[20],pp179[20],pp181[19],pp183[18],pp185[17],pp187[16],pp189[15],pp191[14],pp193[13],pp195[12],pp197[11],pp199[10],s129[146],s130[146],s131[146],s132[146],s133[146],s134[146],s135[146],s136[146],s137[146],s138[146],s139[146],s140[146],pp0[222],pp1[222],pp2[222],pp3[222],pp4[222],pp5[222],pp6[222],pp7[222],pp8[222],pp9[222],pp223[9],pp225[8],pp227[7],pp229[6],pp231[5],pp233[4],pp235[3],pp237[2],pp239[1],pp241[0],s10[105],s11[105],s12[105],s13[105],s14[105],s15[105],s16[105],s17[105],s18[105],s19[105],s20[105],s21[105],s22[105],s23[105],s24[105],s23[107],s22[109],s21[111],s20[113],s19[115],s18[117],s17[119],s16[121],s15[123],s14[125],s13[127],s12[129],s11[131],s10[133],s140[196],s139[198],s138[200],s137[202],s136[204],s135[206],s134[208],s133[210],s132[212],s131[214],s130[216],s129[218],pp255[28],pp254[30],pp253[32],pp252[34],pp251[36],pp250[38],pp249[40],pp248[42],pp247[44],pp246[46],pp245[48],pp244[50],pp243[52],pp242[54],pp241[56],pp240[58],pp239[60],pp238[62],pp237[64],pp236[66],pp235[68],pp234[70],pp233[72],pp232[74],pp231[76],pp230[78],pp229[80],pp228[82],pp227[84],pp226[86],pp225[88],pp224[90],pp223[92],pp222[94],pp221[96],pp220[98],pp99[220],pp97[223],pp95[226],pp93[229],pp91[232],pp89[235],pp87[238],pp85[241],pp83[244],pp81[247],pp79[250],pp77[253],pp231[100],pp229[103],pp227[106],pp225[109],pp223[112],pp221[115],pp219[118],pp217[121],pp215[124],pp213[127],pp211[130],pp209[133],pp207[136],pp205[139],pp203[142],pp201[145],pp199[148],pp197[151],pp195[154],pp193[157],pp191[160],pp189[163],pp187[166],pp185[169],pp183[172],pp182[174],pp181[176],pp180[178],pp179[180],pp178[182],pp177[184],pp176[186],pp175[188],pp174[190],pp173[192],pp172[194],pp171[196],pp170[198],pp169[200],pp168[202],pp167[204],pp166[206],pp165[208],pp164[210],pp163[212],pp162[214],pp161[216],pp160[218],pp159[220],pp158[222],pp157[224],pp156[226],pp155[228],pp154[230],pp155[230],pp156[230],pp157[230],pp158[230],pp159[230],pp160[230],pp161[230],pp162[230],pp163[230],pp164[230],pp165[230],pp166[230],pp167[230],pp168[230],pp169[230],pp170[230],pp171[230],pp172[230],pp173[230],pp174[230],pp175[230],pp176[230],pp177[230],pp178[230],pp179[230],pp180[230],pp181[230],pp182[230],pp183[230],pp184[230],pp185[230],pp186[230],pp187[230],pp188[230],pp189[230],pp190[230],pp191[230],pp192[230],pp193[230],pp194[230],pp195[230],pp196[230],pp197[230],pp198[230],pp199[230],pp200[230],pp201[230],pp202[230],pp203[230],pp204[230],pp205[230]};
    CLA_360 KS_141(s141, c141, in141_1, in141_2);
    wire[357:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp36[41],pp36[42],pp36[43],pp36[44],pp36[45],pp36[46],pp36[47],pp36[48],pp36[49],pp36[50],pp36[51],pp36[52],pp36[53],pp36[54],pp36[55],pp36[56],pp36[57],pp36[58],pp36[59],pp36[60],pp36[61],pp36[62],pp36[63],pp35[65],pp34[67],pp33[69],pp32[71],pp31[73],pp30[75],pp29[77],pp28[79],pp27[81],pp26[83],pp25[85],pp24[87],pp23[89],pp22[91],pp21[93],pp20[95],pp19[97],pp18[99],pp8[110],pp6[113],pp4[116],pp2[119],pp0[122],pp112[11],pp111[13],pp110[15],pp109[17],pp108[19],pp109[19],pp110[19],pp111[19],pp112[19],pp113[19],pp114[19],pp115[19],pp116[19],pp117[19],pp118[19],pp119[19],pp120[19],pp121[19],pp122[19],pp123[19],pp124[19],pp125[19],pp126[19],pp127[19],pp128[19],pp129[19],pp130[19],pp131[19],pp132[19],pp133[19],pp134[19],pp135[19],pp136[19],pp137[19],pp138[19],pp139[19],pp140[19],pp141[19],pp142[19],pp143[19],pp144[19],pp145[19],pp146[19],pp147[19],pp148[19],pp149[19],pp150[19],pp151[19],pp152[19],pp153[19],pp154[19],pp155[19],pp156[19],pp157[19],pp158[19],pp159[19],pp160[19],pp161[19],pp162[19],pp163[19],pp164[19],pp165[19],pp166[19],pp167[19],pp168[19],pp169[19],pp170[19],pp171[19],pp172[19],pp173[19],pp174[19],pp175[19],pp176[19],pp177[19],pp178[19],pp179[19],pp180[19],pp182[18],pp184[17],pp186[16],pp188[15],pp190[14],pp192[13],pp194[12],pp196[11],pp198[10],s129[145],s130[145],s131[145],s132[145],s133[145],s134[145],s135[145],s136[145],s137[145],s138[145],s139[145],s140[145],s141[145],s141[146],s141[147],s141[148],s141[149],s141[150],s141[151],s141[152],s141[153],s141[154],s141[155],s141[156],s141[157],s141[158],s141[159],s141[160],s141[161],s141[162],s141[163],s141[164],s141[165],s141[166],s141[167],s141[168],s141[169],s141[170],s141[171],s141[172],s141[173],s141[174],s141[175],s141[176],s141[177],s141[178],s141[179],s141[180],s141[181],s141[182],s141[183],s141[184],s141[185],s141[186],s141[187],s141[188],s141[189],s141[190],s141[191],s141[192],s141[193],s141[194],s141[195],s140[197],s139[199],s138[201],s137[203],s136[205],s135[207],s134[209],s133[211],s132[213],s131[215],s130[217],s129[219],pp255[29],pp254[31],pp253[33],pp252[35],pp251[37],pp250[39],pp249[41],pp248[43],pp247[45],pp246[47],pp245[49],pp244[51],pp243[53],pp242[55],pp241[57],pp240[59],pp239[61],pp238[63],pp237[65],pp236[67],pp235[69],pp234[71],pp233[73],pp232[75],pp231[77],pp230[79],pp229[81],pp228[83],pp227[85],pp226[87],pp225[89],pp224[91],pp223[93],pp222[95],pp221[97],pp220[99],pp98[222],pp96[225],pp94[228],pp92[231],pp90[234],pp88[237],pp86[240],pp84[243],pp82[246],pp80[249],pp78[252],pp76[255],pp230[102],pp228[105],pp226[108],pp224[111],pp222[114],pp220[117],pp218[120],pp216[123],pp214[126],pp212[129],pp210[132],pp208[135],pp206[138],pp204[141],pp202[144],pp200[147],pp198[150],pp196[153],pp194[156],pp192[159],pp190[162],pp188[165],pp186[168],pp184[171],pp183[173],pp182[175],pp181[177],pp180[179],pp179[181],pp178[183],pp177[185],pp176[187],pp175[189],pp174[191],pp173[193],pp172[195],pp171[197],pp170[199],pp169[201],pp168[203],pp167[205],pp166[207],pp165[209],pp164[211],pp163[213],pp162[215],pp161[217],pp160[219],pp159[221],pp158[223],pp157[225],pp156[227],pp155[229],pp156[229],pp157[229],pp158[229],pp159[229],pp160[229],pp161[229],pp162[229],pp163[229],pp164[229],pp165[229],pp166[229],pp167[229],pp168[229],pp169[229],pp170[229],pp171[229],pp172[229],pp173[229],pp174[229],pp175[229],pp176[229],pp177[229],pp178[229],pp179[229],pp180[229],pp181[229],pp182[229],pp183[229],pp184[229],pp185[229],pp186[229],pp187[229],pp188[229],pp189[229],pp190[229],pp191[229],pp192[229],pp193[229],pp194[229],pp195[229],pp196[229],pp197[229],pp198[229],pp199[229],pp200[229],pp201[229],pp202[229],pp203[229],pp204[229],pp205[229]};
    assign in142_2 = {pp37[40],pp37[41],pp37[42],pp37[43],pp37[44],pp37[45],pp37[46],pp37[47],pp37[48],pp37[49],pp37[50],pp37[51],pp37[52],pp37[53],pp37[54],pp37[55],pp37[56],pp37[57],pp37[58],pp37[59],pp37[60],pp37[61],pp37[62],pp36[64],pp35[66],pp34[68],pp33[70],pp32[72],pp31[74],pp30[76],pp29[78],pp28[80],pp27[82],pp26[84],pp25[86],pp24[88],pp23[90],pp22[92],pp21[94],pp20[96],pp19[98],pp9[109],pp7[112],pp5[115],pp3[118],pp1[121],pp113[10],pp112[12],pp111[14],pp110[16],pp109[18],pp110[18],pp111[18],pp112[18],pp113[18],pp114[18],pp115[18],pp116[18],pp117[18],pp118[18],pp119[18],pp120[18],pp121[18],pp122[18],pp123[18],pp124[18],pp125[18],pp126[18],pp127[18],pp128[18],pp129[18],pp130[18],pp131[18],pp132[18],pp133[18],pp134[18],pp135[18],pp136[18],pp137[18],pp138[18],pp139[18],pp140[18],pp141[18],pp142[18],pp143[18],pp144[18],pp145[18],pp146[18],pp147[18],pp148[18],pp149[18],pp150[18],pp151[18],pp152[18],pp153[18],pp154[18],pp155[18],pp156[18],pp157[18],pp158[18],pp159[18],pp160[18],pp161[18],pp162[18],pp163[18],pp164[18],pp165[18],pp166[18],pp167[18],pp168[18],pp169[18],pp170[18],pp171[18],pp172[18],pp173[18],pp174[18],pp175[18],pp176[18],pp177[18],pp178[18],pp179[18],pp180[18],pp181[18],pp183[17],pp185[16],pp187[15],pp189[14],pp191[13],pp193[12],pp195[11],pp197[10],s129[144],s130[144],s131[144],s132[144],s133[144],s134[144],s135[144],s136[144],s137[144],s138[144],s139[144],s140[144],s141[144],pp0[221],pp1[221],pp2[221],pp3[221],pp4[221],pp5[221],pp6[221],pp7[221],pp8[221],pp9[221],pp222[9],pp224[8],pp226[7],pp228[6],pp230[5],pp232[4],pp234[3],pp236[2],pp238[1],pp240[0],s10[104],s11[104],s12[104],s13[104],s14[104],s15[104],s16[104],s17[104],s18[104],s19[104],s20[104],s21[104],s22[104],s23[104],s24[104],s25[104],s24[106],s23[108],s22[110],s21[112],s20[114],s19[116],s18[118],s17[120],s16[122],s15[124],s14[126],s13[128],s12[130],s11[132],s10[134],s141[196],s140[198],s139[200],s138[202],s137[204],s136[206],s135[208],s134[210],s133[212],s132[214],s131[216],s130[218],s129[220],pp255[30],pp254[32],pp253[34],pp252[36],pp251[38],pp250[40],pp249[42],pp248[44],pp247[46],pp246[48],pp245[50],pp244[52],pp243[54],pp242[56],pp241[58],pp240[60],pp239[62],pp238[64],pp237[66],pp236[68],pp235[70],pp234[72],pp233[74],pp232[76],pp231[78],pp230[80],pp229[82],pp228[84],pp227[86],pp226[88],pp225[90],pp224[92],pp223[94],pp222[96],pp221[98],pp99[221],pp97[224],pp95[227],pp93[230],pp91[233],pp89[236],pp87[239],pp85[242],pp83[245],pp81[248],pp79[251],pp77[254],pp231[101],pp229[104],pp227[107],pp225[110],pp223[113],pp221[116],pp219[119],pp217[122],pp215[125],pp213[128],pp211[131],pp209[134],pp207[137],pp205[140],pp203[143],pp201[146],pp199[149],pp197[152],pp195[155],pp193[158],pp191[161],pp189[164],pp187[167],pp185[170],pp184[172],pp183[174],pp182[176],pp181[178],pp180[180],pp179[182],pp178[184],pp177[186],pp176[188],pp175[190],pp174[192],pp173[194],pp172[196],pp171[198],pp170[200],pp169[202],pp168[204],pp167[206],pp166[208],pp165[210],pp164[212],pp163[214],pp162[216],pp161[218],pp160[220],pp159[222],pp158[224],pp157[226],pp156[228],pp157[228],pp158[228],pp159[228],pp160[228],pp161[228],pp162[228],pp163[228],pp164[228],pp165[228],pp166[228],pp167[228],pp168[228],pp169[228],pp170[228],pp171[228],pp172[228],pp173[228],pp174[228],pp175[228],pp176[228],pp177[228],pp178[228],pp179[228],pp180[228],pp181[228],pp182[228],pp183[228],pp184[228],pp185[228],pp186[228],pp187[228],pp188[228],pp189[228],pp190[228],pp191[228],pp192[228],pp193[228],pp194[228],pp195[228],pp196[228],pp197[228],pp198[228],pp199[228],pp200[228],pp201[228],pp202[228],pp203[228],pp204[228],pp205[228],pp206[228]};
    CLA_358 KS_142(s142, c142, in142_1, in142_2);
    wire[355:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp38[40],pp38[41],pp38[42],pp38[43],pp38[44],pp38[45],pp38[46],pp38[47],pp38[48],pp38[49],pp38[50],pp38[51],pp38[52],pp38[53],pp38[54],pp38[55],pp38[56],pp38[57],pp38[58],pp38[59],pp38[60],pp38[61],pp37[63],pp36[65],pp35[67],pp34[69],pp33[71],pp32[73],pp31[75],pp30[77],pp29[79],pp28[81],pp27[83],pp26[85],pp25[87],pp24[89],pp23[91],pp22[93],pp21[95],pp20[97],pp19[99],pp8[111],pp6[114],pp4[117],pp2[120],pp0[123],pp113[11],pp112[13],pp111[15],pp110[17],pp111[17],pp112[17],pp113[17],pp114[17],pp115[17],pp116[17],pp117[17],pp118[17],pp119[17],pp120[17],pp121[17],pp122[17],pp123[17],pp124[17],pp125[17],pp126[17],pp127[17],pp128[17],pp129[17],pp130[17],pp131[17],pp132[17],pp133[17],pp134[17],pp135[17],pp136[17],pp137[17],pp138[17],pp139[17],pp140[17],pp141[17],pp142[17],pp143[17],pp144[17],pp145[17],pp146[17],pp147[17],pp148[17],pp149[17],pp150[17],pp151[17],pp152[17],pp153[17],pp154[17],pp155[17],pp156[17],pp157[17],pp158[17],pp159[17],pp160[17],pp161[17],pp162[17],pp163[17],pp164[17],pp165[17],pp166[17],pp167[17],pp168[17],pp169[17],pp170[17],pp171[17],pp172[17],pp173[17],pp174[17],pp175[17],pp176[17],pp177[17],pp178[17],pp179[17],pp180[17],pp181[17],pp182[17],pp184[16],pp186[15],pp188[14],pp190[13],pp192[12],pp194[11],pp196[10],s129[143],s130[143],s131[143],s132[143],s133[143],s134[143],s135[143],s136[143],s137[143],s138[143],s139[143],s140[143],s141[143],s142[143],s142[144],s142[145],s142[146],s142[147],s142[148],s142[149],s142[150],s142[151],s142[152],s142[153],s142[154],s142[155],s142[156],s142[157],s142[158],s142[159],s142[160],s142[161],s142[162],s142[163],s142[164],s142[165],s142[166],s142[167],s142[168],s142[169],s142[170],s142[171],s142[172],s142[173],s142[174],s142[175],s142[176],s142[177],s142[178],s142[179],s142[180],s142[181],s142[182],s142[183],s142[184],s142[185],s142[186],s142[187],s142[188],s142[189],s142[190],s142[191],s142[192],s142[193],s142[194],s142[195],s141[197],s140[199],s139[201],s138[203],s137[205],s136[207],s135[209],s134[211],s133[213],s132[215],s131[217],s130[219],s129[221],pp255[31],pp254[33],pp253[35],pp252[37],pp251[39],pp250[41],pp249[43],pp248[45],pp247[47],pp246[49],pp245[51],pp244[53],pp243[55],pp242[57],pp241[59],pp240[61],pp239[63],pp238[65],pp237[67],pp236[69],pp235[71],pp234[73],pp233[75],pp232[77],pp231[79],pp230[81],pp229[83],pp228[85],pp227[87],pp226[89],pp225[91],pp224[93],pp223[95],pp222[97],pp221[99],pp98[223],pp96[226],pp94[229],pp92[232],pp90[235],pp88[238],pp86[241],pp84[244],pp82[247],pp80[250],pp78[253],pp232[100],pp230[103],pp228[106],pp226[109],pp224[112],pp222[115],pp220[118],pp218[121],pp216[124],pp214[127],pp212[130],pp210[133],pp208[136],pp206[139],pp204[142],pp202[145],pp200[148],pp198[151],pp196[154],pp194[157],pp192[160],pp190[163],pp188[166],pp186[169],pp185[171],pp184[173],pp183[175],pp182[177],pp181[179],pp180[181],pp179[183],pp178[185],pp177[187],pp176[189],pp175[191],pp174[193],pp173[195],pp172[197],pp171[199],pp170[201],pp169[203],pp168[205],pp167[207],pp166[209],pp165[211],pp164[213],pp163[215],pp162[217],pp161[219],pp160[221],pp159[223],pp158[225],pp157[227],pp158[227],pp159[227],pp160[227],pp161[227],pp162[227],pp163[227],pp164[227],pp165[227],pp166[227],pp167[227],pp168[227],pp169[227],pp170[227],pp171[227],pp172[227],pp173[227],pp174[227],pp175[227],pp176[227],pp177[227],pp178[227],pp179[227],pp180[227],pp181[227],pp182[227],pp183[227],pp184[227],pp185[227],pp186[227],pp187[227],pp188[227],pp189[227],pp190[227],pp191[227],pp192[227],pp193[227],pp194[227],pp195[227],pp196[227],pp197[227],pp198[227],pp199[227],pp200[227],pp201[227],pp202[227],pp203[227],pp204[227],pp205[227],pp206[227]};
    assign in143_2 = {pp39[39],pp39[40],pp39[41],pp39[42],pp39[43],pp39[44],pp39[45],pp39[46],pp39[47],pp39[48],pp39[49],pp39[50],pp39[51],pp39[52],pp39[53],pp39[54],pp39[55],pp39[56],pp39[57],pp39[58],pp39[59],pp39[60],pp38[62],pp37[64],pp36[66],pp35[68],pp34[70],pp33[72],pp32[74],pp31[76],pp30[78],pp29[80],pp28[82],pp27[84],pp26[86],pp25[88],pp24[90],pp23[92],pp22[94],pp21[96],pp20[98],pp9[110],pp7[113],pp5[116],pp3[119],pp1[122],pp114[10],pp113[12],pp112[14],pp111[16],pp112[16],pp113[16],pp114[16],pp115[16],pp116[16],pp117[16],pp118[16],pp119[16],pp120[16],pp121[16],pp122[16],pp123[16],pp124[16],pp125[16],pp126[16],pp127[16],pp128[16],pp129[16],pp130[16],pp131[16],pp132[16],pp133[16],pp134[16],pp135[16],pp136[16],pp137[16],pp138[16],pp139[16],pp140[16],pp141[16],pp142[16],pp143[16],pp144[16],pp145[16],pp146[16],pp147[16],pp148[16],pp149[16],pp150[16],pp151[16],pp152[16],pp153[16],pp154[16],pp155[16],pp156[16],pp157[16],pp158[16],pp159[16],pp160[16],pp161[16],pp162[16],pp163[16],pp164[16],pp165[16],pp166[16],pp167[16],pp168[16],pp169[16],pp170[16],pp171[16],pp172[16],pp173[16],pp174[16],pp175[16],pp176[16],pp177[16],pp178[16],pp179[16],pp180[16],pp181[16],pp182[16],pp183[16],pp185[15],pp187[14],pp189[13],pp191[12],pp193[11],pp195[10],s129[142],s130[142],s131[142],s132[142],s133[142],s134[142],s135[142],s136[142],s137[142],s138[142],s139[142],s140[142],s141[142],s142[142],pp0[220],pp1[220],pp2[220],pp3[220],pp4[220],pp5[220],pp6[220],pp7[220],pp8[220],pp9[220],pp221[9],pp223[8],pp225[7],pp227[6],pp229[5],pp231[4],pp233[3],pp235[2],pp237[1],pp239[0],s10[103],s11[103],s12[103],s13[103],s14[103],s15[103],s16[103],s17[103],s18[103],s19[103],s20[103],s21[103],s22[103],s23[103],s24[103],s25[103],s26[103],s25[105],s24[107],s23[109],s22[111],s21[113],s20[115],s19[117],s18[119],s17[121],s16[123],s15[125],s14[127],s13[129],s12[131],s11[133],s10[135],s142[196],s141[198],s140[200],s139[202],s138[204],s137[206],s136[208],s135[210],s134[212],s133[214],s132[216],s131[218],s130[220],s129[222],pp255[32],pp254[34],pp253[36],pp252[38],pp251[40],pp250[42],pp249[44],pp248[46],pp247[48],pp246[50],pp245[52],pp244[54],pp243[56],pp242[58],pp241[60],pp240[62],pp239[64],pp238[66],pp237[68],pp236[70],pp235[72],pp234[74],pp233[76],pp232[78],pp231[80],pp230[82],pp229[84],pp228[86],pp227[88],pp226[90],pp225[92],pp224[94],pp223[96],pp222[98],pp99[222],pp97[225],pp95[228],pp93[231],pp91[234],pp89[237],pp87[240],pp85[243],pp83[246],pp81[249],pp79[252],pp77[255],pp231[102],pp229[105],pp227[108],pp225[111],pp223[114],pp221[117],pp219[120],pp217[123],pp215[126],pp213[129],pp211[132],pp209[135],pp207[138],pp205[141],pp203[144],pp201[147],pp199[150],pp197[153],pp195[156],pp193[159],pp191[162],pp189[165],pp187[168],pp186[170],pp185[172],pp184[174],pp183[176],pp182[178],pp181[180],pp180[182],pp179[184],pp178[186],pp177[188],pp176[190],pp175[192],pp174[194],pp173[196],pp172[198],pp171[200],pp170[202],pp169[204],pp168[206],pp167[208],pp166[210],pp165[212],pp164[214],pp163[216],pp162[218],pp161[220],pp160[222],pp159[224],pp158[226],pp159[226],pp160[226],pp161[226],pp162[226],pp163[226],pp164[226],pp165[226],pp166[226],pp167[226],pp168[226],pp169[226],pp170[226],pp171[226],pp172[226],pp173[226],pp174[226],pp175[226],pp176[226],pp177[226],pp178[226],pp179[226],pp180[226],pp181[226],pp182[226],pp183[226],pp184[226],pp185[226],pp186[226],pp187[226],pp188[226],pp189[226],pp190[226],pp191[226],pp192[226],pp193[226],pp194[226],pp195[226],pp196[226],pp197[226],pp198[226],pp199[226],pp200[226],pp201[226],pp202[226],pp203[226],pp204[226],pp205[226],pp206[226],pp207[226]};
    CLA_356 KS_143(s143, c143, in143_1, in143_2);
    wire[353:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp40[39],pp40[40],pp40[41],pp40[42],pp40[43],pp40[44],pp40[45],pp40[46],pp40[47],pp40[48],pp40[49],pp40[50],pp40[51],pp40[52],pp40[53],pp40[54],pp40[55],pp40[56],pp40[57],pp40[58],pp40[59],pp39[61],pp38[63],pp37[65],pp36[67],pp35[69],pp34[71],pp33[73],pp32[75],pp31[77],pp30[79],pp29[81],pp28[83],pp27[85],pp26[87],pp25[89],pp24[91],pp23[93],pp22[95],pp21[97],pp20[99],pp8[112],pp6[115],pp4[118],pp2[121],pp0[124],pp114[11],pp113[13],pp112[15],pp113[15],pp114[15],pp115[15],pp116[15],pp117[15],pp118[15],pp119[15],pp120[15],pp121[15],pp122[15],pp123[15],pp124[15],pp125[15],pp126[15],pp127[15],pp128[15],pp129[15],pp130[15],pp131[15],pp132[15],pp133[15],pp134[15],pp135[15],pp136[15],pp137[15],pp138[15],pp139[15],pp140[15],pp141[15],pp142[15],pp143[15],pp144[15],pp145[15],pp146[15],pp147[15],pp148[15],pp149[15],pp150[15],pp151[15],pp152[15],pp153[15],pp154[15],pp155[15],pp156[15],pp157[15],pp158[15],pp159[15],pp160[15],pp161[15],pp162[15],pp163[15],pp164[15],pp165[15],pp166[15],pp167[15],pp168[15],pp169[15],pp170[15],pp171[15],pp172[15],pp173[15],pp174[15],pp175[15],pp176[15],pp177[15],pp178[15],pp179[15],pp180[15],pp181[15],pp182[15],pp183[15],pp184[15],pp186[14],pp188[13],pp190[12],pp192[11],pp194[10],s129[141],s130[141],s131[141],s132[141],s133[141],s134[141],s135[141],s136[141],s137[141],s138[141],s139[141],s140[141],s141[141],s142[141],s143[141],s143[142],s143[143],s143[144],s143[145],s143[146],s143[147],s143[148],s143[149],s143[150],s143[151],s143[152],s143[153],s143[154],s143[155],s143[156],s143[157],s143[158],s143[159],s143[160],s143[161],s143[162],s143[163],s143[164],s143[165],s143[166],s143[167],s143[168],s143[169],s143[170],s143[171],s143[172],s143[173],s143[174],s143[175],s143[176],s143[177],s143[178],s143[179],s143[180],s143[181],s143[182],s143[183],s143[184],s143[185],s143[186],s143[187],s143[188],s143[189],s143[190],s143[191],s143[192],s143[193],s143[194],s143[195],s142[197],s141[199],s140[201],s139[203],s138[205],s137[207],s136[209],s135[211],s134[213],s133[215],s132[217],s131[219],s130[221],s129[223],pp255[33],pp254[35],pp253[37],pp252[39],pp251[41],pp250[43],pp249[45],pp248[47],pp247[49],pp246[51],pp245[53],pp244[55],pp243[57],pp242[59],pp241[61],pp240[63],pp239[65],pp238[67],pp237[69],pp236[71],pp235[73],pp234[75],pp233[77],pp232[79],pp231[81],pp230[83],pp229[85],pp228[87],pp227[89],pp226[91],pp225[93],pp224[95],pp223[97],pp222[99],pp98[224],pp96[227],pp94[230],pp92[233],pp90[236],pp88[239],pp86[242],pp84[245],pp82[248],pp80[251],pp78[254],pp232[101],pp230[104],pp228[107],pp226[110],pp224[113],pp222[116],pp220[119],pp218[122],pp216[125],pp214[128],pp212[131],pp210[134],pp208[137],pp206[140],pp204[143],pp202[146],pp200[149],pp198[152],pp196[155],pp194[158],pp192[161],pp190[164],pp188[167],pp187[169],pp186[171],pp185[173],pp184[175],pp183[177],pp182[179],pp181[181],pp180[183],pp179[185],pp178[187],pp177[189],pp176[191],pp175[193],pp174[195],pp173[197],pp172[199],pp171[201],pp170[203],pp169[205],pp168[207],pp167[209],pp166[211],pp165[213],pp164[215],pp163[217],pp162[219],pp161[221],pp160[223],pp159[225],pp160[225],pp161[225],pp162[225],pp163[225],pp164[225],pp165[225],pp166[225],pp167[225],pp168[225],pp169[225],pp170[225],pp171[225],pp172[225],pp173[225],pp174[225],pp175[225],pp176[225],pp177[225],pp178[225],pp179[225],pp180[225],pp181[225],pp182[225],pp183[225],pp184[225],pp185[225],pp186[225],pp187[225],pp188[225],pp189[225],pp190[225],pp191[225],pp192[225],pp193[225],pp194[225],pp195[225],pp196[225],pp197[225],pp198[225],pp199[225],pp200[225],pp201[225],pp202[225],pp203[225],pp204[225],pp205[225],pp206[225],pp207[225]};
    assign in144_2 = {pp41[38],pp41[39],pp41[40],pp41[41],pp41[42],pp41[43],pp41[44],pp41[45],pp41[46],pp41[47],pp41[48],pp41[49],pp41[50],pp41[51],pp41[52],pp41[53],pp41[54],pp41[55],pp41[56],pp41[57],pp41[58],pp40[60],pp39[62],pp38[64],pp37[66],pp36[68],pp35[70],pp34[72],pp33[74],pp32[76],pp31[78],pp30[80],pp29[82],pp28[84],pp27[86],pp26[88],pp25[90],pp24[92],pp23[94],pp22[96],pp21[98],pp9[111],pp7[114],pp5[117],pp3[120],pp1[123],pp115[10],pp114[12],pp113[14],pp114[14],pp115[14],pp116[14],pp117[14],pp118[14],pp119[14],pp120[14],pp121[14],pp122[14],pp123[14],pp124[14],pp125[14],pp126[14],pp127[14],pp128[14],pp129[14],pp130[14],pp131[14],pp132[14],pp133[14],pp134[14],pp135[14],pp136[14],pp137[14],pp138[14],pp139[14],pp140[14],pp141[14],pp142[14],pp143[14],pp144[14],pp145[14],pp146[14],pp147[14],pp148[14],pp149[14],pp150[14],pp151[14],pp152[14],pp153[14],pp154[14],pp155[14],pp156[14],pp157[14],pp158[14],pp159[14],pp160[14],pp161[14],pp162[14],pp163[14],pp164[14],pp165[14],pp166[14],pp167[14],pp168[14],pp169[14],pp170[14],pp171[14],pp172[14],pp173[14],pp174[14],pp175[14],pp176[14],pp177[14],pp178[14],pp179[14],pp180[14],pp181[14],pp182[14],pp183[14],pp184[14],pp185[14],pp187[13],pp189[12],pp191[11],pp193[10],s129[140],s130[140],s131[140],s132[140],s133[140],s134[140],s135[140],s136[140],s137[140],s138[140],s139[140],s140[140],s141[140],s142[140],s143[140],pp0[219],pp1[219],pp2[219],pp3[219],pp4[219],pp5[219],pp6[219],pp7[219],pp8[219],pp9[219],pp220[9],pp222[8],pp224[7],pp226[6],pp228[5],pp230[4],pp232[3],pp234[2],pp236[1],pp238[0],s10[102],s11[102],s12[102],s13[102],s14[102],s15[102],s16[102],s17[102],s18[102],s19[102],s20[102],s21[102],s22[102],s23[102],s24[102],s25[102],s26[102],s27[102],s26[104],s25[106],s24[108],s23[110],s22[112],s21[114],s20[116],s19[118],s18[120],s17[122],s16[124],s15[126],s14[128],s13[130],s12[132],s11[134],s10[136],s143[196],s142[198],s141[200],s140[202],s139[204],s138[206],s137[208],s136[210],s135[212],s134[214],s133[216],s132[218],s131[220],s130[222],s129[224],pp255[34],pp254[36],pp253[38],pp252[40],pp251[42],pp250[44],pp249[46],pp248[48],pp247[50],pp246[52],pp245[54],pp244[56],pp243[58],pp242[60],pp241[62],pp240[64],pp239[66],pp238[68],pp237[70],pp236[72],pp235[74],pp234[76],pp233[78],pp232[80],pp231[82],pp230[84],pp229[86],pp228[88],pp227[90],pp226[92],pp225[94],pp224[96],pp223[98],pp99[223],pp97[226],pp95[229],pp93[232],pp91[235],pp89[238],pp87[241],pp85[244],pp83[247],pp81[250],pp79[253],pp233[100],pp231[103],pp229[106],pp227[109],pp225[112],pp223[115],pp221[118],pp219[121],pp217[124],pp215[127],pp213[130],pp211[133],pp209[136],pp207[139],pp205[142],pp203[145],pp201[148],pp199[151],pp197[154],pp195[157],pp193[160],pp191[163],pp189[166],pp188[168],pp187[170],pp186[172],pp185[174],pp184[176],pp183[178],pp182[180],pp181[182],pp180[184],pp179[186],pp178[188],pp177[190],pp176[192],pp175[194],pp174[196],pp173[198],pp172[200],pp171[202],pp170[204],pp169[206],pp168[208],pp167[210],pp166[212],pp165[214],pp164[216],pp163[218],pp162[220],pp161[222],pp160[224],pp161[224],pp162[224],pp163[224],pp164[224],pp165[224],pp166[224],pp167[224],pp168[224],pp169[224],pp170[224],pp171[224],pp172[224],pp173[224],pp174[224],pp175[224],pp176[224],pp177[224],pp178[224],pp179[224],pp180[224],pp181[224],pp182[224],pp183[224],pp184[224],pp185[224],pp186[224],pp187[224],pp188[224],pp189[224],pp190[224],pp191[224],pp192[224],pp193[224],pp194[224],pp195[224],pp196[224],pp197[224],pp198[224],pp199[224],pp200[224],pp201[224],pp202[224],pp203[224],pp204[224],pp205[224],pp206[224],pp207[224],pp208[224]};
    CLA_354 KS_144(s144, c144, in144_1, in144_2);
    wire[351:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp42[38],pp42[39],pp42[40],pp42[41],pp42[42],pp42[43],pp42[44],pp42[45],pp42[46],pp42[47],pp42[48],pp42[49],pp42[50],pp42[51],pp42[52],pp42[53],pp42[54],pp42[55],pp42[56],pp42[57],pp41[59],pp40[61],pp39[63],pp38[65],pp37[67],pp36[69],pp35[71],pp34[73],pp33[75],pp32[77],pp31[79],pp30[81],pp29[83],pp28[85],pp27[87],pp26[89],pp25[91],pp24[93],pp23[95],pp22[97],pp21[99],pp8[113],pp6[116],pp4[119],pp2[122],pp0[125],pp115[11],pp114[13],pp115[13],pp116[13],pp117[13],pp118[13],pp119[13],pp120[13],pp121[13],pp122[13],pp123[13],pp124[13],pp125[13],pp126[13],pp127[13],pp128[13],pp129[13],pp130[13],pp131[13],pp132[13],pp133[13],pp134[13],pp135[13],pp136[13],pp137[13],pp138[13],pp139[13],pp140[13],pp141[13],pp142[13],pp143[13],pp144[13],pp145[13],pp146[13],pp147[13],pp148[13],pp149[13],pp150[13],pp151[13],pp152[13],pp153[13],pp154[13],pp155[13],pp156[13],pp157[13],pp158[13],pp159[13],pp160[13],pp161[13],pp162[13],pp163[13],pp164[13],pp165[13],pp166[13],pp167[13],pp168[13],pp169[13],pp170[13],pp171[13],pp172[13],pp173[13],pp174[13],pp175[13],pp176[13],pp177[13],pp178[13],pp179[13],pp180[13],pp181[13],pp182[13],pp183[13],pp184[13],pp185[13],pp186[13],pp188[12],pp190[11],pp192[10],s129[139],s130[139],s131[139],s132[139],s133[139],s134[139],s135[139],s136[139],s137[139],s138[139],s139[139],s140[139],s141[139],s142[139],s143[139],s144[139],s144[140],s144[141],s144[142],s144[143],s144[144],s144[145],s144[146],s144[147],s144[148],s144[149],s144[150],s144[151],s144[152],s144[153],s144[154],s144[155],s144[156],s144[157],s144[158],s144[159],s144[160],s144[161],s144[162],s144[163],s144[164],s144[165],s144[166],s144[167],s144[168],s144[169],s144[170],s144[171],s144[172],s144[173],s144[174],s144[175],s144[176],s144[177],s144[178],s144[179],s144[180],s144[181],s144[182],s144[183],s144[184],s144[185],s144[186],s144[187],s144[188],s144[189],s144[190],s144[191],s144[192],s144[193],s144[194],s144[195],s143[197],s142[199],s141[201],s140[203],s139[205],s138[207],s137[209],s136[211],s135[213],s134[215],s133[217],s132[219],s131[221],s130[223],s129[225],pp255[35],pp254[37],pp253[39],pp252[41],pp251[43],pp250[45],pp249[47],pp248[49],pp247[51],pp246[53],pp245[55],pp244[57],pp243[59],pp242[61],pp241[63],pp240[65],pp239[67],pp238[69],pp237[71],pp236[73],pp235[75],pp234[77],pp233[79],pp232[81],pp231[83],pp230[85],pp229[87],pp228[89],pp227[91],pp226[93],pp225[95],pp224[97],pp223[99],pp98[225],pp96[228],pp94[231],pp92[234],pp90[237],pp88[240],pp86[243],pp84[246],pp82[249],pp80[252],pp78[255],pp232[102],pp230[105],pp228[108],pp226[111],pp224[114],pp222[117],pp220[120],pp218[123],pp216[126],pp214[129],pp212[132],pp210[135],pp208[138],pp206[141],pp204[144],pp202[147],pp200[150],pp198[153],pp196[156],pp194[159],pp192[162],pp190[165],pp189[167],pp188[169],pp187[171],pp186[173],pp185[175],pp184[177],pp183[179],pp182[181],pp181[183],pp180[185],pp179[187],pp178[189],pp177[191],pp176[193],pp175[195],pp174[197],pp173[199],pp172[201],pp171[203],pp170[205],pp169[207],pp168[209],pp167[211],pp166[213],pp165[215],pp164[217],pp163[219],pp162[221],pp161[223],pp162[223],pp163[223],pp164[223],pp165[223],pp166[223],pp167[223],pp168[223],pp169[223],pp170[223],pp171[223],pp172[223],pp173[223],pp174[223],pp175[223],pp176[223],pp177[223],pp178[223],pp179[223],pp180[223],pp181[223],pp182[223],pp183[223],pp184[223],pp185[223],pp186[223],pp187[223],pp188[223],pp189[223],pp190[223],pp191[223],pp192[223],pp193[223],pp194[223],pp195[223],pp196[223],pp197[223],pp198[223],pp199[223],pp200[223],pp201[223],pp202[223],pp203[223],pp204[223],pp205[223],pp206[223],pp207[223],pp208[223]};
    assign in145_2 = {pp43[37],pp43[38],pp43[39],pp43[40],pp43[41],pp43[42],pp43[43],pp43[44],pp43[45],pp43[46],pp43[47],pp43[48],pp43[49],pp43[50],pp43[51],pp43[52],pp43[53],pp43[54],pp43[55],pp43[56],pp42[58],pp41[60],pp40[62],pp39[64],pp38[66],pp37[68],pp36[70],pp35[72],pp34[74],pp33[76],pp32[78],pp31[80],pp30[82],pp29[84],pp28[86],pp27[88],pp26[90],pp25[92],pp24[94],pp23[96],pp22[98],pp9[112],pp7[115],pp5[118],pp3[121],pp1[124],pp116[10],pp115[12],pp116[12],pp117[12],pp118[12],pp119[12],pp120[12],pp121[12],pp122[12],pp123[12],pp124[12],pp125[12],pp126[12],pp127[12],pp128[12],pp129[12],pp130[12],pp131[12],pp132[12],pp133[12],pp134[12],pp135[12],pp136[12],pp137[12],pp138[12],pp139[12],pp140[12],pp141[12],pp142[12],pp143[12],pp144[12],pp145[12],pp146[12],pp147[12],pp148[12],pp149[12],pp150[12],pp151[12],pp152[12],pp153[12],pp154[12],pp155[12],pp156[12],pp157[12],pp158[12],pp159[12],pp160[12],pp161[12],pp162[12],pp163[12],pp164[12],pp165[12],pp166[12],pp167[12],pp168[12],pp169[12],pp170[12],pp171[12],pp172[12],pp173[12],pp174[12],pp175[12],pp176[12],pp177[12],pp178[12],pp179[12],pp180[12],pp181[12],pp182[12],pp183[12],pp184[12],pp185[12],pp186[12],pp187[12],pp189[11],pp191[10],s129[138],s130[138],s131[138],s132[138],s133[138],s134[138],s135[138],s136[138],s137[138],s138[138],s139[138],s140[138],s141[138],s142[138],s143[138],s144[138],pp0[218],pp1[218],pp2[218],pp3[218],pp4[218],pp5[218],pp6[218],pp7[218],pp8[218],pp9[218],pp219[9],pp221[8],pp223[7],pp225[6],pp227[5],pp229[4],pp231[3],pp233[2],pp235[1],pp237[0],s10[101],s11[101],s12[101],s13[101],s14[101],s15[101],s16[101],s17[101],s18[101],s19[101],s20[101],s21[101],s22[101],s23[101],s24[101],s25[101],s26[101],s27[101],s28[101],s27[103],s26[105],s25[107],s24[109],s23[111],s22[113],s21[115],s20[117],s19[119],s18[121],s17[123],s16[125],s15[127],s14[129],s13[131],s12[133],s11[135],s10[137],s144[196],s143[198],s142[200],s141[202],s140[204],s139[206],s138[208],s137[210],s136[212],s135[214],s134[216],s133[218],s132[220],s131[222],s130[224],s129[226],pp255[36],pp254[38],pp253[40],pp252[42],pp251[44],pp250[46],pp249[48],pp248[50],pp247[52],pp246[54],pp245[56],pp244[58],pp243[60],pp242[62],pp241[64],pp240[66],pp239[68],pp238[70],pp237[72],pp236[74],pp235[76],pp234[78],pp233[80],pp232[82],pp231[84],pp230[86],pp229[88],pp228[90],pp227[92],pp226[94],pp225[96],pp224[98],pp99[224],pp97[227],pp95[230],pp93[233],pp91[236],pp89[239],pp87[242],pp85[245],pp83[248],pp81[251],pp79[254],pp233[101],pp231[104],pp229[107],pp227[110],pp225[113],pp223[116],pp221[119],pp219[122],pp217[125],pp215[128],pp213[131],pp211[134],pp209[137],pp207[140],pp205[143],pp203[146],pp201[149],pp199[152],pp197[155],pp195[158],pp193[161],pp191[164],pp190[166],pp189[168],pp188[170],pp187[172],pp186[174],pp185[176],pp184[178],pp183[180],pp182[182],pp181[184],pp180[186],pp179[188],pp178[190],pp177[192],pp176[194],pp175[196],pp174[198],pp173[200],pp172[202],pp171[204],pp170[206],pp169[208],pp168[210],pp167[212],pp166[214],pp165[216],pp164[218],pp163[220],pp162[222],pp163[222],pp164[222],pp165[222],pp166[222],pp167[222],pp168[222],pp169[222],pp170[222],pp171[222],pp172[222],pp173[222],pp174[222],pp175[222],pp176[222],pp177[222],pp178[222],pp179[222],pp180[222],pp181[222],pp182[222],pp183[222],pp184[222],pp185[222],pp186[222],pp187[222],pp188[222],pp189[222],pp190[222],pp191[222],pp192[222],pp193[222],pp194[222],pp195[222],pp196[222],pp197[222],pp198[222],pp199[222],pp200[222],pp201[222],pp202[222],pp203[222],pp204[222],pp205[222],pp206[222],pp207[222],pp208[222],pp209[222]};
    CLA_352 KS_145(s145, c145, in145_1, in145_2);
    wire[349:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp44[37],pp44[38],pp44[39],pp44[40],pp44[41],pp44[42],pp44[43],pp44[44],pp44[45],pp44[46],pp44[47],pp44[48],pp44[49],pp44[50],pp44[51],pp44[52],pp44[53],pp44[54],pp44[55],pp43[57],pp42[59],pp41[61],pp40[63],pp39[65],pp38[67],pp37[69],pp36[71],pp35[73],pp34[75],pp33[77],pp32[79],pp31[81],pp30[83],pp29[85],pp28[87],pp27[89],pp26[91],pp25[93],pp24[95],pp23[97],pp22[99],pp8[114],pp6[117],pp4[120],pp2[123],pp0[126],pp116[11],pp117[11],pp118[11],pp119[11],pp120[11],pp121[11],pp122[11],pp123[11],pp124[11],pp125[11],pp126[11],pp127[11],pp128[11],pp129[11],pp130[11],pp131[11],pp132[11],pp133[11],pp134[11],pp135[11],pp136[11],pp137[11],pp138[11],pp139[11],pp140[11],pp141[11],pp142[11],pp143[11],pp144[11],pp145[11],pp146[11],pp147[11],pp148[11],pp149[11],pp150[11],pp151[11],pp152[11],pp153[11],pp154[11],pp155[11],pp156[11],pp157[11],pp158[11],pp159[11],pp160[11],pp161[11],pp162[11],pp163[11],pp164[11],pp165[11],pp166[11],pp167[11],pp168[11],pp169[11],pp170[11],pp171[11],pp172[11],pp173[11],pp174[11],pp175[11],pp176[11],pp177[11],pp178[11],pp179[11],pp180[11],pp181[11],pp182[11],pp183[11],pp184[11],pp185[11],pp186[11],pp187[11],pp188[11],pp190[10],s129[137],s130[137],s131[137],s132[137],s133[137],s134[137],s135[137],s136[137],s137[137],s138[137],s139[137],s140[137],s141[137],s142[137],s143[137],s144[137],s145[137],s145[138],s145[139],s145[140],s145[141],s145[142],s145[143],s145[144],s145[145],s145[146],s145[147],s145[148],s145[149],s145[150],s145[151],s145[152],s145[153],s145[154],s145[155],s145[156],s145[157],s145[158],s145[159],s145[160],s145[161],s145[162],s145[163],s145[164],s145[165],s145[166],s145[167],s145[168],s145[169],s145[170],s145[171],s145[172],s145[173],s145[174],s145[175],s145[176],s145[177],s145[178],s145[179],s145[180],s145[181],s145[182],s145[183],s145[184],s145[185],s145[186],s145[187],s145[188],s145[189],s145[190],s145[191],s145[192],s145[193],s145[194],s145[195],s144[197],s143[199],s142[201],s141[203],s140[205],s139[207],s138[209],s137[211],s136[213],s135[215],s134[217],s133[219],s132[221],s131[223],s130[225],s129[227],pp255[37],pp254[39],pp253[41],pp252[43],pp251[45],pp250[47],pp249[49],pp248[51],pp247[53],pp246[55],pp245[57],pp244[59],pp243[61],pp242[63],pp241[65],pp240[67],pp239[69],pp238[71],pp237[73],pp236[75],pp235[77],pp234[79],pp233[81],pp232[83],pp231[85],pp230[87],pp229[89],pp228[91],pp227[93],pp226[95],pp225[97],pp224[99],pp98[226],pp96[229],pp94[232],pp92[235],pp90[238],pp88[241],pp86[244],pp84[247],pp82[250],pp80[253],pp234[100],pp232[103],pp230[106],pp228[109],pp226[112],pp224[115],pp222[118],pp220[121],pp218[124],pp216[127],pp214[130],pp212[133],pp210[136],pp208[139],pp206[142],pp204[145],pp202[148],pp200[151],pp198[154],pp196[157],pp194[160],pp192[163],pp191[165],pp190[167],pp189[169],pp188[171],pp187[173],pp186[175],pp185[177],pp184[179],pp183[181],pp182[183],pp181[185],pp180[187],pp179[189],pp178[191],pp177[193],pp176[195],pp175[197],pp174[199],pp173[201],pp172[203],pp171[205],pp170[207],pp169[209],pp168[211],pp167[213],pp166[215],pp165[217],pp164[219],pp163[221],pp164[221],pp165[221],pp166[221],pp167[221],pp168[221],pp169[221],pp170[221],pp171[221],pp172[221],pp173[221],pp174[221],pp175[221],pp176[221],pp177[221],pp178[221],pp179[221],pp180[221],pp181[221],pp182[221],pp183[221],pp184[221],pp185[221],pp186[221],pp187[221],pp188[221],pp189[221],pp190[221],pp191[221],pp192[221],pp193[221],pp194[221],pp195[221],pp196[221],pp197[221],pp198[221],pp199[221],pp200[221],pp201[221],pp202[221],pp203[221],pp204[221],pp205[221],pp206[221],pp207[221],pp208[221],pp209[221]};
    assign in146_2 = {pp45[36],pp45[37],pp45[38],pp45[39],pp45[40],pp45[41],pp45[42],pp45[43],pp45[44],pp45[45],pp45[46],pp45[47],pp45[48],pp45[49],pp45[50],pp45[51],pp45[52],pp45[53],pp45[54],pp44[56],pp43[58],pp42[60],pp41[62],pp40[64],pp39[66],pp38[68],pp37[70],pp36[72],pp35[74],pp34[76],pp33[78],pp32[80],pp31[82],pp30[84],pp29[86],pp28[88],pp27[90],pp26[92],pp25[94],pp24[96],pp23[98],pp9[113],pp7[116],pp5[119],pp3[122],pp1[125],pp117[10],pp118[10],pp119[10],pp120[10],pp121[10],pp122[10],pp123[10],pp124[10],pp125[10],pp126[10],pp127[10],pp128[10],pp129[10],pp130[10],pp131[10],pp132[10],pp133[10],pp134[10],pp135[10],pp136[10],pp137[10],pp138[10],pp139[10],pp140[10],pp141[10],pp142[10],pp143[10],pp144[10],pp145[10],pp146[10],pp147[10],pp148[10],pp149[10],pp150[10],pp151[10],pp152[10],pp153[10],pp154[10],pp155[10],pp156[10],pp157[10],pp158[10],pp159[10],pp160[10],pp161[10],pp162[10],pp163[10],pp164[10],pp165[10],pp166[10],pp167[10],pp168[10],pp169[10],pp170[10],pp171[10],pp172[10],pp173[10],pp174[10],pp175[10],pp176[10],pp177[10],pp178[10],pp179[10],pp180[10],pp181[10],pp182[10],pp183[10],pp184[10],pp185[10],pp186[10],pp187[10],pp188[10],pp189[10],s129[136],s130[136],s131[136],s132[136],s133[136],s134[136],s135[136],s136[136],s137[136],s138[136],s139[136],s140[136],s141[136],s142[136],s143[136],s144[136],s145[136],pp0[217],pp1[217],pp2[217],pp3[217],pp4[217],pp5[217],pp6[217],pp7[217],pp8[217],pp9[217],pp218[9],pp220[8],pp222[7],pp224[6],pp226[5],pp228[4],pp230[3],pp232[2],pp234[1],pp236[0],s10[100],s11[100],s12[100],s13[100],s14[100],s15[100],s16[100],s17[100],s18[100],s19[100],s20[100],s21[100],s22[100],s23[100],s24[100],s25[100],s26[100],s27[100],s28[100],s29[100],s28[102],s27[104],s26[106],s25[108],s24[110],s23[112],s22[114],s21[116],s20[118],s19[120],s18[122],s17[124],s16[126],s15[128],s14[130],s13[132],s12[134],s11[136],s10[138],s145[196],s144[198],s143[200],s142[202],s141[204],s140[206],s139[208],s138[210],s137[212],s136[214],s135[216],s134[218],s133[220],s132[222],s131[224],s130[226],s129[228],pp255[38],pp254[40],pp253[42],pp252[44],pp251[46],pp250[48],pp249[50],pp248[52],pp247[54],pp246[56],pp245[58],pp244[60],pp243[62],pp242[64],pp241[66],pp240[68],pp239[70],pp238[72],pp237[74],pp236[76],pp235[78],pp234[80],pp233[82],pp232[84],pp231[86],pp230[88],pp229[90],pp228[92],pp227[94],pp226[96],pp225[98],pp99[225],pp97[228],pp95[231],pp93[234],pp91[237],pp89[240],pp87[243],pp85[246],pp83[249],pp81[252],pp79[255],pp233[102],pp231[105],pp229[108],pp227[111],pp225[114],pp223[117],pp221[120],pp219[123],pp217[126],pp215[129],pp213[132],pp211[135],pp209[138],pp207[141],pp205[144],pp203[147],pp201[150],pp199[153],pp197[156],pp195[159],pp193[162],pp192[164],pp191[166],pp190[168],pp189[170],pp188[172],pp187[174],pp186[176],pp185[178],pp184[180],pp183[182],pp182[184],pp181[186],pp180[188],pp179[190],pp178[192],pp177[194],pp176[196],pp175[198],pp174[200],pp173[202],pp172[204],pp171[206],pp170[208],pp169[210],pp168[212],pp167[214],pp166[216],pp165[218],pp164[220],pp165[220],pp166[220],pp167[220],pp168[220],pp169[220],pp170[220],pp171[220],pp172[220],pp173[220],pp174[220],pp175[220],pp176[220],pp177[220],pp178[220],pp179[220],pp180[220],pp181[220],pp182[220],pp183[220],pp184[220],pp185[220],pp186[220],pp187[220],pp188[220],pp189[220],pp190[220],pp191[220],pp192[220],pp193[220],pp194[220],pp195[220],pp196[220],pp197[220],pp198[220],pp199[220],pp200[220],pp201[220],pp202[220],pp203[220],pp204[220],pp205[220],pp206[220],pp207[220],pp208[220],pp209[220],pp210[220]};
    CLA_350 KS_146(s146, c146, in146_1, in146_2);
    wire[347:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp46[36],pp46[37],pp46[38],pp46[39],pp46[40],pp46[41],pp46[42],pp46[43],pp46[44],pp46[45],pp46[46],pp46[47],pp46[48],pp46[49],pp46[50],pp46[51],pp46[52],pp46[53],pp45[55],pp44[57],pp43[59],pp42[61],pp41[63],pp40[65],pp39[67],pp38[69],pp37[71],pp36[73],pp35[75],pp34[77],pp33[79],pp32[81],pp31[83],pp30[85],pp29[87],pp28[89],pp27[91],pp26[93],pp25[95],pp24[97],pp23[99],pp8[115],pp6[118],pp4[121],pp2[124],pp0[127],pp0[128],pp0[129],pp0[130],pp0[131],pp0[132],pp0[133],pp0[134],pp0[135],pp0[136],pp0[137],pp0[138],pp0[139],pp0[140],pp0[141],pp0[142],pp0[143],pp0[144],pp0[145],pp0[146],pp0[147],pp0[148],pp0[149],pp0[150],pp0[151],pp0[152],pp0[153],pp0[154],pp0[155],pp0[156],pp0[157],pp0[158],pp0[159],pp0[160],pp0[161],pp0[162],pp0[163],s129[100],s129[101],s129[102],s129[103],s129[104],s129[105],s129[106],s129[107],s129[108],s129[109],s129[110],s129[111],s129[112],s129[113],s129[114],s129[115],s129[116],s129[117],s129[118],s129[119],s129[120],s129[121],s129[122],s129[123],s129[124],s129[125],s129[126],s129[127],s129[128],s129[129],s129[130],s129[131],s129[132],s129[133],s129[134],s129[135],s130[135],s131[135],s132[135],s133[135],s134[135],s135[135],s136[135],s137[135],s138[135],s139[135],s140[135],s141[135],s142[135],s143[135],s144[135],s145[135],s146[135],s146[136],s146[137],s146[138],s146[139],s146[140],s146[141],s146[142],s146[143],s146[144],s146[145],s146[146],s146[147],s146[148],s146[149],s146[150],s146[151],s146[152],s146[153],s146[154],s146[155],s146[156],s146[157],s146[158],s146[159],s146[160],s146[161],s146[162],s146[163],s146[164],s146[165],s146[166],s146[167],s146[168],s146[169],s146[170],s146[171],s146[172],s146[173],s146[174],s146[175],s146[176],s146[177],s146[178],s146[179],s146[180],s146[181],s146[182],s146[183],s146[184],s146[185],s146[186],s146[187],s146[188],s146[189],s146[190],s146[191],s146[192],s146[193],s146[194],s146[195],s145[197],s144[199],s143[201],s142[203],s141[205],s140[207],s139[209],s138[211],s137[213],s136[215],s135[217],s134[219],s133[221],s132[223],s131[225],s130[227],s129[229],pp255[39],pp254[41],pp253[43],pp252[45],pp251[47],pp250[49],pp249[51],pp248[53],pp247[55],pp246[57],pp245[59],pp244[61],pp243[63],pp242[65],pp241[67],pp240[69],pp239[71],pp238[73],pp237[75],pp236[77],pp235[79],pp234[81],pp233[83],pp232[85],pp231[87],pp230[89],pp229[91],pp228[93],pp227[95],pp226[97],pp225[99],pp98[227],pp96[230],pp94[233],pp92[236],pp90[239],pp88[242],pp86[245],pp84[248],pp82[251],pp80[254],pp234[101],pp232[104],pp230[107],pp228[110],pp226[113],pp224[116],pp222[119],pp220[122],pp218[125],pp216[128],pp214[131],pp212[134],pp210[137],pp208[140],pp206[143],pp204[146],pp202[149],pp200[152],pp198[155],pp196[158],pp194[161],pp193[163],pp192[165],pp191[167],pp190[169],pp189[171],pp188[173],pp187[175],pp186[177],pp185[179],pp184[181],pp183[183],pp182[185],pp181[187],pp180[189],pp179[191],pp178[193],pp177[195],pp176[197],pp175[199],pp174[201],pp173[203],pp172[205],pp171[207],pp170[209],pp169[211],pp168[213],pp167[215],pp166[217],pp165[219],pp166[219],pp167[219],pp168[219],pp169[219],pp170[219],pp171[219],pp172[219],pp173[219],pp174[219],pp175[219],pp176[219],pp177[219],pp178[219],pp179[219],pp180[219],pp181[219],pp182[219],pp183[219],pp184[219],pp185[219],pp186[219],pp187[219],pp188[219],pp189[219],pp190[219],pp191[219],pp192[219],pp193[219],pp194[219],pp195[219],pp196[219],pp197[219],pp198[219],pp199[219],pp200[219],pp201[219],pp202[219],pp203[219],pp204[219],pp205[219],pp206[219],pp207[219],pp208[219],pp209[219],pp210[219]};
    assign in147_2 = {pp47[35],pp47[36],pp47[37],pp47[38],pp47[39],pp47[40],pp47[41],pp47[42],pp47[43],pp47[44],pp47[45],pp47[46],pp47[47],pp47[48],pp47[49],pp47[50],pp47[51],pp47[52],pp46[54],pp45[56],pp44[58],pp43[60],pp42[62],pp41[64],pp40[66],pp39[68],pp38[70],pp37[72],pp36[74],pp35[76],pp34[78],pp33[80],pp32[82],pp31[84],pp30[86],pp29[88],pp28[90],pp27[92],pp26[94],pp25[96],pp24[98],pp9[114],pp7[117],pp5[120],pp3[123],pp1[126],pp1[127],pp1[128],pp1[129],pp1[130],pp1[131],pp1[132],pp1[133],pp1[134],pp1[135],pp1[136],pp1[137],pp1[138],pp1[139],pp1[140],pp1[141],pp1[142],pp1[143],pp1[144],pp1[145],pp1[146],pp1[147],pp1[148],pp1[149],pp1[150],pp1[151],pp1[152],pp1[153],pp1[154],pp1[155],pp1[156],pp1[157],pp1[158],pp1[159],pp1[160],pp1[161],pp1[162],pp0[164],s130[100],s130[101],s130[102],s130[103],s130[104],s130[105],s130[106],s130[107],s130[108],s130[109],s130[110],s130[111],s130[112],s130[113],s130[114],s130[115],s130[116],s130[117],s130[118],s130[119],s130[120],s130[121],s130[122],s130[123],s130[124],s130[125],s130[126],s130[127],s130[128],s130[129],s130[130],s130[131],s130[132],s130[133],s130[134],s131[134],s132[134],s133[134],s134[134],s135[134],s136[134],s137[134],s138[134],s139[134],s140[134],s141[134],s142[134],s143[134],s144[134],s145[134],s146[134],pp0[216],pp1[216],pp2[216],pp3[216],pp4[216],pp5[216],pp6[216],pp7[216],pp8[216],pp9[216],pp217[9],pp219[8],pp221[7],pp223[6],pp225[5],pp227[4],pp229[3],pp231[2],pp233[1],pp235[0],s1[108],s100[10],s100[11],s100[12],s100[13],s100[14],s100[15],s100[16],s100[17],s100[18],s100[19],s100[20],s100[21],s100[22],s100[23],s100[24],s100[25],s100[26],s100[27],s100[28],s100[29],s29[101],s28[103],s27[105],s26[107],s25[109],s24[111],s23[113],s22[115],s21[117],s20[119],s19[121],s18[123],s17[125],s16[127],s15[129],s14[131],s13[133],s12[135],s11[137],s10[139],s146[196],s145[198],s144[200],s143[202],s142[204],s141[206],s140[208],s139[210],s138[212],s137[214],s136[216],s135[218],s134[220],s133[222],s132[224],s131[226],s130[228],s129[230],pp255[40],pp254[42],pp253[44],pp252[46],pp251[48],pp250[50],pp249[52],pp248[54],pp247[56],pp246[58],pp245[60],pp244[62],pp243[64],pp242[66],pp241[68],pp240[70],pp239[72],pp238[74],pp237[76],pp236[78],pp235[80],pp234[82],pp233[84],pp232[86],pp231[88],pp230[90],pp229[92],pp228[94],pp227[96],pp226[98],pp99[226],pp97[229],pp95[232],pp93[235],pp91[238],pp89[241],pp87[244],pp85[247],pp83[250],pp81[253],pp235[100],pp233[103],pp231[106],pp229[109],pp227[112],pp225[115],pp223[118],pp221[121],pp219[124],pp217[127],pp215[130],pp213[133],pp211[136],pp209[139],pp207[142],pp205[145],pp203[148],pp201[151],pp199[154],pp197[157],pp195[160],pp194[162],pp193[164],pp192[166],pp191[168],pp190[170],pp189[172],pp188[174],pp187[176],pp186[178],pp185[180],pp184[182],pp183[184],pp182[186],pp181[188],pp180[190],pp179[192],pp178[194],pp177[196],pp176[198],pp175[200],pp174[202],pp173[204],pp172[206],pp171[208],pp170[210],pp169[212],pp168[214],pp167[216],pp166[218],pp167[218],pp168[218],pp169[218],pp170[218],pp171[218],pp172[218],pp173[218],pp174[218],pp175[218],pp176[218],pp177[218],pp178[218],pp179[218],pp180[218],pp181[218],pp182[218],pp183[218],pp184[218],pp185[218],pp186[218],pp187[218],pp188[218],pp189[218],pp190[218],pp191[218],pp192[218],pp193[218],pp194[218],pp195[218],pp196[218],pp197[218],pp198[218],pp199[218],pp200[218],pp201[218],pp202[218],pp203[218],pp204[218],pp205[218],pp206[218],pp207[218],pp208[218],pp209[218],pp210[218],pp211[218]};
    CLA_348 KS_147(s147, c147, in147_1, in147_2);
    wire[345:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp48[35],pp48[36],pp48[37],pp48[38],pp48[39],pp48[40],pp48[41],pp48[42],pp48[43],pp48[44],pp48[45],pp48[46],pp48[47],pp48[48],pp48[49],pp48[50],pp48[51],pp47[53],pp46[55],pp45[57],pp44[59],pp43[61],pp42[63],pp41[65],pp40[67],pp39[69],pp38[71],pp37[73],pp36[75],pp35[77],pp34[79],pp33[81],pp32[83],pp31[85],pp30[87],pp29[89],pp28[91],pp27[93],pp26[95],pp25[97],pp24[99],pp8[116],pp6[119],pp4[122],pp2[125],pp2[126],pp2[127],pp2[128],pp2[129],pp2[130],pp2[131],pp2[132],pp2[133],pp2[134],pp2[135],pp2[136],pp2[137],pp2[138],pp2[139],pp2[140],pp2[141],pp2[142],pp2[143],pp2[144],pp2[145],pp2[146],pp2[147],pp2[148],pp2[149],pp2[150],pp2[151],pp2[152],pp2[153],pp2[154],pp2[155],pp2[156],pp2[157],pp2[158],pp2[159],pp2[160],pp2[161],pp1[163],pp0[165],s131[100],s131[101],s131[102],s131[103],s131[104],s131[105],s131[106],s131[107],s131[108],s131[109],s131[110],s131[111],s131[112],s131[113],s131[114],s131[115],s131[116],s131[117],s131[118],s131[119],s131[120],s131[121],s131[122],s131[123],s131[124],s131[125],s131[126],s131[127],s131[128],s131[129],s131[130],s131[131],s131[132],s131[133],s132[133],s133[133],s134[133],s135[133],s136[133],s137[133],s138[133],s139[133],s140[133],s141[133],s142[133],s143[133],s144[133],s145[133],s146[133],s147[133],s147[134],s147[135],s147[136],s147[137],s147[138],s147[139],s147[140],s147[141],s147[142],s147[143],s147[144],s147[145],s147[146],s147[147],s147[148],s147[149],s147[150],s147[151],s147[152],s147[153],s147[154],s147[155],s147[156],s147[157],s147[158],s147[159],s147[160],s147[161],s147[162],s147[163],s147[164],s147[165],s147[166],s147[167],s147[168],s147[169],s147[170],s147[171],s147[172],s147[173],s147[174],s147[175],s147[176],s147[177],s147[178],s147[179],s147[180],s147[181],s147[182],s147[183],s147[184],s147[185],s147[186],s147[187],s147[188],s147[189],s147[190],s147[191],s147[192],s147[193],s147[194],s147[195],s146[197],s145[199],s144[201],s143[203],s142[205],s141[207],s140[209],s139[211],s138[213],s137[215],s136[217],s135[219],s134[221],s133[223],s132[225],s131[227],s130[229],s129[231],pp255[41],pp254[43],pp253[45],pp252[47],pp251[49],pp250[51],pp249[53],pp248[55],pp247[57],pp246[59],pp245[61],pp244[63],pp243[65],pp242[67],pp241[69],pp240[71],pp239[73],pp238[75],pp237[77],pp236[79],pp235[81],pp234[83],pp233[85],pp232[87],pp231[89],pp230[91],pp229[93],pp228[95],pp227[97],pp226[99],pp98[228],pp96[231],pp94[234],pp92[237],pp90[240],pp88[243],pp86[246],pp84[249],pp82[252],pp80[255],pp234[102],pp232[105],pp230[108],pp228[111],pp226[114],pp224[117],pp222[120],pp220[123],pp218[126],pp216[129],pp214[132],pp212[135],pp210[138],pp208[141],pp206[144],pp204[147],pp202[150],pp200[153],pp198[156],pp196[159],pp195[161],pp194[163],pp193[165],pp192[167],pp191[169],pp190[171],pp189[173],pp188[175],pp187[177],pp186[179],pp185[181],pp184[183],pp183[185],pp182[187],pp181[189],pp180[191],pp179[193],pp178[195],pp177[197],pp176[199],pp175[201],pp174[203],pp173[205],pp172[207],pp171[209],pp170[211],pp169[213],pp168[215],pp167[217],pp168[217],pp169[217],pp170[217],pp171[217],pp172[217],pp173[217],pp174[217],pp175[217],pp176[217],pp177[217],pp178[217],pp179[217],pp180[217],pp181[217],pp182[217],pp183[217],pp184[217],pp185[217],pp186[217],pp187[217],pp188[217],pp189[217],pp190[217],pp191[217],pp192[217],pp193[217],pp194[217],pp195[217],pp196[217],pp197[217],pp198[217],pp199[217],pp200[217],pp201[217],pp202[217],pp203[217],pp204[217],pp205[217],pp206[217],pp207[217],pp208[217],pp209[217],pp210[217],pp211[217]};
    assign in148_2 = {pp49[34],pp49[35],pp49[36],pp49[37],pp49[38],pp49[39],pp49[40],pp49[41],pp49[42],pp49[43],pp49[44],pp49[45],pp49[46],pp49[47],pp49[48],pp49[49],pp49[50],pp48[52],pp47[54],pp46[56],pp45[58],pp44[60],pp43[62],pp42[64],pp41[66],pp40[68],pp39[70],pp38[72],pp37[74],pp36[76],pp35[78],pp34[80],pp33[82],pp32[84],pp31[86],pp30[88],pp29[90],pp28[92],pp27[94],pp26[96],pp25[98],pp9[115],pp7[118],pp5[121],pp3[124],pp3[125],pp3[126],pp3[127],pp3[128],pp3[129],pp3[130],pp3[131],pp3[132],pp3[133],pp3[134],pp3[135],pp3[136],pp3[137],pp3[138],pp3[139],pp3[140],pp3[141],pp3[142],pp3[143],pp3[144],pp3[145],pp3[146],pp3[147],pp3[148],pp3[149],pp3[150],pp3[151],pp3[152],pp3[153],pp3[154],pp3[155],pp3[156],pp3[157],pp3[158],pp3[159],pp3[160],pp2[162],pp1[164],pp0[166],s132[100],s132[101],s132[102],s132[103],s132[104],s132[105],s132[106],s132[107],s132[108],s132[109],s132[110],s132[111],s132[112],s132[113],s132[114],s132[115],s132[116],s132[117],s132[118],s132[119],s132[120],s132[121],s132[122],s132[123],s132[124],s132[125],s132[126],s132[127],s132[128],s132[129],s132[130],s132[131],s132[132],s133[132],s134[132],s135[132],s136[132],s137[132],s138[132],s139[132],s140[132],s141[132],s142[132],s143[132],s144[132],s145[132],s146[132],s147[132],pp0[215],pp1[215],pp2[215],pp3[215],pp4[215],pp5[215],pp6[215],pp7[215],pp8[215],pp9[215],pp216[9],pp218[8],pp220[7],pp222[6],pp224[5],pp226[4],pp228[3],pp230[2],pp232[1],pp234[0],s1[107],s2[107],s1[109],s101[10],s101[11],s101[12],s101[13],s101[14],s101[15],s101[16],s101[17],s101[18],s101[19],s101[20],s101[21],s101[22],s101[23],s101[24],s101[25],s101[26],s101[27],s101[28],s30[100],s29[102],s28[104],s27[106],s26[108],s25[110],s24[112],s23[114],s22[116],s21[118],s20[120],s19[122],s18[124],s17[126],s16[128],s15[130],s14[132],s13[134],s12[136],s11[138],s10[140],s147[196],s146[198],s145[200],s144[202],s143[204],s142[206],s141[208],s140[210],s139[212],s138[214],s137[216],s136[218],s135[220],s134[222],s133[224],s132[226],s131[228],s130[230],s129[232],pp255[42],pp254[44],pp253[46],pp252[48],pp251[50],pp250[52],pp249[54],pp248[56],pp247[58],pp246[60],pp245[62],pp244[64],pp243[66],pp242[68],pp241[70],pp240[72],pp239[74],pp238[76],pp237[78],pp236[80],pp235[82],pp234[84],pp233[86],pp232[88],pp231[90],pp230[92],pp229[94],pp228[96],pp227[98],pp99[227],pp97[230],pp95[233],pp93[236],pp91[239],pp89[242],pp87[245],pp85[248],pp83[251],pp81[254],pp235[101],pp233[104],pp231[107],pp229[110],pp227[113],pp225[116],pp223[119],pp221[122],pp219[125],pp217[128],pp215[131],pp213[134],pp211[137],pp209[140],pp207[143],pp205[146],pp203[149],pp201[152],pp199[155],pp197[158],pp196[160],pp195[162],pp194[164],pp193[166],pp192[168],pp191[170],pp190[172],pp189[174],pp188[176],pp187[178],pp186[180],pp185[182],pp184[184],pp183[186],pp182[188],pp181[190],pp180[192],pp179[194],pp178[196],pp177[198],pp176[200],pp175[202],pp174[204],pp173[206],pp172[208],pp171[210],pp170[212],pp169[214],pp168[216],pp169[216],pp170[216],pp171[216],pp172[216],pp173[216],pp174[216],pp175[216],pp176[216],pp177[216],pp178[216],pp179[216],pp180[216],pp181[216],pp182[216],pp183[216],pp184[216],pp185[216],pp186[216],pp187[216],pp188[216],pp189[216],pp190[216],pp191[216],pp192[216],pp193[216],pp194[216],pp195[216],pp196[216],pp197[216],pp198[216],pp199[216],pp200[216],pp201[216],pp202[216],pp203[216],pp204[216],pp205[216],pp206[216],pp207[216],pp208[216],pp209[216],pp210[216],pp211[216],pp212[216]};
    CLA_346 KS_148(s148, c148, in148_1, in148_2);
    wire[343:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp50[34],pp50[35],pp50[36],pp50[37],pp50[38],pp50[39],pp50[40],pp50[41],pp50[42],pp50[43],pp50[44],pp50[45],pp50[46],pp50[47],pp50[48],pp50[49],pp49[51],pp48[53],pp47[55],pp46[57],pp45[59],pp44[61],pp43[63],pp42[65],pp41[67],pp40[69],pp39[71],pp38[73],pp37[75],pp36[77],pp35[79],pp34[81],pp33[83],pp32[85],pp31[87],pp30[89],pp29[91],pp28[93],pp27[95],pp26[97],pp25[99],pp8[117],pp6[120],pp4[123],pp4[124],pp4[125],pp4[126],pp4[127],pp4[128],pp4[129],pp4[130],pp4[131],pp4[132],pp4[133],pp4[134],pp4[135],pp4[136],pp4[137],pp4[138],pp4[139],pp4[140],pp4[141],pp4[142],pp4[143],pp4[144],pp4[145],pp4[146],pp4[147],pp4[148],pp4[149],pp4[150],pp4[151],pp4[152],pp4[153],pp4[154],pp4[155],pp4[156],pp4[157],pp4[158],pp4[159],pp3[161],pp2[163],pp1[165],pp0[167],s133[100],s133[101],s133[102],s133[103],s133[104],s133[105],s133[106],s133[107],s133[108],s133[109],s133[110],s133[111],s133[112],s133[113],s133[114],s133[115],s133[116],s133[117],s133[118],s133[119],s133[120],s133[121],s133[122],s133[123],s133[124],s133[125],s133[126],s133[127],s133[128],s133[129],s133[130],s133[131],s134[131],s135[131],s136[131],s137[131],s138[131],s139[131],s140[131],s141[131],s142[131],s143[131],s144[131],s145[131],s146[131],s147[131],s148[131],s148[132],s148[133],s148[134],s148[135],s148[136],s148[137],s148[138],s148[139],s148[140],s148[141],s148[142],s148[143],s148[144],s148[145],s148[146],s148[147],s148[148],s148[149],s148[150],s148[151],s148[152],s148[153],s148[154],s148[155],s148[156],s148[157],s148[158],s148[159],s148[160],s148[161],s148[162],s148[163],s148[164],s148[165],s148[166],s148[167],s148[168],s148[169],s148[170],s148[171],s148[172],s148[173],s148[174],s148[175],s148[176],s148[177],s148[178],s148[179],s148[180],s148[181],s148[182],s148[183],s148[184],s148[185],s148[186],s148[187],s148[188],s148[189],s148[190],s148[191],s148[192],s148[193],s148[194],s148[195],s147[197],s146[199],s145[201],s144[203],s143[205],s142[207],s141[209],s140[211],s139[213],s138[215],s137[217],s136[219],s135[221],s134[223],s133[225],s132[227],s131[229],s130[231],s129[233],pp255[43],pp254[45],pp253[47],pp252[49],pp251[51],pp250[53],pp249[55],pp248[57],pp247[59],pp246[61],pp245[63],pp244[65],pp243[67],pp242[69],pp241[71],pp240[73],pp239[75],pp238[77],pp237[79],pp236[81],pp235[83],pp234[85],pp233[87],pp232[89],pp231[91],pp230[93],pp229[95],pp228[97],pp227[99],pp98[229],pp96[232],pp94[235],pp92[238],pp90[241],pp88[244],pp86[247],pp84[250],pp82[253],pp236[100],pp234[103],pp232[106],pp230[109],pp228[112],pp226[115],pp224[118],pp222[121],pp220[124],pp218[127],pp216[130],pp214[133],pp212[136],pp210[139],pp208[142],pp206[145],pp204[148],pp202[151],pp200[154],pp198[157],pp197[159],pp196[161],pp195[163],pp194[165],pp193[167],pp192[169],pp191[171],pp190[173],pp189[175],pp188[177],pp187[179],pp186[181],pp185[183],pp184[185],pp183[187],pp182[189],pp181[191],pp180[193],pp179[195],pp178[197],pp177[199],pp176[201],pp175[203],pp174[205],pp173[207],pp172[209],pp171[211],pp170[213],pp169[215],pp170[215],pp171[215],pp172[215],pp173[215],pp174[215],pp175[215],pp176[215],pp177[215],pp178[215],pp179[215],pp180[215],pp181[215],pp182[215],pp183[215],pp184[215],pp185[215],pp186[215],pp187[215],pp188[215],pp189[215],pp190[215],pp191[215],pp192[215],pp193[215],pp194[215],pp195[215],pp196[215],pp197[215],pp198[215],pp199[215],pp200[215],pp201[215],pp202[215],pp203[215],pp204[215],pp205[215],pp206[215],pp207[215],pp208[215],pp209[215],pp210[215],pp211[215],pp212[215]};
    assign in149_2 = {pp51[33],pp51[34],pp51[35],pp51[36],pp51[37],pp51[38],pp51[39],pp51[40],pp51[41],pp51[42],pp51[43],pp51[44],pp51[45],pp51[46],pp51[47],pp51[48],pp50[50],pp49[52],pp48[54],pp47[56],pp46[58],pp45[60],pp44[62],pp43[64],pp42[66],pp41[68],pp40[70],pp39[72],pp38[74],pp37[76],pp36[78],pp35[80],pp34[82],pp33[84],pp32[86],pp31[88],pp30[90],pp29[92],pp28[94],pp27[96],pp26[98],pp9[116],pp7[119],pp5[122],pp5[123],pp5[124],pp5[125],pp5[126],pp5[127],pp5[128],pp5[129],pp5[130],pp5[131],pp5[132],pp5[133],pp5[134],pp5[135],pp5[136],pp5[137],pp5[138],pp5[139],pp5[140],pp5[141],pp5[142],pp5[143],pp5[144],pp5[145],pp5[146],pp5[147],pp5[148],pp5[149],pp5[150],pp5[151],pp5[152],pp5[153],pp5[154],pp5[155],pp5[156],pp5[157],pp5[158],pp4[160],pp3[162],pp2[164],pp1[166],pp0[168],s134[100],s134[101],s134[102],s134[103],s134[104],s134[105],s134[106],s134[107],s134[108],s134[109],s134[110],s134[111],s134[112],s134[113],s134[114],s134[115],s134[116],s134[117],s134[118],s134[119],s134[120],s134[121],s134[122],s134[123],s134[124],s134[125],s134[126],s134[127],s134[128],s134[129],s134[130],s135[130],s136[130],s137[130],s138[130],s139[130],s140[130],s141[130],s142[130],s143[130],s144[130],s145[130],s146[130],s147[130],s148[130],pp0[214],pp1[214],pp2[214],pp3[214],pp4[214],pp5[214],pp6[214],pp7[214],pp8[214],pp9[214],pp215[9],pp217[8],pp219[7],pp221[6],pp223[5],pp225[4],pp227[3],pp229[2],pp231[1],pp233[0],s1[106],s2[106],s3[106],s2[108],s1[110],s102[10],s102[11],s102[12],s102[13],s102[14],s102[15],s102[16],s102[17],s102[18],s102[19],s102[20],s102[21],s102[22],s102[23],s102[24],s102[25],s102[26],s102[27],s100[30],s30[101],s29[103],s28[105],s27[107],s26[109],s25[111],s24[113],s23[115],s22[117],s21[119],s20[121],s19[123],s18[125],s17[127],s16[129],s15[131],s14[133],s13[135],s12[137],s11[139],s10[141],s148[196],s147[198],s146[200],s145[202],s144[204],s143[206],s142[208],s141[210],s140[212],s139[214],s138[216],s137[218],s136[220],s135[222],s134[224],s133[226],s132[228],s131[230],s130[232],s129[234],pp255[44],pp254[46],pp253[48],pp252[50],pp251[52],pp250[54],pp249[56],pp248[58],pp247[60],pp246[62],pp245[64],pp244[66],pp243[68],pp242[70],pp241[72],pp240[74],pp239[76],pp238[78],pp237[80],pp236[82],pp235[84],pp234[86],pp233[88],pp232[90],pp231[92],pp230[94],pp229[96],pp228[98],pp99[228],pp97[231],pp95[234],pp93[237],pp91[240],pp89[243],pp87[246],pp85[249],pp83[252],pp81[255],pp235[102],pp233[105],pp231[108],pp229[111],pp227[114],pp225[117],pp223[120],pp221[123],pp219[126],pp217[129],pp215[132],pp213[135],pp211[138],pp209[141],pp207[144],pp205[147],pp203[150],pp201[153],pp199[156],pp198[158],pp197[160],pp196[162],pp195[164],pp194[166],pp193[168],pp192[170],pp191[172],pp190[174],pp189[176],pp188[178],pp187[180],pp186[182],pp185[184],pp184[186],pp183[188],pp182[190],pp181[192],pp180[194],pp179[196],pp178[198],pp177[200],pp176[202],pp175[204],pp174[206],pp173[208],pp172[210],pp171[212],pp170[214],pp171[214],pp172[214],pp173[214],pp174[214],pp175[214],pp176[214],pp177[214],pp178[214],pp179[214],pp180[214],pp181[214],pp182[214],pp183[214],pp184[214],pp185[214],pp186[214],pp187[214],pp188[214],pp189[214],pp190[214],pp191[214],pp192[214],pp193[214],pp194[214],pp195[214],pp196[214],pp197[214],pp198[214],pp199[214],pp200[214],pp201[214],pp202[214],pp203[214],pp204[214],pp205[214],pp206[214],pp207[214],pp208[214],pp209[214],pp210[214],pp211[214],pp212[214],pp213[214]};
    CLA_344 KS_149(s149, c149, in149_1, in149_2);
    wire[341:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp52[33],pp52[34],pp52[35],pp52[36],pp52[37],pp52[38],pp52[39],pp52[40],pp52[41],pp52[42],pp52[43],pp52[44],pp52[45],pp52[46],pp52[47],pp51[49],pp50[51],pp49[53],pp48[55],pp47[57],pp46[59],pp45[61],pp44[63],pp43[65],pp42[67],pp41[69],pp40[71],pp39[73],pp38[75],pp37[77],pp36[79],pp35[81],pp34[83],pp33[85],pp32[87],pp31[89],pp30[91],pp29[93],pp28[95],pp27[97],pp26[99],pp8[118],pp6[121],pp6[122],pp6[123],pp6[124],pp6[125],pp6[126],pp6[127],pp6[128],pp6[129],pp6[130],pp6[131],pp6[132],pp6[133],pp6[134],pp6[135],pp6[136],pp6[137],pp6[138],pp6[139],pp6[140],pp6[141],pp6[142],pp6[143],pp6[144],pp6[145],pp6[146],pp6[147],pp6[148],pp6[149],pp6[150],pp6[151],pp6[152],pp6[153],pp6[154],pp6[155],pp6[156],pp6[157],pp5[159],pp4[161],pp3[163],pp2[165],pp1[167],pp0[169],s135[100],s135[101],s135[102],s135[103],s135[104],s135[105],s135[106],s135[107],s135[108],s135[109],s135[110],s135[111],s135[112],s135[113],s135[114],s135[115],s135[116],s135[117],s135[118],s135[119],s135[120],s135[121],s135[122],s135[123],s135[124],s135[125],s135[126],s135[127],s135[128],s135[129],s136[129],s137[129],s138[129],s139[129],s140[129],s141[129],s142[129],s143[129],s144[129],s145[129],s146[129],s147[129],s148[129],s149[129],s149[130],s149[131],s149[132],s149[133],s149[134],s149[135],s149[136],s149[137],s149[138],s149[139],s149[140],s149[141],s149[142],s149[143],s149[144],s149[145],s149[146],s149[147],s149[148],s149[149],s149[150],s149[151],s149[152],s149[153],s149[154],s149[155],s149[156],s149[157],s149[158],s149[159],s149[160],s149[161],s149[162],s149[163],s149[164],s149[165],s149[166],s149[167],s149[168],s149[169],s149[170],s149[171],s149[172],s149[173],s149[174],s149[175],s149[176],s149[177],s149[178],s149[179],s149[180],s149[181],s149[182],s149[183],s149[184],s149[185],s149[186],s149[187],s149[188],s149[189],s149[190],s149[191],s149[192],s149[193],s149[194],s149[195],s148[197],s147[199],s146[201],s145[203],s144[205],s143[207],s142[209],s141[211],s140[213],s139[215],s138[217],s137[219],s136[221],s135[223],s134[225],s133[227],s132[229],s131[231],s130[233],s129[235],pp255[45],pp254[47],pp253[49],pp252[51],pp251[53],pp250[55],pp249[57],pp248[59],pp247[61],pp246[63],pp245[65],pp244[67],pp243[69],pp242[71],pp241[73],pp240[75],pp239[77],pp238[79],pp237[81],pp236[83],pp235[85],pp234[87],pp233[89],pp232[91],pp231[93],pp230[95],pp229[97],pp228[99],pp98[230],pp96[233],pp94[236],pp92[239],pp90[242],pp88[245],pp86[248],pp84[251],pp82[254],pp236[101],pp234[104],pp232[107],pp230[110],pp228[113],pp226[116],pp224[119],pp222[122],pp220[125],pp218[128],pp216[131],pp214[134],pp212[137],pp210[140],pp208[143],pp206[146],pp204[149],pp202[152],pp200[155],pp199[157],pp198[159],pp197[161],pp196[163],pp195[165],pp194[167],pp193[169],pp192[171],pp191[173],pp190[175],pp189[177],pp188[179],pp187[181],pp186[183],pp185[185],pp184[187],pp183[189],pp182[191],pp181[193],pp180[195],pp179[197],pp178[199],pp177[201],pp176[203],pp175[205],pp174[207],pp173[209],pp172[211],pp171[213],pp172[213],pp173[213],pp174[213],pp175[213],pp176[213],pp177[213],pp178[213],pp179[213],pp180[213],pp181[213],pp182[213],pp183[213],pp184[213],pp185[213],pp186[213],pp187[213],pp188[213],pp189[213],pp190[213],pp191[213],pp192[213],pp193[213],pp194[213],pp195[213],pp196[213],pp197[213],pp198[213],pp199[213],pp200[213],pp201[213],pp202[213],pp203[213],pp204[213],pp205[213],pp206[213],pp207[213],pp208[213],pp209[213],pp210[213],pp211[213],pp212[213],pp213[213]};
    assign in150_2 = {pp53[32],pp53[33],pp53[34],pp53[35],pp53[36],pp53[37],pp53[38],pp53[39],pp53[40],pp53[41],pp53[42],pp53[43],pp53[44],pp53[45],pp53[46],pp52[48],pp51[50],pp50[52],pp49[54],pp48[56],pp47[58],pp46[60],pp45[62],pp44[64],pp43[66],pp42[68],pp41[70],pp40[72],pp39[74],pp38[76],pp37[78],pp36[80],pp35[82],pp34[84],pp33[86],pp32[88],pp31[90],pp30[92],pp29[94],pp28[96],pp27[98],pp9[117],pp7[120],pp7[121],pp7[122],pp7[123],pp7[124],pp7[125],pp7[126],pp7[127],pp7[128],pp7[129],pp7[130],pp7[131],pp7[132],pp7[133],pp7[134],pp7[135],pp7[136],pp7[137],pp7[138],pp7[139],pp7[140],pp7[141],pp7[142],pp7[143],pp7[144],pp7[145],pp7[146],pp7[147],pp7[148],pp7[149],pp7[150],pp7[151],pp7[152],pp7[153],pp7[154],pp7[155],pp7[156],pp6[158],pp5[160],pp4[162],pp3[164],pp2[166],pp1[168],pp0[170],s136[100],s136[101],s136[102],s136[103],s136[104],s136[105],s136[106],s136[107],s136[108],s136[109],s136[110],s136[111],s136[112],s136[113],s136[114],s136[115],s136[116],s136[117],s136[118],s136[119],s136[120],s136[121],s136[122],s136[123],s136[124],s136[125],s136[126],s136[127],s136[128],s137[128],s138[128],s139[128],s140[128],s141[128],s142[128],s143[128],s144[128],s145[128],s146[128],s147[128],s148[128],s149[128],pp0[213],pp1[213],pp2[213],pp3[213],pp4[213],pp5[213],pp6[213],pp7[213],pp8[213],pp9[213],pp214[9],pp216[8],pp218[7],pp220[6],pp222[5],pp224[4],pp226[3],pp228[2],pp230[1],pp232[0],s1[105],s2[105],s3[105],s4[105],s3[107],s2[109],s1[111],s103[10],s103[11],s103[12],s103[13],s103[14],s103[15],s103[16],s103[17],s103[18],s103[19],s103[20],s103[21],s103[22],s103[23],s103[24],s103[25],s103[26],s101[29],s31[100],s30[102],s29[104],s28[106],s27[108],s26[110],s25[112],s24[114],s23[116],s22[118],s21[120],s20[122],s19[124],s18[126],s17[128],s16[130],s15[132],s14[134],s13[136],s12[138],s11[140],s10[142],s149[196],s148[198],s147[200],s146[202],s145[204],s144[206],s143[208],s142[210],s141[212],s140[214],s139[216],s138[218],s137[220],s136[222],s135[224],s134[226],s133[228],s132[230],s131[232],s130[234],s129[236],pp255[46],pp254[48],pp253[50],pp252[52],pp251[54],pp250[56],pp249[58],pp248[60],pp247[62],pp246[64],pp245[66],pp244[68],pp243[70],pp242[72],pp241[74],pp240[76],pp239[78],pp238[80],pp237[82],pp236[84],pp235[86],pp234[88],pp233[90],pp232[92],pp231[94],pp230[96],pp229[98],pp99[229],pp97[232],pp95[235],pp93[238],pp91[241],pp89[244],pp87[247],pp85[250],pp83[253],pp237[100],pp235[103],pp233[106],pp231[109],pp229[112],pp227[115],pp225[118],pp223[121],pp221[124],pp219[127],pp217[130],pp215[133],pp213[136],pp211[139],pp209[142],pp207[145],pp205[148],pp203[151],pp201[154],pp200[156],pp199[158],pp198[160],pp197[162],pp196[164],pp195[166],pp194[168],pp193[170],pp192[172],pp191[174],pp190[176],pp189[178],pp188[180],pp187[182],pp186[184],pp185[186],pp184[188],pp183[190],pp182[192],pp181[194],pp180[196],pp179[198],pp178[200],pp177[202],pp176[204],pp175[206],pp174[208],pp173[210],pp172[212],pp173[212],pp174[212],pp175[212],pp176[212],pp177[212],pp178[212],pp179[212],pp180[212],pp181[212],pp182[212],pp183[212],pp184[212],pp185[212],pp186[212],pp187[212],pp188[212],pp189[212],pp190[212],pp191[212],pp192[212],pp193[212],pp194[212],pp195[212],pp196[212],pp197[212],pp198[212],pp199[212],pp200[212],pp201[212],pp202[212],pp203[212],pp204[212],pp205[212],pp206[212],pp207[212],pp208[212],pp209[212],pp210[212],pp211[212],pp212[212],pp213[212],pp214[212]};
    CLA_342 KS_150(s150, c150, in150_1, in150_2);
    wire[339:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp54[32],pp54[33],pp54[34],pp54[35],pp54[36],pp54[37],pp54[38],pp54[39],pp54[40],pp54[41],pp54[42],pp54[43],pp54[44],pp54[45],pp53[47],pp52[49],pp51[51],pp50[53],pp49[55],pp48[57],pp47[59],pp46[61],pp45[63],pp44[65],pp43[67],pp42[69],pp41[71],pp40[73],pp39[75],pp38[77],pp37[79],pp36[81],pp35[83],pp34[85],pp33[87],pp32[89],pp31[91],pp30[93],pp29[95],pp28[97],pp27[99],pp8[119],pp8[120],pp8[121],pp8[122],pp8[123],pp8[124],pp8[125],pp8[126],pp8[127],pp8[128],pp8[129],pp8[130],pp8[131],pp8[132],pp8[133],pp8[134],pp8[135],pp8[136],pp8[137],pp8[138],pp8[139],pp8[140],pp8[141],pp8[142],pp8[143],pp8[144],pp8[145],pp8[146],pp8[147],pp8[148],pp8[149],pp8[150],pp8[151],pp8[152],pp8[153],pp8[154],pp8[155],pp7[157],pp6[159],pp5[161],pp4[163],pp3[165],pp2[167],pp1[169],pp0[171],s137[100],s137[101],s137[102],s137[103],s137[104],s137[105],s137[106],s137[107],s137[108],s137[109],s137[110],s137[111],s137[112],s137[113],s137[114],s137[115],s137[116],s137[117],s137[118],s137[119],s137[120],s137[121],s137[122],s137[123],s137[124],s137[125],s137[126],s137[127],s138[127],s139[127],s140[127],s141[127],s142[127],s143[127],s144[127],s145[127],s146[127],s147[127],s148[127],s149[127],s150[127],s150[128],s150[129],s150[130],s150[131],s150[132],s150[133],s150[134],s150[135],s150[136],s150[137],s150[138],s150[139],s150[140],s150[141],s150[142],s150[143],s150[144],s150[145],s150[146],s150[147],s150[148],s150[149],s150[150],s150[151],s150[152],s150[153],s150[154],s150[155],s150[156],s150[157],s150[158],s150[159],s150[160],s150[161],s150[162],s150[163],s150[164],s150[165],s150[166],s150[167],s150[168],s150[169],s150[170],s150[171],s150[172],s150[173],s150[174],s150[175],s150[176],s150[177],s150[178],s150[179],s150[180],s150[181],s150[182],s150[183],s150[184],s150[185],s150[186],s150[187],s150[188],s150[189],s150[190],s150[191],s150[192],s150[193],s150[194],s150[195],s149[197],s148[199],s147[201],s146[203],s145[205],s144[207],s143[209],s142[211],s141[213],s140[215],s139[217],s138[219],s137[221],s136[223],s135[225],s134[227],s133[229],s132[231],s131[233],s130[235],s129[237],pp255[47],pp254[49],pp253[51],pp252[53],pp251[55],pp250[57],pp249[59],pp248[61],pp247[63],pp246[65],pp245[67],pp244[69],pp243[71],pp242[73],pp241[75],pp240[77],pp239[79],pp238[81],pp237[83],pp236[85],pp235[87],pp234[89],pp233[91],pp232[93],pp231[95],pp230[97],pp229[99],pp98[231],pp96[234],pp94[237],pp92[240],pp90[243],pp88[246],pp86[249],pp84[252],pp82[255],pp236[102],pp234[105],pp232[108],pp230[111],pp228[114],pp226[117],pp224[120],pp222[123],pp220[126],pp218[129],pp216[132],pp214[135],pp212[138],pp210[141],pp208[144],pp206[147],pp204[150],pp202[153],pp201[155],pp200[157],pp199[159],pp198[161],pp197[163],pp196[165],pp195[167],pp194[169],pp193[171],pp192[173],pp191[175],pp190[177],pp189[179],pp188[181],pp187[183],pp186[185],pp185[187],pp184[189],pp183[191],pp182[193],pp181[195],pp180[197],pp179[199],pp178[201],pp177[203],pp176[205],pp175[207],pp174[209],pp173[211],pp174[211],pp175[211],pp176[211],pp177[211],pp178[211],pp179[211],pp180[211],pp181[211],pp182[211],pp183[211],pp184[211],pp185[211],pp186[211],pp187[211],pp188[211],pp189[211],pp190[211],pp191[211],pp192[211],pp193[211],pp194[211],pp195[211],pp196[211],pp197[211],pp198[211],pp199[211],pp200[211],pp201[211],pp202[211],pp203[211],pp204[211],pp205[211],pp206[211],pp207[211],pp208[211],pp209[211],pp210[211],pp211[211],pp212[211],pp213[211],pp214[211]};
    assign in151_2 = {pp55[31],pp55[32],pp55[33],pp55[34],pp55[35],pp55[36],pp55[37],pp55[38],pp55[39],pp55[40],pp55[41],pp55[42],pp55[43],pp55[44],pp54[46],pp53[48],pp52[50],pp51[52],pp50[54],pp49[56],pp48[58],pp47[60],pp46[62],pp45[64],pp44[66],pp43[68],pp42[70],pp41[72],pp40[74],pp39[76],pp38[78],pp37[80],pp36[82],pp35[84],pp34[86],pp33[88],pp32[90],pp31[92],pp30[94],pp29[96],pp28[98],pp9[118],pp9[119],pp9[120],pp9[121],pp9[122],pp9[123],pp9[124],pp9[125],pp9[126],pp9[127],pp9[128],pp9[129],pp9[130],pp9[131],pp9[132],pp9[133],pp9[134],pp9[135],pp9[136],pp9[137],pp9[138],pp9[139],pp9[140],pp9[141],pp9[142],pp9[143],pp9[144],pp9[145],pp9[146],pp9[147],pp9[148],pp9[149],pp9[150],pp9[151],pp9[152],pp9[153],pp9[154],pp8[156],pp7[158],pp6[160],pp5[162],pp4[164],pp3[166],pp2[168],pp1[170],pp0[172],s138[100],s138[101],s138[102],s138[103],s138[104],s138[105],s138[106],s138[107],s138[108],s138[109],s138[110],s138[111],s138[112],s138[113],s138[114],s138[115],s138[116],s138[117],s138[118],s138[119],s138[120],s138[121],s138[122],s138[123],s138[124],s138[125],s138[126],s139[126],s140[126],s141[126],s142[126],s143[126],s144[126],s145[126],s146[126],s147[126],s148[126],s149[126],s150[126],pp0[212],pp1[212],pp2[212],pp3[212],pp4[212],pp5[212],pp6[212],pp7[212],pp8[212],pp9[212],pp213[9],pp215[8],pp217[7],pp219[6],pp221[5],pp223[4],pp225[3],pp227[2],pp229[1],pp231[0],s1[104],s2[104],s3[104],s4[104],s5[104],s4[106],s3[108],s2[110],s1[112],s104[10],s104[11],s104[12],s104[13],s104[14],s104[15],s104[16],s104[17],s104[18],s104[19],s104[20],s104[21],s104[22],s104[23],s104[24],s104[25],s102[28],s100[31],s31[101],s30[103],s29[105],s28[107],s27[109],s26[111],s25[113],s24[115],s23[117],s22[119],s21[121],s20[123],s19[125],s18[127],s17[129],s16[131],s15[133],s14[135],s13[137],s12[139],s11[141],s10[143],s150[196],s149[198],s148[200],s147[202],s146[204],s145[206],s144[208],s143[210],s142[212],s141[214],s140[216],s139[218],s138[220],s137[222],s136[224],s135[226],s134[228],s133[230],s132[232],s131[234],s130[236],s129[238],pp255[48],pp254[50],pp253[52],pp252[54],pp251[56],pp250[58],pp249[60],pp248[62],pp247[64],pp246[66],pp245[68],pp244[70],pp243[72],pp242[74],pp241[76],pp240[78],pp239[80],pp238[82],pp237[84],pp236[86],pp235[88],pp234[90],pp233[92],pp232[94],pp231[96],pp230[98],pp99[230],pp97[233],pp95[236],pp93[239],pp91[242],pp89[245],pp87[248],pp85[251],pp83[254],pp237[101],pp235[104],pp233[107],pp231[110],pp229[113],pp227[116],pp225[119],pp223[122],pp221[125],pp219[128],pp217[131],pp215[134],pp213[137],pp211[140],pp209[143],pp207[146],pp205[149],pp203[152],pp202[154],pp201[156],pp200[158],pp199[160],pp198[162],pp197[164],pp196[166],pp195[168],pp194[170],pp193[172],pp192[174],pp191[176],pp190[178],pp189[180],pp188[182],pp187[184],pp186[186],pp185[188],pp184[190],pp183[192],pp182[194],pp181[196],pp180[198],pp179[200],pp178[202],pp177[204],pp176[206],pp175[208],pp174[210],pp175[210],pp176[210],pp177[210],pp178[210],pp179[210],pp180[210],pp181[210],pp182[210],pp183[210],pp184[210],pp185[210],pp186[210],pp187[210],pp188[210],pp189[210],pp190[210],pp191[210],pp192[210],pp193[210],pp194[210],pp195[210],pp196[210],pp197[210],pp198[210],pp199[210],pp200[210],pp201[210],pp202[210],pp203[210],pp204[210],pp205[210],pp206[210],pp207[210],pp208[210],pp209[210],pp210[210],pp211[210],pp212[210],pp213[210],pp214[210],pp215[210]};
    CLA_340 KS_151(s151, c151, in151_1, in151_2);
    wire[337:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp56[31],pp56[32],pp56[33],pp56[34],pp56[35],pp56[36],pp56[37],pp56[38],pp56[39],pp56[40],pp56[41],pp56[42],pp56[43],pp55[45],pp54[47],pp53[49],pp52[51],pp51[53],pp50[55],pp49[57],pp48[59],pp47[61],pp46[63],pp45[65],pp44[67],pp43[69],pp42[71],pp41[73],pp40[75],pp39[77],pp38[79],pp37[81],pp36[83],pp35[85],pp34[87],pp33[89],pp32[91],pp31[93],pp30[95],pp29[97],pp28[99],pp29[99],pp30[99],pp31[99],pp32[99],pp33[99],pp34[99],pp35[99],pp36[99],pp37[99],pp38[99],pp39[99],pp40[99],pp41[99],pp42[99],pp43[99],pp44[99],pp45[99],pp46[99],pp47[99],pp48[99],pp49[99],pp50[99],pp51[99],pp52[99],pp53[99],pp54[99],pp55[99],pp56[99],pp57[99],pp58[99],pp59[99],pp60[99],pp61[99],pp62[99],pp63[99],pp64[99],pp9[155],pp8[157],pp7[159],pp6[161],pp5[163],pp4[165],pp3[167],pp2[169],pp1[171],pp0[173],s139[100],s139[101],s139[102],s139[103],s139[104],s139[105],s139[106],s139[107],s139[108],s139[109],s139[110],s139[111],s139[112],s139[113],s139[114],s139[115],s139[116],s139[117],s139[118],s139[119],s139[120],s139[121],s139[122],s139[123],s139[124],s139[125],s140[125],s141[125],s142[125],s143[125],s144[125],s145[125],s146[125],s147[125],s148[125],s149[125],s150[125],s151[125],s151[126],s151[127],s151[128],s151[129],s151[130],s151[131],s151[132],s151[133],s151[134],s151[135],s151[136],s151[137],s151[138],s151[139],s151[140],s151[141],s151[142],s151[143],s151[144],s151[145],s151[146],s151[147],s151[148],s151[149],s151[150],s151[151],s151[152],s151[153],s151[154],s151[155],s151[156],s151[157],s151[158],s151[159],s151[160],s151[161],s151[162],s151[163],s151[164],s151[165],s151[166],s151[167],s151[168],s151[169],s151[170],s151[171],s151[172],s151[173],s151[174],s151[175],s151[176],s151[177],s151[178],s151[179],s151[180],s151[181],s151[182],s151[183],s151[184],s151[185],s151[186],s151[187],s151[188],s151[189],s151[190],s151[191],s151[192],s151[193],s151[194],s151[195],s150[197],s149[199],s148[201],s147[203],s146[205],s145[207],s144[209],s143[211],s142[213],s141[215],s140[217],s139[219],s138[221],s137[223],s136[225],s135[227],s134[229],s133[231],s132[233],s131[235],s130[237],s129[239],pp255[49],pp254[51],pp253[53],pp252[55],pp251[57],pp250[59],pp249[61],pp248[63],pp247[65],pp246[67],pp245[69],pp244[71],pp243[73],pp242[75],pp241[77],pp240[79],pp239[81],pp238[83],pp237[85],pp236[87],pp235[89],pp234[91],pp233[93],pp232[95],pp231[97],pp230[99],pp98[232],pp96[235],pp94[238],pp92[241],pp90[244],pp88[247],pp86[250],pp84[253],pp238[100],pp236[103],pp234[106],pp232[109],pp230[112],pp228[115],pp226[118],pp224[121],pp222[124],pp220[127],pp218[130],pp216[133],pp214[136],pp212[139],pp210[142],pp208[145],pp206[148],pp204[151],pp203[153],pp202[155],pp201[157],pp200[159],pp199[161],pp198[163],pp197[165],pp196[167],pp195[169],pp194[171],pp193[173],pp192[175],pp191[177],pp190[179],pp189[181],pp188[183],pp187[185],pp186[187],pp185[189],pp184[191],pp183[193],pp182[195],pp181[197],pp180[199],pp179[201],pp178[203],pp177[205],pp176[207],pp175[209],pp176[209],pp177[209],pp178[209],pp179[209],pp180[209],pp181[209],pp182[209],pp183[209],pp184[209],pp185[209],pp186[209],pp187[209],pp188[209],pp189[209],pp190[209],pp191[209],pp192[209],pp193[209],pp194[209],pp195[209],pp196[209],pp197[209],pp198[209],pp199[209],pp200[209],pp201[209],pp202[209],pp203[209],pp204[209],pp205[209],pp206[209],pp207[209],pp208[209],pp209[209],pp210[209],pp211[209],pp212[209],pp213[209],pp214[209],pp215[209]};
    assign in152_2 = {pp57[30],pp57[31],pp57[32],pp57[33],pp57[34],pp57[35],pp57[36],pp57[37],pp57[38],pp57[39],pp57[40],pp57[41],pp57[42],pp56[44],pp55[46],pp54[48],pp53[50],pp52[52],pp51[54],pp50[56],pp49[58],pp48[60],pp47[62],pp46[64],pp45[66],pp44[68],pp43[70],pp42[72],pp41[74],pp40[76],pp39[78],pp38[80],pp37[82],pp36[84],pp35[86],pp34[88],pp33[90],pp32[92],pp31[94],pp30[96],pp29[98],pp30[98],pp31[98],pp32[98],pp33[98],pp34[98],pp35[98],pp36[98],pp37[98],pp38[98],pp39[98],pp40[98],pp41[98],pp42[98],pp43[98],pp44[98],pp45[98],pp46[98],pp47[98],pp48[98],pp49[98],pp50[98],pp51[98],pp52[98],pp53[98],pp54[98],pp55[98],pp56[98],pp57[98],pp58[98],pp59[98],pp60[98],pp61[98],pp62[98],pp63[98],pp64[98],pp65[98],pp65[99],pp9[156],pp8[158],pp7[160],pp6[162],pp5[164],pp4[166],pp3[168],pp2[170],pp1[172],pp0[174],s140[100],s140[101],s140[102],s140[103],s140[104],s140[105],s140[106],s140[107],s140[108],s140[109],s140[110],s140[111],s140[112],s140[113],s140[114],s140[115],s140[116],s140[117],s140[118],s140[119],s140[120],s140[121],s140[122],s140[123],s140[124],s141[124],s142[124],s143[124],s144[124],s145[124],s146[124],s147[124],s148[124],s149[124],s150[124],s151[124],pp0[211],pp1[211],pp2[211],pp3[211],pp4[211],pp5[211],pp6[211],pp7[211],pp8[211],pp9[211],pp212[9],pp214[8],pp216[7],pp218[6],pp220[5],pp222[4],pp224[3],pp226[2],pp228[1],pp230[0],s1[103],s2[103],s3[103],s4[103],s5[103],s6[103],s5[105],s4[107],s3[109],s2[111],s1[113],s105[10],s105[11],s105[12],s105[13],s105[14],s105[15],s105[16],s105[17],s105[18],s105[19],s105[20],s105[21],s105[22],s105[23],s105[24],s103[27],s101[30],s32[100],s31[102],s30[104],s29[106],s28[108],s27[110],s26[112],s25[114],s24[116],s23[118],s22[120],s21[122],s20[124],s19[126],s18[128],s17[130],s16[132],s15[134],s14[136],s13[138],s12[140],s11[142],s10[144],s151[196],s150[198],s149[200],s148[202],s147[204],s146[206],s145[208],s144[210],s143[212],s142[214],s141[216],s140[218],s139[220],s138[222],s137[224],s136[226],s135[228],s134[230],s133[232],s132[234],s131[236],s130[238],s129[240],pp255[50],pp254[52],pp253[54],pp252[56],pp251[58],pp250[60],pp249[62],pp248[64],pp247[66],pp246[68],pp245[70],pp244[72],pp243[74],pp242[76],pp241[78],pp240[80],pp239[82],pp238[84],pp237[86],pp236[88],pp235[90],pp234[92],pp233[94],pp232[96],pp231[98],pp99[231],pp97[234],pp95[237],pp93[240],pp91[243],pp89[246],pp87[249],pp85[252],pp83[255],pp237[102],pp235[105],pp233[108],pp231[111],pp229[114],pp227[117],pp225[120],pp223[123],pp221[126],pp219[129],pp217[132],pp215[135],pp213[138],pp211[141],pp209[144],pp207[147],pp205[150],pp204[152],pp203[154],pp202[156],pp201[158],pp200[160],pp199[162],pp198[164],pp197[166],pp196[168],pp195[170],pp194[172],pp193[174],pp192[176],pp191[178],pp190[180],pp189[182],pp188[184],pp187[186],pp186[188],pp185[190],pp184[192],pp183[194],pp182[196],pp181[198],pp180[200],pp179[202],pp178[204],pp177[206],pp176[208],pp177[208],pp178[208],pp179[208],pp180[208],pp181[208],pp182[208],pp183[208],pp184[208],pp185[208],pp186[208],pp187[208],pp188[208],pp189[208],pp190[208],pp191[208],pp192[208],pp193[208],pp194[208],pp195[208],pp196[208],pp197[208],pp198[208],pp199[208],pp200[208],pp201[208],pp202[208],pp203[208],pp204[208],pp205[208],pp206[208],pp207[208],pp208[208],pp209[208],pp210[208],pp211[208],pp212[208],pp213[208],pp214[208],pp215[208],pp216[208]};
    CLA_338 KS_152(s152, c152, in152_1, in152_2);
    wire[335:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp58[30],pp58[31],pp58[32],pp58[33],pp58[34],pp58[35],pp58[36],pp58[37],pp58[38],pp58[39],pp58[40],pp58[41],pp57[43],pp56[45],pp55[47],pp54[49],pp53[51],pp52[53],pp51[55],pp50[57],pp49[59],pp48[61],pp47[63],pp46[65],pp45[67],pp44[69],pp43[71],pp42[73],pp41[75],pp40[77],pp39[79],pp38[81],pp37[83],pp36[85],pp35[87],pp34[89],pp33[91],pp32[93],pp31[95],pp30[97],pp31[97],pp32[97],pp33[97],pp34[97],pp35[97],pp36[97],pp37[97],pp38[97],pp39[97],pp40[97],pp41[97],pp42[97],pp43[97],pp44[97],pp45[97],pp46[97],pp47[97],pp48[97],pp49[97],pp50[97],pp51[97],pp52[97],pp53[97],pp54[97],pp55[97],pp56[97],pp57[97],pp58[97],pp59[97],pp60[97],pp61[97],pp62[97],pp63[97],pp64[97],pp65[97],pp66[97],pp66[98],pp66[99],pp9[157],pp8[159],pp7[161],pp6[163],pp5[165],pp4[167],pp3[169],pp2[171],pp1[173],pp0[175],s141[100],s141[101],s141[102],s141[103],s141[104],s141[105],s141[106],s141[107],s141[108],s141[109],s141[110],s141[111],s141[112],s141[113],s141[114],s141[115],s141[116],s141[117],s141[118],s141[119],s141[120],s141[121],s141[122],s141[123],s142[123],s143[123],s144[123],s145[123],s146[123],s147[123],s148[123],s149[123],s150[123],s151[123],s152[123],s152[124],s152[125],s152[126],s152[127],s152[128],s152[129],s152[130],s152[131],s152[132],s152[133],s152[134],s152[135],s152[136],s152[137],s152[138],s152[139],s152[140],s152[141],s152[142],s152[143],s152[144],s152[145],s152[146],s152[147],s152[148],s152[149],s152[150],s152[151],s152[152],s152[153],s152[154],s152[155],s152[156],s152[157],s152[158],s152[159],s152[160],s152[161],s152[162],s152[163],s152[164],s152[165],s152[166],s152[167],s152[168],s152[169],s152[170],s152[171],s152[172],s152[173],s152[174],s152[175],s152[176],s152[177],s152[178],s152[179],s152[180],s152[181],s152[182],s152[183],s152[184],s152[185],s152[186],s152[187],s152[188],s152[189],s152[190],s152[191],s152[192],s152[193],s152[194],s152[195],s151[197],s150[199],s149[201],s148[203],s147[205],s146[207],s145[209],s144[211],s143[213],s142[215],s141[217],s140[219],s139[221],s138[223],s137[225],s136[227],s135[229],s134[231],s133[233],s132[235],s131[237],s130[239],s129[241],pp255[51],pp254[53],pp253[55],pp252[57],pp251[59],pp250[61],pp249[63],pp248[65],pp247[67],pp246[69],pp245[71],pp244[73],pp243[75],pp242[77],pp241[79],pp240[81],pp239[83],pp238[85],pp237[87],pp236[89],pp235[91],pp234[93],pp233[95],pp232[97],pp231[99],pp98[233],pp96[236],pp94[239],pp92[242],pp90[245],pp88[248],pp86[251],pp84[254],pp238[101],pp236[104],pp234[107],pp232[110],pp230[113],pp228[116],pp226[119],pp224[122],pp222[125],pp220[128],pp218[131],pp216[134],pp214[137],pp212[140],pp210[143],pp208[146],pp206[149],pp205[151],pp204[153],pp203[155],pp202[157],pp201[159],pp200[161],pp199[163],pp198[165],pp197[167],pp196[169],pp195[171],pp194[173],pp193[175],pp192[177],pp191[179],pp190[181],pp189[183],pp188[185],pp187[187],pp186[189],pp185[191],pp184[193],pp183[195],pp182[197],pp181[199],pp180[201],pp179[203],pp178[205],pp177[207],pp178[207],pp179[207],pp180[207],pp181[207],pp182[207],pp183[207],pp184[207],pp185[207],pp186[207],pp187[207],pp188[207],pp189[207],pp190[207],pp191[207],pp192[207],pp193[207],pp194[207],pp195[207],pp196[207],pp197[207],pp198[207],pp199[207],pp200[207],pp201[207],pp202[207],pp203[207],pp204[207],pp205[207],pp206[207],pp207[207],pp208[207],pp209[207],pp210[207],pp211[207],pp212[207],pp213[207],pp214[207],pp215[207],pp216[207]};
    assign in153_2 = {pp59[29],pp59[30],pp59[31],pp59[32],pp59[33],pp59[34],pp59[35],pp59[36],pp59[37],pp59[38],pp59[39],pp59[40],pp58[42],pp57[44],pp56[46],pp55[48],pp54[50],pp53[52],pp52[54],pp51[56],pp50[58],pp49[60],pp48[62],pp47[64],pp46[66],pp45[68],pp44[70],pp43[72],pp42[74],pp41[76],pp40[78],pp39[80],pp38[82],pp37[84],pp36[86],pp35[88],pp34[90],pp33[92],pp32[94],pp31[96],pp32[96],pp33[96],pp34[96],pp35[96],pp36[96],pp37[96],pp38[96],pp39[96],pp40[96],pp41[96],pp42[96],pp43[96],pp44[96],pp45[96],pp46[96],pp47[96],pp48[96],pp49[96],pp50[96],pp51[96],pp52[96],pp53[96],pp54[96],pp55[96],pp56[96],pp57[96],pp58[96],pp59[96],pp60[96],pp61[96],pp62[96],pp63[96],pp64[96],pp65[96],pp66[96],pp67[96],pp67[97],pp67[98],pp67[99],pp9[158],pp8[160],pp7[162],pp6[164],pp5[166],pp4[168],pp3[170],pp2[172],pp1[174],pp0[176],s142[100],s142[101],s142[102],s142[103],s142[104],s142[105],s142[106],s142[107],s142[108],s142[109],s142[110],s142[111],s142[112],s142[113],s142[114],s142[115],s142[116],s142[117],s142[118],s142[119],s142[120],s142[121],s142[122],s143[122],s144[122],s145[122],s146[122],s147[122],s148[122],s149[122],s150[122],s151[122],s152[122],pp0[210],pp1[210],pp2[210],pp3[210],pp4[210],pp5[210],pp6[210],pp7[210],pp8[210],pp9[210],pp211[9],pp213[8],pp215[7],pp217[6],pp219[5],pp221[4],pp223[3],pp225[2],pp227[1],pp229[0],s1[102],s2[102],s3[102],s4[102],s5[102],s6[102],s7[102],s6[104],s5[106],s4[108],s3[110],s2[112],s1[114],s106[10],s106[11],s106[12],s106[13],s106[14],s106[15],s106[16],s106[17],s106[18],s106[19],s106[20],s106[21],s106[22],s106[23],s104[26],s102[29],s100[32],s32[101],s31[103],s30[105],s29[107],s28[109],s27[111],s26[113],s25[115],s24[117],s23[119],s22[121],s21[123],s20[125],s19[127],s18[129],s17[131],s16[133],s15[135],s14[137],s13[139],s12[141],s11[143],s10[145],s152[196],s151[198],s150[200],s149[202],s148[204],s147[206],s146[208],s145[210],s144[212],s143[214],s142[216],s141[218],s140[220],s139[222],s138[224],s137[226],s136[228],s135[230],s134[232],s133[234],s132[236],s131[238],s130[240],s129[242],pp255[52],pp254[54],pp253[56],pp252[58],pp251[60],pp250[62],pp249[64],pp248[66],pp247[68],pp246[70],pp245[72],pp244[74],pp243[76],pp242[78],pp241[80],pp240[82],pp239[84],pp238[86],pp237[88],pp236[90],pp235[92],pp234[94],pp233[96],pp232[98],pp99[232],pp97[235],pp95[238],pp93[241],pp91[244],pp89[247],pp87[250],pp85[253],pp239[100],pp237[103],pp235[106],pp233[109],pp231[112],pp229[115],pp227[118],pp225[121],pp223[124],pp221[127],pp219[130],pp217[133],pp215[136],pp213[139],pp211[142],pp209[145],pp207[148],pp206[150],pp205[152],pp204[154],pp203[156],pp202[158],pp201[160],pp200[162],pp199[164],pp198[166],pp197[168],pp196[170],pp195[172],pp194[174],pp193[176],pp192[178],pp191[180],pp190[182],pp189[184],pp188[186],pp187[188],pp186[190],pp185[192],pp184[194],pp183[196],pp182[198],pp181[200],pp180[202],pp179[204],pp178[206],pp179[206],pp180[206],pp181[206],pp182[206],pp183[206],pp184[206],pp185[206],pp186[206],pp187[206],pp188[206],pp189[206],pp190[206],pp191[206],pp192[206],pp193[206],pp194[206],pp195[206],pp196[206],pp197[206],pp198[206],pp199[206],pp200[206],pp201[206],pp202[206],pp203[206],pp204[206],pp205[206],pp206[206],pp207[206],pp208[206],pp209[206],pp210[206],pp211[206],pp212[206],pp213[206],pp214[206],pp215[206],pp216[206],pp217[206]};
    CLA_336 KS_153(s153, c153, in153_1, in153_2);
    wire[333:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp60[29],pp60[30],pp60[31],pp60[32],pp60[33],pp60[34],pp60[35],pp60[36],pp60[37],pp60[38],pp60[39],pp59[41],pp58[43],pp57[45],pp56[47],pp55[49],pp54[51],pp53[53],pp52[55],pp51[57],pp50[59],pp49[61],pp48[63],pp47[65],pp46[67],pp45[69],pp44[71],pp43[73],pp42[75],pp41[77],pp40[79],pp39[81],pp38[83],pp37[85],pp36[87],pp35[89],pp34[91],pp33[93],pp32[95],pp33[95],pp34[95],pp35[95],pp36[95],pp37[95],pp38[95],pp39[95],pp40[95],pp41[95],pp42[95],pp43[95],pp44[95],pp45[95],pp46[95],pp47[95],pp48[95],pp49[95],pp50[95],pp51[95],pp52[95],pp53[95],pp54[95],pp55[95],pp56[95],pp57[95],pp58[95],pp59[95],pp60[95],pp61[95],pp62[95],pp63[95],pp64[95],pp65[95],pp66[95],pp67[95],pp68[95],pp68[96],pp68[97],pp68[98],pp68[99],pp9[159],pp8[161],pp7[163],pp6[165],pp5[167],pp4[169],pp3[171],pp2[173],pp1[175],pp0[177],s143[100],s143[101],s143[102],s143[103],s143[104],s143[105],s143[106],s143[107],s143[108],s143[109],s143[110],s143[111],s143[112],s143[113],s143[114],s143[115],s143[116],s143[117],s143[118],s143[119],s143[120],s143[121],s144[121],s145[121],s146[121],s147[121],s148[121],s149[121],s150[121],s151[121],s152[121],s153[121],s153[122],s153[123],s153[124],s153[125],s153[126],s153[127],s153[128],s153[129],s153[130],s153[131],s153[132],s153[133],s153[134],s153[135],s153[136],s153[137],s153[138],s153[139],s153[140],s153[141],s153[142],s153[143],s153[144],s153[145],s153[146],s153[147],s153[148],s153[149],s153[150],s153[151],s153[152],s153[153],s153[154],s153[155],s153[156],s153[157],s153[158],s153[159],s153[160],s153[161],s153[162],s153[163],s153[164],s153[165],s153[166],s153[167],s153[168],s153[169],s153[170],s153[171],s153[172],s153[173],s153[174],s153[175],s153[176],s153[177],s153[178],s153[179],s153[180],s153[181],s153[182],s153[183],s153[184],s153[185],s153[186],s153[187],s153[188],s153[189],s153[190],s153[191],s153[192],s153[193],s153[194],s153[195],s152[197],s151[199],s150[201],s149[203],s148[205],s147[207],s146[209],s145[211],s144[213],s143[215],s142[217],s141[219],s140[221],s139[223],s138[225],s137[227],s136[229],s135[231],s134[233],s133[235],s132[237],s131[239],s130[241],s129[243],pp255[53],pp254[55],pp253[57],pp252[59],pp251[61],pp250[63],pp249[65],pp248[67],pp247[69],pp246[71],pp245[73],pp244[75],pp243[77],pp242[79],pp241[81],pp240[83],pp239[85],pp238[87],pp237[89],pp236[91],pp235[93],pp234[95],pp233[97],pp232[99],pp98[234],pp96[237],pp94[240],pp92[243],pp90[246],pp88[249],pp86[252],pp84[255],pp238[102],pp236[105],pp234[108],pp232[111],pp230[114],pp228[117],pp226[120],pp224[123],pp222[126],pp220[129],pp218[132],pp216[135],pp214[138],pp212[141],pp210[144],pp208[147],pp207[149],pp206[151],pp205[153],pp204[155],pp203[157],pp202[159],pp201[161],pp200[163],pp199[165],pp198[167],pp197[169],pp196[171],pp195[173],pp194[175],pp193[177],pp192[179],pp191[181],pp190[183],pp189[185],pp188[187],pp187[189],pp186[191],pp185[193],pp184[195],pp183[197],pp182[199],pp181[201],pp180[203],pp179[205],pp180[205],pp181[205],pp182[205],pp183[205],pp184[205],pp185[205],pp186[205],pp187[205],pp188[205],pp189[205],pp190[205],pp191[205],pp192[205],pp193[205],pp194[205],pp195[205],pp196[205],pp197[205],pp198[205],pp199[205],pp200[205],pp201[205],pp202[205],pp203[205],pp204[205],pp205[205],pp206[205],pp207[205],pp208[205],pp209[205],pp210[205],pp211[205],pp212[205],pp213[205],pp214[205],pp215[205],pp216[205],pp217[205]};
    assign in154_2 = {pp61[28],pp61[29],pp61[30],pp61[31],pp61[32],pp61[33],pp61[34],pp61[35],pp61[36],pp61[37],pp61[38],pp60[40],pp59[42],pp58[44],pp57[46],pp56[48],pp55[50],pp54[52],pp53[54],pp52[56],pp51[58],pp50[60],pp49[62],pp48[64],pp47[66],pp46[68],pp45[70],pp44[72],pp43[74],pp42[76],pp41[78],pp40[80],pp39[82],pp38[84],pp37[86],pp36[88],pp35[90],pp34[92],pp33[94],pp34[94],pp35[94],pp36[94],pp37[94],pp38[94],pp39[94],pp40[94],pp41[94],pp42[94],pp43[94],pp44[94],pp45[94],pp46[94],pp47[94],pp48[94],pp49[94],pp50[94],pp51[94],pp52[94],pp53[94],pp54[94],pp55[94],pp56[94],pp57[94],pp58[94],pp59[94],pp60[94],pp61[94],pp62[94],pp63[94],pp64[94],pp65[94],pp66[94],pp67[94],pp68[94],pp69[94],pp69[95],pp69[96],pp69[97],pp69[98],pp69[99],pp9[160],pp8[162],pp7[164],pp6[166],pp5[168],pp4[170],pp3[172],pp2[174],pp1[176],pp0[178],s144[100],s144[101],s144[102],s144[103],s144[104],s144[105],s144[106],s144[107],s144[108],s144[109],s144[110],s144[111],s144[112],s144[113],s144[114],s144[115],s144[116],s144[117],s144[118],s144[119],s144[120],s145[120],s146[120],s147[120],s148[120],s149[120],s150[120],s151[120],s152[120],s153[120],pp0[209],pp1[209],pp2[209],pp3[209],pp4[209],pp5[209],pp6[209],pp7[209],pp8[209],pp9[209],pp210[9],pp212[8],pp214[7],pp216[6],pp218[5],pp220[4],pp222[3],pp224[2],pp226[1],pp228[0],s1[101],s2[101],s3[101],s4[101],s5[101],s6[101],s7[101],s8[101],s7[103],s6[105],s5[107],s4[109],s3[111],s2[113],s1[115],s107[10],s107[11],s107[12],s107[13],s107[14],s107[15],s107[16],s107[17],s107[18],s107[19],s107[20],s107[21],s107[22],s105[25],s103[28],s101[31],s33[100],s32[102],s31[104],s30[106],s29[108],s28[110],s27[112],s26[114],s25[116],s24[118],s23[120],s22[122],s21[124],s20[126],s19[128],s18[130],s17[132],s16[134],s15[136],s14[138],s13[140],s12[142],s11[144],s10[146],s153[196],s152[198],s151[200],s150[202],s149[204],s148[206],s147[208],s146[210],s145[212],s144[214],s143[216],s142[218],s141[220],s140[222],s139[224],s138[226],s137[228],s136[230],s135[232],s134[234],s133[236],s132[238],s131[240],s130[242],s129[244],pp255[54],pp254[56],pp253[58],pp252[60],pp251[62],pp250[64],pp249[66],pp248[68],pp247[70],pp246[72],pp245[74],pp244[76],pp243[78],pp242[80],pp241[82],pp240[84],pp239[86],pp238[88],pp237[90],pp236[92],pp235[94],pp234[96],pp233[98],pp99[233],pp97[236],pp95[239],pp93[242],pp91[245],pp89[248],pp87[251],pp85[254],pp239[101],pp237[104],pp235[107],pp233[110],pp231[113],pp229[116],pp227[119],pp225[122],pp223[125],pp221[128],pp219[131],pp217[134],pp215[137],pp213[140],pp211[143],pp209[146],pp208[148],pp207[150],pp206[152],pp205[154],pp204[156],pp203[158],pp202[160],pp201[162],pp200[164],pp199[166],pp198[168],pp197[170],pp196[172],pp195[174],pp194[176],pp193[178],pp192[180],pp191[182],pp190[184],pp189[186],pp188[188],pp187[190],pp186[192],pp185[194],pp184[196],pp183[198],pp182[200],pp181[202],pp180[204],pp181[204],pp182[204],pp183[204],pp184[204],pp185[204],pp186[204],pp187[204],pp188[204],pp189[204],pp190[204],pp191[204],pp192[204],pp193[204],pp194[204],pp195[204],pp196[204],pp197[204],pp198[204],pp199[204],pp200[204],pp201[204],pp202[204],pp203[204],pp204[204],pp205[204],pp206[204],pp207[204],pp208[204],pp209[204],pp210[204],pp211[204],pp212[204],pp213[204],pp214[204],pp215[204],pp216[204],pp217[204],pp218[204]};
    CLA_334 KS_154(s154, c154, in154_1, in154_2);
    wire[331:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp62[28],pp62[29],pp62[30],pp62[31],pp62[32],pp62[33],pp62[34],pp62[35],pp62[36],pp62[37],pp61[39],pp60[41],pp59[43],pp58[45],pp57[47],pp56[49],pp55[51],pp54[53],pp53[55],pp52[57],pp51[59],pp50[61],pp49[63],pp48[65],pp47[67],pp46[69],pp45[71],pp44[73],pp43[75],pp42[77],pp41[79],pp40[81],pp39[83],pp38[85],pp37[87],pp36[89],pp35[91],pp34[93],pp35[93],pp36[93],pp37[93],pp38[93],pp39[93],pp40[93],pp41[93],pp42[93],pp43[93],pp44[93],pp45[93],pp46[93],pp47[93],pp48[93],pp49[93],pp50[93],pp51[93],pp52[93],pp53[93],pp54[93],pp55[93],pp56[93],pp57[93],pp58[93],pp59[93],pp60[93],pp61[93],pp62[93],pp63[93],pp64[93],pp65[93],pp66[93],pp67[93],pp68[93],pp69[93],pp70[93],pp70[94],pp70[95],pp70[96],pp70[97],pp70[98],pp70[99],pp9[161],pp8[163],pp7[165],pp6[167],pp5[169],pp4[171],pp3[173],pp2[175],pp1[177],pp0[179],s145[100],s145[101],s145[102],s145[103],s145[104],s145[105],s145[106],s145[107],s145[108],s145[109],s145[110],s145[111],s145[112],s145[113],s145[114],s145[115],s145[116],s145[117],s145[118],s145[119],s146[119],s147[119],s148[119],s149[119],s150[119],s151[119],s152[119],s153[119],s154[119],s154[120],s154[121],s154[122],s154[123],s154[124],s154[125],s154[126],s154[127],s154[128],s154[129],s154[130],s154[131],s154[132],s154[133],s154[134],s154[135],s154[136],s154[137],s154[138],s154[139],s154[140],s154[141],s154[142],s154[143],s154[144],s154[145],s154[146],s154[147],s154[148],s154[149],s154[150],s154[151],s154[152],s154[153],s154[154],s154[155],s154[156],s154[157],s154[158],s154[159],s154[160],s154[161],s154[162],s154[163],s154[164],s154[165],s154[166],s154[167],s154[168],s154[169],s154[170],s154[171],s154[172],s154[173],s154[174],s154[175],s154[176],s154[177],s154[178],s154[179],s154[180],s154[181],s154[182],s154[183],s154[184],s154[185],s154[186],s154[187],s154[188],s154[189],s154[190],s154[191],s154[192],s154[193],s154[194],s154[195],s153[197],s152[199],s151[201],s150[203],s149[205],s148[207],s147[209],s146[211],s145[213],s144[215],s143[217],s142[219],s141[221],s140[223],s139[225],s138[227],s137[229],s136[231],s135[233],s134[235],s133[237],s132[239],s131[241],s130[243],s129[245],pp255[55],pp254[57],pp253[59],pp252[61],pp251[63],pp250[65],pp249[67],pp248[69],pp247[71],pp246[73],pp245[75],pp244[77],pp243[79],pp242[81],pp241[83],pp240[85],pp239[87],pp238[89],pp237[91],pp236[93],pp235[95],pp234[97],pp233[99],pp98[235],pp96[238],pp94[241],pp92[244],pp90[247],pp88[250],pp86[253],pp240[100],pp238[103],pp236[106],pp234[109],pp232[112],pp230[115],pp228[118],pp226[121],pp224[124],pp222[127],pp220[130],pp218[133],pp216[136],pp214[139],pp212[142],pp210[145],pp209[147],pp208[149],pp207[151],pp206[153],pp205[155],pp204[157],pp203[159],pp202[161],pp201[163],pp200[165],pp199[167],pp198[169],pp197[171],pp196[173],pp195[175],pp194[177],pp193[179],pp192[181],pp191[183],pp190[185],pp189[187],pp188[189],pp187[191],pp186[193],pp185[195],pp184[197],pp183[199],pp182[201],pp181[203],pp182[203],pp183[203],pp184[203],pp185[203],pp186[203],pp187[203],pp188[203],pp189[203],pp190[203],pp191[203],pp192[203],pp193[203],pp194[203],pp195[203],pp196[203],pp197[203],pp198[203],pp199[203],pp200[203],pp201[203],pp202[203],pp203[203],pp204[203],pp205[203],pp206[203],pp207[203],pp208[203],pp209[203],pp210[203],pp211[203],pp212[203],pp213[203],pp214[203],pp215[203],pp216[203],pp217[203],pp218[203]};
    assign in155_2 = {pp63[27],pp63[28],pp63[29],pp63[30],pp63[31],pp63[32],pp63[33],pp63[34],pp63[35],pp63[36],pp62[38],pp61[40],pp60[42],pp59[44],pp58[46],pp57[48],pp56[50],pp55[52],pp54[54],pp53[56],pp52[58],pp51[60],pp50[62],pp49[64],pp48[66],pp47[68],pp46[70],pp45[72],pp44[74],pp43[76],pp42[78],pp41[80],pp40[82],pp39[84],pp38[86],pp37[88],pp36[90],pp35[92],pp36[92],pp37[92],pp38[92],pp39[92],pp40[92],pp41[92],pp42[92],pp43[92],pp44[92],pp45[92],pp46[92],pp47[92],pp48[92],pp49[92],pp50[92],pp51[92],pp52[92],pp53[92],pp54[92],pp55[92],pp56[92],pp57[92],pp58[92],pp59[92],pp60[92],pp61[92],pp62[92],pp63[92],pp64[92],pp65[92],pp66[92],pp67[92],pp68[92],pp69[92],pp70[92],pp71[92],pp71[93],pp71[94],pp71[95],pp71[96],pp71[97],pp71[98],pp71[99],pp9[162],pp8[164],pp7[166],pp6[168],pp5[170],pp4[172],pp3[174],pp2[176],pp1[178],pp0[180],s146[100],s146[101],s146[102],s146[103],s146[104],s146[105],s146[106],s146[107],s146[108],s146[109],s146[110],s146[111],s146[112],s146[113],s146[114],s146[115],s146[116],s146[117],s146[118],s147[118],s148[118],s149[118],s150[118],s151[118],s152[118],s153[118],s154[118],pp0[208],pp1[208],pp2[208],pp3[208],pp4[208],pp5[208],pp6[208],pp7[208],pp8[208],pp9[208],pp209[9],pp211[8],pp213[7],pp215[6],pp217[5],pp219[4],pp221[3],pp223[2],pp225[1],pp227[0],s1[100],s2[100],s3[100],s4[100],s5[100],s6[100],s7[100],s8[100],s9[100],s8[102],s7[104],s6[106],s5[108],s4[110],s3[112],s2[114],s1[116],s108[10],s108[11],s108[12],s108[13],s108[14],s108[15],s108[16],s108[17],s108[18],s108[19],s108[20],s108[21],s106[24],s104[27],s102[30],s100[33],s33[101],s32[103],s31[105],s30[107],s29[109],s28[111],s27[113],s26[115],s25[117],s24[119],s23[121],s22[123],s21[125],s20[127],s19[129],s18[131],s17[133],s16[135],s15[137],s14[139],s13[141],s12[143],s11[145],s10[147],s154[196],s153[198],s152[200],s151[202],s150[204],s149[206],s148[208],s147[210],s146[212],s145[214],s144[216],s143[218],s142[220],s141[222],s140[224],s139[226],s138[228],s137[230],s136[232],s135[234],s134[236],s133[238],s132[240],s131[242],s130[244],s129[246],pp255[56],pp254[58],pp253[60],pp252[62],pp251[64],pp250[66],pp249[68],pp248[70],pp247[72],pp246[74],pp245[76],pp244[78],pp243[80],pp242[82],pp241[84],pp240[86],pp239[88],pp238[90],pp237[92],pp236[94],pp235[96],pp234[98],pp99[234],pp97[237],pp95[240],pp93[243],pp91[246],pp89[249],pp87[252],pp85[255],pp239[102],pp237[105],pp235[108],pp233[111],pp231[114],pp229[117],pp227[120],pp225[123],pp223[126],pp221[129],pp219[132],pp217[135],pp215[138],pp213[141],pp211[144],pp210[146],pp209[148],pp208[150],pp207[152],pp206[154],pp205[156],pp204[158],pp203[160],pp202[162],pp201[164],pp200[166],pp199[168],pp198[170],pp197[172],pp196[174],pp195[176],pp194[178],pp193[180],pp192[182],pp191[184],pp190[186],pp189[188],pp188[190],pp187[192],pp186[194],pp185[196],pp184[198],pp183[200],pp182[202],pp183[202],pp184[202],pp185[202],pp186[202],pp187[202],pp188[202],pp189[202],pp190[202],pp191[202],pp192[202],pp193[202],pp194[202],pp195[202],pp196[202],pp197[202],pp198[202],pp199[202],pp200[202],pp201[202],pp202[202],pp203[202],pp204[202],pp205[202],pp206[202],pp207[202],pp208[202],pp209[202],pp210[202],pp211[202],pp212[202],pp213[202],pp214[202],pp215[202],pp216[202],pp217[202],pp218[202],pp219[202]};
    CLA_332 KS_155(s155, c155, in155_1, in155_2);
    wire[329:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp64[27],pp64[28],pp64[29],pp64[30],pp64[31],pp64[32],pp64[33],pp64[34],pp64[35],pp63[37],pp62[39],pp61[41],pp60[43],pp59[45],pp58[47],pp57[49],pp56[51],pp55[53],pp54[55],pp53[57],pp52[59],pp51[61],pp50[63],pp49[65],pp48[67],pp47[69],pp46[71],pp45[73],pp44[75],pp43[77],pp42[79],pp41[81],pp40[83],pp39[85],pp38[87],pp37[89],pp36[91],pp37[91],pp38[91],pp39[91],pp40[91],pp41[91],pp42[91],pp43[91],pp44[91],pp45[91],pp46[91],pp47[91],pp48[91],pp49[91],pp50[91],pp51[91],pp52[91],pp53[91],pp54[91],pp55[91],pp56[91],pp57[91],pp58[91],pp59[91],pp60[91],pp61[91],pp62[91],pp63[91],pp64[91],pp65[91],pp66[91],pp67[91],pp68[91],pp69[91],pp70[91],pp71[91],pp72[91],pp72[92],pp72[93],pp72[94],pp72[95],pp72[96],pp72[97],pp72[98],pp72[99],pp9[163],pp8[165],pp7[167],pp6[169],pp5[171],pp4[173],pp3[175],pp2[177],pp1[179],pp0[181],s147[100],s147[101],s147[102],s147[103],s147[104],s147[105],s147[106],s147[107],s147[108],s147[109],s147[110],s147[111],s147[112],s147[113],s147[114],s147[115],s147[116],s147[117],s148[117],s149[117],s150[117],s151[117],s152[117],s153[117],s154[117],s155[117],s155[118],s155[119],s155[120],s155[121],s155[122],s155[123],s155[124],s155[125],s155[126],s155[127],s155[128],s155[129],s155[130],s155[131],s155[132],s155[133],s155[134],s155[135],s155[136],s155[137],s155[138],s155[139],s155[140],s155[141],s155[142],s155[143],s155[144],s155[145],s155[146],s155[147],s155[148],s155[149],s155[150],s155[151],s155[152],s155[153],s155[154],s155[155],s155[156],s155[157],s155[158],s155[159],s155[160],s155[161],s155[162],s155[163],s155[164],s155[165],s155[166],s155[167],s155[168],s155[169],s155[170],s155[171],s155[172],s155[173],s155[174],s155[175],s155[176],s155[177],s155[178],s155[179],s155[180],s155[181],s155[182],s155[183],s155[184],s155[185],s155[186],s155[187],s155[188],s155[189],s155[190],s155[191],s155[192],s155[193],s155[194],s155[195],s154[197],s153[199],s152[201],s151[203],s150[205],s149[207],s148[209],s147[211],s146[213],s145[215],s144[217],s143[219],s142[221],s141[223],s140[225],s139[227],s138[229],s137[231],s136[233],s135[235],s134[237],s133[239],s132[241],s131[243],s130[245],s129[247],pp255[57],pp254[59],pp253[61],pp252[63],pp251[65],pp250[67],pp249[69],pp248[71],pp247[73],pp246[75],pp245[77],pp244[79],pp243[81],pp242[83],pp241[85],pp240[87],pp239[89],pp238[91],pp237[93],pp236[95],pp235[97],pp234[99],pp98[236],pp96[239],pp94[242],pp92[245],pp90[248],pp88[251],pp86[254],pp240[101],pp238[104],pp236[107],pp234[110],pp232[113],pp230[116],pp228[119],pp226[122],pp224[125],pp222[128],pp220[131],pp218[134],pp216[137],pp214[140],pp212[143],pp211[145],pp210[147],pp209[149],pp208[151],pp207[153],pp206[155],pp205[157],pp204[159],pp203[161],pp202[163],pp201[165],pp200[167],pp199[169],pp198[171],pp197[173],pp196[175],pp195[177],pp194[179],pp193[181],pp192[183],pp191[185],pp190[187],pp189[189],pp188[191],pp187[193],pp186[195],pp185[197],pp184[199],pp183[201],pp184[201],pp185[201],pp186[201],pp187[201],pp188[201],pp189[201],pp190[201],pp191[201],pp192[201],pp193[201],pp194[201],pp195[201],pp196[201],pp197[201],pp198[201],pp199[201],pp200[201],pp201[201],pp202[201],pp203[201],pp204[201],pp205[201],pp206[201],pp207[201],pp208[201],pp209[201],pp210[201],pp211[201],pp212[201],pp213[201],pp214[201],pp215[201],pp216[201],pp217[201],pp218[201],pp219[201]};
    assign in156_2 = {pp65[26],pp65[27],pp65[28],pp65[29],pp65[30],pp65[31],pp65[32],pp65[33],pp65[34],pp64[36],pp63[38],pp62[40],pp61[42],pp60[44],pp59[46],pp58[48],pp57[50],pp56[52],pp55[54],pp54[56],pp53[58],pp52[60],pp51[62],pp50[64],pp49[66],pp48[68],pp47[70],pp46[72],pp45[74],pp44[76],pp43[78],pp42[80],pp41[82],pp40[84],pp39[86],pp38[88],pp37[90],pp38[90],pp39[90],pp40[90],pp41[90],pp42[90],pp43[90],pp44[90],pp45[90],pp46[90],pp47[90],pp48[90],pp49[90],pp50[90],pp51[90],pp52[90],pp53[90],pp54[90],pp55[90],pp56[90],pp57[90],pp58[90],pp59[90],pp60[90],pp61[90],pp62[90],pp63[90],pp64[90],pp65[90],pp66[90],pp67[90],pp68[90],pp69[90],pp70[90],pp71[90],pp72[90],pp73[90],pp73[91],pp73[92],pp73[93],pp73[94],pp73[95],pp73[96],pp73[97],pp73[98],pp73[99],pp9[164],pp8[166],pp7[168],pp6[170],pp5[172],pp4[174],pp3[176],pp2[178],pp1[180],pp0[182],s148[100],s148[101],s148[102],s148[103],s148[104],s148[105],s148[106],s148[107],s148[108],s148[109],s148[110],s148[111],s148[112],s148[113],s148[114],s148[115],s148[116],s149[116],s150[116],s151[116],s152[116],s153[116],s154[116],s155[116],pp0[207],pp1[207],pp2[207],pp3[207],pp4[207],pp5[207],pp6[207],pp7[207],pp8[207],pp9[207],pp208[9],pp210[8],pp212[7],pp214[6],pp216[5],pp218[4],pp220[3],pp222[2],pp224[1],pp226[0],s10[90],s10[91],s10[92],s10[93],s10[94],s10[95],s10[96],s10[97],s10[98],s10[99],s9[101],s8[103],s7[105],s6[107],s5[109],s4[111],s3[113],s2[115],s1[117],s109[10],s109[11],s109[12],s109[13],s109[14],s109[15],s109[16],s109[17],s109[18],s109[19],s109[20],s107[23],s105[26],s103[29],s101[32],s34[100],s33[102],s32[104],s31[106],s30[108],s29[110],s28[112],s27[114],s26[116],s25[118],s24[120],s23[122],s22[124],s21[126],s20[128],s19[130],s18[132],s17[134],s16[136],s15[138],s14[140],s13[142],s12[144],s11[146],s10[148],s155[196],s154[198],s153[200],s152[202],s151[204],s150[206],s149[208],s148[210],s147[212],s146[214],s145[216],s144[218],s143[220],s142[222],s141[224],s140[226],s139[228],s138[230],s137[232],s136[234],s135[236],s134[238],s133[240],s132[242],s131[244],s130[246],s129[248],pp255[58],pp254[60],pp253[62],pp252[64],pp251[66],pp250[68],pp249[70],pp248[72],pp247[74],pp246[76],pp245[78],pp244[80],pp243[82],pp242[84],pp241[86],pp240[88],pp239[90],pp238[92],pp237[94],pp236[96],pp235[98],pp99[235],pp97[238],pp95[241],pp93[244],pp91[247],pp89[250],pp87[253],pp241[100],pp239[103],pp237[106],pp235[109],pp233[112],pp231[115],pp229[118],pp227[121],pp225[124],pp223[127],pp221[130],pp219[133],pp217[136],pp215[139],pp213[142],pp212[144],pp211[146],pp210[148],pp209[150],pp208[152],pp207[154],pp206[156],pp205[158],pp204[160],pp203[162],pp202[164],pp201[166],pp200[168],pp199[170],pp198[172],pp197[174],pp196[176],pp195[178],pp194[180],pp193[182],pp192[184],pp191[186],pp190[188],pp189[190],pp188[192],pp187[194],pp186[196],pp185[198],pp184[200],pp185[200],pp186[200],pp187[200],pp188[200],pp189[200],pp190[200],pp191[200],pp192[200],pp193[200],pp194[200],pp195[200],pp196[200],pp197[200],pp198[200],pp199[200],pp200[200],pp201[200],pp202[200],pp203[200],pp204[200],pp205[200],pp206[200],pp207[200],pp208[200],pp209[200],pp210[200],pp211[200],pp212[200],pp213[200],pp214[200],pp215[200],pp216[200],pp217[200],pp218[200],pp219[200],pp220[200]};
    CLA_330 KS_156(s156, c156, in156_1, in156_2);
    wire[327:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp66[26],pp66[27],pp66[28],pp66[29],pp66[30],pp66[31],pp66[32],pp66[33],pp65[35],pp64[37],pp63[39],pp62[41],pp61[43],pp60[45],pp59[47],pp58[49],pp57[51],pp56[53],pp55[55],pp54[57],pp53[59],pp52[61],pp51[63],pp50[65],pp49[67],pp48[69],pp47[71],pp46[73],pp45[75],pp44[77],pp43[79],pp42[81],pp41[83],pp40[85],pp39[87],pp38[89],pp39[89],pp40[89],pp41[89],pp42[89],pp43[89],pp44[89],pp45[89],pp46[89],pp47[89],pp48[89],pp49[89],pp50[89],pp51[89],pp52[89],pp53[89],pp54[89],pp55[89],pp56[89],pp57[89],pp58[89],pp59[89],pp60[89],pp61[89],pp62[89],pp63[89],pp64[89],pp65[89],pp66[89],pp67[89],pp68[89],pp69[89],pp70[89],pp71[89],pp72[89],pp73[89],pp74[89],pp74[90],pp74[91],pp74[92],pp74[93],pp74[94],pp74[95],pp74[96],pp74[97],pp74[98],pp74[99],pp9[165],pp8[167],pp7[169],pp6[171],pp5[173],pp4[175],pp3[177],pp2[179],pp1[181],pp0[183],s149[100],s149[101],s149[102],s149[103],s149[104],s149[105],s149[106],s149[107],s149[108],s149[109],s149[110],s149[111],s149[112],s149[113],s149[114],s149[115],s150[115],s151[115],s152[115],s153[115],s154[115],s155[115],s156[115],s156[116],s156[117],s156[118],s156[119],s156[120],s156[121],s156[122],s156[123],s156[124],s156[125],s156[126],s156[127],s156[128],s156[129],s156[130],s156[131],s156[132],s156[133],s156[134],s156[135],s156[136],s156[137],s156[138],s156[139],s156[140],s156[141],s156[142],s156[143],s156[144],s156[145],s156[146],s156[147],s156[148],s156[149],s156[150],s156[151],s156[152],s156[153],s156[154],s156[155],s156[156],s156[157],s156[158],s156[159],s156[160],s156[161],s156[162],s156[163],s156[164],s156[165],s156[166],s156[167],s156[168],s156[169],s156[170],s156[171],s156[172],s156[173],s156[174],s156[175],s156[176],s156[177],s156[178],s156[179],s156[180],s156[181],s156[182],s156[183],s156[184],s156[185],s156[186],s156[187],s156[188],s156[189],s156[190],s156[191],s156[192],s156[193],s156[194],s156[195],s155[197],s154[199],s153[201],s152[203],s151[205],s150[207],s149[209],s148[211],s147[213],s146[215],s145[217],s144[219],s143[221],s142[223],s141[225],s140[227],s139[229],s138[231],s137[233],s136[235],s135[237],s134[239],s133[241],s132[243],s131[245],s130[247],s129[249],pp255[59],pp254[61],pp253[63],pp252[65],pp251[67],pp250[69],pp249[71],pp248[73],pp247[75],pp246[77],pp245[79],pp244[81],pp243[83],pp242[85],pp241[87],pp240[89],pp239[91],pp238[93],pp237[95],pp236[97],pp235[99],pp98[237],pp96[240],pp94[243],pp92[246],pp90[249],pp88[252],pp86[255],pp240[102],pp238[105],pp236[108],pp234[111],pp232[114],pp230[117],pp228[120],pp226[123],pp224[126],pp222[129],pp220[132],pp218[135],pp216[138],pp214[141],pp213[143],pp212[145],pp211[147],pp210[149],pp209[151],pp208[153],pp207[155],pp206[157],pp205[159],pp204[161],pp203[163],pp202[165],pp201[167],pp200[169],pp199[171],pp198[173],pp197[175],pp196[177],pp195[179],pp194[181],pp193[183],pp192[185],pp191[187],pp190[189],pp189[191],pp188[193],pp187[195],pp186[197],pp185[199],pp186[199],pp187[199],pp188[199],pp189[199],pp190[199],pp191[199],pp192[199],pp193[199],pp194[199],pp195[199],pp196[199],pp197[199],pp198[199],pp199[199],pp200[199],pp201[199],pp202[199],pp203[199],pp204[199],pp205[199],pp206[199],pp207[199],pp208[199],pp209[199],pp210[199],pp211[199],pp212[199],pp213[199],pp214[199],pp215[199],pp216[199],pp217[199],pp218[199],pp219[199],pp220[199]};
    assign in157_2 = {pp67[25],pp67[26],pp67[27],pp67[28],pp67[29],pp67[30],pp67[31],pp67[32],pp66[34],pp65[36],pp64[38],pp63[40],pp62[42],pp61[44],pp60[46],pp59[48],pp58[50],pp57[52],pp56[54],pp55[56],pp54[58],pp53[60],pp52[62],pp51[64],pp50[66],pp49[68],pp48[70],pp47[72],pp46[74],pp45[76],pp44[78],pp43[80],pp42[82],pp41[84],pp40[86],pp39[88],pp40[88],pp41[88],pp42[88],pp43[88],pp44[88],pp45[88],pp46[88],pp47[88],pp48[88],pp49[88],pp50[88],pp51[88],pp52[88],pp53[88],pp54[88],pp55[88],pp56[88],pp57[88],pp58[88],pp59[88],pp60[88],pp61[88],pp62[88],pp63[88],pp64[88],pp65[88],pp66[88],pp67[88],pp68[88],pp69[88],pp70[88],pp71[88],pp72[88],pp73[88],pp74[88],pp75[88],pp75[89],pp75[90],pp75[91],pp75[92],pp75[93],pp75[94],pp75[95],pp75[96],pp75[97],pp75[98],pp75[99],pp9[166],pp8[168],pp7[170],pp6[172],pp5[174],pp4[176],pp3[178],pp2[180],pp1[182],pp0[184],s150[100],s150[101],s150[102],s150[103],s150[104],s150[105],s150[106],s150[107],s150[108],s150[109],s150[110],s150[111],s150[112],s150[113],s150[114],s151[114],s152[114],s153[114],s154[114],s155[114],s156[114],pp0[206],pp1[206],pp2[206],pp3[206],pp4[206],pp5[206],pp6[206],pp7[206],pp8[206],pp9[206],pp207[9],pp209[8],pp211[7],pp213[6],pp215[5],pp217[4],pp219[3],pp221[2],pp223[1],pp225[0],s10[89],s11[89],s11[90],s11[91],s11[92],s11[93],s11[94],s11[95],s11[96],s11[97],s11[98],s11[99],s9[102],s8[104],s7[106],s6[108],s5[110],s4[112],s3[114],s2[116],s1[118],s110[10],s110[11],s110[12],s110[13],s110[14],s110[15],s110[16],s110[17],s110[18],s110[19],s108[22],s106[25],s104[28],s102[31],s100[34],s34[101],s33[103],s32[105],s31[107],s30[109],s29[111],s28[113],s27[115],s26[117],s25[119],s24[121],s23[123],s22[125],s21[127],s20[129],s19[131],s18[133],s17[135],s16[137],s15[139],s14[141],s13[143],s12[145],s11[147],s10[149],s156[196],s155[198],s154[200],s153[202],s152[204],s151[206],s150[208],s149[210],s148[212],s147[214],s146[216],s145[218],s144[220],s143[222],s142[224],s141[226],s140[228],s139[230],s138[232],s137[234],s136[236],s135[238],s134[240],s133[242],s132[244],s131[246],s130[248],s129[250],pp255[60],pp254[62],pp253[64],pp252[66],pp251[68],pp250[70],pp249[72],pp248[74],pp247[76],pp246[78],pp245[80],pp244[82],pp243[84],pp242[86],pp241[88],pp240[90],pp239[92],pp238[94],pp237[96],pp236[98],pp99[236],pp97[239],pp95[242],pp93[245],pp91[248],pp89[251],pp87[254],pp241[101],pp239[104],pp237[107],pp235[110],pp233[113],pp231[116],pp229[119],pp227[122],pp225[125],pp223[128],pp221[131],pp219[134],pp217[137],pp215[140],pp214[142],pp213[144],pp212[146],pp211[148],pp210[150],pp209[152],pp208[154],pp207[156],pp206[158],pp205[160],pp204[162],pp203[164],pp202[166],pp201[168],pp200[170],pp199[172],pp198[174],pp197[176],pp196[178],pp195[180],pp194[182],pp193[184],pp192[186],pp191[188],pp190[190],pp189[192],pp188[194],pp187[196],pp186[198],pp187[198],pp188[198],pp189[198],pp190[198],pp191[198],pp192[198],pp193[198],pp194[198],pp195[198],pp196[198],pp197[198],pp198[198],pp199[198],pp200[198],pp201[198],pp202[198],pp203[198],pp204[198],pp205[198],pp206[198],pp207[198],pp208[198],pp209[198],pp210[198],pp211[198],pp212[198],pp213[198],pp214[198],pp215[198],pp216[198],pp217[198],pp218[198],pp219[198],pp220[198],pp221[198]};
    CLA_328 KS_157(s157, c157, in157_1, in157_2);
    wire[325:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp68[25],pp68[26],pp68[27],pp68[28],pp68[29],pp68[30],pp68[31],pp67[33],pp66[35],pp65[37],pp64[39],pp63[41],pp62[43],pp61[45],pp60[47],pp59[49],pp58[51],pp57[53],pp56[55],pp55[57],pp54[59],pp53[61],pp52[63],pp51[65],pp50[67],pp49[69],pp48[71],pp47[73],pp46[75],pp45[77],pp44[79],pp43[81],pp42[83],pp41[85],pp40[87],pp41[87],pp42[87],pp43[87],pp44[87],pp45[87],pp46[87],pp47[87],pp48[87],pp49[87],pp50[87],pp51[87],pp52[87],pp53[87],pp54[87],pp55[87],pp56[87],pp57[87],pp58[87],pp59[87],pp60[87],pp61[87],pp62[87],pp63[87],pp64[87],pp65[87],pp66[87],pp67[87],pp68[87],pp69[87],pp70[87],pp71[87],pp72[87],pp73[87],pp74[87],pp75[87],pp76[87],pp76[88],pp76[89],pp76[90],pp76[91],pp76[92],pp76[93],pp76[94],pp76[95],pp76[96],pp76[97],pp76[98],pp76[99],pp9[167],pp8[169],pp7[171],pp6[173],pp5[175],pp4[177],pp3[179],pp2[181],pp1[183],pp0[185],s151[100],s151[101],s151[102],s151[103],s151[104],s151[105],s151[106],s151[107],s151[108],s151[109],s151[110],s151[111],s151[112],s151[113],s152[113],s153[113],s154[113],s155[113],s156[113],s157[113],s157[114],s157[115],s157[116],s157[117],s157[118],s157[119],s157[120],s157[121],s157[122],s157[123],s157[124],s157[125],s157[126],s157[127],s157[128],s157[129],s157[130],s157[131],s157[132],s157[133],s157[134],s157[135],s157[136],s157[137],s157[138],s157[139],s157[140],s157[141],s157[142],s157[143],s157[144],s157[145],s157[146],s157[147],s157[148],s157[149],s157[150],s157[151],s157[152],s157[153],s157[154],s157[155],s157[156],s157[157],s157[158],s157[159],s157[160],s157[161],s157[162],s157[163],s157[164],s157[165],s157[166],s157[167],s157[168],s157[169],s157[170],s157[171],s157[172],s157[173],s157[174],s157[175],s157[176],s157[177],s157[178],s157[179],s157[180],s157[181],s157[182],s157[183],s157[184],s157[185],s157[186],s157[187],s157[188],s157[189],s157[190],s157[191],s157[192],s157[193],s157[194],s157[195],s156[197],s155[199],s154[201],s153[203],s152[205],s151[207],s150[209],s149[211],s148[213],s147[215],s146[217],s145[219],s144[221],s143[223],s142[225],s141[227],s140[229],s139[231],s138[233],s137[235],s136[237],s135[239],s134[241],s133[243],s132[245],s131[247],s130[249],s129[251],pp255[61],pp254[63],pp253[65],pp252[67],pp251[69],pp250[71],pp249[73],pp248[75],pp247[77],pp246[79],pp245[81],pp244[83],pp243[85],pp242[87],pp241[89],pp240[91],pp239[93],pp238[95],pp237[97],pp236[99],pp98[238],pp96[241],pp94[244],pp92[247],pp90[250],pp88[253],pp242[100],pp240[103],pp238[106],pp236[109],pp234[112],pp232[115],pp230[118],pp228[121],pp226[124],pp224[127],pp222[130],pp220[133],pp218[136],pp216[139],pp215[141],pp214[143],pp213[145],pp212[147],pp211[149],pp210[151],pp209[153],pp208[155],pp207[157],pp206[159],pp205[161],pp204[163],pp203[165],pp202[167],pp201[169],pp200[171],pp199[173],pp198[175],pp197[177],pp196[179],pp195[181],pp194[183],pp193[185],pp192[187],pp191[189],pp190[191],pp189[193],pp188[195],pp187[197],pp188[197],pp189[197],pp190[197],pp191[197],pp192[197],pp193[197],pp194[197],pp195[197],pp196[197],pp197[197],pp198[197],pp199[197],pp200[197],pp201[197],pp202[197],pp203[197],pp204[197],pp205[197],pp206[197],pp207[197],pp208[197],pp209[197],pp210[197],pp211[197],pp212[197],pp213[197],pp214[197],pp215[197],pp216[197],pp217[197],pp218[197],pp219[197],pp220[197],pp221[197]};
    assign in158_2 = {pp69[24],pp69[25],pp69[26],pp69[27],pp69[28],pp69[29],pp69[30],pp68[32],pp67[34],pp66[36],pp65[38],pp64[40],pp63[42],pp62[44],pp61[46],pp60[48],pp59[50],pp58[52],pp57[54],pp56[56],pp55[58],pp54[60],pp53[62],pp52[64],pp51[66],pp50[68],pp49[70],pp48[72],pp47[74],pp46[76],pp45[78],pp44[80],pp43[82],pp42[84],pp41[86],pp42[86],pp43[86],pp44[86],pp45[86],pp46[86],pp47[86],pp48[86],pp49[86],pp50[86],pp51[86],pp52[86],pp53[86],pp54[86],pp55[86],pp56[86],pp57[86],pp58[86],pp59[86],pp60[86],pp61[86],pp62[86],pp63[86],pp64[86],pp65[86],pp66[86],pp67[86],pp68[86],pp69[86],pp70[86],pp71[86],pp72[86],pp73[86],pp74[86],pp75[86],pp76[86],pp77[86],pp77[87],pp77[88],pp77[89],pp77[90],pp77[91],pp77[92],pp77[93],pp77[94],pp77[95],pp77[96],pp77[97],pp77[98],pp77[99],pp9[168],pp8[170],pp7[172],pp6[174],pp5[176],pp4[178],pp3[180],pp2[182],pp1[184],pp0[186],s152[100],s152[101],s152[102],s152[103],s152[104],s152[105],s152[106],s152[107],s152[108],s152[109],s152[110],s152[111],s152[112],s153[112],s154[112],s155[112],s156[112],s157[112],pp0[205],pp1[205],pp2[205],pp3[205],pp4[205],pp5[205],pp6[205],pp7[205],pp8[205],pp9[205],pp206[9],pp208[8],pp210[7],pp212[6],pp214[5],pp216[4],pp218[3],pp220[2],pp222[1],pp224[0],s10[88],s11[88],s12[88],s12[89],s12[90],s12[91],s12[92],s12[93],s12[94],s12[95],s12[96],s12[97],s12[98],s12[99],s9[103],s8[105],s7[107],s6[109],s5[111],s4[113],s3[115],s2[117],s1[119],s111[10],s111[11],s111[12],s111[13],s111[14],s111[15],s111[16],s111[17],s111[18],s109[21],s107[24],s105[27],s103[30],s101[33],s35[100],s34[102],s33[104],s32[106],s31[108],s30[110],s29[112],s28[114],s27[116],s26[118],s25[120],s24[122],s23[124],s22[126],s21[128],s20[130],s19[132],s18[134],s17[136],s16[138],s15[140],s14[142],s13[144],s12[146],s11[148],s10[150],s157[196],s156[198],s155[200],s154[202],s153[204],s152[206],s151[208],s150[210],s149[212],s148[214],s147[216],s146[218],s145[220],s144[222],s143[224],s142[226],s141[228],s140[230],s139[232],s138[234],s137[236],s136[238],s135[240],s134[242],s133[244],s132[246],s131[248],s130[250],s129[252],pp255[62],pp254[64],pp253[66],pp252[68],pp251[70],pp250[72],pp249[74],pp248[76],pp247[78],pp246[80],pp245[82],pp244[84],pp243[86],pp242[88],pp241[90],pp240[92],pp239[94],pp238[96],pp237[98],pp99[237],pp97[240],pp95[243],pp93[246],pp91[249],pp89[252],pp87[255],pp241[102],pp239[105],pp237[108],pp235[111],pp233[114],pp231[117],pp229[120],pp227[123],pp225[126],pp223[129],pp221[132],pp219[135],pp217[138],pp216[140],pp215[142],pp214[144],pp213[146],pp212[148],pp211[150],pp210[152],pp209[154],pp208[156],pp207[158],pp206[160],pp205[162],pp204[164],pp203[166],pp202[168],pp201[170],pp200[172],pp199[174],pp198[176],pp197[178],pp196[180],pp195[182],pp194[184],pp193[186],pp192[188],pp191[190],pp190[192],pp189[194],pp188[196],pp189[196],pp190[196],pp191[196],pp192[196],pp193[196],pp194[196],pp195[196],pp196[196],pp197[196],pp198[196],pp199[196],pp200[196],pp201[196],pp202[196],pp203[196],pp204[196],pp205[196],pp206[196],pp207[196],pp208[196],pp209[196],pp210[196],pp211[196],pp212[196],pp213[196],pp214[196],pp215[196],pp216[196],pp217[196],pp218[196],pp219[196],pp220[196],pp221[196],pp222[196]};
    CLA_326 KS_158(s158, c158, in158_1, in158_2);
    wire[323:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp70[24],pp70[25],pp70[26],pp70[27],pp70[28],pp70[29],pp69[31],pp68[33],pp67[35],pp66[37],pp65[39],pp64[41],pp63[43],pp62[45],pp61[47],pp60[49],pp59[51],pp58[53],pp57[55],pp56[57],pp55[59],pp54[61],pp53[63],pp52[65],pp51[67],pp50[69],pp49[71],pp48[73],pp47[75],pp46[77],pp45[79],pp44[81],pp43[83],pp42[85],pp43[85],pp44[85],pp45[85],pp46[85],pp47[85],pp48[85],pp49[85],pp50[85],pp51[85],pp52[85],pp53[85],pp54[85],pp55[85],pp56[85],pp57[85],pp58[85],pp59[85],pp60[85],pp61[85],pp62[85],pp63[85],pp64[85],pp65[85],pp66[85],pp67[85],pp68[85],pp69[85],pp70[85],pp71[85],pp72[85],pp73[85],pp74[85],pp75[85],pp76[85],pp77[85],pp78[85],pp78[86],pp78[87],pp78[88],pp78[89],pp78[90],pp78[91],pp78[92],pp78[93],pp78[94],pp78[95],pp78[96],pp78[97],pp78[98],pp78[99],pp9[169],pp8[171],pp7[173],pp6[175],pp5[177],pp4[179],pp3[181],pp2[183],pp1[185],pp0[187],s153[100],s153[101],s153[102],s153[103],s153[104],s153[105],s153[106],s153[107],s153[108],s153[109],s153[110],s153[111],s154[111],s155[111],s156[111],s157[111],s158[111],s158[112],s158[113],s158[114],s158[115],s158[116],s158[117],s158[118],s158[119],s158[120],s158[121],s158[122],s158[123],s158[124],s158[125],s158[126],s158[127],s158[128],s158[129],s158[130],s158[131],s158[132],s158[133],s158[134],s158[135],s158[136],s158[137],s158[138],s158[139],s158[140],s158[141],s158[142],s158[143],s158[144],s158[145],s158[146],s158[147],s158[148],s158[149],s158[150],s158[151],s158[152],s158[153],s158[154],s158[155],s158[156],s158[157],s158[158],s158[159],s158[160],s158[161],s158[162],s158[163],s158[164],s158[165],s158[166],s158[167],s158[168],s158[169],s158[170],s158[171],s158[172],s158[173],s158[174],s158[175],s158[176],s158[177],s158[178],s158[179],s158[180],s158[181],s158[182],s158[183],s158[184],s158[185],s158[186],s158[187],s158[188],s158[189],s158[190],s158[191],s158[192],s158[193],s158[194],s158[195],s157[197],s156[199],s155[201],s154[203],s153[205],s152[207],s151[209],s150[211],s149[213],s148[215],s147[217],s146[219],s145[221],s144[223],s143[225],s142[227],s141[229],s140[231],s139[233],s138[235],s137[237],s136[239],s135[241],s134[243],s133[245],s132[247],s131[249],s130[251],s129[253],pp255[63],pp254[65],pp253[67],pp252[69],pp251[71],pp250[73],pp249[75],pp248[77],pp247[79],pp246[81],pp245[83],pp244[85],pp243[87],pp242[89],pp241[91],pp240[93],pp239[95],pp238[97],pp237[99],pp98[239],pp96[242],pp94[245],pp92[248],pp90[251],pp88[254],pp242[101],pp240[104],pp238[107],pp236[110],pp234[113],pp232[116],pp230[119],pp228[122],pp226[125],pp224[128],pp222[131],pp220[134],pp218[137],pp217[139],pp216[141],pp215[143],pp214[145],pp213[147],pp212[149],pp211[151],pp210[153],pp209[155],pp208[157],pp207[159],pp206[161],pp205[163],pp204[165],pp203[167],pp202[169],pp201[171],pp200[173],pp199[175],pp198[177],pp197[179],pp196[181],pp195[183],pp194[185],pp193[187],pp192[189],pp191[191],pp190[193],pp189[195],pp190[195],pp191[195],pp192[195],pp193[195],pp194[195],pp195[195],pp196[195],pp197[195],pp198[195],pp199[195],pp200[195],pp201[195],pp202[195],pp203[195],pp204[195],pp205[195],pp206[195],pp207[195],pp208[195],pp209[195],pp210[195],pp211[195],pp212[195],pp213[195],pp214[195],pp215[195],pp216[195],pp217[195],pp218[195],pp219[195],pp220[195],pp221[195],pp222[195]};
    assign in159_2 = {pp71[23],pp71[24],pp71[25],pp71[26],pp71[27],pp71[28],pp70[30],pp69[32],pp68[34],pp67[36],pp66[38],pp65[40],pp64[42],pp63[44],pp62[46],pp61[48],pp60[50],pp59[52],pp58[54],pp57[56],pp56[58],pp55[60],pp54[62],pp53[64],pp52[66],pp51[68],pp50[70],pp49[72],pp48[74],pp47[76],pp46[78],pp45[80],pp44[82],pp43[84],pp44[84],pp45[84],pp46[84],pp47[84],pp48[84],pp49[84],pp50[84],pp51[84],pp52[84],pp53[84],pp54[84],pp55[84],pp56[84],pp57[84],pp58[84],pp59[84],pp60[84],pp61[84],pp62[84],pp63[84],pp64[84],pp65[84],pp66[84],pp67[84],pp68[84],pp69[84],pp70[84],pp71[84],pp72[84],pp73[84],pp74[84],pp75[84],pp76[84],pp77[84],pp78[84],pp79[84],pp79[85],pp79[86],pp79[87],pp79[88],pp79[89],pp79[90],pp79[91],pp79[92],pp79[93],pp79[94],pp79[95],pp79[96],pp79[97],pp79[98],pp79[99],pp9[170],pp8[172],pp7[174],pp6[176],pp5[178],pp4[180],pp3[182],pp2[184],pp1[186],pp0[188],s154[100],s154[101],s154[102],s154[103],s154[104],s154[105],s154[106],s154[107],s154[108],s154[109],s154[110],s155[110],s156[110],s157[110],s158[110],pp0[204],pp1[204],pp2[204],pp3[204],pp4[204],pp5[204],pp6[204],pp7[204],pp8[204],pp9[204],pp205[9],pp207[8],pp209[7],pp211[6],pp213[5],pp215[4],pp217[3],pp219[2],pp221[1],pp223[0],s10[87],s11[87],s12[87],s13[87],s13[88],s13[89],s13[90],s13[91],s13[92],s13[93],s13[94],s13[95],s13[96],s13[97],s13[98],s13[99],s9[104],s8[106],s7[108],s6[110],s5[112],s4[114],s3[116],s2[118],s1[120],s112[10],s112[11],s112[12],s112[13],s112[14],s112[15],s112[16],s112[17],s110[20],s108[23],s106[26],s104[29],s102[32],s100[35],s35[101],s34[103],s33[105],s32[107],s31[109],s30[111],s29[113],s28[115],s27[117],s26[119],s25[121],s24[123],s23[125],s22[127],s21[129],s20[131],s19[133],s18[135],s17[137],s16[139],s15[141],s14[143],s13[145],s12[147],s11[149],s10[151],s158[196],s157[198],s156[200],s155[202],s154[204],s153[206],s152[208],s151[210],s150[212],s149[214],s148[216],s147[218],s146[220],s145[222],s144[224],s143[226],s142[228],s141[230],s140[232],s139[234],s138[236],s137[238],s136[240],s135[242],s134[244],s133[246],s132[248],s131[250],s130[252],s129[254],pp255[64],pp254[66],pp253[68],pp252[70],pp251[72],pp250[74],pp249[76],pp248[78],pp247[80],pp246[82],pp245[84],pp244[86],pp243[88],pp242[90],pp241[92],pp240[94],pp239[96],pp238[98],pp99[238],pp97[241],pp95[244],pp93[247],pp91[250],pp89[253],pp243[100],pp241[103],pp239[106],pp237[109],pp235[112],pp233[115],pp231[118],pp229[121],pp227[124],pp225[127],pp223[130],pp221[133],pp219[136],pp218[138],pp217[140],pp216[142],pp215[144],pp214[146],pp213[148],pp212[150],pp211[152],pp210[154],pp209[156],pp208[158],pp207[160],pp206[162],pp205[164],pp204[166],pp203[168],pp202[170],pp201[172],pp200[174],pp199[176],pp198[178],pp197[180],pp196[182],pp195[184],pp194[186],pp193[188],pp192[190],pp191[192],pp190[194],pp191[194],pp192[194],pp193[194],pp194[194],pp195[194],pp196[194],pp197[194],pp198[194],pp199[194],pp200[194],pp201[194],pp202[194],pp203[194],pp204[194],pp205[194],pp206[194],pp207[194],pp208[194],pp209[194],pp210[194],pp211[194],pp212[194],pp213[194],pp214[194],pp215[194],pp216[194],pp217[194],pp218[194],pp219[194],pp220[194],pp221[194],pp222[194],pp223[194]};
    CLA_324 KS_159(s159, c159, in159_1, in159_2);
    wire[321:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp72[23],pp72[24],pp72[25],pp72[26],pp72[27],pp71[29],pp70[31],pp69[33],pp68[35],pp67[37],pp66[39],pp65[41],pp64[43],pp63[45],pp62[47],pp61[49],pp60[51],pp59[53],pp58[55],pp57[57],pp56[59],pp55[61],pp54[63],pp53[65],pp52[67],pp51[69],pp50[71],pp49[73],pp48[75],pp47[77],pp46[79],pp45[81],pp44[83],pp45[83],pp46[83],pp47[83],pp48[83],pp49[83],pp50[83],pp51[83],pp52[83],pp53[83],pp54[83],pp55[83],pp56[83],pp57[83],pp58[83],pp59[83],pp60[83],pp61[83],pp62[83],pp63[83],pp64[83],pp65[83],pp66[83],pp67[83],pp68[83],pp69[83],pp70[83],pp71[83],pp72[83],pp73[83],pp74[83],pp75[83],pp76[83],pp77[83],pp78[83],pp79[83],pp80[83],pp80[84],pp80[85],pp80[86],pp80[87],pp80[88],pp80[89],pp80[90],pp80[91],pp80[92],pp80[93],pp80[94],pp80[95],pp80[96],pp80[97],pp80[98],pp80[99],pp9[171],pp8[173],pp7[175],pp6[177],pp5[179],pp4[181],pp3[183],pp2[185],pp1[187],pp0[189],s155[100],s155[101],s155[102],s155[103],s155[104],s155[105],s155[106],s155[107],s155[108],s155[109],s156[109],s157[109],s158[109],s159[109],s159[110],s159[111],s159[112],s159[113],s159[114],s159[115],s159[116],s159[117],s159[118],s159[119],s159[120],s159[121],s159[122],s159[123],s159[124],s159[125],s159[126],s159[127],s159[128],s159[129],s159[130],s159[131],s159[132],s159[133],s159[134],s159[135],s159[136],s159[137],s159[138],s159[139],s159[140],s159[141],s159[142],s159[143],s159[144],s159[145],s159[146],s159[147],s159[148],s159[149],s159[150],s159[151],s159[152],s159[153],s159[154],s159[155],s159[156],s159[157],s159[158],s159[159],s159[160],s159[161],s159[162],s159[163],s159[164],s159[165],s159[166],s159[167],s159[168],s159[169],s159[170],s159[171],s159[172],s159[173],s159[174],s159[175],s159[176],s159[177],s159[178],s159[179],s159[180],s159[181],s159[182],s159[183],s159[184],s159[185],s159[186],s159[187],s159[188],s159[189],s159[190],s159[191],s159[192],s159[193],s159[194],s159[195],s158[197],s157[199],s156[201],s155[203],s154[205],s153[207],s152[209],s151[211],s150[213],s149[215],s148[217],s147[219],s146[221],s145[223],s144[225],s143[227],s142[229],s141[231],s140[233],s139[235],s138[237],s137[239],s136[241],s135[243],s134[245],s133[247],s132[249],s131[251],s130[253],s129[255],pp255[65],pp254[67],pp253[69],pp252[71],pp251[73],pp250[75],pp249[77],pp248[79],pp247[81],pp246[83],pp245[85],pp244[87],pp243[89],pp242[91],pp241[93],pp240[95],pp239[97],pp238[99],pp98[240],pp96[243],pp94[246],pp92[249],pp90[252],pp88[255],pp242[102],pp240[105],pp238[108],pp236[111],pp234[114],pp232[117],pp230[120],pp228[123],pp226[126],pp224[129],pp222[132],pp220[135],pp219[137],pp218[139],pp217[141],pp216[143],pp215[145],pp214[147],pp213[149],pp212[151],pp211[153],pp210[155],pp209[157],pp208[159],pp207[161],pp206[163],pp205[165],pp204[167],pp203[169],pp202[171],pp201[173],pp200[175],pp199[177],pp198[179],pp197[181],pp196[183],pp195[185],pp194[187],pp193[189],pp192[191],pp191[193],pp192[193],pp193[193],pp194[193],pp195[193],pp196[193],pp197[193],pp198[193],pp199[193],pp200[193],pp201[193],pp202[193],pp203[193],pp204[193],pp205[193],pp206[193],pp207[193],pp208[193],pp209[193],pp210[193],pp211[193],pp212[193],pp213[193],pp214[193],pp215[193],pp216[193],pp217[193],pp218[193],pp219[193],pp220[193],pp221[193],pp222[193],pp223[193]};
    assign in160_2 = {pp73[22],pp73[23],pp73[24],pp73[25],pp73[26],pp72[28],pp71[30],pp70[32],pp69[34],pp68[36],pp67[38],pp66[40],pp65[42],pp64[44],pp63[46],pp62[48],pp61[50],pp60[52],pp59[54],pp58[56],pp57[58],pp56[60],pp55[62],pp54[64],pp53[66],pp52[68],pp51[70],pp50[72],pp49[74],pp48[76],pp47[78],pp46[80],pp45[82],pp46[82],pp47[82],pp48[82],pp49[82],pp50[82],pp51[82],pp52[82],pp53[82],pp54[82],pp55[82],pp56[82],pp57[82],pp58[82],pp59[82],pp60[82],pp61[82],pp62[82],pp63[82],pp64[82],pp65[82],pp66[82],pp67[82],pp68[82],pp69[82],pp70[82],pp71[82],pp72[82],pp73[82],pp74[82],pp75[82],pp76[82],pp77[82],pp78[82],pp79[82],pp80[82],pp81[82],pp81[83],pp81[84],pp81[85],pp81[86],pp81[87],pp81[88],pp81[89],pp81[90],pp81[91],pp81[92],pp81[93],pp81[94],pp81[95],pp81[96],pp81[97],pp81[98],pp81[99],pp9[172],pp8[174],pp7[176],pp6[178],pp5[180],pp4[182],pp3[184],pp2[186],pp1[188],pp0[190],s156[100],s156[101],s156[102],s156[103],s156[104],s156[105],s156[106],s156[107],s156[108],s157[108],s158[108],s159[108],pp0[203],pp1[203],pp2[203],pp3[203],pp4[203],pp5[203],pp6[203],pp7[203],pp8[203],pp9[203],pp204[9],pp206[8],pp208[7],pp210[6],pp212[5],pp214[4],pp216[3],pp218[2],pp220[1],pp222[0],s10[86],s11[86],s12[86],s13[86],s14[86],s14[87],s14[88],s14[89],s14[90],s14[91],s14[92],s14[93],s14[94],s14[95],s14[96],s14[97],s14[98],s14[99],s9[105],s8[107],s7[109],s6[111],s5[113],s4[115],s3[117],s2[119],s1[121],s113[10],s113[11],s113[12],s113[13],s113[14],s113[15],s113[16],s111[19],s109[22],s107[25],s105[28],s103[31],s101[34],s36[100],s35[102],s34[104],s33[106],s32[108],s31[110],s30[112],s29[114],s28[116],s27[118],s26[120],s25[122],s24[124],s23[126],s22[128],s21[130],s20[132],s19[134],s18[136],s17[138],s16[140],s15[142],s14[144],s13[146],s12[148],s11[150],s10[152],s159[196],s158[198],s157[200],s156[202],s155[204],s154[206],s153[208],s152[210],s151[212],s150[214],s149[216],s148[218],s147[220],s146[222],s145[224],s144[226],s143[228],s142[230],s141[232],s140[234],s139[236],s138[238],s137[240],s136[242],s135[244],s134[246],s133[248],s132[250],s131[252],s130[254],s129[256],pp255[66],pp254[68],pp253[70],pp252[72],pp251[74],pp250[76],pp249[78],pp248[80],pp247[82],pp246[84],pp245[86],pp244[88],pp243[90],pp242[92],pp241[94],pp240[96],pp239[98],pp99[239],pp97[242],pp95[245],pp93[248],pp91[251],pp89[254],pp243[101],pp241[104],pp239[107],pp237[110],pp235[113],pp233[116],pp231[119],pp229[122],pp227[125],pp225[128],pp223[131],pp221[134],pp220[136],pp219[138],pp218[140],pp217[142],pp216[144],pp215[146],pp214[148],pp213[150],pp212[152],pp211[154],pp210[156],pp209[158],pp208[160],pp207[162],pp206[164],pp205[166],pp204[168],pp203[170],pp202[172],pp201[174],pp200[176],pp199[178],pp198[180],pp197[182],pp196[184],pp195[186],pp194[188],pp193[190],pp192[192],pp193[192],pp194[192],pp195[192],pp196[192],pp197[192],pp198[192],pp199[192],pp200[192],pp201[192],pp202[192],pp203[192],pp204[192],pp205[192],pp206[192],pp207[192],pp208[192],pp209[192],pp210[192],pp211[192],pp212[192],pp213[192],pp214[192],pp215[192],pp216[192],pp217[192],pp218[192],pp219[192],pp220[192],pp221[192],pp222[192],pp223[192],pp224[192]};
    CLA_322 KS_160(s160, c160, in160_1, in160_2);
    wire[319:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp74[22],pp74[23],pp74[24],pp74[25],pp73[27],pp72[29],pp71[31],pp70[33],pp69[35],pp68[37],pp67[39],pp66[41],pp65[43],pp64[45],pp63[47],pp62[49],pp61[51],pp60[53],pp59[55],pp58[57],pp57[59],pp56[61],pp55[63],pp54[65],pp53[67],pp52[69],pp51[71],pp50[73],pp49[75],pp48[77],pp47[79],pp46[81],pp47[81],pp48[81],pp49[81],pp50[81],pp51[81],pp52[81],pp53[81],pp54[81],pp55[81],pp56[81],pp57[81],pp58[81],pp59[81],pp60[81],pp61[81],pp62[81],pp63[81],pp64[81],pp65[81],pp66[81],pp67[81],pp68[81],pp69[81],pp70[81],pp71[81],pp72[81],pp73[81],pp74[81],pp75[81],pp76[81],pp77[81],pp78[81],pp79[81],pp80[81],pp81[81],pp82[81],pp82[82],pp82[83],pp82[84],pp82[85],pp82[86],pp82[87],pp82[88],pp82[89],pp82[90],pp82[91],pp82[92],pp82[93],pp82[94],pp82[95],pp82[96],pp82[97],pp82[98],pp82[99],pp9[173],pp8[175],pp7[177],pp6[179],pp5[181],pp4[183],pp3[185],pp2[187],pp1[189],pp0[191],s157[100],s157[101],s157[102],s157[103],s157[104],s157[105],s157[106],s157[107],s158[107],s159[107],s160[107],s160[108],s160[109],s160[110],s160[111],s160[112],s160[113],s160[114],s160[115],s160[116],s160[117],s160[118],s160[119],s160[120],s160[121],s160[122],s160[123],s160[124],s160[125],s160[126],s160[127],s160[128],s160[129],s160[130],s160[131],s160[132],s160[133],s160[134],s160[135],s160[136],s160[137],s160[138],s160[139],s160[140],s160[141],s160[142],s160[143],s160[144],s160[145],s160[146],s160[147],s160[148],s160[149],s160[150],s160[151],s160[152],s160[153],s160[154],s160[155],s160[156],s160[157],s160[158],s160[159],s160[160],s160[161],s160[162],s160[163],s160[164],s160[165],s160[166],s160[167],s160[168],s160[169],s160[170],s160[171],s160[172],s160[173],s160[174],s160[175],s160[176],s160[177],s160[178],s160[179],s160[180],s160[181],s160[182],s160[183],s160[184],s160[185],s160[186],s160[187],s160[188],s160[189],s160[190],s160[191],s160[192],s160[193],s160[194],s160[195],s159[197],s158[199],s157[201],s156[203],s155[205],s154[207],s153[209],s152[211],s151[213],s150[215],s149[217],s148[219],s147[221],s146[223],s145[225],s144[227],s143[229],s142[231],s141[233],s140[235],s139[237],s138[239],s137[241],s136[243],s135[245],s134[247],s133[249],s132[251],s131[253],s130[255],s129[257],pp255[67],pp254[69],pp253[71],pp252[73],pp251[75],pp250[77],pp249[79],pp248[81],pp247[83],pp246[85],pp245[87],pp244[89],pp243[91],pp242[93],pp241[95],pp240[97],pp239[99],pp98[241],pp96[244],pp94[247],pp92[250],pp90[253],pp244[100],pp242[103],pp240[106],pp238[109],pp236[112],pp234[115],pp232[118],pp230[121],pp228[124],pp226[127],pp224[130],pp222[133],pp221[135],pp220[137],pp219[139],pp218[141],pp217[143],pp216[145],pp215[147],pp214[149],pp213[151],pp212[153],pp211[155],pp210[157],pp209[159],pp208[161],pp207[163],pp206[165],pp205[167],pp204[169],pp203[171],pp202[173],pp201[175],pp200[177],pp199[179],pp198[181],pp197[183],pp196[185],pp195[187],pp194[189],pp193[191],pp194[191],pp195[191],pp196[191],pp197[191],pp198[191],pp199[191],pp200[191],pp201[191],pp202[191],pp203[191],pp204[191],pp205[191],pp206[191],pp207[191],pp208[191],pp209[191],pp210[191],pp211[191],pp212[191],pp213[191],pp214[191],pp215[191],pp216[191],pp217[191],pp218[191],pp219[191],pp220[191],pp221[191],pp222[191],pp223[191],pp224[191]};
    assign in161_2 = {pp75[21],pp75[22],pp75[23],pp75[24],pp74[26],pp73[28],pp72[30],pp71[32],pp70[34],pp69[36],pp68[38],pp67[40],pp66[42],pp65[44],pp64[46],pp63[48],pp62[50],pp61[52],pp60[54],pp59[56],pp58[58],pp57[60],pp56[62],pp55[64],pp54[66],pp53[68],pp52[70],pp51[72],pp50[74],pp49[76],pp48[78],pp47[80],pp48[80],pp49[80],pp50[80],pp51[80],pp52[80],pp53[80],pp54[80],pp55[80],pp56[80],pp57[80],pp58[80],pp59[80],pp60[80],pp61[80],pp62[80],pp63[80],pp64[80],pp65[80],pp66[80],pp67[80],pp68[80],pp69[80],pp70[80],pp71[80],pp72[80],pp73[80],pp74[80],pp75[80],pp76[80],pp77[80],pp78[80],pp79[80],pp80[80],pp81[80],pp82[80],pp83[80],pp83[81],pp83[82],pp83[83],pp83[84],pp83[85],pp83[86],pp83[87],pp83[88],pp83[89],pp83[90],pp83[91],pp83[92],pp83[93],pp83[94],pp83[95],pp83[96],pp83[97],pp83[98],pp83[99],pp9[174],pp8[176],pp7[178],pp6[180],pp5[182],pp4[184],pp3[186],pp2[188],pp1[190],pp0[192],s158[100],s158[101],s158[102],s158[103],s158[104],s158[105],s158[106],s159[106],s160[106],pp0[202],pp1[202],pp2[202],pp3[202],pp4[202],pp5[202],pp6[202],pp7[202],pp8[202],pp9[202],pp203[9],pp205[8],pp207[7],pp209[6],pp211[5],pp213[4],pp215[3],pp217[2],pp219[1],pp221[0],s10[85],s11[85],s12[85],s13[85],s14[85],s15[85],s15[86],s15[87],s15[88],s15[89],s15[90],s15[91],s15[92],s15[93],s15[94],s15[95],s15[96],s15[97],s15[98],s15[99],s9[106],s8[108],s7[110],s6[112],s5[114],s4[116],s3[118],s2[120],s1[122],s114[10],s114[11],s114[12],s114[13],s114[14],s114[15],s112[18],s110[21],s108[24],s106[27],s104[30],s102[33],s100[36],s36[101],s35[103],s34[105],s33[107],s32[109],s31[111],s30[113],s29[115],s28[117],s27[119],s26[121],s25[123],s24[125],s23[127],s22[129],s21[131],s20[133],s19[135],s18[137],s17[139],s16[141],s15[143],s14[145],s13[147],s12[149],s11[151],s10[153],s160[196],s159[198],s158[200],s157[202],s156[204],s155[206],s154[208],s153[210],s152[212],s151[214],s150[216],s149[218],s148[220],s147[222],s146[224],s145[226],s144[228],s143[230],s142[232],s141[234],s140[236],s139[238],s138[240],s137[242],s136[244],s135[246],s134[248],s133[250],s132[252],s131[254],s130[256],s129[258],pp255[68],pp254[70],pp253[72],pp252[74],pp251[76],pp250[78],pp249[80],pp248[82],pp247[84],pp246[86],pp245[88],pp244[90],pp243[92],pp242[94],pp241[96],pp240[98],pp99[240],pp97[243],pp95[246],pp93[249],pp91[252],pp89[255],pp243[102],pp241[105],pp239[108],pp237[111],pp235[114],pp233[117],pp231[120],pp229[123],pp227[126],pp225[129],pp223[132],pp222[134],pp221[136],pp220[138],pp219[140],pp218[142],pp217[144],pp216[146],pp215[148],pp214[150],pp213[152],pp212[154],pp211[156],pp210[158],pp209[160],pp208[162],pp207[164],pp206[166],pp205[168],pp204[170],pp203[172],pp202[174],pp201[176],pp200[178],pp199[180],pp198[182],pp197[184],pp196[186],pp195[188],pp194[190],pp195[190],pp196[190],pp197[190],pp198[190],pp199[190],pp200[190],pp201[190],pp202[190],pp203[190],pp204[190],pp205[190],pp206[190],pp207[190],pp208[190],pp209[190],pp210[190],pp211[190],pp212[190],pp213[190],pp214[190],pp215[190],pp216[190],pp217[190],pp218[190],pp219[190],pp220[190],pp221[190],pp222[190],pp223[190],pp224[190],pp225[190]};
    CLA_320 KS_161(s161, c161, in161_1, in161_2);
    wire[317:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp76[21],pp76[22],pp76[23],pp75[25],pp74[27],pp73[29],pp72[31],pp71[33],pp70[35],pp69[37],pp68[39],pp67[41],pp66[43],pp65[45],pp64[47],pp63[49],pp62[51],pp61[53],pp60[55],pp59[57],pp58[59],pp57[61],pp56[63],pp55[65],pp54[67],pp53[69],pp52[71],pp51[73],pp50[75],pp49[77],pp48[79],pp49[79],pp50[79],pp51[79],pp52[79],pp53[79],pp54[79],pp55[79],pp56[79],pp57[79],pp58[79],pp59[79],pp60[79],pp61[79],pp62[79],pp63[79],pp64[79],pp65[79],pp66[79],pp67[79],pp68[79],pp69[79],pp70[79],pp71[79],pp72[79],pp73[79],pp74[79],pp75[79],pp76[79],pp77[79],pp78[79],pp79[79],pp80[79],pp81[79],pp82[79],pp83[79],pp84[79],pp84[80],pp84[81],pp84[82],pp84[83],pp84[84],pp84[85],pp84[86],pp84[87],pp84[88],pp84[89],pp84[90],pp84[91],pp84[92],pp84[93],pp84[94],pp84[95],pp84[96],pp84[97],pp84[98],pp84[99],pp9[175],pp8[177],pp7[179],pp6[181],pp5[183],pp4[185],pp3[187],pp2[189],pp1[191],pp0[193],s159[100],s159[101],s159[102],s159[103],s159[104],s159[105],s160[105],s161[105],s161[106],s161[107],s161[108],s161[109],s161[110],s161[111],s161[112],s161[113],s161[114],s161[115],s161[116],s161[117],s161[118],s161[119],s161[120],s161[121],s161[122],s161[123],s161[124],s161[125],s161[126],s161[127],s161[128],s161[129],s161[130],s161[131],s161[132],s161[133],s161[134],s161[135],s161[136],s161[137],s161[138],s161[139],s161[140],s161[141],s161[142],s161[143],s161[144],s161[145],s161[146],s161[147],s161[148],s161[149],s161[150],s161[151],s161[152],s161[153],s161[154],s161[155],s161[156],s161[157],s161[158],s161[159],s161[160],s161[161],s161[162],s161[163],s161[164],s161[165],s161[166],s161[167],s161[168],s161[169],s161[170],s161[171],s161[172],s161[173],s161[174],s161[175],s161[176],s161[177],s161[178],s161[179],s161[180],s161[181],s161[182],s161[183],s161[184],s161[185],s161[186],s161[187],s161[188],s161[189],s161[190],s161[191],s161[192],s161[193],s161[194],s161[195],s160[197],s159[199],s158[201],s157[203],s156[205],s155[207],s154[209],s153[211],s152[213],s151[215],s150[217],s149[219],s148[221],s147[223],s146[225],s145[227],s144[229],s143[231],s142[233],s141[235],s140[237],s139[239],s138[241],s137[243],s136[245],s135[247],s134[249],s133[251],s132[253],s131[255],s130[257],s129[259],pp255[69],pp254[71],pp253[73],pp252[75],pp251[77],pp250[79],pp249[81],pp248[83],pp247[85],pp246[87],pp245[89],pp244[91],pp243[93],pp242[95],pp241[97],pp240[99],pp98[242],pp96[245],pp94[248],pp92[251],pp90[254],pp244[101],pp242[104],pp240[107],pp238[110],pp236[113],pp234[116],pp232[119],pp230[122],pp228[125],pp226[128],pp224[131],pp223[133],pp222[135],pp221[137],pp220[139],pp219[141],pp218[143],pp217[145],pp216[147],pp215[149],pp214[151],pp213[153],pp212[155],pp211[157],pp210[159],pp209[161],pp208[163],pp207[165],pp206[167],pp205[169],pp204[171],pp203[173],pp202[175],pp201[177],pp200[179],pp199[181],pp198[183],pp197[185],pp196[187],pp195[189],pp196[189],pp197[189],pp198[189],pp199[189],pp200[189],pp201[189],pp202[189],pp203[189],pp204[189],pp205[189],pp206[189],pp207[189],pp208[189],pp209[189],pp210[189],pp211[189],pp212[189],pp213[189],pp214[189],pp215[189],pp216[189],pp217[189],pp218[189],pp219[189],pp220[189],pp221[189],pp222[189],pp223[189],pp224[189],pp225[189]};
    assign in162_2 = {pp77[20],pp77[21],pp77[22],pp76[24],pp75[26],pp74[28],pp73[30],pp72[32],pp71[34],pp70[36],pp69[38],pp68[40],pp67[42],pp66[44],pp65[46],pp64[48],pp63[50],pp62[52],pp61[54],pp60[56],pp59[58],pp58[60],pp57[62],pp56[64],pp55[66],pp54[68],pp53[70],pp52[72],pp51[74],pp50[76],pp49[78],pp50[78],pp51[78],pp52[78],pp53[78],pp54[78],pp55[78],pp56[78],pp57[78],pp58[78],pp59[78],pp60[78],pp61[78],pp62[78],pp63[78],pp64[78],pp65[78],pp66[78],pp67[78],pp68[78],pp69[78],pp70[78],pp71[78],pp72[78],pp73[78],pp74[78],pp75[78],pp76[78],pp77[78],pp78[78],pp79[78],pp80[78],pp81[78],pp82[78],pp83[78],pp84[78],pp85[78],pp85[79],pp85[80],pp85[81],pp85[82],pp85[83],pp85[84],pp85[85],pp85[86],pp85[87],pp85[88],pp85[89],pp85[90],pp85[91],pp85[92],pp85[93],pp85[94],pp85[95],pp85[96],pp85[97],pp85[98],pp85[99],pp9[176],pp8[178],pp7[180],pp6[182],pp5[184],pp4[186],pp3[188],pp2[190],pp1[192],pp0[194],s160[100],s160[101],s160[102],s160[103],s160[104],s161[104],pp0[201],pp1[201],pp2[201],pp3[201],pp4[201],pp5[201],pp6[201],pp7[201],pp8[201],pp9[201],pp202[9],pp204[8],pp206[7],pp208[6],pp210[5],pp212[4],pp214[3],pp216[2],pp218[1],pp220[0],s10[84],s11[84],s12[84],s13[84],s14[84],s15[84],s16[84],s16[85],s16[86],s16[87],s16[88],s16[89],s16[90],s16[91],s16[92],s16[93],s16[94],s16[95],s16[96],s16[97],s16[98],s16[99],s9[107],s8[109],s7[111],s6[113],s5[115],s4[117],s3[119],s2[121],s1[123],s115[10],s115[11],s115[12],s115[13],s115[14],s113[17],s111[20],s109[23],s107[26],s105[29],s103[32],s101[35],s37[100],s36[102],s35[104],s34[106],s33[108],s32[110],s31[112],s30[114],s29[116],s28[118],s27[120],s26[122],s25[124],s24[126],s23[128],s22[130],s21[132],s20[134],s19[136],s18[138],s17[140],s16[142],s15[144],s14[146],s13[148],s12[150],s11[152],s10[154],s161[196],s160[198],s159[200],s158[202],s157[204],s156[206],s155[208],s154[210],s153[212],s152[214],s151[216],s150[218],s149[220],s148[222],s147[224],s146[226],s145[228],s144[230],s143[232],s142[234],s141[236],s140[238],s139[240],s138[242],s137[244],s136[246],s135[248],s134[250],s133[252],s132[254],s131[256],s130[258],s129[260],pp255[70],pp254[72],pp253[74],pp252[76],pp251[78],pp250[80],pp249[82],pp248[84],pp247[86],pp246[88],pp245[90],pp244[92],pp243[94],pp242[96],pp241[98],pp99[241],pp97[244],pp95[247],pp93[250],pp91[253],pp245[100],pp243[103],pp241[106],pp239[109],pp237[112],pp235[115],pp233[118],pp231[121],pp229[124],pp227[127],pp225[130],pp224[132],pp223[134],pp222[136],pp221[138],pp220[140],pp219[142],pp218[144],pp217[146],pp216[148],pp215[150],pp214[152],pp213[154],pp212[156],pp211[158],pp210[160],pp209[162],pp208[164],pp207[166],pp206[168],pp205[170],pp204[172],pp203[174],pp202[176],pp201[178],pp200[180],pp199[182],pp198[184],pp197[186],pp196[188],pp197[188],pp198[188],pp199[188],pp200[188],pp201[188],pp202[188],pp203[188],pp204[188],pp205[188],pp206[188],pp207[188],pp208[188],pp209[188],pp210[188],pp211[188],pp212[188],pp213[188],pp214[188],pp215[188],pp216[188],pp217[188],pp218[188],pp219[188],pp220[188],pp221[188],pp222[188],pp223[188],pp224[188],pp225[188],pp226[188]};
    CLA_318 KS_162(s162, c162, in162_1, in162_2);
    wire[315:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp78[20],pp78[21],pp77[23],pp76[25],pp75[27],pp74[29],pp73[31],pp72[33],pp71[35],pp70[37],pp69[39],pp68[41],pp67[43],pp66[45],pp65[47],pp64[49],pp63[51],pp62[53],pp61[55],pp60[57],pp59[59],pp58[61],pp57[63],pp56[65],pp55[67],pp54[69],pp53[71],pp52[73],pp51[75],pp50[77],pp51[77],pp52[77],pp53[77],pp54[77],pp55[77],pp56[77],pp57[77],pp58[77],pp59[77],pp60[77],pp61[77],pp62[77],pp63[77],pp64[77],pp65[77],pp66[77],pp67[77],pp68[77],pp69[77],pp70[77],pp71[77],pp72[77],pp73[77],pp74[77],pp75[77],pp76[77],pp77[77],pp78[77],pp79[77],pp80[77],pp81[77],pp82[77],pp83[77],pp84[77],pp85[77],pp86[77],pp86[78],pp86[79],pp86[80],pp86[81],pp86[82],pp86[83],pp86[84],pp86[85],pp86[86],pp86[87],pp86[88],pp86[89],pp86[90],pp86[91],pp86[92],pp86[93],pp86[94],pp86[95],pp86[96],pp86[97],pp86[98],pp86[99],pp9[177],pp8[179],pp7[181],pp6[183],pp5[185],pp4[187],pp3[189],pp2[191],pp1[193],pp0[195],s161[100],s161[101],s161[102],s161[103],s162[103],s162[104],s162[105],s162[106],s162[107],s162[108],s162[109],s162[110],s162[111],s162[112],s162[113],s162[114],s162[115],s162[116],s162[117],s162[118],s162[119],s162[120],s162[121],s162[122],s162[123],s162[124],s162[125],s162[126],s162[127],s162[128],s162[129],s162[130],s162[131],s162[132],s162[133],s162[134],s162[135],s162[136],s162[137],s162[138],s162[139],s162[140],s162[141],s162[142],s162[143],s162[144],s162[145],s162[146],s162[147],s162[148],s162[149],s162[150],s162[151],s162[152],s162[153],s162[154],s162[155],s162[156],s162[157],s162[158],s162[159],s162[160],s162[161],s162[162],s162[163],s162[164],s162[165],s162[166],s162[167],s162[168],s162[169],s162[170],s162[171],s162[172],s162[173],s162[174],s162[175],s162[176],s162[177],s162[178],s162[179],s162[180],s162[181],s162[182],s162[183],s162[184],s162[185],s162[186],s162[187],s162[188],s162[189],s162[190],s162[191],s162[192],s162[193],s162[194],s162[195],s161[197],s160[199],s159[201],s158[203],s157[205],s156[207],s155[209],s154[211],s153[213],s152[215],s151[217],s150[219],s149[221],s148[223],s147[225],s146[227],s145[229],s144[231],s143[233],s142[235],s141[237],s140[239],s139[241],s138[243],s137[245],s136[247],s135[249],s134[251],s133[253],s132[255],s131[257],s130[259],s129[261],pp255[71],pp254[73],pp253[75],pp252[77],pp251[79],pp250[81],pp249[83],pp248[85],pp247[87],pp246[89],pp245[91],pp244[93],pp243[95],pp242[97],pp241[99],pp98[243],pp96[246],pp94[249],pp92[252],pp90[255],pp244[102],pp242[105],pp240[108],pp238[111],pp236[114],pp234[117],pp232[120],pp230[123],pp228[126],pp226[129],pp225[131],pp224[133],pp223[135],pp222[137],pp221[139],pp220[141],pp219[143],pp218[145],pp217[147],pp216[149],pp215[151],pp214[153],pp213[155],pp212[157],pp211[159],pp210[161],pp209[163],pp208[165],pp207[167],pp206[169],pp205[171],pp204[173],pp203[175],pp202[177],pp201[179],pp200[181],pp199[183],pp198[185],pp197[187],pp198[187],pp199[187],pp200[187],pp201[187],pp202[187],pp203[187],pp204[187],pp205[187],pp206[187],pp207[187],pp208[187],pp209[187],pp210[187],pp211[187],pp212[187],pp213[187],pp214[187],pp215[187],pp216[187],pp217[187],pp218[187],pp219[187],pp220[187],pp221[187],pp222[187],pp223[187],pp224[187],pp225[187],pp226[187]};
    assign in163_2 = {pp79[19],pp79[20],pp78[22],pp77[24],pp76[26],pp75[28],pp74[30],pp73[32],pp72[34],pp71[36],pp70[38],pp69[40],pp68[42],pp67[44],pp66[46],pp65[48],pp64[50],pp63[52],pp62[54],pp61[56],pp60[58],pp59[60],pp58[62],pp57[64],pp56[66],pp55[68],pp54[70],pp53[72],pp52[74],pp51[76],pp52[76],pp53[76],pp54[76],pp55[76],pp56[76],pp57[76],pp58[76],pp59[76],pp60[76],pp61[76],pp62[76],pp63[76],pp64[76],pp65[76],pp66[76],pp67[76],pp68[76],pp69[76],pp70[76],pp71[76],pp72[76],pp73[76],pp74[76],pp75[76],pp76[76],pp77[76],pp78[76],pp79[76],pp80[76],pp81[76],pp82[76],pp83[76],pp84[76],pp85[76],pp86[76],pp87[76],pp87[77],pp87[78],pp87[79],pp87[80],pp87[81],pp87[82],pp87[83],pp87[84],pp87[85],pp87[86],pp87[87],pp87[88],pp87[89],pp87[90],pp87[91],pp87[92],pp87[93],pp87[94],pp87[95],pp87[96],pp87[97],pp87[98],pp87[99],pp9[178],pp8[180],pp7[182],pp6[184],pp5[186],pp4[188],pp3[190],pp2[192],pp1[194],pp0[196],s162[100],s162[101],s162[102],pp0[200],pp1[200],pp2[200],pp3[200],pp4[200],pp5[200],pp6[200],pp7[200],pp8[200],pp9[200],pp201[9],pp203[8],pp205[7],pp207[6],pp209[5],pp211[4],pp213[3],pp215[2],pp217[1],pp219[0],s10[83],s11[83],s12[83],s13[83],s14[83],s15[83],s16[83],s17[83],s17[84],s17[85],s17[86],s17[87],s17[88],s17[89],s17[90],s17[91],s17[92],s17[93],s17[94],s17[95],s17[96],s17[97],s17[98],s17[99],s9[108],s8[110],s7[112],s6[114],s5[116],s4[118],s3[120],s2[122],s1[124],s116[10],s116[11],s116[12],s116[13],s114[16],s112[19],s110[22],s108[25],s106[28],s104[31],s102[34],s100[37],s37[101],s36[103],s35[105],s34[107],s33[109],s32[111],s31[113],s30[115],s29[117],s28[119],s27[121],s26[123],s25[125],s24[127],s23[129],s22[131],s21[133],s20[135],s19[137],s18[139],s17[141],s16[143],s15[145],s14[147],s13[149],s12[151],s11[153],s10[155],s162[196],s161[198],s160[200],s159[202],s158[204],s157[206],s156[208],s155[210],s154[212],s153[214],s152[216],s151[218],s150[220],s149[222],s148[224],s147[226],s146[228],s145[230],s144[232],s143[234],s142[236],s141[238],s140[240],s139[242],s138[244],s137[246],s136[248],s135[250],s134[252],s133[254],s132[256],s131[258],s130[260],s129[262],pp255[72],pp254[74],pp253[76],pp252[78],pp251[80],pp250[82],pp249[84],pp248[86],pp247[88],pp246[90],pp245[92],pp244[94],pp243[96],pp242[98],pp99[242],pp97[245],pp95[248],pp93[251],pp91[254],pp245[101],pp243[104],pp241[107],pp239[110],pp237[113],pp235[116],pp233[119],pp231[122],pp229[125],pp227[128],pp226[130],pp225[132],pp224[134],pp223[136],pp222[138],pp221[140],pp220[142],pp219[144],pp218[146],pp217[148],pp216[150],pp215[152],pp214[154],pp213[156],pp212[158],pp211[160],pp210[162],pp209[164],pp208[166],pp207[168],pp206[170],pp205[172],pp204[174],pp203[176],pp202[178],pp201[180],pp200[182],pp199[184],pp198[186],pp199[186],pp200[186],pp201[186],pp202[186],pp203[186],pp204[186],pp205[186],pp206[186],pp207[186],pp208[186],pp209[186],pp210[186],pp211[186],pp212[186],pp213[186],pp214[186],pp215[186],pp216[186],pp217[186],pp218[186],pp219[186],pp220[186],pp221[186],pp222[186],pp223[186],pp224[186],pp225[186],pp226[186],pp227[186]};
    CLA_316 KS_163(s163, c163, in163_1, in163_2);
    wire[313:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp80[19],pp79[21],pp78[23],pp77[25],pp76[27],pp75[29],pp74[31],pp73[33],pp72[35],pp71[37],pp70[39],pp69[41],pp68[43],pp67[45],pp66[47],pp65[49],pp64[51],pp63[53],pp62[55],pp61[57],pp60[59],pp59[61],pp58[63],pp57[65],pp56[67],pp55[69],pp54[71],pp53[73],pp52[75],pp53[75],pp54[75],pp55[75],pp56[75],pp57[75],pp58[75],pp59[75],pp60[75],pp61[75],pp62[75],pp63[75],pp64[75],pp65[75],pp66[75],pp67[75],pp68[75],pp69[75],pp70[75],pp71[75],pp72[75],pp73[75],pp74[75],pp75[75],pp76[75],pp77[75],pp78[75],pp79[75],pp80[75],pp81[75],pp82[75],pp83[75],pp84[75],pp85[75],pp86[75],pp87[75],pp88[75],pp88[76],pp88[77],pp88[78],pp88[79],pp88[80],pp88[81],pp88[82],pp88[83],pp88[84],pp88[85],pp88[86],pp88[87],pp88[88],pp88[89],pp88[90],pp88[91],pp88[92],pp88[93],pp88[94],pp88[95],pp88[96],pp88[97],pp88[98],pp88[99],pp9[179],pp8[181],pp7[183],pp6[185],pp5[187],pp4[189],pp3[191],pp2[193],pp1[195],pp0[197],s163[100],s163[101],s163[102],s163[103],s163[104],s163[105],s163[106],s163[107],s163[108],s163[109],s163[110],s163[111],s163[112],s163[113],s163[114],s163[115],s163[116],s163[117],s163[118],s163[119],s163[120],s163[121],s163[122],s163[123],s163[124],s163[125],s163[126],s163[127],s163[128],s163[129],s163[130],s163[131],s163[132],s163[133],s163[134],s163[135],s163[136],s163[137],s163[138],s163[139],s163[140],s163[141],s163[142],s163[143],s163[144],s163[145],s163[146],s163[147],s163[148],s163[149],s163[150],s163[151],s163[152],s163[153],s163[154],s163[155],s163[156],s163[157],s163[158],s163[159],s163[160],s163[161],s163[162],s163[163],s163[164],s163[165],s163[166],s163[167],s163[168],s163[169],s163[170],s163[171],s163[172],s163[173],s163[174],s163[175],s163[176],s163[177],s163[178],s163[179],s163[180],s163[181],s163[182],s163[183],s163[184],s163[185],s163[186],s163[187],s163[188],s163[189],s163[190],s163[191],s163[192],s163[193],s163[194],s163[195],s162[197],s161[199],s160[201],s159[203],s158[205],s157[207],s156[209],s155[211],s154[213],s153[215],s152[217],s151[219],s150[221],s149[223],s148[225],s147[227],s146[229],s145[231],s144[233],s143[235],s142[237],s141[239],s140[241],s139[243],s138[245],s137[247],s136[249],s135[251],s134[253],s133[255],s132[257],s131[259],s130[261],s129[263],pp255[73],pp254[75],pp253[77],pp252[79],pp251[81],pp250[83],pp249[85],pp248[87],pp247[89],pp246[91],pp245[93],pp244[95],pp243[97],pp242[99],pp98[244],pp96[247],pp94[250],pp92[253],pp246[100],pp244[103],pp242[106],pp240[109],pp238[112],pp236[115],pp234[118],pp232[121],pp230[124],pp228[127],pp227[129],pp226[131],pp225[133],pp224[135],pp223[137],pp222[139],pp221[141],pp220[143],pp219[145],pp218[147],pp217[149],pp216[151],pp215[153],pp214[155],pp213[157],pp212[159],pp211[161],pp210[163],pp209[165],pp208[167],pp207[169],pp206[171],pp205[173],pp204[175],pp203[177],pp202[179],pp201[181],pp200[183],pp199[185],pp200[185],pp201[185],pp202[185],pp203[185],pp204[185],pp205[185],pp206[185],pp207[185],pp208[185],pp209[185],pp210[185],pp211[185],pp212[185],pp213[185],pp214[185],pp215[185],pp216[185],pp217[185],pp218[185],pp219[185],pp220[185],pp221[185],pp222[185],pp223[185],pp224[185],pp225[185],pp226[185],pp227[185]};
    assign in164_2 = {pp81[18],pp80[20],pp79[22],pp78[24],pp77[26],pp76[28],pp75[30],pp74[32],pp73[34],pp72[36],pp71[38],pp70[40],pp69[42],pp68[44],pp67[46],pp66[48],pp65[50],pp64[52],pp63[54],pp62[56],pp61[58],pp60[60],pp59[62],pp58[64],pp57[66],pp56[68],pp55[70],pp54[72],pp53[74],pp54[74],pp55[74],pp56[74],pp57[74],pp58[74],pp59[74],pp60[74],pp61[74],pp62[74],pp63[74],pp64[74],pp65[74],pp66[74],pp67[74],pp68[74],pp69[74],pp70[74],pp71[74],pp72[74],pp73[74],pp74[74],pp75[74],pp76[74],pp77[74],pp78[74],pp79[74],pp80[74],pp81[74],pp82[74],pp83[74],pp84[74],pp85[74],pp86[74],pp87[74],pp88[74],pp89[74],pp89[75],pp89[76],pp89[77],pp89[78],pp89[79],pp89[80],pp89[81],pp89[82],pp89[83],pp89[84],pp89[85],pp89[86],pp89[87],pp89[88],pp89[89],pp89[90],pp89[91],pp89[92],pp89[93],pp89[94],pp89[95],pp89[96],pp89[97],pp89[98],pp89[99],pp9[180],pp8[182],pp7[184],pp6[186],pp5[188],pp4[190],pp3[192],pp2[194],pp1[196],pp0[198],pp0[199],pp1[199],pp2[199],pp3[199],pp4[199],pp5[199],pp6[199],pp7[199],pp8[199],pp9[199],pp200[9],pp202[8],pp204[7],pp206[6],pp208[5],pp210[4],pp212[3],pp214[2],pp216[1],pp218[0],s10[82],s11[82],s12[82],s13[82],s14[82],s15[82],s16[82],s17[82],s18[82],s18[83],s18[84],s18[85],s18[86],s18[87],s18[88],s18[89],s18[90],s18[91],s18[92],s18[93],s18[94],s18[95],s18[96],s18[97],s18[98],s18[99],s9[109],s8[111],s7[113],s6[115],s5[117],s4[119],s3[121],s2[123],s1[125],s117[10],s117[11],s117[12],s115[15],s113[18],s111[21],s109[24],s107[27],s105[30],s103[33],s101[36],s38[100],s37[102],s36[104],s35[106],s34[108],s33[110],s32[112],s31[114],s30[116],s29[118],s28[120],s27[122],s26[124],s25[126],s24[128],s23[130],s22[132],s21[134],s20[136],s19[138],s18[140],s17[142],s16[144],s15[146],s14[148],s13[150],s12[152],s11[154],s10[156],s163[196],s162[198],s161[200],s160[202],s159[204],s158[206],s157[208],s156[210],s155[212],s154[214],s153[216],s152[218],s151[220],s150[222],s149[224],s148[226],s147[228],s146[230],s145[232],s144[234],s143[236],s142[238],s141[240],s140[242],s139[244],s138[246],s137[248],s136[250],s135[252],s134[254],s133[256],s132[258],s131[260],s130[262],s129[264],pp255[74],pp254[76],pp253[78],pp252[80],pp251[82],pp250[84],pp249[86],pp248[88],pp247[90],pp246[92],pp245[94],pp244[96],pp243[98],pp99[243],pp97[246],pp95[249],pp93[252],pp91[255],pp245[102],pp243[105],pp241[108],pp239[111],pp237[114],pp235[117],pp233[120],pp231[123],pp229[126],pp228[128],pp227[130],pp226[132],pp225[134],pp224[136],pp223[138],pp222[140],pp221[142],pp220[144],pp219[146],pp218[148],pp217[150],pp216[152],pp215[154],pp214[156],pp213[158],pp212[160],pp211[162],pp210[164],pp209[166],pp208[168],pp207[170],pp206[172],pp205[174],pp204[176],pp203[178],pp202[180],pp201[182],pp200[184],pp201[184],pp202[184],pp203[184],pp204[184],pp205[184],pp206[184],pp207[184],pp208[184],pp209[184],pp210[184],pp211[184],pp212[184],pp213[184],pp214[184],pp215[184],pp216[184],pp217[184],pp218[184],pp219[184],pp220[184],pp221[184],pp222[184],pp223[184],pp224[184],pp225[184],pp226[184],pp227[184],pp228[184]};
    CLA_314 KS_164(s164, c164, in164_1, in164_2);
    wire[311:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {pp81[19],pp80[21],pp79[23],pp78[25],pp77[27],pp76[29],pp75[31],pp74[33],pp73[35],pp72[37],pp71[39],pp70[41],pp69[43],pp68[45],pp67[47],pp66[49],pp65[51],pp64[53],pp63[55],pp62[57],pp61[59],pp60[61],pp59[63],pp58[65],pp57[67],pp56[69],pp55[71],pp54[73],pp55[73],pp56[73],pp57[73],pp58[73],pp59[73],pp60[73],pp61[73],pp62[73],pp63[73],pp64[73],pp65[73],pp66[73],pp67[73],pp68[73],pp69[73],pp70[73],pp71[73],pp72[73],pp73[73],pp74[73],pp75[73],pp76[73],pp77[73],pp78[73],pp79[73],pp80[73],pp81[73],pp82[73],pp83[73],pp84[73],pp85[73],pp86[73],pp87[73],pp88[73],pp89[73],pp90[73],pp90[74],pp90[75],pp90[76],pp90[77],pp90[78],pp90[79],pp90[80],pp90[81],pp90[82],pp90[83],pp90[84],pp90[85],pp90[86],pp90[87],pp90[88],pp90[89],pp90[90],pp90[91],pp90[92],pp90[93],pp90[94],pp90[95],pp90[96],pp90[97],pp90[98],pp90[99],pp9[181],pp8[183],pp7[185],pp6[187],pp5[189],pp4[191],pp3[193],pp2[195],pp1[197],s164[100],s164[101],s164[102],s164[103],s164[104],s164[105],s164[106],s164[107],s164[108],s164[109],s164[110],s164[111],s164[112],s164[113],s164[114],s164[115],s164[116],s164[117],s164[118],s164[119],s164[120],s164[121],s164[122],s164[123],s164[124],s164[125],s164[126],s164[127],s164[128],s164[129],s164[130],s164[131],s164[132],s164[133],s164[134],s164[135],s164[136],s164[137],s164[138],s164[139],s164[140],s164[141],s164[142],s164[143],s164[144],s164[145],s164[146],s164[147],s164[148],s164[149],s164[150],s164[151],s164[152],s164[153],s164[154],s164[155],s164[156],s164[157],s164[158],s164[159],s164[160],s164[161],s164[162],s164[163],s164[164],s164[165],s164[166],s164[167],s164[168],s164[169],s164[170],s164[171],s164[172],s164[173],s164[174],s164[175],s164[176],s164[177],s164[178],s164[179],s164[180],s164[181],s164[182],s164[183],s164[184],s164[185],s164[186],s164[187],s164[188],s164[189],s164[190],s164[191],s164[192],s164[193],s164[194],s164[195],s163[197],s162[199],s161[201],s160[203],s159[205],s158[207],s157[209],s156[211],s155[213],s154[215],s153[217],s152[219],s151[221],s150[223],s149[225],s148[227],s147[229],s146[231],s145[233],s144[235],s143[237],s142[239],s141[241],s140[243],s139[245],s138[247],s137[249],s136[251],s135[253],s134[255],s133[257],s132[259],s131[261],s130[263],s129[265],pp255[75],pp254[77],pp253[79],pp252[81],pp251[83],pp250[85],pp249[87],pp248[89],pp247[91],pp246[93],pp245[95],pp244[97],pp243[99],pp98[245],pp96[248],pp94[251],pp92[254],pp246[101],pp244[104],pp242[107],pp240[110],pp238[113],pp236[116],pp234[119],pp232[122],pp230[125],pp229[127],pp228[129],pp227[131],pp226[133],pp225[135],pp224[137],pp223[139],pp222[141],pp221[143],pp220[145],pp219[147],pp218[149],pp217[151],pp216[153],pp215[155],pp214[157],pp213[159],pp212[161],pp211[163],pp210[165],pp209[167],pp208[169],pp207[171],pp206[173],pp205[175],pp204[177],pp203[179],pp202[181],pp201[183],pp202[183],pp203[183],pp204[183],pp205[183],pp206[183],pp207[183],pp208[183],pp209[183],pp210[183],pp211[183],pp212[183],pp213[183],pp214[183],pp215[183],pp216[183],pp217[183],pp218[183],pp219[183],pp220[183],pp221[183],pp222[183],pp223[183],pp224[183],pp225[183],pp226[183],pp227[183],pp228[183]};
    assign in165_2 = {pp82[18],pp81[20],pp80[22],pp79[24],pp78[26],pp77[28],pp76[30],pp75[32],pp74[34],pp73[36],pp72[38],pp71[40],pp70[42],pp69[44],pp68[46],pp67[48],pp66[50],pp65[52],pp64[54],pp63[56],pp62[58],pp61[60],pp60[62],pp59[64],pp58[66],pp57[68],pp56[70],pp55[72],pp56[72],pp57[72],pp58[72],pp59[72],pp60[72],pp61[72],pp62[72],pp63[72],pp64[72],pp65[72],pp66[72],pp67[72],pp68[72],pp69[72],pp70[72],pp71[72],pp72[72],pp73[72],pp74[72],pp75[72],pp76[72],pp77[72],pp78[72],pp79[72],pp80[72],pp81[72],pp82[72],pp83[72],pp84[72],pp85[72],pp86[72],pp87[72],pp88[72],pp89[72],pp90[72],pp91[72],pp91[73],pp91[74],pp91[75],pp91[76],pp91[77],pp91[78],pp91[79],pp91[80],pp91[81],pp91[82],pp91[83],pp91[84],pp91[85],pp91[86],pp91[87],pp91[88],pp91[89],pp91[90],pp91[91],pp91[92],pp91[93],pp91[94],pp91[95],pp91[96],pp91[97],pp91[98],pp91[99],pp9[182],pp8[184],pp7[186],pp6[188],pp5[190],pp4[192],pp3[194],pp2[196],pp1[198],pp2[198],pp3[198],pp4[198],pp5[198],pp6[198],pp7[198],pp8[198],pp9[198],pp199[9],pp201[8],pp203[7],pp205[6],pp207[5],pp209[4],pp211[3],pp213[2],pp215[1],pp217[0],s10[81],s11[81],s12[81],s13[81],s14[81],s15[81],s16[81],s17[81],s18[81],s19[81],s19[82],s19[83],s19[84],s19[85],s19[86],s19[87],s19[88],s19[89],s19[90],s19[91],s19[92],s19[93],s19[94],s19[95],s19[96],s19[97],s19[98],s19[99],s9[110],s8[112],s7[114],s6[116],s5[118],s4[120],s3[122],s2[124],s1[126],s118[10],s118[11],s116[14],s114[17],s112[20],s110[23],s108[26],s106[29],s104[32],s102[35],s100[38],s38[101],s37[103],s36[105],s35[107],s34[109],s33[111],s32[113],s31[115],s30[117],s29[119],s28[121],s27[123],s26[125],s25[127],s24[129],s23[131],s22[133],s21[135],s20[137],s19[139],s18[141],s17[143],s16[145],s15[147],s14[149],s13[151],s12[153],s11[155],s10[157],s164[196],s163[198],s162[200],s161[202],s160[204],s159[206],s158[208],s157[210],s156[212],s155[214],s154[216],s153[218],s152[220],s151[222],s150[224],s149[226],s148[228],s147[230],s146[232],s145[234],s144[236],s143[238],s142[240],s141[242],s140[244],s139[246],s138[248],s137[250],s136[252],s135[254],s134[256],s133[258],s132[260],s131[262],s130[264],s129[266],pp255[76],pp254[78],pp253[80],pp252[82],pp251[84],pp250[86],pp249[88],pp248[90],pp247[92],pp246[94],pp245[96],pp244[98],pp99[244],pp97[247],pp95[250],pp93[253],pp247[100],pp245[103],pp243[106],pp241[109],pp239[112],pp237[115],pp235[118],pp233[121],pp231[124],pp230[126],pp229[128],pp228[130],pp227[132],pp226[134],pp225[136],pp224[138],pp223[140],pp222[142],pp221[144],pp220[146],pp219[148],pp218[150],pp217[152],pp216[154],pp215[156],pp214[158],pp213[160],pp212[162],pp211[164],pp210[166],pp209[168],pp208[170],pp207[172],pp206[174],pp205[176],pp204[178],pp203[180],pp202[182],pp203[182],pp204[182],pp205[182],pp206[182],pp207[182],pp208[182],pp209[182],pp210[182],pp211[182],pp212[182],pp213[182],pp214[182],pp215[182],pp216[182],pp217[182],pp218[182],pp219[182],pp220[182],pp221[182],pp222[182],pp223[182],pp224[182],pp225[182],pp226[182],pp227[182],pp228[182],pp229[182]};
    CLA_312 KS_165(s165, c165, in165_1, in165_2);
    wire[309:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {pp82[19],pp81[21],pp80[23],pp79[25],pp78[27],pp77[29],pp76[31],pp75[33],pp74[35],pp73[37],pp72[39],pp71[41],pp70[43],pp69[45],pp68[47],pp67[49],pp66[51],pp65[53],pp64[55],pp63[57],pp62[59],pp61[61],pp60[63],pp59[65],pp58[67],pp57[69],pp56[71],pp57[71],pp58[71],pp59[71],pp60[71],pp61[71],pp62[71],pp63[71],pp64[71],pp65[71],pp66[71],pp67[71],pp68[71],pp69[71],pp70[71],pp71[71],pp72[71],pp73[71],pp74[71],pp75[71],pp76[71],pp77[71],pp78[71],pp79[71],pp80[71],pp81[71],pp82[71],pp83[71],pp84[71],pp85[71],pp86[71],pp87[71],pp88[71],pp89[71],pp90[71],pp91[71],pp92[71],pp92[72],pp92[73],pp92[74],pp92[75],pp92[76],pp92[77],pp92[78],pp92[79],pp92[80],pp92[81],pp92[82],pp92[83],pp92[84],pp92[85],pp92[86],pp92[87],pp92[88],pp92[89],pp92[90],pp92[91],pp92[92],pp92[93],pp92[94],pp92[95],pp92[96],pp92[97],pp92[98],pp92[99],pp9[183],pp8[185],pp7[187],pp6[189],pp5[191],pp4[193],pp3[195],pp2[197],s165[100],s165[101],s165[102],s165[103],s165[104],s165[105],s165[106],s165[107],s165[108],s165[109],s165[110],s165[111],s165[112],s165[113],s165[114],s165[115],s165[116],s165[117],s165[118],s165[119],s165[120],s165[121],s165[122],s165[123],s165[124],s165[125],s165[126],s165[127],s165[128],s165[129],s165[130],s165[131],s165[132],s165[133],s165[134],s165[135],s165[136],s165[137],s165[138],s165[139],s165[140],s165[141],s165[142],s165[143],s165[144],s165[145],s165[146],s165[147],s165[148],s165[149],s165[150],s165[151],s165[152],s165[153],s165[154],s165[155],s165[156],s165[157],s165[158],s165[159],s165[160],s165[161],s165[162],s165[163],s165[164],s165[165],s165[166],s165[167],s165[168],s165[169],s165[170],s165[171],s165[172],s165[173],s165[174],s165[175],s165[176],s165[177],s165[178],s165[179],s165[180],s165[181],s165[182],s165[183],s165[184],s165[185],s165[186],s165[187],s165[188],s165[189],s165[190],s165[191],s165[192],s165[193],s165[194],s165[195],s164[197],s163[199],s162[201],s161[203],s160[205],s159[207],s158[209],s157[211],s156[213],s155[215],s154[217],s153[219],s152[221],s151[223],s150[225],s149[227],s148[229],s147[231],s146[233],s145[235],s144[237],s143[239],s142[241],s141[243],s140[245],s139[247],s138[249],s137[251],s136[253],s135[255],s134[257],s133[259],s132[261],s131[263],s130[265],s129[267],pp255[77],pp254[79],pp253[81],pp252[83],pp251[85],pp250[87],pp249[89],pp248[91],pp247[93],pp246[95],pp245[97],pp244[99],pp98[246],pp96[249],pp94[252],pp92[255],pp246[102],pp244[105],pp242[108],pp240[111],pp238[114],pp236[117],pp234[120],pp232[123],pp231[125],pp230[127],pp229[129],pp228[131],pp227[133],pp226[135],pp225[137],pp224[139],pp223[141],pp222[143],pp221[145],pp220[147],pp219[149],pp218[151],pp217[153],pp216[155],pp215[157],pp214[159],pp213[161],pp212[163],pp211[165],pp210[167],pp209[169],pp208[171],pp207[173],pp206[175],pp205[177],pp204[179],pp203[181],pp204[181],pp205[181],pp206[181],pp207[181],pp208[181],pp209[181],pp210[181],pp211[181],pp212[181],pp213[181],pp214[181],pp215[181],pp216[181],pp217[181],pp218[181],pp219[181],pp220[181],pp221[181],pp222[181],pp223[181],pp224[181],pp225[181],pp226[181],pp227[181],pp228[181],pp229[181]};
    assign in166_2 = {pp83[18],pp82[20],pp81[22],pp80[24],pp79[26],pp78[28],pp77[30],pp76[32],pp75[34],pp74[36],pp73[38],pp72[40],pp71[42],pp70[44],pp69[46],pp68[48],pp67[50],pp66[52],pp65[54],pp64[56],pp63[58],pp62[60],pp61[62],pp60[64],pp59[66],pp58[68],pp57[70],pp58[70],pp59[70],pp60[70],pp61[70],pp62[70],pp63[70],pp64[70],pp65[70],pp66[70],pp67[70],pp68[70],pp69[70],pp70[70],pp71[70],pp72[70],pp73[70],pp74[70],pp75[70],pp76[70],pp77[70],pp78[70],pp79[70],pp80[70],pp81[70],pp82[70],pp83[70],pp84[70],pp85[70],pp86[70],pp87[70],pp88[70],pp89[70],pp90[70],pp91[70],pp92[70],pp93[70],pp93[71],pp93[72],pp93[73],pp93[74],pp93[75],pp93[76],pp93[77],pp93[78],pp93[79],pp93[80],pp93[81],pp93[82],pp93[83],pp93[84],pp93[85],pp93[86],pp93[87],pp93[88],pp93[89],pp93[90],pp93[91],pp93[92],pp93[93],pp93[94],pp93[95],pp93[96],pp93[97],pp93[98],pp93[99],pp9[184],pp8[186],pp7[188],pp6[190],pp5[192],pp4[194],pp3[196],pp3[197],pp4[197],pp5[197],pp6[197],pp7[197],pp8[197],pp9[197],pp198[9],pp200[8],pp202[7],pp204[6],pp206[5],pp208[4],pp210[3],pp212[2],pp214[1],pp216[0],s10[80],s11[80],s12[80],s13[80],s14[80],s15[80],s16[80],s17[80],s18[80],s19[80],s20[80],s20[81],s20[82],s20[83],s20[84],s20[85],s20[86],s20[87],s20[88],s20[89],s20[90],s20[91],s20[92],s20[93],s20[94],s20[95],s20[96],s20[97],s20[98],s20[99],s9[111],s8[113],s7[115],s6[117],s5[119],s4[121],s3[123],s2[125],s1[127],s119[10],s117[13],s115[16],s113[19],s111[22],s109[25],s107[28],s105[31],s103[34],s101[37],s39[100],s38[102],s37[104],s36[106],s35[108],s34[110],s33[112],s32[114],s31[116],s30[118],s29[120],s28[122],s27[124],s26[126],s25[128],s24[130],s23[132],s22[134],s21[136],s20[138],s19[140],s18[142],s17[144],s16[146],s15[148],s14[150],s13[152],s12[154],s11[156],s10[158],s165[196],s164[198],s163[200],s162[202],s161[204],s160[206],s159[208],s158[210],s157[212],s156[214],s155[216],s154[218],s153[220],s152[222],s151[224],s150[226],s149[228],s148[230],s147[232],s146[234],s145[236],s144[238],s143[240],s142[242],s141[244],s140[246],s139[248],s138[250],s137[252],s136[254],s135[256],s134[258],s133[260],s132[262],s131[264],s130[266],s129[268],pp255[78],pp254[80],pp253[82],pp252[84],pp251[86],pp250[88],pp249[90],pp248[92],pp247[94],pp246[96],pp245[98],pp99[245],pp97[248],pp95[251],pp93[254],pp247[101],pp245[104],pp243[107],pp241[110],pp239[113],pp237[116],pp235[119],pp233[122],pp232[124],pp231[126],pp230[128],pp229[130],pp228[132],pp227[134],pp226[136],pp225[138],pp224[140],pp223[142],pp222[144],pp221[146],pp220[148],pp219[150],pp218[152],pp217[154],pp216[156],pp215[158],pp214[160],pp213[162],pp212[164],pp211[166],pp210[168],pp209[170],pp208[172],pp207[174],pp206[176],pp205[178],pp204[180],pp205[180],pp206[180],pp207[180],pp208[180],pp209[180],pp210[180],pp211[180],pp212[180],pp213[180],pp214[180],pp215[180],pp216[180],pp217[180],pp218[180],pp219[180],pp220[180],pp221[180],pp222[180],pp223[180],pp224[180],pp225[180],pp226[180],pp227[180],pp228[180],pp229[180],pp230[180]};
    CLA_310 KS_166(s166, c166, in166_1, in166_2);
    wire[307:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {pp83[19],pp82[21],pp81[23],pp80[25],pp79[27],pp78[29],pp77[31],pp76[33],pp75[35],pp74[37],pp73[39],pp72[41],pp71[43],pp70[45],pp69[47],pp68[49],pp67[51],pp66[53],pp65[55],pp64[57],pp63[59],pp62[61],pp61[63],pp60[65],pp59[67],pp58[69],pp59[69],pp60[69],pp61[69],pp62[69],pp63[69],pp64[69],pp65[69],pp66[69],pp67[69],pp68[69],pp69[69],pp70[69],pp71[69],pp72[69],pp73[69],pp74[69],pp75[69],pp76[69],pp77[69],pp78[69],pp79[69],pp80[69],pp81[69],pp82[69],pp83[69],pp84[69],pp85[69],pp86[69],pp87[69],pp88[69],pp89[69],pp90[69],pp91[69],pp92[69],pp93[69],pp94[69],pp94[70],pp94[71],pp94[72],pp94[73],pp94[74],pp94[75],pp94[76],pp94[77],pp94[78],pp94[79],pp94[80],pp94[81],pp94[82],pp94[83],pp94[84],pp94[85],pp94[86],pp94[87],pp94[88],pp94[89],pp94[90],pp94[91],pp94[92],pp94[93],pp94[94],pp94[95],pp94[96],pp94[97],pp94[98],pp94[99],pp9[185],pp8[187],pp7[189],pp6[191],pp5[193],pp4[195],pp4[196],s166[100],s166[101],s166[102],s166[103],s166[104],s166[105],s166[106],s166[107],s166[108],s166[109],s166[110],s166[111],s166[112],s166[113],s166[114],s166[115],s166[116],s166[117],s166[118],s166[119],s166[120],s166[121],s166[122],s166[123],s166[124],s166[125],s166[126],s166[127],s166[128],s166[129],s166[130],s166[131],s166[132],s166[133],s166[134],s166[135],s166[136],s166[137],s166[138],s166[139],s166[140],s166[141],s166[142],s166[143],s166[144],s166[145],s166[146],s166[147],s166[148],s166[149],s166[150],s166[151],s166[152],s166[153],s166[154],s166[155],s166[156],s166[157],s166[158],s166[159],s166[160],s166[161],s166[162],s166[163],s166[164],s166[165],s166[166],s166[167],s166[168],s166[169],s166[170],s166[171],s166[172],s166[173],s166[174],s166[175],s166[176],s166[177],s166[178],s166[179],s166[180],s166[181],s166[182],s166[183],s166[184],s166[185],s166[186],s166[187],s166[188],s166[189],s166[190],s166[191],s166[192],s166[193],s166[194],s166[195],s165[197],s164[199],s163[201],s162[203],s161[205],s160[207],s159[209],s158[211],s157[213],s156[215],s155[217],s154[219],s153[221],s152[223],s151[225],s150[227],s149[229],s148[231],s147[233],s146[235],s145[237],s144[239],s143[241],s142[243],s141[245],s140[247],s139[249],s138[251],s137[253],s136[255],s135[257],s134[259],s133[261],s132[263],s131[265],s130[267],s129[269],pp255[79],pp254[81],pp253[83],pp252[85],pp251[87],pp250[89],pp249[91],pp248[93],pp247[95],pp246[97],pp245[99],pp98[247],pp96[250],pp94[253],pp248[100],pp246[103],pp244[106],pp242[109],pp240[112],pp238[115],pp236[118],pp234[121],pp233[123],pp232[125],pp231[127],pp230[129],pp229[131],pp228[133],pp227[135],pp226[137],pp225[139],pp224[141],pp223[143],pp222[145],pp221[147],pp220[149],pp219[151],pp218[153],pp217[155],pp216[157],pp215[159],pp214[161],pp213[163],pp212[165],pp211[167],pp210[169],pp209[171],pp208[173],pp207[175],pp206[177],pp205[179],pp206[179],pp207[179],pp208[179],pp209[179],pp210[179],pp211[179],pp212[179],pp213[179],pp214[179],pp215[179],pp216[179],pp217[179],pp218[179],pp219[179],pp220[179],pp221[179],pp222[179],pp223[179],pp224[179],pp225[179],pp226[179],pp227[179],pp228[179],pp229[179],pp230[179]};
    assign in167_2 = {pp84[18],pp83[20],pp82[22],pp81[24],pp80[26],pp79[28],pp78[30],pp77[32],pp76[34],pp75[36],pp74[38],pp73[40],pp72[42],pp71[44],pp70[46],pp69[48],pp68[50],pp67[52],pp66[54],pp65[56],pp64[58],pp63[60],pp62[62],pp61[64],pp60[66],pp59[68],pp60[68],pp61[68],pp62[68],pp63[68],pp64[68],pp65[68],pp66[68],pp67[68],pp68[68],pp69[68],pp70[68],pp71[68],pp72[68],pp73[68],pp74[68],pp75[68],pp76[68],pp77[68],pp78[68],pp79[68],pp80[68],pp81[68],pp82[68],pp83[68],pp84[68],pp85[68],pp86[68],pp87[68],pp88[68],pp89[68],pp90[68],pp91[68],pp92[68],pp93[68],pp94[68],pp95[68],pp95[69],pp95[70],pp95[71],pp95[72],pp95[73],pp95[74],pp95[75],pp95[76],pp95[77],pp95[78],pp95[79],pp95[80],pp95[81],pp95[82],pp95[83],pp95[84],pp95[85],pp95[86],pp95[87],pp95[88],pp95[89],pp95[90],pp95[91],pp95[92],pp95[93],pp95[94],pp95[95],pp95[96],pp95[97],pp95[98],pp95[99],pp9[186],pp8[188],pp7[190],pp6[192],pp5[194],pp5[195],pp5[196],pp6[196],pp7[196],pp8[196],pp9[196],pp197[9],pp199[8],pp201[7],pp203[6],pp205[5],pp207[4],pp209[3],pp211[2],pp213[1],pp215[0],s10[79],s11[79],s12[79],s13[79],s14[79],s15[79],s16[79],s17[79],s18[79],s19[79],s20[79],s21[79],s21[80],s21[81],s21[82],s21[83],s21[84],s21[85],s21[86],s21[87],s21[88],s21[89],s21[90],s21[91],s21[92],s21[93],s21[94],s21[95],s21[96],s21[97],s21[98],s21[99],s9[112],s8[114],s7[116],s6[118],s5[120],s4[122],s3[124],s2[126],s1[128],s118[12],s116[15],s114[18],s112[21],s110[24],s108[27],s106[30],s104[33],s102[36],s100[39],s39[101],s38[103],s37[105],s36[107],s35[109],s34[111],s33[113],s32[115],s31[117],s30[119],s29[121],s28[123],s27[125],s26[127],s25[129],s24[131],s23[133],s22[135],s21[137],s20[139],s19[141],s18[143],s17[145],s16[147],s15[149],s14[151],s13[153],s12[155],s11[157],s10[159],s166[196],s165[198],s164[200],s163[202],s162[204],s161[206],s160[208],s159[210],s158[212],s157[214],s156[216],s155[218],s154[220],s153[222],s152[224],s151[226],s150[228],s149[230],s148[232],s147[234],s146[236],s145[238],s144[240],s143[242],s142[244],s141[246],s140[248],s139[250],s138[252],s137[254],s136[256],s135[258],s134[260],s133[262],s132[264],s131[266],s130[268],s129[270],pp255[80],pp254[82],pp253[84],pp252[86],pp251[88],pp250[90],pp249[92],pp248[94],pp247[96],pp246[98],pp99[246],pp97[249],pp95[252],pp93[255],pp247[102],pp245[105],pp243[108],pp241[111],pp239[114],pp237[117],pp235[120],pp234[122],pp233[124],pp232[126],pp231[128],pp230[130],pp229[132],pp228[134],pp227[136],pp226[138],pp225[140],pp224[142],pp223[144],pp222[146],pp221[148],pp220[150],pp219[152],pp218[154],pp217[156],pp216[158],pp215[160],pp214[162],pp213[164],pp212[166],pp211[168],pp210[170],pp209[172],pp208[174],pp207[176],pp206[178],pp207[178],pp208[178],pp209[178],pp210[178],pp211[178],pp212[178],pp213[178],pp214[178],pp215[178],pp216[178],pp217[178],pp218[178],pp219[178],pp220[178],pp221[178],pp222[178],pp223[178],pp224[178],pp225[178],pp226[178],pp227[178],pp228[178],pp229[178],pp230[178],pp231[178]};
    CLA_308 KS_167(s167, c167, in167_1, in167_2);
    wire[305:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {pp84[19],pp83[21],pp82[23],pp81[25],pp80[27],pp79[29],pp78[31],pp77[33],pp76[35],pp75[37],pp74[39],pp73[41],pp72[43],pp71[45],pp70[47],pp69[49],pp68[51],pp67[53],pp66[55],pp65[57],pp64[59],pp63[61],pp62[63],pp61[65],pp60[67],pp61[67],pp62[67],pp63[67],pp64[67],pp65[67],pp66[67],pp67[67],pp68[67],pp69[67],pp70[67],pp71[67],pp72[67],pp73[67],pp74[67],pp75[67],pp76[67],pp77[67],pp78[67],pp79[67],pp80[67],pp81[67],pp82[67],pp83[67],pp84[67],pp85[67],pp86[67],pp87[67],pp88[67],pp89[67],pp90[67],pp91[67],pp92[67],pp93[67],pp94[67],pp95[67],pp96[67],pp96[68],pp96[69],pp96[70],pp96[71],pp96[72],pp96[73],pp96[74],pp96[75],pp96[76],pp96[77],pp96[78],pp96[79],pp96[80],pp96[81],pp96[82],pp96[83],pp96[84],pp96[85],pp96[86],pp96[87],pp96[88],pp96[89],pp96[90],pp96[91],pp96[92],pp96[93],pp96[94],pp96[95],pp96[96],pp96[97],pp96[98],pp96[99],pp9[187],pp8[189],pp7[191],pp6[193],pp6[194],pp6[195],s167[100],s167[101],s167[102],s167[103],s167[104],s167[105],s167[106],s167[107],s167[108],s167[109],s167[110],s167[111],s167[112],s167[113],s167[114],s167[115],s167[116],s167[117],s167[118],s167[119],s167[120],s167[121],s167[122],s167[123],s167[124],s167[125],s167[126],s167[127],s167[128],s167[129],s167[130],s167[131],s167[132],s167[133],s167[134],s167[135],s167[136],s167[137],s167[138],s167[139],s167[140],s167[141],s167[142],s167[143],s167[144],s167[145],s167[146],s167[147],s167[148],s167[149],s167[150],s167[151],s167[152],s167[153],s167[154],s167[155],s167[156],s167[157],s167[158],s167[159],s167[160],s167[161],s167[162],s167[163],s167[164],s167[165],s167[166],s167[167],s167[168],s167[169],s167[170],s167[171],s167[172],s167[173],s167[174],s167[175],s167[176],s167[177],s167[178],s167[179],s167[180],s167[181],s167[182],s167[183],s167[184],s167[185],s167[186],s167[187],s167[188],s167[189],s167[190],s167[191],s167[192],s167[193],s167[194],s167[195],s166[197],s165[199],s164[201],s163[203],s162[205],s161[207],s160[209],s159[211],s158[213],s157[215],s156[217],s155[219],s154[221],s153[223],s152[225],s151[227],s150[229],s149[231],s148[233],s147[235],s146[237],s145[239],s144[241],s143[243],s142[245],s141[247],s140[249],s139[251],s138[253],s137[255],s136[257],s135[259],s134[261],s133[263],s132[265],s131[267],s130[269],s129[271],pp255[81],pp254[83],pp253[85],pp252[87],pp251[89],pp250[91],pp249[93],pp248[95],pp247[97],pp246[99],pp98[248],pp96[251],pp94[254],pp248[101],pp246[104],pp244[107],pp242[110],pp240[113],pp238[116],pp236[119],pp235[121],pp234[123],pp233[125],pp232[127],pp231[129],pp230[131],pp229[133],pp228[135],pp227[137],pp226[139],pp225[141],pp224[143],pp223[145],pp222[147],pp221[149],pp220[151],pp219[153],pp218[155],pp217[157],pp216[159],pp215[161],pp214[163],pp213[165],pp212[167],pp211[169],pp210[171],pp209[173],pp208[175],pp207[177],pp208[177],pp209[177],pp210[177],pp211[177],pp212[177],pp213[177],pp214[177],pp215[177],pp216[177],pp217[177],pp218[177],pp219[177],pp220[177],pp221[177],pp222[177],pp223[177],pp224[177],pp225[177],pp226[177],pp227[177],pp228[177],pp229[177],pp230[177],pp231[177]};
    assign in168_2 = {pp85[18],pp84[20],pp83[22],pp82[24],pp81[26],pp80[28],pp79[30],pp78[32],pp77[34],pp76[36],pp75[38],pp74[40],pp73[42],pp72[44],pp71[46],pp70[48],pp69[50],pp68[52],pp67[54],pp66[56],pp65[58],pp64[60],pp63[62],pp62[64],pp61[66],pp62[66],pp63[66],pp64[66],pp65[66],pp66[66],pp67[66],pp68[66],pp69[66],pp70[66],pp71[66],pp72[66],pp73[66],pp74[66],pp75[66],pp76[66],pp77[66],pp78[66],pp79[66],pp80[66],pp81[66],pp82[66],pp83[66],pp84[66],pp85[66],pp86[66],pp87[66],pp88[66],pp89[66],pp90[66],pp91[66],pp92[66],pp93[66],pp94[66],pp95[66],pp96[66],pp97[66],pp97[67],pp97[68],pp97[69],pp97[70],pp97[71],pp97[72],pp97[73],pp97[74],pp97[75],pp97[76],pp97[77],pp97[78],pp97[79],pp97[80],pp97[81],pp97[82],pp97[83],pp97[84],pp97[85],pp97[86],pp97[87],pp97[88],pp97[89],pp97[90],pp97[91],pp97[92],pp97[93],pp97[94],pp97[95],pp97[96],pp97[97],pp97[98],pp97[99],pp9[188],pp8[190],pp7[192],pp7[193],pp7[194],pp7[195],pp8[195],pp9[195],pp196[9],pp198[8],pp200[7],pp202[6],pp204[5],pp206[4],pp208[3],pp210[2],pp212[1],pp214[0],s10[78],s11[78],s12[78],s13[78],s14[78],s15[78],s16[78],s17[78],s18[78],s19[78],s20[78],s21[78],s22[78],s22[79],s22[80],s22[81],s22[82],s22[83],s22[84],s22[85],s22[86],s22[87],s22[88],s22[89],s22[90],s22[91],s22[92],s22[93],s22[94],s22[95],s22[96],s22[97],s22[98],s22[99],s9[113],s8[115],s7[117],s6[119],s5[121],s4[123],s3[125],s2[127],s119[11],s117[14],s115[17],s113[20],s111[23],s109[26],s107[29],s105[32],s103[35],s101[38],s40[100],s39[102],s38[104],s37[106],s36[108],s35[110],s34[112],s33[114],s32[116],s31[118],s30[120],s29[122],s28[124],s27[126],s26[128],s25[130],s24[132],s23[134],s22[136],s21[138],s20[140],s19[142],s18[144],s17[146],s16[148],s15[150],s14[152],s13[154],s12[156],s11[158],s10[160],s167[196],s166[198],s165[200],s164[202],s163[204],s162[206],s161[208],s160[210],s159[212],s158[214],s157[216],s156[218],s155[220],s154[222],s153[224],s152[226],s151[228],s150[230],s149[232],s148[234],s147[236],s146[238],s145[240],s144[242],s143[244],s142[246],s141[248],s140[250],s139[252],s138[254],s137[256],s136[258],s135[260],s134[262],s133[264],s132[266],s131[268],s130[270],s129[272],pp255[82],pp254[84],pp253[86],pp252[88],pp251[90],pp250[92],pp249[94],pp248[96],pp247[98],pp99[247],pp97[250],pp95[253],pp249[100],pp247[103],pp245[106],pp243[109],pp241[112],pp239[115],pp237[118],pp236[120],pp235[122],pp234[124],pp233[126],pp232[128],pp231[130],pp230[132],pp229[134],pp228[136],pp227[138],pp226[140],pp225[142],pp224[144],pp223[146],pp222[148],pp221[150],pp220[152],pp219[154],pp218[156],pp217[158],pp216[160],pp215[162],pp214[164],pp213[166],pp212[168],pp211[170],pp210[172],pp209[174],pp208[176],pp209[176],pp210[176],pp211[176],pp212[176],pp213[176],pp214[176],pp215[176],pp216[176],pp217[176],pp218[176],pp219[176],pp220[176],pp221[176],pp222[176],pp223[176],pp224[176],pp225[176],pp226[176],pp227[176],pp228[176],pp229[176],pp230[176],pp231[176],pp232[176]};
    CLA_306 KS_168(s168, c168, in168_1, in168_2);
    wire[303:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {pp85[19],pp84[21],pp83[23],pp82[25],pp81[27],pp80[29],pp79[31],pp78[33],pp77[35],pp76[37],pp75[39],pp74[41],pp73[43],pp72[45],pp71[47],pp70[49],pp69[51],pp68[53],pp67[55],pp66[57],pp65[59],pp64[61],pp63[63],pp62[65],pp63[65],pp64[65],pp65[65],pp66[65],pp67[65],pp68[65],pp69[65],pp70[65],pp71[65],pp72[65],pp73[65],pp74[65],pp75[65],pp76[65],pp77[65],pp78[65],pp79[65],pp80[65],pp81[65],pp82[65],pp83[65],pp84[65],pp85[65],pp86[65],pp87[65],pp88[65],pp89[65],pp90[65],pp91[65],pp92[65],pp93[65],pp94[65],pp95[65],pp96[65],pp97[65],pp98[65],pp98[66],pp98[67],pp98[68],pp98[69],pp98[70],pp98[71],pp98[72],pp98[73],pp98[74],pp98[75],pp98[76],pp98[77],pp98[78],pp98[79],pp98[80],pp98[81],pp98[82],pp98[83],pp98[84],pp98[85],pp98[86],pp98[87],pp98[88],pp98[89],pp98[90],pp98[91],pp98[92],pp98[93],pp98[94],pp98[95],pp98[96],pp98[97],pp98[98],pp98[99],pp9[189],pp8[191],pp8[192],pp8[193],pp8[194],s168[100],s168[101],s168[102],s168[103],s168[104],s168[105],s168[106],s168[107],s168[108],s168[109],s168[110],s168[111],s168[112],s168[113],s168[114],s168[115],s168[116],s168[117],s168[118],s168[119],s168[120],s168[121],s168[122],s168[123],s168[124],s168[125],s168[126],s168[127],s168[128],s168[129],s168[130],s168[131],s168[132],s168[133],s168[134],s168[135],s168[136],s168[137],s168[138],s168[139],s168[140],s168[141],s168[142],s168[143],s168[144],s168[145],s168[146],s168[147],s168[148],s168[149],s168[150],s168[151],s168[152],s168[153],s168[154],s168[155],s168[156],s168[157],s168[158],s168[159],s168[160],s168[161],s168[162],s168[163],s168[164],s168[165],s168[166],s168[167],s168[168],s168[169],s168[170],s168[171],s168[172],s168[173],s168[174],s168[175],s168[176],s168[177],s168[178],s168[179],s168[180],s168[181],s168[182],s168[183],s168[184],s168[185],s168[186],s168[187],s168[188],s168[189],s168[190],s168[191],s168[192],s168[193],s168[194],s168[195],s167[197],s166[199],s165[201],s164[203],s163[205],s162[207],s161[209],s160[211],s159[213],s158[215],s157[217],s156[219],s155[221],s154[223],s153[225],s152[227],s151[229],s150[231],s149[233],s148[235],s147[237],s146[239],s145[241],s144[243],s143[245],s142[247],s141[249],s140[251],s139[253],s138[255],s137[257],s136[259],s135[261],s134[263],s133[265],s132[267],s131[269],s130[271],s129[273],pp255[83],pp254[85],pp253[87],pp252[89],pp251[91],pp250[93],pp249[95],pp248[97],pp247[99],pp98[249],pp96[252],pp94[255],pp248[102],pp246[105],pp244[108],pp242[111],pp240[114],pp238[117],pp237[119],pp236[121],pp235[123],pp234[125],pp233[127],pp232[129],pp231[131],pp230[133],pp229[135],pp228[137],pp227[139],pp226[141],pp225[143],pp224[145],pp223[147],pp222[149],pp221[151],pp220[153],pp219[155],pp218[157],pp217[159],pp216[161],pp215[163],pp214[165],pp213[167],pp212[169],pp211[171],pp210[173],pp209[175],pp210[175],pp211[175],pp212[175],pp213[175],pp214[175],pp215[175],pp216[175],pp217[175],pp218[175],pp219[175],pp220[175],pp221[175],pp222[175],pp223[175],pp224[175],pp225[175],pp226[175],pp227[175],pp228[175],pp229[175],pp230[175],pp231[175],pp232[175]};
    assign in169_2 = {pp86[18],pp85[20],pp84[22],pp83[24],pp82[26],pp81[28],pp80[30],pp79[32],pp78[34],pp77[36],pp76[38],pp75[40],pp74[42],pp73[44],pp72[46],pp71[48],pp70[50],pp69[52],pp68[54],pp67[56],pp66[58],pp65[60],pp64[62],pp63[64],pp64[64],pp65[64],pp66[64],pp67[64],pp68[64],pp69[64],pp70[64],pp71[64],pp72[64],pp73[64],pp74[64],pp75[64],pp76[64],pp77[64],pp78[64],pp79[64],pp80[64],pp81[64],pp82[64],pp83[64],pp84[64],pp85[64],pp86[64],pp87[64],pp88[64],pp89[64],pp90[64],pp91[64],pp92[64],pp93[64],pp94[64],pp95[64],pp96[64],pp97[64],pp98[64],pp99[64],pp99[65],pp99[66],pp99[67],pp99[68],pp99[69],pp99[70],pp99[71],pp99[72],pp99[73],pp99[74],pp99[75],pp99[76],pp99[77],pp99[78],pp99[79],pp99[80],pp99[81],pp99[82],pp99[83],pp99[84],pp99[85],pp99[86],pp99[87],pp99[88],pp99[89],pp99[90],pp99[91],pp99[92],pp99[93],pp99[94],pp99[95],pp99[96],pp99[97],pp99[98],pp99[99],pp9[190],pp9[191],pp9[192],pp9[193],pp9[194],pp195[9],pp197[8],pp199[7],pp201[6],pp203[5],pp205[4],pp207[3],pp209[2],pp211[1],pp213[0],s10[77],s11[77],s12[77],s13[77],s14[77],s15[77],s16[77],s17[77],s18[77],s19[77],s20[77],s21[77],s22[77],s23[77],s23[78],s23[79],s23[80],s23[81],s23[82],s23[83],s23[84],s23[85],s23[86],s23[87],s23[88],s23[89],s23[90],s23[91],s23[92],s23[93],s23[94],s23[95],s23[96],s23[97],s23[98],s23[99],s9[114],s8[116],s7[118],s6[120],s5[122],s4[124],s3[126],s120[10],s118[13],s116[16],s114[19],s112[22],s110[25],s108[28],s106[31],s104[34],s102[37],s100[40],s40[101],s39[103],s38[105],s37[107],s36[109],s35[111],s34[113],s33[115],s32[117],s31[119],s30[121],s29[123],s28[125],s27[127],s26[129],s25[131],s24[133],s23[135],s22[137],s21[139],s20[141],s19[143],s18[145],s17[147],s16[149],s15[151],s14[153],s13[155],s12[157],s11[159],s10[161],s168[196],s167[198],s166[200],s165[202],s164[204],s163[206],s162[208],s161[210],s160[212],s159[214],s158[216],s157[218],s156[220],s155[222],s154[224],s153[226],s152[228],s151[230],s150[232],s149[234],s148[236],s147[238],s146[240],s145[242],s144[244],s143[246],s142[248],s141[250],s140[252],s139[254],s138[256],s137[258],s136[260],s135[262],s134[264],s133[266],s132[268],s131[270],s130[272],s129[274],pp255[84],pp254[86],pp253[88],pp252[90],pp251[92],pp250[94],pp249[96],pp248[98],pp99[248],pp97[251],pp95[254],pp249[101],pp247[104],pp245[107],pp243[110],pp241[113],pp239[116],pp238[118],pp237[120],pp236[122],pp235[124],pp234[126],pp233[128],pp232[130],pp231[132],pp230[134],pp229[136],pp228[138],pp227[140],pp226[142],pp225[144],pp224[146],pp223[148],pp222[150],pp221[152],pp220[154],pp219[156],pp218[158],pp217[160],pp216[162],pp215[164],pp214[166],pp213[168],pp212[170],pp211[172],pp210[174],pp211[174],pp212[174],pp213[174],pp214[174],pp215[174],pp216[174],pp217[174],pp218[174],pp219[174],pp220[174],pp221[174],pp222[174],pp223[174],pp224[174],pp225[174],pp226[174],pp227[174],pp228[174],pp229[174],pp230[174],pp231[174],pp232[174],pp233[174]};
    CLA_304 KS_169(s169, c169, in169_1, in169_2);
    wire[301:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {pp86[19],pp85[21],pp84[23],pp83[25],pp82[27],pp81[29],pp80[31],pp79[33],pp78[35],pp77[37],pp76[39],pp75[41],pp74[43],pp73[45],pp72[47],pp71[49],pp70[51],pp69[53],pp68[55],pp67[57],pp66[59],pp65[61],pp64[63],pp65[63],pp66[63],pp67[63],pp68[63],pp69[63],pp70[63],pp71[63],pp72[63],pp73[63],pp74[63],pp75[63],pp76[63],pp77[63],pp78[63],pp79[63],pp80[63],pp81[63],pp82[63],pp83[63],pp84[63],pp85[63],pp86[63],pp87[63],pp88[63],pp89[63],pp90[63],pp91[63],pp92[63],pp93[63],pp94[63],pp95[63],pp96[63],pp97[63],pp98[63],pp99[63],pp154[9],pp155[9],pp156[9],pp157[9],pp158[9],pp159[9],pp160[9],pp161[9],pp162[9],pp163[9],pp164[9],pp165[9],pp166[9],pp167[9],pp168[9],pp169[9],pp170[9],pp171[9],pp172[9],pp173[9],pp174[9],pp175[9],pp176[9],pp177[9],pp178[9],pp179[9],pp180[9],pp181[9],pp182[9],pp183[9],pp184[9],pp185[9],pp186[9],pp187[9],pp188[9],pp189[9],pp190[9],pp191[9],pp192[9],pp193[9],pp194[9],s169[100],s169[101],s169[102],s169[103],s169[104],s169[105],s169[106],s169[107],s169[108],s169[109],s169[110],s169[111],s169[112],s169[113],s169[114],s169[115],s169[116],s169[117],s169[118],s169[119],s169[120],s169[121],s169[122],s169[123],s169[124],s169[125],s169[126],s169[127],s169[128],s169[129],s169[130],s169[131],s169[132],s169[133],s169[134],s169[135],s169[136],s169[137],s169[138],s169[139],s169[140],s169[141],s169[142],s169[143],s169[144],s169[145],s169[146],s169[147],s169[148],s169[149],s169[150],s169[151],s169[152],s169[153],s169[154],s169[155],s169[156],s169[157],s169[158],s169[159],s169[160],s169[161],s169[162],s169[163],s169[164],s169[165],s169[166],s169[167],s169[168],s169[169],s169[170],s169[171],s169[172],s169[173],s169[174],s169[175],s169[176],s169[177],s169[178],s169[179],s169[180],s169[181],s169[182],s169[183],s169[184],s169[185],s169[186],s169[187],s169[188],s169[189],s169[190],s169[191],s169[192],s169[193],s169[194],s169[195],s168[197],s167[199],s166[201],s165[203],s164[205],s163[207],s162[209],s161[211],s160[213],s159[215],s158[217],s157[219],s156[221],s155[223],s154[225],s153[227],s152[229],s151[231],s150[233],s149[235],s148[237],s147[239],s146[241],s145[243],s144[245],s143[247],s142[249],s141[251],s140[253],s139[255],s138[257],s137[259],s136[261],s135[263],s134[265],s133[267],s132[269],s131[271],s130[273],s129[275],pp255[85],pp254[87],pp253[89],pp252[91],pp251[93],pp250[95],pp249[97],pp248[99],pp98[250],pp96[253],pp250[100],pp248[103],pp246[106],pp244[109],pp242[112],pp240[115],pp239[117],pp238[119],pp237[121],pp236[123],pp235[125],pp234[127],pp233[129],pp232[131],pp231[133],pp230[135],pp229[137],pp228[139],pp227[141],pp226[143],pp225[145],pp224[147],pp223[149],pp222[151],pp221[153],pp220[155],pp219[157],pp218[159],pp217[161],pp216[163],pp215[165],pp214[167],pp213[169],pp212[171],pp211[173],pp212[173],pp213[173],pp214[173],pp215[173],pp216[173],pp217[173],pp218[173],pp219[173],pp220[173],pp221[173],pp222[173],pp223[173],pp224[173],pp225[173],pp226[173],pp227[173],pp228[173],pp229[173],pp230[173],pp231[173],pp232[173],pp233[173]};
    assign in170_2 = {pp87[18],pp86[20],pp85[22],pp84[24],pp83[26],pp82[28],pp81[30],pp80[32],pp79[34],pp78[36],pp77[38],pp76[40],pp75[42],pp74[44],pp73[46],pp72[48],pp71[50],pp70[52],pp69[54],pp68[56],pp67[58],pp66[60],pp65[62],pp66[62],pp67[62],pp68[62],pp69[62],pp70[62],pp71[62],pp72[62],pp73[62],pp74[62],pp75[62],pp76[62],pp77[62],pp78[62],pp79[62],pp80[62],pp81[62],pp82[62],pp83[62],pp84[62],pp85[62],pp86[62],pp87[62],pp88[62],pp89[62],pp90[62],pp91[62],pp92[62],pp93[62],pp94[62],pp95[62],pp96[62],pp97[62],pp98[62],pp99[62],pp153[9],pp155[8],pp156[8],pp157[8],pp158[8],pp159[8],pp160[8],pp161[8],pp162[8],pp163[8],pp164[8],pp165[8],pp166[8],pp167[8],pp168[8],pp169[8],pp170[8],pp171[8],pp172[8],pp173[8],pp174[8],pp175[8],pp176[8],pp177[8],pp178[8],pp179[8],pp180[8],pp181[8],pp182[8],pp183[8],pp184[8],pp185[8],pp186[8],pp187[8],pp188[8],pp189[8],pp190[8],pp191[8],pp192[8],pp193[8],pp194[8],pp195[8],pp196[8],pp198[7],pp200[6],pp202[5],pp204[4],pp206[3],pp208[2],pp210[1],pp212[0],s10[76],s11[76],s12[76],s13[76],s14[76],s15[76],s16[76],s17[76],s18[76],s19[76],s20[76],s21[76],s22[76],s23[76],s24[76],s24[77],s24[78],s24[79],s24[80],s24[81],s24[82],s24[83],s24[84],s24[85],s24[86],s24[87],s24[88],s24[89],s24[90],s24[91],s24[92],s24[93],s24[94],s24[95],s24[96],s24[97],s24[98],s24[99],s9[115],s8[117],s7[119],s6[121],s5[123],s4[125],s1[129],s119[12],s117[15],s115[18],s113[21],s111[24],s109[27],s107[30],s105[33],s103[36],s101[39],s41[100],s40[102],s39[104],s38[106],s37[108],s36[110],s35[112],s34[114],s33[116],s32[118],s31[120],s30[122],s29[124],s28[126],s27[128],s26[130],s25[132],s24[134],s23[136],s22[138],s21[140],s20[142],s19[144],s18[146],s17[148],s16[150],s15[152],s14[154],s13[156],s12[158],s11[160],s10[162],s169[196],s168[198],s167[200],s166[202],s165[204],s164[206],s163[208],s162[210],s161[212],s160[214],s159[216],s158[218],s157[220],s156[222],s155[224],s154[226],s153[228],s152[230],s151[232],s150[234],s149[236],s148[238],s147[240],s146[242],s145[244],s144[246],s143[248],s142[250],s141[252],s140[254],s139[256],s138[258],s137[260],s136[262],s135[264],s134[266],s133[268],s132[270],s131[272],s130[274],s129[276],pp255[86],pp254[88],pp253[90],pp252[92],pp251[94],pp250[96],pp249[98],pp99[249],pp97[252],pp95[255],pp249[102],pp247[105],pp245[108],pp243[111],pp241[114],pp240[116],pp239[118],pp238[120],pp237[122],pp236[124],pp235[126],pp234[128],pp233[130],pp232[132],pp231[134],pp230[136],pp229[138],pp228[140],pp227[142],pp226[144],pp225[146],pp224[148],pp223[150],pp222[152],pp221[154],pp220[156],pp219[158],pp218[160],pp217[162],pp216[164],pp215[166],pp214[168],pp213[170],pp212[172],pp213[172],pp214[172],pp215[172],pp216[172],pp217[172],pp218[172],pp219[172],pp220[172],pp221[172],pp222[172],pp223[172],pp224[172],pp225[172],pp226[172],pp227[172],pp228[172],pp229[172],pp230[172],pp231[172],pp232[172],pp233[172],pp234[172]};
    CLA_302 KS_170(s170, c170, in170_1, in170_2);
    wire[299:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {pp87[19],pp86[21],pp85[23],pp84[25],pp83[27],pp82[29],pp81[31],pp80[33],pp79[35],pp78[37],pp77[39],pp76[41],pp75[43],pp74[45],pp73[47],pp72[49],pp71[51],pp70[53],pp69[55],pp68[57],pp67[59],pp66[61],pp67[61],pp68[61],pp69[61],pp70[61],pp71[61],pp72[61],pp73[61],pp74[61],pp75[61],pp76[61],pp77[61],pp78[61],pp79[61],pp80[61],pp81[61],pp82[61],pp83[61],pp84[61],pp85[61],pp86[61],pp87[61],pp88[61],pp89[61],pp90[61],pp91[61],pp92[61],pp93[61],pp94[61],pp95[61],pp96[61],pp97[61],pp98[61],pp99[61],pp152[9],pp154[8],pp156[7],pp157[7],pp158[7],pp159[7],pp160[7],pp161[7],pp162[7],pp163[7],pp164[7],pp165[7],pp166[7],pp167[7],pp168[7],pp169[7],pp170[7],pp171[7],pp172[7],pp173[7],pp174[7],pp175[7],pp176[7],pp177[7],pp178[7],pp179[7],pp180[7],pp181[7],pp182[7],pp183[7],pp184[7],pp185[7],pp186[7],pp187[7],pp188[7],pp189[7],pp190[7],pp191[7],pp192[7],pp193[7],pp194[7],pp195[7],pp196[7],pp197[7],s170[100],s170[101],s170[102],s170[103],s170[104],s170[105],s170[106],s170[107],s170[108],s170[109],s170[110],s170[111],s170[112],s170[113],s170[114],s170[115],s170[116],s170[117],s170[118],s170[119],s170[120],s170[121],s170[122],s170[123],s170[124],s170[125],s170[126],s170[127],s170[128],s170[129],s170[130],s170[131],s170[132],s170[133],s170[134],s170[135],s170[136],s170[137],s170[138],s170[139],s170[140],s170[141],s170[142],s170[143],s170[144],s170[145],s170[146],s170[147],s170[148],s170[149],s170[150],s170[151],s170[152],s170[153],s170[154],s170[155],s170[156],s170[157],s170[158],s170[159],s170[160],s170[161],s170[162],s170[163],s170[164],s170[165],s170[166],s170[167],s170[168],s170[169],s170[170],s170[171],s170[172],s170[173],s170[174],s170[175],s170[176],s170[177],s170[178],s170[179],s170[180],s170[181],s170[182],s170[183],s170[184],s170[185],s170[186],s170[187],s170[188],s170[189],s170[190],s170[191],s170[192],s170[193],s170[194],s170[195],s169[197],s168[199],s167[201],s166[203],s165[205],s164[207],s163[209],s162[211],s161[213],s160[215],s159[217],s158[219],s157[221],s156[223],s155[225],s154[227],s153[229],s152[231],s151[233],s150[235],s149[237],s148[239],s147[241],s146[243],s145[245],s144[247],s143[249],s142[251],s141[253],s140[255],s139[257],s138[259],s137[261],s136[263],s135[265],s134[267],s133[269],s132[271],s131[273],s130[275],s129[277],pp255[87],pp254[89],pp253[91],pp252[93],pp251[95],pp250[97],pp249[99],pp98[251],pp96[254],pp250[101],pp248[104],pp246[107],pp244[110],pp242[113],pp241[115],pp240[117],pp239[119],pp238[121],pp237[123],pp236[125],pp235[127],pp234[129],pp233[131],pp232[133],pp231[135],pp230[137],pp229[139],pp228[141],pp227[143],pp226[145],pp225[147],pp224[149],pp223[151],pp222[153],pp221[155],pp220[157],pp219[159],pp218[161],pp217[163],pp216[165],pp215[167],pp214[169],pp213[171],pp214[171],pp215[171],pp216[171],pp217[171],pp218[171],pp219[171],pp220[171],pp221[171],pp222[171],pp223[171],pp224[171],pp225[171],pp226[171],pp227[171],pp228[171],pp229[171],pp230[171],pp231[171],pp232[171],pp233[171],pp234[171]};
    assign in171_2 = {pp88[18],pp87[20],pp86[22],pp85[24],pp84[26],pp83[28],pp82[30],pp81[32],pp80[34],pp79[36],pp78[38],pp77[40],pp76[42],pp75[44],pp74[46],pp73[48],pp72[50],pp71[52],pp70[54],pp69[56],pp68[58],pp67[60],pp68[60],pp69[60],pp70[60],pp71[60],pp72[60],pp73[60],pp74[60],pp75[60],pp76[60],pp77[60],pp78[60],pp79[60],pp80[60],pp81[60],pp82[60],pp83[60],pp84[60],pp85[60],pp86[60],pp87[60],pp88[60],pp89[60],pp90[60],pp91[60],pp92[60],pp93[60],pp94[60],pp95[60],pp96[60],pp97[60],pp98[60],pp99[60],pp151[9],pp153[8],pp155[7],pp157[6],pp158[6],pp159[6],pp160[6],pp161[6],pp162[6],pp163[6],pp164[6],pp165[6],pp166[6],pp167[6],pp168[6],pp169[6],pp170[6],pp171[6],pp172[6],pp173[6],pp174[6],pp175[6],pp176[6],pp177[6],pp178[6],pp179[6],pp180[6],pp181[6],pp182[6],pp183[6],pp184[6],pp185[6],pp186[6],pp187[6],pp188[6],pp189[6],pp190[6],pp191[6],pp192[6],pp193[6],pp194[6],pp195[6],pp196[6],pp197[6],pp198[6],pp199[6],pp201[5],pp203[4],pp205[3],pp207[2],pp209[1],pp211[0],s10[75],s11[75],s12[75],s13[75],s14[75],s15[75],s16[75],s17[75],s18[75],s19[75],s20[75],s21[75],s22[75],s23[75],s24[75],s25[75],s25[76],s25[77],s25[78],s25[79],s25[80],s25[81],s25[82],s25[83],s25[84],s25[85],s25[86],s25[87],s25[88],s25[89],s25[90],s25[91],s25[92],s25[93],s25[94],s25[95],s25[96],s25[97],s25[98],s25[99],s9[116],s8[118],s7[120],s6[122],s5[124],s2[128],s120[11],s118[14],s116[17],s114[20],s112[23],s110[26],s108[29],s106[32],s104[35],s102[38],s100[41],s41[101],s40[103],s39[105],s38[107],s37[109],s36[111],s35[113],s34[115],s33[117],s32[119],s31[121],s30[123],s29[125],s28[127],s27[129],s26[131],s25[133],s24[135],s23[137],s22[139],s21[141],s20[143],s19[145],s18[147],s17[149],s16[151],s15[153],s14[155],s13[157],s12[159],s11[161],s10[163],s170[196],s169[198],s168[200],s167[202],s166[204],s165[206],s164[208],s163[210],s162[212],s161[214],s160[216],s159[218],s158[220],s157[222],s156[224],s155[226],s154[228],s153[230],s152[232],s151[234],s150[236],s149[238],s148[240],s147[242],s146[244],s145[246],s144[248],s143[250],s142[252],s141[254],s140[256],s139[258],s138[260],s137[262],s136[264],s135[266],s134[268],s133[270],s132[272],s131[274],s130[276],s129[278],pp255[88],pp254[90],pp253[92],pp252[94],pp251[96],pp250[98],pp99[250],pp97[253],pp251[100],pp249[103],pp247[106],pp245[109],pp243[112],pp242[114],pp241[116],pp240[118],pp239[120],pp238[122],pp237[124],pp236[126],pp235[128],pp234[130],pp233[132],pp232[134],pp231[136],pp230[138],pp229[140],pp228[142],pp227[144],pp226[146],pp225[148],pp224[150],pp223[152],pp222[154],pp221[156],pp220[158],pp219[160],pp218[162],pp217[164],pp216[166],pp215[168],pp214[170],pp215[170],pp216[170],pp217[170],pp218[170],pp219[170],pp220[170],pp221[170],pp222[170],pp223[170],pp224[170],pp225[170],pp226[170],pp227[170],pp228[170],pp229[170],pp230[170],pp231[170],pp232[170],pp233[170],pp234[170],pp235[170]};
    CLA_300 KS_171(s171, c171, in171_1, in171_2);
    wire[297:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {pp88[19],pp87[21],pp86[23],pp85[25],pp84[27],pp83[29],pp82[31],pp81[33],pp80[35],pp79[37],pp78[39],pp77[41],pp76[43],pp75[45],pp74[47],pp73[49],pp72[51],pp71[53],pp70[55],pp69[57],pp68[59],pp69[59],pp70[59],pp71[59],pp72[59],pp73[59],pp74[59],pp75[59],pp76[59],pp77[59],pp78[59],pp79[59],pp80[59],pp81[59],pp82[59],pp83[59],pp84[59],pp85[59],pp86[59],pp87[59],pp88[59],pp89[59],pp90[59],pp91[59],pp92[59],pp93[59],pp94[59],pp95[59],pp96[59],pp97[59],pp98[59],pp99[59],pp150[9],pp152[8],pp154[7],pp156[6],pp158[5],pp159[5],pp160[5],pp161[5],pp162[5],pp163[5],pp164[5],pp165[5],pp166[5],pp167[5],pp168[5],pp169[5],pp170[5],pp171[5],pp172[5],pp173[5],pp174[5],pp175[5],pp176[5],pp177[5],pp178[5],pp179[5],pp180[5],pp181[5],pp182[5],pp183[5],pp184[5],pp185[5],pp186[5],pp187[5],pp188[5],pp189[5],pp190[5],pp191[5],pp192[5],pp193[5],pp194[5],pp195[5],pp196[5],pp197[5],pp198[5],pp199[5],pp200[5],s171[100],s171[101],s171[102],s171[103],s171[104],s171[105],s171[106],s171[107],s171[108],s171[109],s171[110],s171[111],s171[112],s171[113],s171[114],s171[115],s171[116],s171[117],s171[118],s171[119],s171[120],s171[121],s171[122],s171[123],s171[124],s171[125],s171[126],s171[127],s171[128],s171[129],s171[130],s171[131],s171[132],s171[133],s171[134],s171[135],s171[136],s171[137],s171[138],s171[139],s171[140],s171[141],s171[142],s171[143],s171[144],s171[145],s171[146],s171[147],s171[148],s171[149],s171[150],s171[151],s171[152],s171[153],s171[154],s171[155],s171[156],s171[157],s171[158],s171[159],s171[160],s171[161],s171[162],s171[163],s171[164],s171[165],s171[166],s171[167],s171[168],s171[169],s171[170],s171[171],s171[172],s171[173],s171[174],s171[175],s171[176],s171[177],s171[178],s171[179],s171[180],s171[181],s171[182],s171[183],s171[184],s171[185],s171[186],s171[187],s171[188],s171[189],s171[190],s171[191],s171[192],s171[193],s171[194],s171[195],s170[197],s169[199],s168[201],s167[203],s166[205],s165[207],s164[209],s163[211],s162[213],s161[215],s160[217],s159[219],s158[221],s157[223],s156[225],s155[227],s154[229],s153[231],s152[233],s151[235],s150[237],s149[239],s148[241],s147[243],s146[245],s145[247],s144[249],s143[251],s142[253],s141[255],s140[257],s139[259],s138[261],s137[263],s136[265],s135[267],s134[269],s133[271],s132[273],s131[275],s130[277],s129[279],pp255[89],pp254[91],pp253[93],pp252[95],pp251[97],pp250[99],pp98[252],pp96[255],pp250[102],pp248[105],pp246[108],pp244[111],pp243[113],pp242[115],pp241[117],pp240[119],pp239[121],pp238[123],pp237[125],pp236[127],pp235[129],pp234[131],pp233[133],pp232[135],pp231[137],pp230[139],pp229[141],pp228[143],pp227[145],pp226[147],pp225[149],pp224[151],pp223[153],pp222[155],pp221[157],pp220[159],pp219[161],pp218[163],pp217[165],pp216[167],pp215[169],pp216[169],pp217[169],pp218[169],pp219[169],pp220[169],pp221[169],pp222[169],pp223[169],pp224[169],pp225[169],pp226[169],pp227[169],pp228[169],pp229[169],pp230[169],pp231[169],pp232[169],pp233[169],pp234[169],pp235[169]};
    assign in172_2 = {pp89[18],pp88[20],pp87[22],pp86[24],pp85[26],pp84[28],pp83[30],pp82[32],pp81[34],pp80[36],pp79[38],pp78[40],pp77[42],pp76[44],pp75[46],pp74[48],pp73[50],pp72[52],pp71[54],pp70[56],pp69[58],pp70[58],pp71[58],pp72[58],pp73[58],pp74[58],pp75[58],pp76[58],pp77[58],pp78[58],pp79[58],pp80[58],pp81[58],pp82[58],pp83[58],pp84[58],pp85[58],pp86[58],pp87[58],pp88[58],pp89[58],pp90[58],pp91[58],pp92[58],pp93[58],pp94[58],pp95[58],pp96[58],pp97[58],pp98[58],pp99[58],pp149[9],pp151[8],pp153[7],pp155[6],pp157[5],pp159[4],pp160[4],pp161[4],pp162[4],pp163[4],pp164[4],pp165[4],pp166[4],pp167[4],pp168[4],pp169[4],pp170[4],pp171[4],pp172[4],pp173[4],pp174[4],pp175[4],pp176[4],pp177[4],pp178[4],pp179[4],pp180[4],pp181[4],pp182[4],pp183[4],pp184[4],pp185[4],pp186[4],pp187[4],pp188[4],pp189[4],pp190[4],pp191[4],pp192[4],pp193[4],pp194[4],pp195[4],pp196[4],pp197[4],pp198[4],pp199[4],pp200[4],pp201[4],pp202[4],pp204[3],pp206[2],pp208[1],pp210[0],s10[74],s11[74],s12[74],s13[74],s14[74],s15[74],s16[74],s17[74],s18[74],s19[74],s20[74],s21[74],s22[74],s23[74],s24[74],s25[74],s26[74],s26[75],s26[76],s26[77],s26[78],s26[79],s26[80],s26[81],s26[82],s26[83],s26[84],s26[85],s26[86],s26[87],s26[88],s26[89],s26[90],s26[91],s26[92],s26[93],s26[94],s26[95],s26[96],s26[97],s26[98],s26[99],s9[117],s8[119],s7[121],s6[123],s3[127],s121[10],s119[13],s117[16],s115[19],s113[22],s111[25],s109[28],s107[31],s105[34],s103[37],s101[40],s42[100],s41[102],s40[104],s39[106],s38[108],s37[110],s36[112],s35[114],s34[116],s33[118],s32[120],s31[122],s30[124],s29[126],s28[128],s27[130],s26[132],s25[134],s24[136],s23[138],s22[140],s21[142],s20[144],s19[146],s18[148],s17[150],s16[152],s15[154],s14[156],s13[158],s12[160],s11[162],s10[164],s171[196],s170[198],s169[200],s168[202],s167[204],s166[206],s165[208],s164[210],s163[212],s162[214],s161[216],s160[218],s159[220],s158[222],s157[224],s156[226],s155[228],s154[230],s153[232],s152[234],s151[236],s150[238],s149[240],s148[242],s147[244],s146[246],s145[248],s144[250],s143[252],s142[254],s141[256],s140[258],s139[260],s138[262],s137[264],s136[266],s135[268],s134[270],s133[272],s132[274],s131[276],s130[278],s129[280],pp255[90],pp254[92],pp253[94],pp252[96],pp251[98],pp99[251],pp97[254],pp251[101],pp249[104],pp247[107],pp245[110],pp244[112],pp243[114],pp242[116],pp241[118],pp240[120],pp239[122],pp238[124],pp237[126],pp236[128],pp235[130],pp234[132],pp233[134],pp232[136],pp231[138],pp230[140],pp229[142],pp228[144],pp227[146],pp226[148],pp225[150],pp224[152],pp223[154],pp222[156],pp221[158],pp220[160],pp219[162],pp218[164],pp217[166],pp216[168],pp217[168],pp218[168],pp219[168],pp220[168],pp221[168],pp222[168],pp223[168],pp224[168],pp225[168],pp226[168],pp227[168],pp228[168],pp229[168],pp230[168],pp231[168],pp232[168],pp233[168],pp234[168],pp235[168],pp236[168]};
    CLA_298 KS_172(s172, c172, in172_1, in172_2);
    wire[295:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {pp89[19],pp88[21],pp87[23],pp86[25],pp85[27],pp84[29],pp83[31],pp82[33],pp81[35],pp80[37],pp79[39],pp78[41],pp77[43],pp76[45],pp75[47],pp74[49],pp73[51],pp72[53],pp71[55],pp70[57],pp71[57],pp72[57],pp73[57],pp74[57],pp75[57],pp76[57],pp77[57],pp78[57],pp79[57],pp80[57],pp81[57],pp82[57],pp83[57],pp84[57],pp85[57],pp86[57],pp87[57],pp88[57],pp89[57],pp90[57],pp91[57],pp92[57],pp93[57],pp94[57],pp95[57],pp96[57],pp97[57],pp98[57],pp99[57],pp148[9],pp150[8],pp152[7],pp154[6],pp156[5],pp158[4],pp160[3],pp161[3],pp162[3],pp163[3],pp164[3],pp165[3],pp166[3],pp167[3],pp168[3],pp169[3],pp170[3],pp171[3],pp172[3],pp173[3],pp174[3],pp175[3],pp176[3],pp177[3],pp178[3],pp179[3],pp180[3],pp181[3],pp182[3],pp183[3],pp184[3],pp185[3],pp186[3],pp187[3],pp188[3],pp189[3],pp190[3],pp191[3],pp192[3],pp193[3],pp194[3],pp195[3],pp196[3],pp197[3],pp198[3],pp199[3],pp200[3],pp201[3],pp202[3],pp203[3],s172[100],s172[101],s172[102],s172[103],s172[104],s172[105],s172[106],s172[107],s172[108],s172[109],s172[110],s172[111],s172[112],s172[113],s172[114],s172[115],s172[116],s172[117],s172[118],s172[119],s172[120],s172[121],s172[122],s172[123],s172[124],s172[125],s172[126],s172[127],s172[128],s172[129],s172[130],s172[131],s172[132],s172[133],s172[134],s172[135],s172[136],s172[137],s172[138],s172[139],s172[140],s172[141],s172[142],s172[143],s172[144],s172[145],s172[146],s172[147],s172[148],s172[149],s172[150],s172[151],s172[152],s172[153],s172[154],s172[155],s172[156],s172[157],s172[158],s172[159],s172[160],s172[161],s172[162],s172[163],s172[164],s172[165],s172[166],s172[167],s172[168],s172[169],s172[170],s172[171],s172[172],s172[173],s172[174],s172[175],s172[176],s172[177],s172[178],s172[179],s172[180],s172[181],s172[182],s172[183],s172[184],s172[185],s172[186],s172[187],s172[188],s172[189],s172[190],s172[191],s172[192],s172[193],s172[194],s172[195],s171[197],s170[199],s169[201],s168[203],s167[205],s166[207],s165[209],s164[211],s163[213],s162[215],s161[217],s160[219],s159[221],s158[223],s157[225],s156[227],s155[229],s154[231],s153[233],s152[235],s151[237],s150[239],s149[241],s148[243],s147[245],s146[247],s145[249],s144[251],s143[253],s142[255],s141[257],s140[259],s139[261],s138[263],s137[265],s136[267],s135[269],s134[271],s133[273],s132[275],s131[277],s130[279],s129[281],pp255[91],pp254[93],pp253[95],pp252[97],pp251[99],pp98[253],pp252[100],pp250[103],pp248[106],pp246[109],pp245[111],pp244[113],pp243[115],pp242[117],pp241[119],pp240[121],pp239[123],pp238[125],pp237[127],pp236[129],pp235[131],pp234[133],pp233[135],pp232[137],pp231[139],pp230[141],pp229[143],pp228[145],pp227[147],pp226[149],pp225[151],pp224[153],pp223[155],pp222[157],pp221[159],pp220[161],pp219[163],pp218[165],pp217[167],pp218[167],pp219[167],pp220[167],pp221[167],pp222[167],pp223[167],pp224[167],pp225[167],pp226[167],pp227[167],pp228[167],pp229[167],pp230[167],pp231[167],pp232[167],pp233[167],pp234[167],pp235[167],pp236[167]};
    assign in173_2 = {pp90[18],pp89[20],pp88[22],pp87[24],pp86[26],pp85[28],pp84[30],pp83[32],pp82[34],pp81[36],pp80[38],pp79[40],pp78[42],pp77[44],pp76[46],pp75[48],pp74[50],pp73[52],pp72[54],pp71[56],pp72[56],pp73[56],pp74[56],pp75[56],pp76[56],pp77[56],pp78[56],pp79[56],pp80[56],pp81[56],pp82[56],pp83[56],pp84[56],pp85[56],pp86[56],pp87[56],pp88[56],pp89[56],pp90[56],pp91[56],pp92[56],pp93[56],pp94[56],pp95[56],pp96[56],pp97[56],pp98[56],pp99[56],pp147[9],pp149[8],pp151[7],pp153[6],pp155[5],pp157[4],pp159[3],pp161[2],pp162[2],pp163[2],pp164[2],pp165[2],pp166[2],pp167[2],pp168[2],pp169[2],pp170[2],pp171[2],pp172[2],pp173[2],pp174[2],pp175[2],pp176[2],pp177[2],pp178[2],pp179[2],pp180[2],pp181[2],pp182[2],pp183[2],pp184[2],pp185[2],pp186[2],pp187[2],pp188[2],pp189[2],pp190[2],pp191[2],pp192[2],pp193[2],pp194[2],pp195[2],pp196[2],pp197[2],pp198[2],pp199[2],pp200[2],pp201[2],pp202[2],pp203[2],pp204[2],pp205[2],pp207[1],pp209[0],s10[73],s11[73],s12[73],s13[73],s14[73],s15[73],s16[73],s17[73],s18[73],s19[73],s20[73],s21[73],s22[73],s23[73],s24[73],s25[73],s26[73],s27[73],s27[74],s27[75],s27[76],s27[77],s27[78],s27[79],s27[80],s27[81],s27[82],s27[83],s27[84],s27[85],s27[86],s27[87],s27[88],s27[89],s27[90],s27[91],s27[92],s27[93],s27[94],s27[95],s27[96],s27[97],s27[98],s27[99],s9[118],s8[120],s7[122],s4[126],s1[130],s120[12],s118[15],s116[18],s114[21],s112[24],s110[27],s108[30],s106[33],s104[36],s102[39],s100[42],s42[101],s41[103],s40[105],s39[107],s38[109],s37[111],s36[113],s35[115],s34[117],s33[119],s32[121],s31[123],s30[125],s29[127],s28[129],s27[131],s26[133],s25[135],s24[137],s23[139],s22[141],s21[143],s20[145],s19[147],s18[149],s17[151],s16[153],s15[155],s14[157],s13[159],s12[161],s11[163],s10[165],s172[196],s171[198],s170[200],s169[202],s168[204],s167[206],s166[208],s165[210],s164[212],s163[214],s162[216],s161[218],s160[220],s159[222],s158[224],s157[226],s156[228],s155[230],s154[232],s153[234],s152[236],s151[238],s150[240],s149[242],s148[244],s147[246],s146[248],s145[250],s144[252],s143[254],s142[256],s141[258],s140[260],s139[262],s138[264],s137[266],s136[268],s135[270],s134[272],s133[274],s132[276],s131[278],s130[280],s129[282],pp255[92],pp254[94],pp253[96],pp252[98],pp99[252],pp97[255],pp251[102],pp249[105],pp247[108],pp246[110],pp245[112],pp244[114],pp243[116],pp242[118],pp241[120],pp240[122],pp239[124],pp238[126],pp237[128],pp236[130],pp235[132],pp234[134],pp233[136],pp232[138],pp231[140],pp230[142],pp229[144],pp228[146],pp227[148],pp226[150],pp225[152],pp224[154],pp223[156],pp222[158],pp221[160],pp220[162],pp219[164],pp218[166],pp219[166],pp220[166],pp221[166],pp222[166],pp223[166],pp224[166],pp225[166],pp226[166],pp227[166],pp228[166],pp229[166],pp230[166],pp231[166],pp232[166],pp233[166],pp234[166],pp235[166],pp236[166],pp237[166]};
    CLA_296 KS_173(s173, c173, in173_1, in173_2);
    wire[293:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp90[19],pp89[21],pp88[23],pp87[25],pp86[27],pp85[29],pp84[31],pp83[33],pp82[35],pp81[37],pp80[39],pp79[41],pp78[43],pp77[45],pp76[47],pp75[49],pp74[51],pp73[53],pp72[55],pp73[55],pp74[55],pp75[55],pp76[55],pp77[55],pp78[55],pp79[55],pp80[55],pp81[55],pp82[55],pp83[55],pp84[55],pp85[55],pp86[55],pp87[55],pp88[55],pp89[55],pp90[55],pp91[55],pp92[55],pp93[55],pp94[55],pp95[55],pp96[55],pp97[55],pp98[55],pp99[55],pp146[9],pp148[8],pp150[7],pp152[6],pp154[5],pp156[4],pp158[3],pp160[2],pp162[1],pp163[1],pp164[1],pp165[1],pp166[1],pp167[1],pp168[1],pp169[1],pp170[1],pp171[1],pp172[1],pp173[1],pp174[1],pp175[1],pp176[1],pp177[1],pp178[1],pp179[1],pp180[1],pp181[1],pp182[1],pp183[1],pp184[1],pp185[1],pp186[1],pp187[1],pp188[1],pp189[1],pp190[1],pp191[1],pp192[1],pp193[1],pp194[1],pp195[1],pp196[1],pp197[1],pp198[1],pp199[1],pp200[1],pp201[1],pp202[1],pp203[1],pp204[1],pp205[1],pp206[1],s173[100],s173[101],s173[102],s173[103],s173[104],s173[105],s173[106],s173[107],s173[108],s173[109],s173[110],s173[111],s173[112],s173[113],s173[114],s173[115],s173[116],s173[117],s173[118],s173[119],s173[120],s173[121],s173[122],s173[123],s173[124],s173[125],s173[126],s173[127],s173[128],s173[129],s173[130],s173[131],s173[132],s173[133],s173[134],s173[135],s173[136],s173[137],s173[138],s173[139],s173[140],s173[141],s173[142],s173[143],s173[144],s173[145],s173[146],s173[147],s173[148],s173[149],s173[150],s173[151],s173[152],s173[153],s173[154],s173[155],s173[156],s173[157],s173[158],s173[159],s173[160],s173[161],s173[162],s173[163],s173[164],s173[165],s173[166],s173[167],s173[168],s173[169],s173[170],s173[171],s173[172],s173[173],s173[174],s173[175],s173[176],s173[177],s173[178],s173[179],s173[180],s173[181],s173[182],s173[183],s173[184],s173[185],s173[186],s173[187],s173[188],s173[189],s173[190],s173[191],s173[192],s173[193],s173[194],s173[195],s172[197],s171[199],s170[201],s169[203],s168[205],s167[207],s166[209],s165[211],s164[213],s163[215],s162[217],s161[219],s160[221],s159[223],s158[225],s157[227],s156[229],s155[231],s154[233],s153[235],s152[237],s151[239],s150[241],s149[243],s148[245],s147[247],s146[249],s145[251],s144[253],s143[255],s142[257],s141[259],s140[261],s139[263],s138[265],s137[267],s136[269],s135[271],s134[273],s133[275],s132[277],s131[279],s130[281],s129[283],pp255[93],pp254[95],pp253[97],pp252[99],pp98[254],pp252[101],pp250[104],pp248[107],pp247[109],pp246[111],pp245[113],pp244[115],pp243[117],pp242[119],pp241[121],pp240[123],pp239[125],pp238[127],pp237[129],pp236[131],pp235[133],pp234[135],pp233[137],pp232[139],pp231[141],pp230[143],pp229[145],pp228[147],pp227[149],pp226[151],pp225[153],pp224[155],pp223[157],pp222[159],pp221[161],pp220[163],pp219[165],pp220[165],pp221[165],pp222[165],pp223[165],pp224[165],pp225[165],pp226[165],pp227[165],pp228[165],pp229[165],pp230[165],pp231[165],pp232[165],pp233[165],pp234[165],pp235[165],pp236[165],pp237[165]};
    assign in174_2 = {pp91[18],pp90[20],pp89[22],pp88[24],pp87[26],pp86[28],pp85[30],pp84[32],pp83[34],pp82[36],pp81[38],pp80[40],pp79[42],pp78[44],pp77[46],pp76[48],pp75[50],pp74[52],pp73[54],pp74[54],pp75[54],pp76[54],pp77[54],pp78[54],pp79[54],pp80[54],pp81[54],pp82[54],pp83[54],pp84[54],pp85[54],pp86[54],pp87[54],pp88[54],pp89[54],pp90[54],pp91[54],pp92[54],pp93[54],pp94[54],pp95[54],pp96[54],pp97[54],pp98[54],pp99[54],pp145[9],pp147[8],pp149[7],pp151[6],pp153[5],pp155[4],pp157[3],pp159[2],pp161[1],pp163[0],pp164[0],pp165[0],pp166[0],pp167[0],pp168[0],pp169[0],pp170[0],pp171[0],pp172[0],pp173[0],pp174[0],pp175[0],pp176[0],pp177[0],pp178[0],pp179[0],pp180[0],pp181[0],pp182[0],pp183[0],pp184[0],pp185[0],pp186[0],pp187[0],pp188[0],pp189[0],pp190[0],pp191[0],pp192[0],pp193[0],pp194[0],pp195[0],pp196[0],pp197[0],pp198[0],pp199[0],pp200[0],pp201[0],pp202[0],pp203[0],pp204[0],pp205[0],pp206[0],pp207[0],pp208[0],s10[72],s11[72],s12[72],s13[72],s14[72],s15[72],s16[72],s17[72],s18[72],s19[72],s20[72],s21[72],s22[72],s23[72],s24[72],s25[72],s26[72],s27[72],s28[72],s28[73],s28[74],s28[75],s28[76],s28[77],s28[78],s28[79],s28[80],s28[81],s28[82],s28[83],s28[84],s28[85],s28[86],s28[87],s28[88],s28[89],s28[90],s28[91],s28[92],s28[93],s28[94],s28[95],s28[96],s28[97],s28[98],s28[99],s9[119],s8[121],s5[125],s2[129],s121[11],s119[14],s117[17],s115[20],s113[23],s111[26],s109[29],s107[32],s105[35],s103[38],s101[41],s43[100],s42[102],s41[104],s40[106],s39[108],s38[110],s37[112],s36[114],s35[116],s34[118],s33[120],s32[122],s31[124],s30[126],s29[128],s28[130],s27[132],s26[134],s25[136],s24[138],s23[140],s22[142],s21[144],s20[146],s19[148],s18[150],s17[152],s16[154],s15[156],s14[158],s13[160],s12[162],s11[164],s10[166],s173[196],s172[198],s171[200],s170[202],s169[204],s168[206],s167[208],s166[210],s165[212],s164[214],s163[216],s162[218],s161[220],s160[222],s159[224],s158[226],s157[228],s156[230],s155[232],s154[234],s153[236],s152[238],s151[240],s150[242],s149[244],s148[246],s147[248],s146[250],s145[252],s144[254],s143[256],s142[258],s141[260],s140[262],s139[264],s138[266],s137[268],s136[270],s135[272],s134[274],s133[276],s132[278],s131[280],s130[282],s129[284],pp255[94],pp254[96],pp253[98],pp99[253],pp253[100],pp251[103],pp249[106],pp248[108],pp247[110],pp246[112],pp245[114],pp244[116],pp243[118],pp242[120],pp241[122],pp240[124],pp239[126],pp238[128],pp237[130],pp236[132],pp235[134],pp234[136],pp233[138],pp232[140],pp231[142],pp230[144],pp229[146],pp228[148],pp227[150],pp226[152],pp225[154],pp224[156],pp223[158],pp222[160],pp221[162],pp220[164],pp221[164],pp222[164],pp223[164],pp224[164],pp225[164],pp226[164],pp227[164],pp228[164],pp229[164],pp230[164],pp231[164],pp232[164],pp233[164],pp234[164],pp235[164],pp236[164],pp237[164],pp238[164]};
    CLA_294 KS_174(s174, c174, in174_1, in174_2);
    wire[291:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp91[19],pp90[21],pp89[23],pp88[25],pp87[27],pp86[29],pp85[31],pp84[33],pp83[35],pp82[37],pp81[39],pp80[41],pp79[43],pp78[45],pp77[47],pp76[49],pp75[51],pp74[53],pp75[53],pp76[53],pp77[53],pp78[53],pp79[53],pp80[53],pp81[53],pp82[53],pp83[53],pp84[53],pp85[53],pp86[53],pp87[53],pp88[53],pp89[53],pp90[53],pp91[53],pp92[53],pp93[53],pp94[53],pp95[53],pp96[53],pp97[53],pp98[53],pp99[53],pp144[9],pp146[8],pp148[7],pp150[6],pp152[5],pp154[4],pp156[3],pp158[2],pp160[1],pp162[0],s129[99],s130[99],s131[99],s132[99],s133[99],s134[99],s135[99],s136[99],s137[99],s138[99],s139[99],s140[99],s141[99],s142[99],s143[99],s144[99],s145[99],s146[99],s147[99],s148[99],s149[99],s150[99],s151[99],s152[99],s153[99],s154[99],s155[99],s156[99],s157[99],s158[99],s159[99],s160[99],s161[99],s162[99],s163[99],s164[99],s165[99],s166[99],s167[99],s168[99],s169[99],s170[99],s171[99],s172[99],s173[99],s174[99],s174[100],s174[101],s174[102],s174[103],s174[104],s174[105],s174[106],s174[107],s174[108],s174[109],s174[110],s174[111],s174[112],s174[113],s174[114],s174[115],s174[116],s174[117],s174[118],s174[119],s174[120],s174[121],s174[122],s174[123],s174[124],s174[125],s174[126],s174[127],s174[128],s174[129],s174[130],s174[131],s174[132],s174[133],s174[134],s174[135],s174[136],s174[137],s174[138],s174[139],s174[140],s174[141],s174[142],s174[143],s174[144],s174[145],s174[146],s174[147],s174[148],s174[149],s174[150],s174[151],s174[152],s174[153],s174[154],s174[155],s174[156],s174[157],s174[158],s174[159],s174[160],s174[161],s174[162],s174[163],s174[164],s174[165],s174[166],s174[167],s174[168],s174[169],s174[170],s174[171],s174[172],s174[173],s174[174],s174[175],s174[176],s174[177],s174[178],s174[179],s174[180],s174[181],s174[182],s174[183],s174[184],s174[185],s174[186],s174[187],s174[188],s174[189],s174[190],s174[191],s174[192],s174[193],s174[194],s174[195],s173[197],s172[199],s171[201],s170[203],s169[205],s168[207],s167[209],s166[211],s165[213],s164[215],s163[217],s162[219],s161[221],s160[223],s159[225],s158[227],s157[229],s156[231],s155[233],s154[235],s153[237],s152[239],s151[241],s150[243],s149[245],s148[247],s147[249],s146[251],s145[253],s144[255],s143[257],s142[259],s141[261],s140[263],s139[265],s138[267],s137[269],s136[271],s135[273],s134[275],s133[277],s132[279],s131[281],s130[283],s129[285],pp255[95],pp254[97],pp253[99],pp98[255],pp252[102],pp250[105],pp249[107],pp248[109],pp247[111],pp246[113],pp245[115],pp244[117],pp243[119],pp242[121],pp241[123],pp240[125],pp239[127],pp238[129],pp237[131],pp236[133],pp235[135],pp234[137],pp233[139],pp232[141],pp231[143],pp230[145],pp229[147],pp228[149],pp227[151],pp226[153],pp225[155],pp224[157],pp223[159],pp222[161],pp221[163],pp222[163],pp223[163],pp224[163],pp225[163],pp226[163],pp227[163],pp228[163],pp229[163],pp230[163],pp231[163],pp232[163],pp233[163],pp234[163],pp235[163],pp236[163],pp237[163],pp238[163]};
    assign in175_2 = {pp92[18],pp91[20],pp90[22],pp89[24],pp88[26],pp87[28],pp86[30],pp85[32],pp84[34],pp83[36],pp82[38],pp81[40],pp80[42],pp79[44],pp78[46],pp77[48],pp76[50],pp75[52],pp76[52],pp77[52],pp78[52],pp79[52],pp80[52],pp81[52],pp82[52],pp83[52],pp84[52],pp85[52],pp86[52],pp87[52],pp88[52],pp89[52],pp90[52],pp91[52],pp92[52],pp93[52],pp94[52],pp95[52],pp96[52],pp97[52],pp98[52],pp99[52],pp143[9],pp145[8],pp147[7],pp149[6],pp151[5],pp153[4],pp155[3],pp157[2],pp159[1],pp161[0],s129[98],s130[98],s131[98],s132[98],s133[98],s134[98],s135[98],s136[98],s137[98],s138[98],s139[98],s140[98],s141[98],s142[98],s143[98],s144[98],s145[98],s146[98],s147[98],s148[98],s149[98],s150[98],s151[98],s152[98],s153[98],s154[98],s155[98],s156[98],s157[98],s158[98],s159[98],s160[98],s161[98],s162[98],s163[98],s164[98],s165[98],s166[98],s167[98],s168[98],s169[98],s170[98],s171[98],s172[98],s173[98],s174[98],s10[71],s11[71],s12[71],s13[71],s14[71],s15[71],s16[71],s17[71],s18[71],s19[71],s20[71],s21[71],s22[71],s23[71],s24[71],s25[71],s26[71],s27[71],s28[71],s29[71],s29[72],s29[73],s29[74],s29[75],s29[76],s29[77],s29[78],s29[79],s29[80],s29[81],s29[82],s29[83],s29[84],s29[85],s29[86],s29[87],s29[88],s29[89],s29[90],s29[91],s29[92],s29[93],s29[94],s29[95],s29[96],s29[97],s29[98],s29[99],s9[120],s6[124],s3[128],s122[10],s120[13],s118[16],s116[19],s114[22],s112[25],s110[28],s108[31],s106[34],s104[37],s102[40],s100[43],s43[101],s42[103],s41[105],s40[107],s39[109],s38[111],s37[113],s36[115],s35[117],s34[119],s33[121],s32[123],s31[125],s30[127],s29[129],s28[131],s27[133],s26[135],s25[137],s24[139],s23[141],s22[143],s21[145],s20[147],s19[149],s18[151],s17[153],s16[155],s15[157],s14[159],s13[161],s12[163],s11[165],s10[167],s174[196],s173[198],s172[200],s171[202],s170[204],s169[206],s168[208],s167[210],s166[212],s165[214],s164[216],s163[218],s162[220],s161[222],s160[224],s159[226],s158[228],s157[230],s156[232],s155[234],s154[236],s153[238],s152[240],s151[242],s150[244],s149[246],s148[248],s147[250],s146[252],s145[254],s144[256],s143[258],s142[260],s141[262],s140[264],s139[266],s138[268],s137[270],s136[272],s135[274],s134[276],s133[278],s132[280],s131[282],s130[284],s129[286],pp255[96],pp254[98],pp99[254],pp253[101],pp251[104],pp250[106],pp249[108],pp248[110],pp247[112],pp246[114],pp245[116],pp244[118],pp243[120],pp242[122],pp241[124],pp240[126],pp239[128],pp238[130],pp237[132],pp236[134],pp235[136],pp234[138],pp233[140],pp232[142],pp231[144],pp230[146],pp229[148],pp228[150],pp227[152],pp226[154],pp225[156],pp224[158],pp223[160],pp222[162],pp223[162],pp224[162],pp225[162],pp226[162],pp227[162],pp228[162],pp229[162],pp230[162],pp231[162],pp232[162],pp233[162],pp234[162],pp235[162],pp236[162],pp237[162],pp238[162],pp239[162]};
    CLA_292 KS_175(s175, c175, in175_1, in175_2);
    wire[289:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp92[19],pp91[21],pp90[23],pp89[25],pp88[27],pp87[29],pp86[31],pp85[33],pp84[35],pp83[37],pp82[39],pp81[41],pp80[43],pp79[45],pp78[47],pp77[49],pp76[51],pp77[51],pp78[51],pp79[51],pp80[51],pp81[51],pp82[51],pp83[51],pp84[51],pp85[51],pp86[51],pp87[51],pp88[51],pp89[51],pp90[51],pp91[51],pp92[51],pp93[51],pp94[51],pp95[51],pp96[51],pp97[51],pp98[51],pp99[51],pp142[9],pp144[8],pp146[7],pp148[6],pp150[5],pp152[4],pp154[3],pp156[2],pp158[1],pp160[0],s129[97],s130[97],s131[97],s132[97],s133[97],s134[97],s135[97],s136[97],s137[97],s138[97],s139[97],s140[97],s141[97],s142[97],s143[97],s144[97],s145[97],s146[97],s147[97],s148[97],s149[97],s150[97],s151[97],s152[97],s153[97],s154[97],s155[97],s156[97],s157[97],s158[97],s159[97],s160[97],s161[97],s162[97],s163[97],s164[97],s165[97],s166[97],s167[97],s168[97],s169[97],s170[97],s171[97],s172[97],s173[97],s174[97],s175[97],s175[98],s175[99],s175[100],s175[101],s175[102],s175[103],s175[104],s175[105],s175[106],s175[107],s175[108],s175[109],s175[110],s175[111],s175[112],s175[113],s175[114],s175[115],s175[116],s175[117],s175[118],s175[119],s175[120],s175[121],s175[122],s175[123],s175[124],s175[125],s175[126],s175[127],s175[128],s175[129],s175[130],s175[131],s175[132],s175[133],s175[134],s175[135],s175[136],s175[137],s175[138],s175[139],s175[140],s175[141],s175[142],s175[143],s175[144],s175[145],s175[146],s175[147],s175[148],s175[149],s175[150],s175[151],s175[152],s175[153],s175[154],s175[155],s175[156],s175[157],s175[158],s175[159],s175[160],s175[161],s175[162],s175[163],s175[164],s175[165],s175[166],s175[167],s175[168],s175[169],s175[170],s175[171],s175[172],s175[173],s175[174],s175[175],s175[176],s175[177],s175[178],s175[179],s175[180],s175[181],s175[182],s175[183],s175[184],s175[185],s175[186],s175[187],s175[188],s175[189],s175[190],s175[191],s175[192],s175[193],s175[194],s175[195],s174[197],s173[199],s172[201],s171[203],s170[205],s169[207],s168[209],s167[211],s166[213],s165[215],s164[217],s163[219],s162[221],s161[223],s160[225],s159[227],s158[229],s157[231],s156[233],s155[235],s154[237],s153[239],s152[241],s151[243],s150[245],s149[247],s148[249],s147[251],s146[253],s145[255],s144[257],s143[259],s142[261],s141[263],s140[265],s139[267],s138[269],s137[271],s136[273],s135[275],s134[277],s133[279],s132[281],s131[283],s130[285],s129[287],pp255[97],pp254[99],pp254[100],pp252[103],pp251[105],pp250[107],pp249[109],pp248[111],pp247[113],pp246[115],pp245[117],pp244[119],pp243[121],pp242[123],pp241[125],pp240[127],pp239[129],pp238[131],pp237[133],pp236[135],pp235[137],pp234[139],pp233[141],pp232[143],pp231[145],pp230[147],pp229[149],pp228[151],pp227[153],pp226[155],pp225[157],pp224[159],pp223[161],pp224[161],pp225[161],pp226[161],pp227[161],pp228[161],pp229[161],pp230[161],pp231[161],pp232[161],pp233[161],pp234[161],pp235[161],pp236[161],pp237[161],pp238[161],pp239[161]};
    assign in176_2 = {pp93[18],pp92[20],pp91[22],pp90[24],pp89[26],pp88[28],pp87[30],pp86[32],pp85[34],pp84[36],pp83[38],pp82[40],pp81[42],pp80[44],pp79[46],pp78[48],pp77[50],pp78[50],pp79[50],pp80[50],pp81[50],pp82[50],pp83[50],pp84[50],pp85[50],pp86[50],pp87[50],pp88[50],pp89[50],pp90[50],pp91[50],pp92[50],pp93[50],pp94[50],pp95[50],pp96[50],pp97[50],pp98[50],pp99[50],pp141[9],pp143[8],pp145[7],pp147[6],pp149[5],pp151[4],pp153[3],pp155[2],pp157[1],pp159[0],s129[96],s130[96],s131[96],s132[96],s133[96],s134[96],s135[96],s136[96],s137[96],s138[96],s139[96],s140[96],s141[96],s142[96],s143[96],s144[96],s145[96],s146[96],s147[96],s148[96],s149[96],s150[96],s151[96],s152[96],s153[96],s154[96],s155[96],s156[96],s157[96],s158[96],s159[96],s160[96],s161[96],s162[96],s163[96],s164[96],s165[96],s166[96],s167[96],s168[96],s169[96],s170[96],s171[96],s172[96],s173[96],s174[96],s175[96],s10[70],s11[70],s12[70],s13[70],s14[70],s15[70],s16[70],s17[70],s18[70],s19[70],s20[70],s21[70],s22[70],s23[70],s24[70],s25[70],s26[70],s27[70],s28[70],s29[70],s30[70],s30[71],s30[72],s30[73],s30[74],s30[75],s30[76],s30[77],s30[78],s30[79],s30[80],s30[81],s30[82],s30[83],s30[84],s30[85],s30[86],s30[87],s30[88],s30[89],s30[90],s30[91],s30[92],s30[93],s30[94],s30[95],s30[96],s30[97],s30[98],s30[99],s7[123],s4[127],s1[131],s121[12],s119[15],s117[18],s115[21],s113[24],s111[27],s109[30],s107[33],s105[36],s103[39],s101[42],s44[100],s43[102],s42[104],s41[106],s40[108],s39[110],s38[112],s37[114],s36[116],s35[118],s34[120],s33[122],s32[124],s31[126],s30[128],s29[130],s28[132],s27[134],s26[136],s25[138],s24[140],s23[142],s22[144],s21[146],s20[148],s19[150],s18[152],s17[154],s16[156],s15[158],s14[160],s13[162],s12[164],s11[166],s10[168],s175[196],s174[198],s173[200],s172[202],s171[204],s170[206],s169[208],s168[210],s167[212],s166[214],s165[216],s164[218],s163[220],s162[222],s161[224],s160[226],s159[228],s158[230],s157[232],s156[234],s155[236],s154[238],s153[240],s152[242],s151[244],s150[246],s149[248],s148[250],s147[252],s146[254],s145[256],s144[258],s143[260],s142[262],s141[264],s140[266],s139[268],s138[270],s137[272],s136[274],s135[276],s134[278],s133[280],s132[282],s131[284],s130[286],s129[288],pp255[98],pp99[255],pp253[102],pp252[104],pp251[106],pp250[108],pp249[110],pp248[112],pp247[114],pp246[116],pp245[118],pp244[120],pp243[122],pp242[124],pp241[126],pp240[128],pp239[130],pp238[132],pp237[134],pp236[136],pp235[138],pp234[140],pp233[142],pp232[144],pp231[146],pp230[148],pp229[150],pp228[152],pp227[154],pp226[156],pp225[158],pp224[160],pp225[160],pp226[160],pp227[160],pp228[160],pp229[160],pp230[160],pp231[160],pp232[160],pp233[160],pp234[160],pp235[160],pp236[160],pp237[160],pp238[160],pp239[160],pp240[160]};
    CLA_290 KS_176(s176, c176, in176_1, in176_2);
    wire[287:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp93[19],pp92[21],pp91[23],pp90[25],pp89[27],pp88[29],pp87[31],pp86[33],pp85[35],pp84[37],pp83[39],pp82[41],pp81[43],pp80[45],pp79[47],pp78[49],pp79[49],pp80[49],pp81[49],pp82[49],pp83[49],pp84[49],pp85[49],pp86[49],pp87[49],pp88[49],pp89[49],pp90[49],pp91[49],pp92[49],pp93[49],pp94[49],pp95[49],pp96[49],pp97[49],pp98[49],pp99[49],pp140[9],pp142[8],pp144[7],pp146[6],pp148[5],pp150[4],pp152[3],pp154[2],pp156[1],pp158[0],s129[95],s130[95],s131[95],s132[95],s133[95],s134[95],s135[95],s136[95],s137[95],s138[95],s139[95],s140[95],s141[95],s142[95],s143[95],s144[95],s145[95],s146[95],s147[95],s148[95],s149[95],s150[95],s151[95],s152[95],s153[95],s154[95],s155[95],s156[95],s157[95],s158[95],s159[95],s160[95],s161[95],s162[95],s163[95],s164[95],s165[95],s166[95],s167[95],s168[95],s169[95],s170[95],s171[95],s172[95],s173[95],s174[95],s175[95],s176[95],s176[96],s176[97],s176[98],s176[99],s176[100],s176[101],s176[102],s176[103],s176[104],s176[105],s176[106],s176[107],s176[108],s176[109],s176[110],s176[111],s176[112],s176[113],s176[114],s176[115],s176[116],s176[117],s176[118],s176[119],s176[120],s176[121],s176[122],s176[123],s176[124],s176[125],s176[126],s176[127],s176[128],s176[129],s176[130],s176[131],s176[132],s176[133],s176[134],s176[135],s176[136],s176[137],s176[138],s176[139],s176[140],s176[141],s176[142],s176[143],s176[144],s176[145],s176[146],s176[147],s176[148],s176[149],s176[150],s176[151],s176[152],s176[153],s176[154],s176[155],s176[156],s176[157],s176[158],s176[159],s176[160],s176[161],s176[162],s176[163],s176[164],s176[165],s176[166],s176[167],s176[168],s176[169],s176[170],s176[171],s176[172],s176[173],s176[174],s176[175],s176[176],s176[177],s176[178],s176[179],s176[180],s176[181],s176[182],s176[183],s176[184],s176[185],s176[186],s176[187],s176[188],s176[189],s176[190],s176[191],s176[192],s176[193],s176[194],s176[195],s175[197],s174[199],s173[201],s172[203],s171[205],s170[207],s169[209],s168[211],s167[213],s166[215],s165[217],s164[219],s163[221],s162[223],s161[225],s160[227],s159[229],s158[231],s157[233],s156[235],s155[237],s154[239],s153[241],s152[243],s151[245],s150[247],s149[249],s148[251],s147[253],s146[255],s145[257],s144[259],s143[261],s142[263],s141[265],s140[267],s139[269],s138[271],s137[273],s136[275],s135[277],s134[279],s133[281],s132[283],s131[285],s130[287],s129[289],pp255[99],pp254[101],pp253[103],pp252[105],pp251[107],pp250[109],pp249[111],pp248[113],pp247[115],pp246[117],pp245[119],pp244[121],pp243[123],pp242[125],pp241[127],pp240[129],pp239[131],pp238[133],pp237[135],pp236[137],pp235[139],pp234[141],pp233[143],pp232[145],pp231[147],pp230[149],pp229[151],pp228[153],pp227[155],pp226[157],pp225[159],pp226[159],pp227[159],pp228[159],pp229[159],pp230[159],pp231[159],pp232[159],pp233[159],pp234[159],pp235[159],pp236[159],pp237[159],pp238[159],pp239[159],pp240[159]};
    assign in177_2 = {pp94[18],pp93[20],pp92[22],pp91[24],pp90[26],pp89[28],pp88[30],pp87[32],pp86[34],pp85[36],pp84[38],pp83[40],pp82[42],pp81[44],pp80[46],pp79[48],pp80[48],pp81[48],pp82[48],pp83[48],pp84[48],pp85[48],pp86[48],pp87[48],pp88[48],pp89[48],pp90[48],pp91[48],pp92[48],pp93[48],pp94[48],pp95[48],pp96[48],pp97[48],pp98[48],pp99[48],pp139[9],pp141[8],pp143[7],pp145[6],pp147[5],pp149[4],pp151[3],pp153[2],pp155[1],pp157[0],s129[94],s130[94],s131[94],s132[94],s133[94],s134[94],s135[94],s136[94],s137[94],s138[94],s139[94],s140[94],s141[94],s142[94],s143[94],s144[94],s145[94],s146[94],s147[94],s148[94],s149[94],s150[94],s151[94],s152[94],s153[94],s154[94],s155[94],s156[94],s157[94],s158[94],s159[94],s160[94],s161[94],s162[94],s163[94],s164[94],s165[94],s166[94],s167[94],s168[94],s169[94],s170[94],s171[94],s172[94],s173[94],s174[94],s175[94],s176[94],s10[69],s11[69],s12[69],s13[69],s14[69],s15[69],s16[69],s17[69],s18[69],s19[69],s20[69],s21[69],s22[69],s23[69],s24[69],s25[69],s26[69],s27[69],s28[69],s29[69],s30[69],s31[69],s31[70],s31[71],s31[72],s31[73],s31[74],s31[75],s31[76],s31[77],s31[78],s31[79],s31[80],s31[81],s31[82],s31[83],s31[84],s31[85],s31[86],s31[87],s31[88],s31[89],s31[90],s31[91],s31[92],s31[93],s31[94],s31[95],s31[96],s31[97],s31[98],s8[122],s5[126],s2[130],s122[11],s120[14],s118[17],s116[20],s114[23],s112[26],s110[29],s108[32],s106[35],s104[38],s102[41],s100[44],s44[101],s43[103],s42[105],s41[107],s40[109],s39[111],s38[113],s37[115],s36[117],s35[119],s34[121],s33[123],s32[125],s31[127],s30[129],s29[131],s28[133],s27[135],s26[137],s25[139],s24[141],s23[143],s22[145],s21[147],s20[149],s19[151],s18[153],s17[155],s16[157],s15[159],s14[161],s13[163],s12[165],s11[167],s10[169],s176[196],s175[198],s174[200],s173[202],s172[204],s171[206],s170[208],s169[210],s168[212],s167[214],s166[216],s165[218],s164[220],s163[222],s162[224],s161[226],s160[228],s159[230],s158[232],s157[234],s156[236],s155[238],s154[240],s153[242],s152[244],s151[246],s150[248],s149[250],s148[252],s147[254],s146[256],s145[258],s144[260],s143[262],s142[264],s141[266],s140[268],s139[270],s138[272],s137[274],s136[276],s135[278],s134[280],s133[282],s132[284],s131[286],s130[288],s129[290],pp255[100],pp254[102],pp253[104],pp252[106],pp251[108],pp250[110],pp249[112],pp248[114],pp247[116],pp246[118],pp245[120],pp244[122],pp243[124],pp242[126],pp241[128],pp240[130],pp239[132],pp238[134],pp237[136],pp236[138],pp235[140],pp234[142],pp233[144],pp232[146],pp231[148],pp230[150],pp229[152],pp228[154],pp227[156],pp226[158],pp227[158],pp228[158],pp229[158],pp230[158],pp231[158],pp232[158],pp233[158],pp234[158],pp235[158],pp236[158],pp237[158],pp238[158],pp239[158],pp240[158],pp241[158]};
    CLA_288 KS_177(s177, c177, in177_1, in177_2);
    wire[285:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {pp94[19],pp93[21],pp92[23],pp91[25],pp90[27],pp89[29],pp88[31],pp87[33],pp86[35],pp85[37],pp84[39],pp83[41],pp82[43],pp81[45],pp80[47],pp81[47],pp82[47],pp83[47],pp84[47],pp85[47],pp86[47],pp87[47],pp88[47],pp89[47],pp90[47],pp91[47],pp92[47],pp93[47],pp94[47],pp95[47],pp96[47],pp97[47],pp98[47],pp99[47],pp138[9],pp140[8],pp142[7],pp144[6],pp146[5],pp148[4],pp150[3],pp152[2],pp154[1],pp156[0],s129[93],s130[93],s131[93],s132[93],s133[93],s134[93],s135[93],s136[93],s137[93],s138[93],s139[93],s140[93],s141[93],s142[93],s143[93],s144[93],s145[93],s146[93],s147[93],s148[93],s149[93],s150[93],s151[93],s152[93],s153[93],s154[93],s155[93],s156[93],s157[93],s158[93],s159[93],s160[93],s161[93],s162[93],s163[93],s164[93],s165[93],s166[93],s167[93],s168[93],s169[93],s170[93],s171[93],s172[93],s173[93],s174[93],s175[93],s176[93],s177[93],s177[94],s177[95],s177[96],s177[97],s177[98],s177[99],s177[100],s177[101],s177[102],s177[103],s177[104],s177[105],s177[106],s177[107],s177[108],s177[109],s177[110],s177[111],s177[112],s177[113],s177[114],s177[115],s177[116],s177[117],s177[118],s177[119],s177[120],s177[121],s177[122],s177[123],s177[124],s177[125],s177[126],s177[127],s177[128],s177[129],s177[130],s177[131],s177[132],s177[133],s177[134],s177[135],s177[136],s177[137],s177[138],s177[139],s177[140],s177[141],s177[142],s177[143],s177[144],s177[145],s177[146],s177[147],s177[148],s177[149],s177[150],s177[151],s177[152],s177[153],s177[154],s177[155],s177[156],s177[157],s177[158],s177[159],s177[160],s177[161],s177[162],s177[163],s177[164],s177[165],s177[166],s177[167],s177[168],s177[169],s177[170],s177[171],s177[172],s177[173],s177[174],s177[175],s177[176],s177[177],s177[178],s177[179],s177[180],s177[181],s177[182],s177[183],s177[184],s177[185],s177[186],s177[187],s177[188],s177[189],s177[190],s177[191],s177[192],s177[193],s177[194],s177[195],s176[197],s175[199],s174[201],s173[203],s172[205],s171[207],s170[209],s169[211],s168[213],s167[215],s166[217],s165[219],s164[221],s163[223],s162[225],s161[227],s160[229],s159[231],s158[233],s157[235],s156[237],s155[239],s154[241],s153[243],s152[245],s151[247],s150[249],s149[251],s148[253],s147[255],s146[257],s145[259],s144[261],s143[263],s142[265],s141[267],s140[269],s139[271],s138[273],s137[275],s136[277],s135[279],s134[281],s133[283],s132[285],s131[287],s130[289],s129[291],pp255[101],pp254[103],pp253[105],pp252[107],pp251[109],pp250[111],pp249[113],pp248[115],pp247[117],pp246[119],pp245[121],pp244[123],pp243[125],pp242[127],pp241[129],pp240[131],pp239[133],pp238[135],pp237[137],pp236[139],pp235[141],pp234[143],pp233[145],pp232[147],pp231[149],pp230[151],pp229[153],pp228[155],pp227[157],pp228[157],pp229[157],pp230[157],pp231[157],pp232[157],pp233[157],pp234[157],pp235[157],pp236[157],pp237[157],pp238[157],pp239[157],pp240[157],pp241[157]};
    assign in178_2 = {pp95[18],pp94[20],pp93[22],pp92[24],pp91[26],pp90[28],pp89[30],pp88[32],pp87[34],pp86[36],pp85[38],pp84[40],pp83[42],pp82[44],pp81[46],pp82[46],pp83[46],pp84[46],pp85[46],pp86[46],pp87[46],pp88[46],pp89[46],pp90[46],pp91[46],pp92[46],pp93[46],pp94[46],pp95[46],pp96[46],pp97[46],pp98[46],pp99[46],pp137[9],pp139[8],pp141[7],pp143[6],pp145[5],pp147[4],pp149[3],pp151[2],pp153[1],pp155[0],s129[92],s130[92],s131[92],s132[92],s133[92],s134[92],s135[92],s136[92],s137[92],s138[92],s139[92],s140[92],s141[92],s142[92],s143[92],s144[92],s145[92],s146[92],s147[92],s148[92],s149[92],s150[92],s151[92],s152[92],s153[92],s154[92],s155[92],s156[92],s157[92],s158[92],s159[92],s160[92],s161[92],s162[92],s163[92],s164[92],s165[92],s166[92],s167[92],s168[92],s169[92],s170[92],s171[92],s172[92],s173[92],s174[92],s175[92],s176[92],s177[92],s10[68],s11[68],s12[68],s13[68],s14[68],s15[68],s16[68],s17[68],s18[68],s19[68],s20[68],s21[68],s22[68],s23[68],s24[68],s25[68],s26[68],s27[68],s28[68],s29[68],s30[68],s31[68],s32[68],s32[69],s32[70],s32[71],s32[72],s32[73],s32[74],s32[75],s32[76],s32[77],s32[78],s32[79],s32[80],s32[81],s32[82],s32[83],s32[84],s32[85],s32[86],s32[87],s32[88],s32[89],s32[90],s32[91],s32[92],s32[93],s32[94],s32[95],s32[96],s32[97],s9[121],s6[125],s3[129],s123[10],s121[13],s119[16],s117[19],s115[22],s113[25],s111[28],s109[31],s107[34],s105[37],s103[40],s101[43],s45[100],s44[102],s43[104],s42[106],s41[108],s40[110],s39[112],s38[114],s37[116],s36[118],s35[120],s34[122],s33[124],s32[126],s31[128],s30[130],s29[132],s28[134],s27[136],s26[138],s25[140],s24[142],s23[144],s22[146],s21[148],s20[150],s19[152],s18[154],s17[156],s16[158],s15[160],s14[162],s13[164],s12[166],s11[168],s10[170],s177[196],s176[198],s175[200],s174[202],s173[204],s172[206],s171[208],s170[210],s169[212],s168[214],s167[216],s166[218],s165[220],s164[222],s163[224],s162[226],s161[228],s160[230],s159[232],s158[234],s157[236],s156[238],s155[240],s154[242],s153[244],s152[246],s151[248],s150[250],s149[252],s148[254],s147[256],s146[258],s145[260],s144[262],s143[264],s142[266],s141[268],s140[270],s139[272],s138[274],s137[276],s136[278],s135[280],s134[282],s133[284],s132[286],s131[288],s130[290],s129[292],pp255[102],pp254[104],pp253[106],pp252[108],pp251[110],pp250[112],pp249[114],pp248[116],pp247[118],pp246[120],pp245[122],pp244[124],pp243[126],pp242[128],pp241[130],pp240[132],pp239[134],pp238[136],pp237[138],pp236[140],pp235[142],pp234[144],pp233[146],pp232[148],pp231[150],pp230[152],pp229[154],pp228[156],pp229[156],pp230[156],pp231[156],pp232[156],pp233[156],pp234[156],pp235[156],pp236[156],pp237[156],pp238[156],pp239[156],pp240[156],pp241[156],pp242[156]};
    CLA_286 KS_178(s178, c178, in178_1, in178_2);
    wire[283:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {pp95[19],pp94[21],pp93[23],pp92[25],pp91[27],pp90[29],pp89[31],pp88[33],pp87[35],pp86[37],pp85[39],pp84[41],pp83[43],pp82[45],pp83[45],pp84[45],pp85[45],pp86[45],pp87[45],pp88[45],pp89[45],pp90[45],pp91[45],pp92[45],pp93[45],pp94[45],pp95[45],pp96[45],pp97[45],pp98[45],pp99[45],pp136[9],pp138[8],pp140[7],pp142[6],pp144[5],pp146[4],pp148[3],pp150[2],pp152[1],pp154[0],s129[91],s130[91],s131[91],s132[91],s133[91],s134[91],s135[91],s136[91],s137[91],s138[91],s139[91],s140[91],s141[91],s142[91],s143[91],s144[91],s145[91],s146[91],s147[91],s148[91],s149[91],s150[91],s151[91],s152[91],s153[91],s154[91],s155[91],s156[91],s157[91],s158[91],s159[91],s160[91],s161[91],s162[91],s163[91],s164[91],s165[91],s166[91],s167[91],s168[91],s169[91],s170[91],s171[91],s172[91],s173[91],s174[91],s175[91],s176[91],s177[91],s178[91],s178[92],s178[93],s178[94],s178[95],s178[96],s178[97],s178[98],s178[99],s178[100],s178[101],s178[102],s178[103],s178[104],s178[105],s178[106],s178[107],s178[108],s178[109],s178[110],s178[111],s178[112],s178[113],s178[114],s178[115],s178[116],s178[117],s178[118],s178[119],s178[120],s178[121],s178[122],s178[123],s178[124],s178[125],s178[126],s178[127],s178[128],s178[129],s178[130],s178[131],s178[132],s178[133],s178[134],s178[135],s178[136],s178[137],s178[138],s178[139],s178[140],s178[141],s178[142],s178[143],s178[144],s178[145],s178[146],s178[147],s178[148],s178[149],s178[150],s178[151],s178[152],s178[153],s178[154],s178[155],s178[156],s178[157],s178[158],s178[159],s178[160],s178[161],s178[162],s178[163],s178[164],s178[165],s178[166],s178[167],s178[168],s178[169],s178[170],s178[171],s178[172],s178[173],s178[174],s178[175],s178[176],s178[177],s178[178],s178[179],s178[180],s178[181],s178[182],s178[183],s178[184],s178[185],s178[186],s178[187],s178[188],s178[189],s178[190],s178[191],s178[192],s178[193],s178[194],s178[195],s177[197],s176[199],s175[201],s174[203],s173[205],s172[207],s171[209],s170[211],s169[213],s168[215],s167[217],s166[219],s165[221],s164[223],s163[225],s162[227],s161[229],s160[231],s159[233],s158[235],s157[237],s156[239],s155[241],s154[243],s153[245],s152[247],s151[249],s150[251],s149[253],s148[255],s147[257],s146[259],s145[261],s144[263],s143[265],s142[267],s141[269],s140[271],s139[273],s138[275],s137[277],s136[279],s135[281],s134[283],s133[285],s132[287],s131[289],s130[291],s129[293],pp255[103],pp254[105],pp253[107],pp252[109],pp251[111],pp250[113],pp249[115],pp248[117],pp247[119],pp246[121],pp245[123],pp244[125],pp243[127],pp242[129],pp241[131],pp240[133],pp239[135],pp238[137],pp237[139],pp236[141],pp235[143],pp234[145],pp233[147],pp232[149],pp231[151],pp230[153],pp229[155],pp230[155],pp231[155],pp232[155],pp233[155],pp234[155],pp235[155],pp236[155],pp237[155],pp238[155],pp239[155],pp240[155],pp241[155],pp242[155]};
    assign in179_2 = {pp96[18],pp95[20],pp94[22],pp93[24],pp92[26],pp91[28],pp90[30],pp89[32],pp88[34],pp87[36],pp86[38],pp85[40],pp84[42],pp83[44],pp84[44],pp85[44],pp86[44],pp87[44],pp88[44],pp89[44],pp90[44],pp91[44],pp92[44],pp93[44],pp94[44],pp95[44],pp96[44],pp97[44],pp98[44],pp99[44],pp135[9],pp137[8],pp139[7],pp141[6],pp143[5],pp145[4],pp147[3],pp149[2],pp151[1],pp153[0],s129[90],s130[90],s131[90],s132[90],s133[90],s134[90],s135[90],s136[90],s137[90],s138[90],s139[90],s140[90],s141[90],s142[90],s143[90],s144[90],s145[90],s146[90],s147[90],s148[90],s149[90],s150[90],s151[90],s152[90],s153[90],s154[90],s155[90],s156[90],s157[90],s158[90],s159[90],s160[90],s161[90],s162[90],s163[90],s164[90],s165[90],s166[90],s167[90],s168[90],s169[90],s170[90],s171[90],s172[90],s173[90],s174[90],s175[90],s176[90],s177[90],s178[90],s10[67],s11[67],s12[67],s13[67],s14[67],s15[67],s16[67],s17[67],s18[67],s19[67],s20[67],s21[67],s22[67],s23[67],s24[67],s25[67],s26[67],s27[67],s28[67],s29[67],s30[67],s31[67],s32[67],s33[67],s33[68],s33[69],s33[70],s33[71],s33[72],s33[73],s33[74],s33[75],s33[76],s33[77],s33[78],s33[79],s33[80],s33[81],s33[82],s33[83],s33[84],s33[85],s33[86],s33[87],s33[88],s33[89],s33[90],s33[91],s33[92],s33[93],s33[94],s33[95],s33[96],s31[99],s7[124],s4[128],s1[132],s122[12],s120[15],s118[18],s116[21],s114[24],s112[27],s110[30],s108[33],s106[36],s104[39],s102[42],s100[45],s45[101],s44[103],s43[105],s42[107],s41[109],s40[111],s39[113],s38[115],s37[117],s36[119],s35[121],s34[123],s33[125],s32[127],s31[129],s30[131],s29[133],s28[135],s27[137],s26[139],s25[141],s24[143],s23[145],s22[147],s21[149],s20[151],s19[153],s18[155],s17[157],s16[159],s15[161],s14[163],s13[165],s12[167],s11[169],s10[171],s178[196],s177[198],s176[200],s175[202],s174[204],s173[206],s172[208],s171[210],s170[212],s169[214],s168[216],s167[218],s166[220],s165[222],s164[224],s163[226],s162[228],s161[230],s160[232],s159[234],s158[236],s157[238],s156[240],s155[242],s154[244],s153[246],s152[248],s151[250],s150[252],s149[254],s148[256],s147[258],s146[260],s145[262],s144[264],s143[266],s142[268],s141[270],s140[272],s139[274],s138[276],s137[278],s136[280],s135[282],s134[284],s133[286],s132[288],s131[290],s130[292],s129[294],pp255[104],pp254[106],pp253[108],pp252[110],pp251[112],pp250[114],pp249[116],pp248[118],pp247[120],pp246[122],pp245[124],pp244[126],pp243[128],pp242[130],pp241[132],pp240[134],pp239[136],pp238[138],pp237[140],pp236[142],pp235[144],pp234[146],pp233[148],pp232[150],pp231[152],pp230[154],pp231[154],pp232[154],pp233[154],pp234[154],pp235[154],pp236[154],pp237[154],pp238[154],pp239[154],pp240[154],pp241[154],pp242[154],pp243[154]};
    CLA_284 KS_179(s179, c179, in179_1, in179_2);
    wire[281:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {pp96[19],pp95[21],pp94[23],pp93[25],pp92[27],pp91[29],pp90[31],pp89[33],pp88[35],pp87[37],pp86[39],pp85[41],pp84[43],pp85[43],pp86[43],pp87[43],pp88[43],pp89[43],pp90[43],pp91[43],pp92[43],pp93[43],pp94[43],pp95[43],pp96[43],pp97[43],pp98[43],pp99[43],pp134[9],pp136[8],pp138[7],pp140[6],pp142[5],pp144[4],pp146[3],pp148[2],pp150[1],pp152[0],s129[89],s130[89],s131[89],s132[89],s133[89],s134[89],s135[89],s136[89],s137[89],s138[89],s139[89],s140[89],s141[89],s142[89],s143[89],s144[89],s145[89],s146[89],s147[89],s148[89],s149[89],s150[89],s151[89],s152[89],s153[89],s154[89],s155[89],s156[89],s157[89],s158[89],s159[89],s160[89],s161[89],s162[89],s163[89],s164[89],s165[89],s166[89],s167[89],s168[89],s169[89],s170[89],s171[89],s172[89],s173[89],s174[89],s175[89],s176[89],s177[89],s178[89],s179[89],s179[90],s179[91],s179[92],s179[93],s179[94],s179[95],s179[96],s179[97],s179[98],s179[99],s179[100],s179[101],s179[102],s179[103],s179[104],s179[105],s179[106],s179[107],s179[108],s179[109],s179[110],s179[111],s179[112],s179[113],s179[114],s179[115],s179[116],s179[117],s179[118],s179[119],s179[120],s179[121],s179[122],s179[123],s179[124],s179[125],s179[126],s179[127],s179[128],s179[129],s179[130],s179[131],s179[132],s179[133],s179[134],s179[135],s179[136],s179[137],s179[138],s179[139],s179[140],s179[141],s179[142],s179[143],s179[144],s179[145],s179[146],s179[147],s179[148],s179[149],s179[150],s179[151],s179[152],s179[153],s179[154],s179[155],s179[156],s179[157],s179[158],s179[159],s179[160],s179[161],s179[162],s179[163],s179[164],s179[165],s179[166],s179[167],s179[168],s179[169],s179[170],s179[171],s179[172],s179[173],s179[174],s179[175],s179[176],s179[177],s179[178],s179[179],s179[180],s179[181],s179[182],s179[183],s179[184],s179[185],s179[186],s179[187],s179[188],s179[189],s179[190],s179[191],s179[192],s179[193],s179[194],s179[195],s178[197],s177[199],s176[201],s175[203],s174[205],s173[207],s172[209],s171[211],s170[213],s169[215],s168[217],s167[219],s166[221],s165[223],s164[225],s163[227],s162[229],s161[231],s160[233],s159[235],s158[237],s157[239],s156[241],s155[243],s154[245],s153[247],s152[249],s151[251],s150[253],s149[255],s148[257],s147[259],s146[261],s145[263],s144[265],s143[267],s142[269],s141[271],s140[273],s139[275],s138[277],s137[279],s136[281],s135[283],s134[285],s133[287],s132[289],s131[291],s130[293],s129[295],pp255[105],pp254[107],pp253[109],pp252[111],pp251[113],pp250[115],pp249[117],pp248[119],pp247[121],pp246[123],pp245[125],pp244[127],pp243[129],pp242[131],pp241[133],pp240[135],pp239[137],pp238[139],pp237[141],pp236[143],pp235[145],pp234[147],pp233[149],pp232[151],pp231[153],pp232[153],pp233[153],pp234[153],pp235[153],pp236[153],pp237[153],pp238[153],pp239[153],pp240[153],pp241[153],pp242[153],pp243[153]};
    assign in180_2 = {pp97[18],pp96[20],pp95[22],pp94[24],pp93[26],pp92[28],pp91[30],pp90[32],pp89[34],pp88[36],pp87[38],pp86[40],pp85[42],pp86[42],pp87[42],pp88[42],pp89[42],pp90[42],pp91[42],pp92[42],pp93[42],pp94[42],pp95[42],pp96[42],pp97[42],pp98[42],pp99[42],pp133[9],pp135[8],pp137[7],pp139[6],pp141[5],pp143[4],pp145[3],pp147[2],pp149[1],pp151[0],s129[88],s130[88],s131[88],s132[88],s133[88],s134[88],s135[88],s136[88],s137[88],s138[88],s139[88],s140[88],s141[88],s142[88],s143[88],s144[88],s145[88],s146[88],s147[88],s148[88],s149[88],s150[88],s151[88],s152[88],s153[88],s154[88],s155[88],s156[88],s157[88],s158[88],s159[88],s160[88],s161[88],s162[88],s163[88],s164[88],s165[88],s166[88],s167[88],s168[88],s169[88],s170[88],s171[88],s172[88],s173[88],s174[88],s175[88],s176[88],s177[88],s178[88],s179[88],s10[66],s11[66],s12[66],s13[66],s14[66],s15[66],s16[66],s17[66],s18[66],s19[66],s20[66],s21[66],s22[66],s23[66],s24[66],s25[66],s26[66],s27[66],s28[66],s29[66],s30[66],s31[66],s32[66],s33[66],s34[66],s34[67],s34[68],s34[69],s34[70],s34[71],s34[72],s34[73],s34[74],s34[75],s34[76],s34[77],s34[78],s34[79],s34[80],s34[81],s34[82],s34[83],s34[84],s34[85],s34[86],s34[87],s34[88],s34[89],s34[90],s34[91],s34[92],s34[93],s34[94],s34[95],s32[98],s8[123],s5[127],s2[131],s123[11],s121[14],s119[17],s117[20],s115[23],s113[26],s111[29],s109[32],s107[35],s105[38],s103[41],s101[44],s46[100],s45[102],s44[104],s43[106],s42[108],s41[110],s40[112],s39[114],s38[116],s37[118],s36[120],s35[122],s34[124],s33[126],s32[128],s31[130],s30[132],s29[134],s28[136],s27[138],s26[140],s25[142],s24[144],s23[146],s22[148],s21[150],s20[152],s19[154],s18[156],s17[158],s16[160],s15[162],s14[164],s13[166],s12[168],s11[170],s10[172],s179[196],s178[198],s177[200],s176[202],s175[204],s174[206],s173[208],s172[210],s171[212],s170[214],s169[216],s168[218],s167[220],s166[222],s165[224],s164[226],s163[228],s162[230],s161[232],s160[234],s159[236],s158[238],s157[240],s156[242],s155[244],s154[246],s153[248],s152[250],s151[252],s150[254],s149[256],s148[258],s147[260],s146[262],s145[264],s144[266],s143[268],s142[270],s141[272],s140[274],s139[276],s138[278],s137[280],s136[282],s135[284],s134[286],s133[288],s132[290],s131[292],s130[294],s129[296],pp255[106],pp254[108],pp253[110],pp252[112],pp251[114],pp250[116],pp249[118],pp248[120],pp247[122],pp246[124],pp245[126],pp244[128],pp243[130],pp242[132],pp241[134],pp240[136],pp239[138],pp238[140],pp237[142],pp236[144],pp235[146],pp234[148],pp233[150],pp232[152],pp233[152],pp234[152],pp235[152],pp236[152],pp237[152],pp238[152],pp239[152],pp240[152],pp241[152],pp242[152],pp243[152],pp244[152]};
    CLA_282 KS_180(s180, c180, in180_1, in180_2);
    wire[279:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp97[19],pp96[21],pp95[23],pp94[25],pp93[27],pp92[29],pp91[31],pp90[33],pp89[35],pp88[37],pp87[39],pp86[41],pp87[41],pp88[41],pp89[41],pp90[41],pp91[41],pp92[41],pp93[41],pp94[41],pp95[41],pp96[41],pp97[41],pp98[41],pp99[41],pp132[9],pp134[8],pp136[7],pp138[6],pp140[5],pp142[4],pp144[3],pp146[2],pp148[1],pp150[0],s129[87],s130[87],s131[87],s132[87],s133[87],s134[87],s135[87],s136[87],s137[87],s138[87],s139[87],s140[87],s141[87],s142[87],s143[87],s144[87],s145[87],s146[87],s147[87],s148[87],s149[87],s150[87],s151[87],s152[87],s153[87],s154[87],s155[87],s156[87],s157[87],s158[87],s159[87],s160[87],s161[87],s162[87],s163[87],s164[87],s165[87],s166[87],s167[87],s168[87],s169[87],s170[87],s171[87],s172[87],s173[87],s174[87],s175[87],s176[87],s177[87],s178[87],s179[87],s180[87],s180[88],s180[89],s180[90],s180[91],s180[92],s180[93],s180[94],s180[95],s180[96],s180[97],s180[98],s180[99],s180[100],s180[101],s180[102],s180[103],s180[104],s180[105],s180[106],s180[107],s180[108],s180[109],s180[110],s180[111],s180[112],s180[113],s180[114],s180[115],s180[116],s180[117],s180[118],s180[119],s180[120],s180[121],s180[122],s180[123],s180[124],s180[125],s180[126],s180[127],s180[128],s180[129],s180[130],s180[131],s180[132],s180[133],s180[134],s180[135],s180[136],s180[137],s180[138],s180[139],s180[140],s180[141],s180[142],s180[143],s180[144],s180[145],s180[146],s180[147],s180[148],s180[149],s180[150],s180[151],s180[152],s180[153],s180[154],s180[155],s180[156],s180[157],s180[158],s180[159],s180[160],s180[161],s180[162],s180[163],s180[164],s180[165],s180[166],s180[167],s180[168],s180[169],s180[170],s180[171],s180[172],s180[173],s180[174],s180[175],s180[176],s180[177],s180[178],s180[179],s180[180],s180[181],s180[182],s180[183],s180[184],s180[185],s180[186],s180[187],s180[188],s180[189],s180[190],s180[191],s180[192],s180[193],s180[194],s180[195],s179[197],s178[199],s177[201],s176[203],s175[205],s174[207],s173[209],s172[211],s171[213],s170[215],s169[217],s168[219],s167[221],s166[223],s165[225],s164[227],s163[229],s162[231],s161[233],s160[235],s159[237],s158[239],s157[241],s156[243],s155[245],s154[247],s153[249],s152[251],s151[253],s150[255],s149[257],s148[259],s147[261],s146[263],s145[265],s144[267],s143[269],s142[271],s141[273],s140[275],s139[277],s138[279],s137[281],s136[283],s135[285],s134[287],s133[289],s132[291],s131[293],s130[295],s129[297],pp255[107],pp254[109],pp253[111],pp252[113],pp251[115],pp250[117],pp249[119],pp248[121],pp247[123],pp246[125],pp245[127],pp244[129],pp243[131],pp242[133],pp241[135],pp240[137],pp239[139],pp238[141],pp237[143],pp236[145],pp235[147],pp234[149],pp233[151],pp234[151],pp235[151],pp236[151],pp237[151],pp238[151],pp239[151],pp240[151],pp241[151],pp242[151],pp243[151],pp244[151]};
    assign in181_2 = {pp98[18],pp97[20],pp96[22],pp95[24],pp94[26],pp93[28],pp92[30],pp91[32],pp90[34],pp89[36],pp88[38],pp87[40],pp88[40],pp89[40],pp90[40],pp91[40],pp92[40],pp93[40],pp94[40],pp95[40],pp96[40],pp97[40],pp98[40],pp99[40],pp131[9],pp133[8],pp135[7],pp137[6],pp139[5],pp141[4],pp143[3],pp145[2],pp147[1],pp149[0],s129[86],s130[86],s131[86],s132[86],s133[86],s134[86],s135[86],s136[86],s137[86],s138[86],s139[86],s140[86],s141[86],s142[86],s143[86],s144[86],s145[86],s146[86],s147[86],s148[86],s149[86],s150[86],s151[86],s152[86],s153[86],s154[86],s155[86],s156[86],s157[86],s158[86],s159[86],s160[86],s161[86],s162[86],s163[86],s164[86],s165[86],s166[86],s167[86],s168[86],s169[86],s170[86],s171[86],s172[86],s173[86],s174[86],s175[86],s176[86],s177[86],s178[86],s179[86],s180[86],s10[65],s11[65],s12[65],s13[65],s14[65],s15[65],s16[65],s17[65],s18[65],s19[65],s20[65],s21[65],s22[65],s23[65],s24[65],s25[65],s26[65],s27[65],s28[65],s29[65],s30[65],s31[65],s32[65],s33[65],s34[65],s35[65],s35[66],s35[67],s35[68],s35[69],s35[70],s35[71],s35[72],s35[73],s35[74],s35[75],s35[76],s35[77],s35[78],s35[79],s35[80],s35[81],s35[82],s35[83],s35[84],s35[85],s35[86],s35[87],s35[88],s35[89],s35[90],s35[91],s35[92],s35[93],s35[94],s33[97],s9[122],s6[126],s3[130],s1[133],s122[13],s120[16],s118[19],s116[22],s114[25],s112[28],s110[31],s108[34],s106[37],s104[40],s102[43],s100[46],s46[101],s45[103],s44[105],s43[107],s42[109],s41[111],s40[113],s39[115],s38[117],s37[119],s36[121],s35[123],s34[125],s33[127],s32[129],s31[131],s30[133],s29[135],s28[137],s27[139],s26[141],s25[143],s24[145],s23[147],s22[149],s21[151],s20[153],s19[155],s18[157],s17[159],s16[161],s15[163],s14[165],s13[167],s12[169],s11[171],s10[173],s180[196],s179[198],s178[200],s177[202],s176[204],s175[206],s174[208],s173[210],s172[212],s171[214],s170[216],s169[218],s168[220],s167[222],s166[224],s165[226],s164[228],s163[230],s162[232],s161[234],s160[236],s159[238],s158[240],s157[242],s156[244],s155[246],s154[248],s153[250],s152[252],s151[254],s150[256],s149[258],s148[260],s147[262],s146[264],s145[266],s144[268],s143[270],s142[272],s141[274],s140[276],s139[278],s138[280],s137[282],s136[284],s135[286],s134[288],s133[290],s132[292],s131[294],s130[296],s129[298],pp255[108],pp254[110],pp253[112],pp252[114],pp251[116],pp250[118],pp249[120],pp248[122],pp247[124],pp246[126],pp245[128],pp244[130],pp243[132],pp242[134],pp241[136],pp240[138],pp239[140],pp238[142],pp237[144],pp236[146],pp235[148],pp234[150],pp235[150],pp236[150],pp237[150],pp238[150],pp239[150],pp240[150],pp241[150],pp242[150],pp243[150],pp244[150],pp245[150]};
    CLA_280 KS_181(s181, c181, in181_1, in181_2);
    wire[277:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp98[19],pp97[21],pp96[23],pp95[25],pp94[27],pp93[29],pp92[31],pp91[33],pp90[35],pp89[37],pp88[39],pp89[39],pp90[39],pp91[39],pp92[39],pp93[39],pp94[39],pp95[39],pp96[39],pp97[39],pp98[39],pp99[39],pp130[9],pp132[8],pp134[7],pp136[6],pp138[5],pp140[4],pp142[3],pp144[2],pp146[1],pp148[0],s129[85],s130[85],s131[85],s132[85],s133[85],s134[85],s135[85],s136[85],s137[85],s138[85],s139[85],s140[85],s141[85],s142[85],s143[85],s144[85],s145[85],s146[85],s147[85],s148[85],s149[85],s150[85],s151[85],s152[85],s153[85],s154[85],s155[85],s156[85],s157[85],s158[85],s159[85],s160[85],s161[85],s162[85],s163[85],s164[85],s165[85],s166[85],s167[85],s168[85],s169[85],s170[85],s171[85],s172[85],s173[85],s174[85],s175[85],s176[85],s177[85],s178[85],s179[85],s180[85],s181[85],s181[86],s181[87],s181[88],s181[89],s181[90],s181[91],s181[92],s181[93],s181[94],s181[95],s181[96],s181[97],s181[98],s181[99],s181[100],s181[101],s181[102],s181[103],s181[104],s181[105],s181[106],s181[107],s181[108],s181[109],s181[110],s181[111],s181[112],s181[113],s181[114],s181[115],s181[116],s181[117],s181[118],s181[119],s181[120],s181[121],s181[122],s181[123],s181[124],s181[125],s181[126],s181[127],s181[128],s181[129],s181[130],s181[131],s181[132],s181[133],s181[134],s181[135],s181[136],s181[137],s181[138],s181[139],s181[140],s181[141],s181[142],s181[143],s181[144],s181[145],s181[146],s181[147],s181[148],s181[149],s181[150],s181[151],s181[152],s181[153],s181[154],s181[155],s181[156],s181[157],s181[158],s181[159],s181[160],s181[161],s181[162],s181[163],s181[164],s181[165],s181[166],s181[167],s181[168],s181[169],s181[170],s181[171],s181[172],s181[173],s181[174],s181[175],s181[176],s181[177],s181[178],s181[179],s181[180],s181[181],s181[182],s181[183],s181[184],s181[185],s181[186],s181[187],s181[188],s181[189],s181[190],s181[191],s181[192],s181[193],s181[194],s181[195],s180[197],s179[199],s178[201],s177[203],s176[205],s175[207],s174[209],s173[211],s172[213],s171[215],s170[217],s169[219],s168[221],s167[223],s166[225],s165[227],s164[229],s163[231],s162[233],s161[235],s160[237],s159[239],s158[241],s157[243],s156[245],s155[247],s154[249],s153[251],s152[253],s151[255],s150[257],s149[259],s148[261],s147[263],s146[265],s145[267],s144[269],s143[271],s142[273],s141[275],s140[277],s139[279],s138[281],s137[283],s136[285],s135[287],s134[289],s133[291],s132[293],s131[295],s130[297],s129[299],pp255[109],pp254[111],pp253[113],pp252[115],pp251[117],pp250[119],pp249[121],pp248[123],pp247[125],pp246[127],pp245[129],pp244[131],pp243[133],pp242[135],pp241[137],pp240[139],pp239[141],pp238[143],pp237[145],pp236[147],pp235[149],pp236[149],pp237[149],pp238[149],pp239[149],pp240[149],pp241[149],pp242[149],pp243[149],pp244[149],pp245[149]};
    assign in182_2 = {pp99[18],pp98[20],pp97[22],pp96[24],pp95[26],pp94[28],pp93[30],pp92[32],pp91[34],pp90[36],pp89[38],pp90[38],pp91[38],pp92[38],pp93[38],pp94[38],pp95[38],pp96[38],pp97[38],pp98[38],pp99[38],pp129[9],pp131[8],pp133[7],pp135[6],pp137[5],pp139[4],pp141[3],pp143[2],pp145[1],pp147[0],s129[84],s130[84],s131[84],s132[84],s133[84],s134[84],s135[84],s136[84],s137[84],s138[84],s139[84],s140[84],s141[84],s142[84],s143[84],s144[84],s145[84],s146[84],s147[84],s148[84],s149[84],s150[84],s151[84],s152[84],s153[84],s154[84],s155[84],s156[84],s157[84],s158[84],s159[84],s160[84],s161[84],s162[84],s163[84],s164[84],s165[84],s166[84],s167[84],s168[84],s169[84],s170[84],s171[84],s172[84],s173[84],s174[84],s175[84],s176[84],s177[84],s178[84],s179[84],s180[84],s181[84],s10[64],s11[64],s12[64],s13[64],s14[64],s15[64],s16[64],s17[64],s18[64],s19[64],s20[64],s21[64],s22[64],s23[64],s24[64],s25[64],s26[64],s27[64],s28[64],s29[64],s30[64],s31[64],s32[64],s33[64],s34[64],s35[64],s36[64],s36[65],s36[66],s36[67],s36[68],s36[69],s36[70],s36[71],s36[72],s36[73],s36[74],s36[75],s36[76],s36[77],s36[78],s36[79],s36[80],s36[81],s36[82],s36[83],s36[84],s36[85],s36[86],s36[87],s36[88],s36[89],s36[90],s36[91],s36[92],s36[93],s34[96],s32[99],s7[125],s4[129],s2[132],s1[134],s121[15],s119[18],s117[21],s115[24],s113[27],s111[30],s109[33],s107[36],s105[39],s103[42],s101[45],s47[100],s46[102],s45[104],s44[106],s43[108],s42[110],s41[112],s40[114],s39[116],s38[118],s37[120],s36[122],s35[124],s34[126],s33[128],s32[130],s31[132],s30[134],s29[136],s28[138],s27[140],s26[142],s25[144],s24[146],s23[148],s22[150],s21[152],s20[154],s19[156],s18[158],s17[160],s16[162],s15[164],s14[166],s13[168],s12[170],s11[172],s10[174],s181[196],s180[198],s179[200],s178[202],s177[204],s176[206],s175[208],s174[210],s173[212],s172[214],s171[216],s170[218],s169[220],s168[222],s167[224],s166[226],s165[228],s164[230],s163[232],s162[234],s161[236],s160[238],s159[240],s158[242],s157[244],s156[246],s155[248],s154[250],s153[252],s152[254],s151[256],s150[258],s149[260],s148[262],s147[264],s146[266],s145[268],s144[270],s143[272],s142[274],s141[276],s140[278],s139[280],s138[282],s137[284],s136[286],s135[288],s134[290],s133[292],s132[294],s131[296],s130[298],s129[300],pp255[110],pp254[112],pp253[114],pp252[116],pp251[118],pp250[120],pp249[122],pp248[124],pp247[126],pp246[128],pp245[130],pp244[132],pp243[134],pp242[136],pp241[138],pp240[140],pp239[142],pp238[144],pp237[146],pp236[148],pp237[148],pp238[148],pp239[148],pp240[148],pp241[148],pp242[148],pp243[148],pp244[148],pp245[148],pp246[148]};
    CLA_278 KS_182(s182, c182, in182_1, in182_2);
    wire[275:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp99[19],pp98[21],pp97[23],pp96[25],pp95[27],pp94[29],pp93[31],pp92[33],pp91[35],pp90[37],pp91[37],pp92[37],pp93[37],pp94[37],pp95[37],pp96[37],pp97[37],pp98[37],pp99[37],pp128[9],pp130[8],pp132[7],pp134[6],pp136[5],pp138[4],pp140[3],pp142[2],pp144[1],pp146[0],s129[83],s130[83],s131[83],s132[83],s133[83],s134[83],s135[83],s136[83],s137[83],s138[83],s139[83],s140[83],s141[83],s142[83],s143[83],s144[83],s145[83],s146[83],s147[83],s148[83],s149[83],s150[83],s151[83],s152[83],s153[83],s154[83],s155[83],s156[83],s157[83],s158[83],s159[83],s160[83],s161[83],s162[83],s163[83],s164[83],s165[83],s166[83],s167[83],s168[83],s169[83],s170[83],s171[83],s172[83],s173[83],s174[83],s175[83],s176[83],s177[83],s178[83],s179[83],s180[83],s181[83],s182[83],s182[84],s182[85],s182[86],s182[87],s182[88],s182[89],s182[90],s182[91],s182[92],s182[93],s182[94],s182[95],s182[96],s182[97],s182[98],s182[99],s182[100],s182[101],s182[102],s182[103],s182[104],s182[105],s182[106],s182[107],s182[108],s182[109],s182[110],s182[111],s182[112],s182[113],s182[114],s182[115],s182[116],s182[117],s182[118],s182[119],s182[120],s182[121],s182[122],s182[123],s182[124],s182[125],s182[126],s182[127],s182[128],s182[129],s182[130],s182[131],s182[132],s182[133],s182[134],s182[135],s182[136],s182[137],s182[138],s182[139],s182[140],s182[141],s182[142],s182[143],s182[144],s182[145],s182[146],s182[147],s182[148],s182[149],s182[150],s182[151],s182[152],s182[153],s182[154],s182[155],s182[156],s182[157],s182[158],s182[159],s182[160],s182[161],s182[162],s182[163],s182[164],s182[165],s182[166],s182[167],s182[168],s182[169],s182[170],s182[171],s182[172],s182[173],s182[174],s182[175],s182[176],s182[177],s182[178],s182[179],s182[180],s182[181],s182[182],s182[183],s182[184],s182[185],s182[186],s182[187],s182[188],s182[189],s182[190],s182[191],s182[192],s182[193],s182[194],s182[195],s181[197],s180[199],s179[201],s178[203],s177[205],s176[207],s175[209],s174[211],s173[213],s172[215],s171[217],s170[219],s169[221],s168[223],s167[225],s166[227],s165[229],s164[231],s163[233],s162[235],s161[237],s160[239],s159[241],s158[243],s157[245],s156[247],s155[249],s154[251],s153[253],s152[255],s151[257],s150[259],s149[261],s148[263],s147[265],s146[267],s145[269],s144[271],s143[273],s142[275],s141[277],s140[279],s139[281],s138[283],s137[285],s136[287],s135[289],s134[291],s133[293],s132[295],s131[297],s130[299],s129[301],pp255[111],pp254[113],pp253[115],pp252[117],pp251[119],pp250[121],pp249[123],pp248[125],pp247[127],pp246[129],pp245[131],pp244[133],pp243[135],pp242[137],pp241[139],pp240[141],pp239[143],pp238[145],pp237[147],pp238[147],pp239[147],pp240[147],pp241[147],pp242[147],pp243[147],pp244[147],pp245[147],pp246[147]};
    assign in183_2 = {pp109[9],pp99[20],pp98[22],pp97[24],pp96[26],pp95[28],pp94[30],pp93[32],pp92[34],pp91[36],pp92[36],pp93[36],pp94[36],pp95[36],pp96[36],pp97[36],pp98[36],pp99[36],pp127[9],pp129[8],pp131[7],pp133[6],pp135[5],pp137[4],pp139[3],pp141[2],pp143[1],pp145[0],s129[82],s130[82],s131[82],s132[82],s133[82],s134[82],s135[82],s136[82],s137[82],s138[82],s139[82],s140[82],s141[82],s142[82],s143[82],s144[82],s145[82],s146[82],s147[82],s148[82],s149[82],s150[82],s151[82],s152[82],s153[82],s154[82],s155[82],s156[82],s157[82],s158[82],s159[82],s160[82],s161[82],s162[82],s163[82],s164[82],s165[82],s166[82],s167[82],s168[82],s169[82],s170[82],s171[82],s172[82],s173[82],s174[82],s175[82],s176[82],s177[82],s178[82],s179[82],s180[82],s181[82],s182[82],s10[63],s11[63],s12[63],s13[63],s14[63],s15[63],s16[63],s17[63],s18[63],s19[63],s20[63],s21[63],s22[63],s23[63],s24[63],s25[63],s26[63],s27[63],s28[63],s29[63],s30[63],s31[63],s32[63],s33[63],s34[63],s35[63],s36[63],s37[63],s37[64],s37[65],s37[66],s37[67],s37[68],s37[69],s37[70],s37[71],s37[72],s37[73],s37[74],s37[75],s37[76],s37[77],s37[78],s37[79],s37[80],s37[81],s37[82],s37[83],s37[84],s37[85],s37[86],s37[87],s37[88],s37[89],s37[90],s37[91],s37[92],s35[95],s33[98],s8[124],s5[128],s3[131],s2[133],s1[135],s120[17],s118[20],s116[23],s114[26],s112[29],s110[32],s108[35],s106[38],s104[41],s102[44],s100[47],s47[101],s46[103],s45[105],s44[107],s43[109],s42[111],s41[113],s40[115],s39[117],s38[119],s37[121],s36[123],s35[125],s34[127],s33[129],s32[131],s31[133],s30[135],s29[137],s28[139],s27[141],s26[143],s25[145],s24[147],s23[149],s22[151],s21[153],s20[155],s19[157],s18[159],s17[161],s16[163],s15[165],s14[167],s13[169],s12[171],s11[173],s10[175],s182[196],s181[198],s180[200],s179[202],s178[204],s177[206],s176[208],s175[210],s174[212],s173[214],s172[216],s171[218],s170[220],s169[222],s168[224],s167[226],s166[228],s165[230],s164[232],s163[234],s162[236],s161[238],s160[240],s159[242],s158[244],s157[246],s156[248],s155[250],s154[252],s153[254],s152[256],s151[258],s150[260],s149[262],s148[264],s147[266],s146[268],s145[270],s144[272],s143[274],s142[276],s141[278],s140[280],s139[282],s138[284],s137[286],s136[288],s135[290],s134[292],s133[294],s132[296],s131[298],s130[300],s129[302],pp255[112],pp254[114],pp253[116],pp252[118],pp251[120],pp250[122],pp249[124],pp248[126],pp247[128],pp246[130],pp245[132],pp244[134],pp243[136],pp242[138],pp241[140],pp240[142],pp239[144],pp238[146],pp239[146],pp240[146],pp241[146],pp242[146],pp243[146],pp244[146],pp245[146],pp246[146],pp247[146]};
    CLA_276 KS_183(s183, c183, in183_1, in183_2);
    wire[273:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp110[9],pp99[21],pp98[23],pp97[25],pp96[27],pp95[29],pp94[31],pp93[33],pp92[35],pp93[35],pp94[35],pp95[35],pp96[35],pp97[35],pp98[35],pp99[35],pp126[9],pp128[8],pp130[7],pp132[6],pp134[5],pp136[4],pp138[3],pp140[2],pp142[1],pp144[0],s129[81],s130[81],s131[81],s132[81],s133[81],s134[81],s135[81],s136[81],s137[81],s138[81],s139[81],s140[81],s141[81],s142[81],s143[81],s144[81],s145[81],s146[81],s147[81],s148[81],s149[81],s150[81],s151[81],s152[81],s153[81],s154[81],s155[81],s156[81],s157[81],s158[81],s159[81],s160[81],s161[81],s162[81],s163[81],s164[81],s165[81],s166[81],s167[81],s168[81],s169[81],s170[81],s171[81],s172[81],s173[81],s174[81],s175[81],s176[81],s177[81],s178[81],s179[81],s180[81],s181[81],s182[81],s183[81],s183[82],s183[83],s183[84],s183[85],s183[86],s183[87],s183[88],s183[89],s183[90],s183[91],s183[92],s183[93],s183[94],s183[95],s183[96],s183[97],s183[98],s183[99],s183[100],s183[101],s183[102],s183[103],s183[104],s183[105],s183[106],s183[107],s183[108],s183[109],s183[110],s183[111],s183[112],s183[113],s183[114],s183[115],s183[116],s183[117],s183[118],s183[119],s183[120],s183[121],s183[122],s183[123],s183[124],s183[125],s183[126],s183[127],s183[128],s183[129],s183[130],s183[131],s183[132],s183[133],s183[134],s183[135],s183[136],s183[137],s183[138],s183[139],s183[140],s183[141],s183[142],s183[143],s183[144],s183[145],s183[146],s183[147],s183[148],s183[149],s183[150],s183[151],s183[152],s183[153],s183[154],s183[155],s183[156],s183[157],s183[158],s183[159],s183[160],s183[161],s183[162],s183[163],s183[164],s183[165],s183[166],s183[167],s183[168],s183[169],s183[170],s183[171],s183[172],s183[173],s183[174],s183[175],s183[176],s183[177],s183[178],s183[179],s183[180],s183[181],s183[182],s183[183],s183[184],s183[185],s183[186],s183[187],s183[188],s183[189],s183[190],s183[191],s183[192],s183[193],s183[194],s183[195],s182[197],s181[199],s180[201],s179[203],s178[205],s177[207],s176[209],s175[211],s174[213],s173[215],s172[217],s171[219],s170[221],s169[223],s168[225],s167[227],s166[229],s165[231],s164[233],s163[235],s162[237],s161[239],s160[241],s159[243],s158[245],s157[247],s156[249],s155[251],s154[253],s153[255],s152[257],s151[259],s150[261],s149[263],s148[265],s147[267],s146[269],s145[271],s144[273],s143[275],s142[277],s141[279],s140[281],s139[283],s138[285],s137[287],s136[289],s135[291],s134[293],s133[295],s132[297],s131[299],s130[301],s129[303],pp255[113],pp254[115],pp253[117],pp252[119],pp251[121],pp250[123],pp249[125],pp248[127],pp247[129],pp246[131],pp245[133],pp244[135],pp243[137],pp242[139],pp241[141],pp240[143],pp239[145],pp240[145],pp241[145],pp242[145],pp243[145],pp244[145],pp245[145],pp246[145],pp247[145]};
    assign in184_2 = {pp111[8],pp111[9],pp99[22],pp98[24],pp97[26],pp96[28],pp95[30],pp94[32],pp93[34],pp94[34],pp95[34],pp96[34],pp97[34],pp98[34],pp99[34],pp125[9],pp127[8],pp129[7],pp131[6],pp133[5],pp135[4],pp137[3],pp139[2],pp141[1],pp143[0],s129[80],s130[80],s131[80],s132[80],s133[80],s134[80],s135[80],s136[80],s137[80],s138[80],s139[80],s140[80],s141[80],s142[80],s143[80],s144[80],s145[80],s146[80],s147[80],s148[80],s149[80],s150[80],s151[80],s152[80],s153[80],s154[80],s155[80],s156[80],s157[80],s158[80],s159[80],s160[80],s161[80],s162[80],s163[80],s164[80],s165[80],s166[80],s167[80],s168[80],s169[80],s170[80],s171[80],s172[80],s173[80],s174[80],s175[80],s176[80],s177[80],s178[80],s179[80],s180[80],s181[80],s182[80],s183[80],s10[62],s11[62],s12[62],s13[62],s14[62],s15[62],s16[62],s17[62],s18[62],s19[62],s20[62],s21[62],s22[62],s23[62],s24[62],s25[62],s26[62],s27[62],s28[62],s29[62],s30[62],s31[62],s32[62],s33[62],s34[62],s35[62],s36[62],s37[62],s38[62],s38[63],s38[64],s38[65],s38[66],s38[67],s38[68],s38[69],s38[70],s38[71],s38[72],s38[73],s38[74],s38[75],s38[76],s38[77],s38[78],s38[79],s38[80],s38[81],s38[82],s38[83],s38[84],s38[85],s38[86],s38[87],s38[88],s38[89],s38[90],s38[91],s36[94],s34[97],s9[123],s6[127],s4[130],s3[132],s2[134],s1[136],s119[19],s117[22],s115[25],s113[28],s111[31],s109[34],s107[37],s105[40],s103[43],s101[46],s48[100],s47[102],s46[104],s45[106],s44[108],s43[110],s42[112],s41[114],s40[116],s39[118],s38[120],s37[122],s36[124],s35[126],s34[128],s33[130],s32[132],s31[134],s30[136],s29[138],s28[140],s27[142],s26[144],s25[146],s24[148],s23[150],s22[152],s21[154],s20[156],s19[158],s18[160],s17[162],s16[164],s15[166],s14[168],s13[170],s12[172],s11[174],s10[176],s183[196],s182[198],s181[200],s180[202],s179[204],s178[206],s177[208],s176[210],s175[212],s174[214],s173[216],s172[218],s171[220],s170[222],s169[224],s168[226],s167[228],s166[230],s165[232],s164[234],s163[236],s162[238],s161[240],s160[242],s159[244],s158[246],s157[248],s156[250],s155[252],s154[254],s153[256],s152[258],s151[260],s150[262],s149[264],s148[266],s147[268],s146[270],s145[272],s144[274],s143[276],s142[278],s141[280],s140[282],s139[284],s138[286],s137[288],s136[290],s135[292],s134[294],s133[296],s132[298],s131[300],s130[302],s129[304],pp255[114],pp254[116],pp253[118],pp252[120],pp251[122],pp250[124],pp249[126],pp248[128],pp247[130],pp246[132],pp245[134],pp244[136],pp243[138],pp242[140],pp241[142],pp240[144],pp241[144],pp242[144],pp243[144],pp244[144],pp245[144],pp246[144],pp247[144],pp248[144]};
    CLA_274 KS_184(s184, c184, in184_1, in184_2);
    wire[271:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {pp112[8],pp112[9],pp99[23],pp98[25],pp97[27],pp96[29],pp95[31],pp94[33],pp95[33],pp96[33],pp97[33],pp98[33],pp99[33],pp124[9],pp126[8],pp128[7],pp130[6],pp132[5],pp134[4],pp136[3],pp138[2],pp140[1],pp142[0],s129[79],s130[79],s131[79],s132[79],s133[79],s134[79],s135[79],s136[79],s137[79],s138[79],s139[79],s140[79],s141[79],s142[79],s143[79],s144[79],s145[79],s146[79],s147[79],s148[79],s149[79],s150[79],s151[79],s152[79],s153[79],s154[79],s155[79],s156[79],s157[79],s158[79],s159[79],s160[79],s161[79],s162[79],s163[79],s164[79],s165[79],s166[79],s167[79],s168[79],s169[79],s170[79],s171[79],s172[79],s173[79],s174[79],s175[79],s176[79],s177[79],s178[79],s179[79],s180[79],s181[79],s182[79],s183[79],s184[79],s184[80],s184[81],s184[82],s184[83],s184[84],s184[85],s184[86],s184[87],s184[88],s184[89],s184[90],s184[91],s184[92],s184[93],s184[94],s184[95],s184[96],s184[97],s184[98],s184[99],s184[100],s184[101],s184[102],s184[103],s184[104],s184[105],s184[106],s184[107],s184[108],s184[109],s184[110],s184[111],s184[112],s184[113],s184[114],s184[115],s184[116],s184[117],s184[118],s184[119],s184[120],s184[121],s184[122],s184[123],s184[124],s184[125],s184[126],s184[127],s184[128],s184[129],s184[130],s184[131],s184[132],s184[133],s184[134],s184[135],s184[136],s184[137],s184[138],s184[139],s184[140],s184[141],s184[142],s184[143],s184[144],s184[145],s184[146],s184[147],s184[148],s184[149],s184[150],s184[151],s184[152],s184[153],s184[154],s184[155],s184[156],s184[157],s184[158],s184[159],s184[160],s184[161],s184[162],s184[163],s184[164],s184[165],s184[166],s184[167],s184[168],s184[169],s184[170],s184[171],s184[172],s184[173],s184[174],s184[175],s184[176],s184[177],s184[178],s184[179],s184[180],s184[181],s184[182],s184[183],s184[184],s184[185],s184[186],s184[187],s184[188],s184[189],s184[190],s184[191],s184[192],s184[193],s184[194],s184[195],s183[197],s182[199],s181[201],s180[203],s179[205],s178[207],s177[209],s176[211],s175[213],s174[215],s173[217],s172[219],s171[221],s170[223],s169[225],s168[227],s167[229],s166[231],s165[233],s164[235],s163[237],s162[239],s161[241],s160[243],s159[245],s158[247],s157[249],s156[251],s155[253],s154[255],s153[257],s152[259],s151[261],s150[263],s149[265],s148[267],s147[269],s146[271],s145[273],s144[275],s143[277],s142[279],s141[281],s140[283],s139[285],s138[287],s137[289],s136[291],s135[293],s134[295],s133[297],s132[299],s131[301],s130[303],s129[305],pp255[115],pp254[117],pp253[119],pp252[121],pp251[123],pp250[125],pp249[127],pp248[129],pp247[131],pp246[133],pp245[135],pp244[137],pp243[139],pp242[141],pp241[143],pp242[143],pp243[143],pp244[143],pp245[143],pp246[143],pp247[143],pp248[143]};
    assign in185_2 = {pp113[7],pp113[8],pp113[9],pp99[24],pp98[26],pp97[28],pp96[30],pp95[32],pp96[32],pp97[32],pp98[32],pp99[32],pp123[9],pp125[8],pp127[7],pp129[6],pp131[5],pp133[4],pp135[3],pp137[2],pp139[1],pp141[0],s129[78],s130[78],s131[78],s132[78],s133[78],s134[78],s135[78],s136[78],s137[78],s138[78],s139[78],s140[78],s141[78],s142[78],s143[78],s144[78],s145[78],s146[78],s147[78],s148[78],s149[78],s150[78],s151[78],s152[78],s153[78],s154[78],s155[78],s156[78],s157[78],s158[78],s159[78],s160[78],s161[78],s162[78],s163[78],s164[78],s165[78],s166[78],s167[78],s168[78],s169[78],s170[78],s171[78],s172[78],s173[78],s174[78],s175[78],s176[78],s177[78],s178[78],s179[78],s180[78],s181[78],s182[78],s183[78],s184[78],s10[61],s11[61],s12[61],s13[61],s14[61],s15[61],s16[61],s17[61],s18[61],s19[61],s20[61],s21[61],s22[61],s23[61],s24[61],s25[61],s26[61],s27[61],s28[61],s29[61],s30[61],s31[61],s32[61],s33[61],s34[61],s35[61],s36[61],s37[61],s38[61],s39[61],s39[62],s39[63],s39[64],s39[65],s39[66],s39[67],s39[68],s39[69],s39[70],s39[71],s39[72],s39[73],s39[74],s39[75],s39[76],s39[77],s39[78],s39[79],s39[80],s39[81],s39[82],s39[83],s39[84],s39[85],s39[86],s39[87],s39[88],s39[89],s39[90],s37[93],s35[96],s33[99],s7[126],s5[129],s4[131],s3[133],s2[135],s1[137],s118[21],s116[24],s114[27],s112[30],s110[33],s108[36],s106[39],s104[42],s102[45],s100[48],s48[101],s47[103],s46[105],s45[107],s44[109],s43[111],s42[113],s41[115],s40[117],s39[119],s38[121],s37[123],s36[125],s35[127],s34[129],s33[131],s32[133],s31[135],s30[137],s29[139],s28[141],s27[143],s26[145],s25[147],s24[149],s23[151],s22[153],s21[155],s20[157],s19[159],s18[161],s17[163],s16[165],s15[167],s14[169],s13[171],s12[173],s11[175],s10[177],s184[196],s183[198],s182[200],s181[202],s180[204],s179[206],s178[208],s177[210],s176[212],s175[214],s174[216],s173[218],s172[220],s171[222],s170[224],s169[226],s168[228],s167[230],s166[232],s165[234],s164[236],s163[238],s162[240],s161[242],s160[244],s159[246],s158[248],s157[250],s156[252],s155[254],s154[256],s153[258],s152[260],s151[262],s150[264],s149[266],s148[268],s147[270],s146[272],s145[274],s144[276],s143[278],s142[280],s141[282],s140[284],s139[286],s138[288],s137[290],s136[292],s135[294],s134[296],s133[298],s132[300],s131[302],s130[304],s129[306],pp255[116],pp254[118],pp253[120],pp252[122],pp251[124],pp250[126],pp249[128],pp248[130],pp247[132],pp246[134],pp245[136],pp244[138],pp243[140],pp242[142],pp243[142],pp244[142],pp245[142],pp246[142],pp247[142],pp248[142],pp249[142]};
    CLA_272 KS_185(s185, c185, in185_1, in185_2);
    wire[269:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {pp114[7],pp114[8],pp114[9],pp99[25],pp98[27],pp97[29],pp96[31],pp97[31],pp98[31],pp99[31],pp122[9],pp124[8],pp126[7],pp128[6],pp130[5],pp132[4],pp134[3],pp136[2],pp138[1],pp140[0],s129[77],s130[77],s131[77],s132[77],s133[77],s134[77],s135[77],s136[77],s137[77],s138[77],s139[77],s140[77],s141[77],s142[77],s143[77],s144[77],s145[77],s146[77],s147[77],s148[77],s149[77],s150[77],s151[77],s152[77],s153[77],s154[77],s155[77],s156[77],s157[77],s158[77],s159[77],s160[77],s161[77],s162[77],s163[77],s164[77],s165[77],s166[77],s167[77],s168[77],s169[77],s170[77],s171[77],s172[77],s173[77],s174[77],s175[77],s176[77],s177[77],s178[77],s179[77],s180[77],s181[77],s182[77],s183[77],s184[77],s185[77],s185[78],s185[79],s185[80],s185[81],s185[82],s185[83],s185[84],s185[85],s185[86],s185[87],s185[88],s185[89],s185[90],s185[91],s185[92],s185[93],s185[94],s185[95],s185[96],s185[97],s185[98],s185[99],s185[100],s185[101],s185[102],s185[103],s185[104],s185[105],s185[106],s185[107],s185[108],s185[109],s185[110],s185[111],s185[112],s185[113],s185[114],s185[115],s185[116],s185[117],s185[118],s185[119],s185[120],s185[121],s185[122],s185[123],s185[124],s185[125],s185[126],s185[127],s185[128],s185[129],s185[130],s185[131],s185[132],s185[133],s185[134],s185[135],s185[136],s185[137],s185[138],s185[139],s185[140],s185[141],s185[142],s185[143],s185[144],s185[145],s185[146],s185[147],s185[148],s185[149],s185[150],s185[151],s185[152],s185[153],s185[154],s185[155],s185[156],s185[157],s185[158],s185[159],s185[160],s185[161],s185[162],s185[163],s185[164],s185[165],s185[166],s185[167],s185[168],s185[169],s185[170],s185[171],s185[172],s185[173],s185[174],s185[175],s185[176],s185[177],s185[178],s185[179],s185[180],s185[181],s185[182],s185[183],s185[184],s185[185],s185[186],s185[187],s185[188],s185[189],s185[190],s185[191],s185[192],s185[193],s185[194],s185[195],s184[197],s183[199],s182[201],s181[203],s180[205],s179[207],s178[209],s177[211],s176[213],s175[215],s174[217],s173[219],s172[221],s171[223],s170[225],s169[227],s168[229],s167[231],s166[233],s165[235],s164[237],s163[239],s162[241],s161[243],s160[245],s159[247],s158[249],s157[251],s156[253],s155[255],s154[257],s153[259],s152[261],s151[263],s150[265],s149[267],s148[269],s147[271],s146[273],s145[275],s144[277],s143[279],s142[281],s141[283],s140[285],s139[287],s138[289],s137[291],s136[293],s135[295],s134[297],s133[299],s132[301],s131[303],s130[305],s129[307],pp255[117],pp254[119],pp253[121],pp252[123],pp251[125],pp250[127],pp249[129],pp248[131],pp247[133],pp246[135],pp245[137],pp244[139],pp243[141],pp244[141],pp245[141],pp246[141],pp247[141],pp248[141],pp249[141]};
    assign in186_2 = {pp115[6],pp115[7],pp115[8],pp115[9],pp99[26],pp98[28],pp97[30],pp98[30],pp99[30],pp121[9],pp123[8],pp125[7],pp127[6],pp129[5],pp131[4],pp133[3],pp135[2],pp137[1],pp139[0],s129[76],s130[76],s131[76],s132[76],s133[76],s134[76],s135[76],s136[76],s137[76],s138[76],s139[76],s140[76],s141[76],s142[76],s143[76],s144[76],s145[76],s146[76],s147[76],s148[76],s149[76],s150[76],s151[76],s152[76],s153[76],s154[76],s155[76],s156[76],s157[76],s158[76],s159[76],s160[76],s161[76],s162[76],s163[76],s164[76],s165[76],s166[76],s167[76],s168[76],s169[76],s170[76],s171[76],s172[76],s173[76],s174[76],s175[76],s176[76],s177[76],s178[76],s179[76],s180[76],s181[76],s182[76],s183[76],s184[76],s185[76],s10[60],s11[60],s12[60],s13[60],s14[60],s15[60],s16[60],s17[60],s18[60],s19[60],s20[60],s21[60],s22[60],s23[60],s24[60],s25[60],s26[60],s27[60],s28[60],s29[60],s30[60],s31[60],s32[60],s33[60],s34[60],s35[60],s36[60],s37[60],s38[60],s39[60],s40[60],s40[61],s40[62],s40[63],s40[64],s40[65],s40[66],s40[67],s40[68],s40[69],s40[70],s40[71],s40[72],s40[73],s40[74],s40[75],s40[76],s40[77],s40[78],s40[79],s40[80],s40[81],s40[82],s40[83],s40[84],s40[85],s40[86],s40[87],s40[88],s40[89],s38[92],s36[95],s34[98],s8[125],s6[128],s5[130],s4[132],s3[134],s2[136],s1[138],s117[23],s115[26],s113[29],s111[32],s109[35],s107[38],s105[41],s103[44],s101[47],s49[100],s48[102],s47[104],s46[106],s45[108],s44[110],s43[112],s42[114],s41[116],s40[118],s39[120],s38[122],s37[124],s36[126],s35[128],s34[130],s33[132],s32[134],s31[136],s30[138],s29[140],s28[142],s27[144],s26[146],s25[148],s24[150],s23[152],s22[154],s21[156],s20[158],s19[160],s18[162],s17[164],s16[166],s15[168],s14[170],s13[172],s12[174],s11[176],s10[178],s185[196],s184[198],s183[200],s182[202],s181[204],s180[206],s179[208],s178[210],s177[212],s176[214],s175[216],s174[218],s173[220],s172[222],s171[224],s170[226],s169[228],s168[230],s167[232],s166[234],s165[236],s164[238],s163[240],s162[242],s161[244],s160[246],s159[248],s158[250],s157[252],s156[254],s155[256],s154[258],s153[260],s152[262],s151[264],s150[266],s149[268],s148[270],s147[272],s146[274],s145[276],s144[278],s143[280],s142[282],s141[284],s140[286],s139[288],s138[290],s137[292],s136[294],s135[296],s134[298],s133[300],s132[302],s131[304],s130[306],s129[308],pp255[118],pp254[120],pp253[122],pp252[124],pp251[126],pp250[128],pp249[130],pp248[132],pp247[134],pp246[136],pp245[138],pp244[140],pp245[140],pp246[140],pp247[140],pp248[140],pp249[140],pp250[140]};
    CLA_270 KS_186(s186, c186, in186_1, in186_2);
    wire[267:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {pp116[6],pp116[7],pp116[8],pp116[9],pp99[27],pp98[29],pp99[29],pp120[9],pp122[8],pp124[7],pp126[6],pp128[5],pp130[4],pp132[3],pp134[2],pp136[1],pp138[0],s129[75],s130[75],s131[75],s132[75],s133[75],s134[75],s135[75],s136[75],s137[75],s138[75],s139[75],s140[75],s141[75],s142[75],s143[75],s144[75],s145[75],s146[75],s147[75],s148[75],s149[75],s150[75],s151[75],s152[75],s153[75],s154[75],s155[75],s156[75],s157[75],s158[75],s159[75],s160[75],s161[75],s162[75],s163[75],s164[75],s165[75],s166[75],s167[75],s168[75],s169[75],s170[75],s171[75],s172[75],s173[75],s174[75],s175[75],s176[75],s177[75],s178[75],s179[75],s180[75],s181[75],s182[75],s183[75],s184[75],s185[75],s186[75],s186[76],s186[77],s186[78],s186[79],s186[80],s186[81],s186[82],s186[83],s186[84],s186[85],s186[86],s186[87],s186[88],s186[89],s186[90],s186[91],s186[92],s186[93],s186[94],s186[95],s186[96],s186[97],s186[98],s186[99],s186[100],s186[101],s186[102],s186[103],s186[104],s186[105],s186[106],s186[107],s186[108],s186[109],s186[110],s186[111],s186[112],s186[113],s186[114],s186[115],s186[116],s186[117],s186[118],s186[119],s186[120],s186[121],s186[122],s186[123],s186[124],s186[125],s186[126],s186[127],s186[128],s186[129],s186[130],s186[131],s186[132],s186[133],s186[134],s186[135],s186[136],s186[137],s186[138],s186[139],s186[140],s186[141],s186[142],s186[143],s186[144],s186[145],s186[146],s186[147],s186[148],s186[149],s186[150],s186[151],s186[152],s186[153],s186[154],s186[155],s186[156],s186[157],s186[158],s186[159],s186[160],s186[161],s186[162],s186[163],s186[164],s186[165],s186[166],s186[167],s186[168],s186[169],s186[170],s186[171],s186[172],s186[173],s186[174],s186[175],s186[176],s186[177],s186[178],s186[179],s186[180],s186[181],s186[182],s186[183],s186[184],s186[185],s186[186],s186[187],s186[188],s186[189],s186[190],s186[191],s186[192],s186[193],s186[194],s186[195],s185[197],s184[199],s183[201],s182[203],s181[205],s180[207],s179[209],s178[211],s177[213],s176[215],s175[217],s174[219],s173[221],s172[223],s171[225],s170[227],s169[229],s168[231],s167[233],s166[235],s165[237],s164[239],s163[241],s162[243],s161[245],s160[247],s159[249],s158[251],s157[253],s156[255],s155[257],s154[259],s153[261],s152[263],s151[265],s150[267],s149[269],s148[271],s147[273],s146[275],s145[277],s144[279],s143[281],s142[283],s141[285],s140[287],s139[289],s138[291],s137[293],s136[295],s135[297],s134[299],s133[301],s132[303],s131[305],s130[307],s129[309],pp255[119],pp254[121],pp253[123],pp252[125],pp251[127],pp250[129],pp249[131],pp248[133],pp247[135],pp246[137],pp245[139],pp246[139],pp247[139],pp248[139],pp249[139],pp250[139]};
    assign in187_2 = {pp117[5],pp117[6],pp117[7],pp117[8],pp117[9],pp99[28],pp119[9],pp121[8],pp123[7],pp125[6],pp127[5],pp129[4],pp131[3],pp133[2],pp135[1],pp137[0],s129[74],s130[74],s131[74],s132[74],s133[74],s134[74],s135[74],s136[74],s137[74],s138[74],s139[74],s140[74],s141[74],s142[74],s143[74],s144[74],s145[74],s146[74],s147[74],s148[74],s149[74],s150[74],s151[74],s152[74],s153[74],s154[74],s155[74],s156[74],s157[74],s158[74],s159[74],s160[74],s161[74],s162[74],s163[74],s164[74],s165[74],s166[74],s167[74],s168[74],s169[74],s170[74],s171[74],s172[74],s173[74],s174[74],s175[74],s176[74],s177[74],s178[74],s179[74],s180[74],s181[74],s182[74],s183[74],s184[74],s185[74],s186[74],s10[59],s11[59],s12[59],s13[59],s14[59],s15[59],s16[59],s17[59],s18[59],s19[59],s20[59],s21[59],s22[59],s23[59],s24[59],s25[59],s26[59],s27[59],s28[59],s29[59],s30[59],s31[59],s32[59],s33[59],s34[59],s35[59],s36[59],s37[59],s38[59],s39[59],s40[59],s41[59],s41[60],s41[61],s41[62],s41[63],s41[64],s41[65],s41[66],s41[67],s41[68],s41[69],s41[70],s41[71],s41[72],s41[73],s41[74],s41[75],s41[76],s41[77],s41[78],s41[79],s41[80],s41[81],s41[82],s41[83],s41[84],s41[85],s41[86],s41[87],s41[88],s39[91],s37[94],s35[97],s9[124],s7[127],s6[129],s5[131],s4[133],s3[135],s2[137],s1[139],s116[25],s114[28],s112[31],s110[34],s108[37],s106[40],s104[43],s102[46],s100[49],s49[101],s48[103],s47[105],s46[107],s45[109],s44[111],s43[113],s42[115],s41[117],s40[119],s39[121],s38[123],s37[125],s36[127],s35[129],s34[131],s33[133],s32[135],s31[137],s30[139],s29[141],s28[143],s27[145],s26[147],s25[149],s24[151],s23[153],s22[155],s21[157],s20[159],s19[161],s18[163],s17[165],s16[167],s15[169],s14[171],s13[173],s12[175],s11[177],s10[179],s186[196],s185[198],s184[200],s183[202],s182[204],s181[206],s180[208],s179[210],s178[212],s177[214],s176[216],s175[218],s174[220],s173[222],s172[224],s171[226],s170[228],s169[230],s168[232],s167[234],s166[236],s165[238],s164[240],s163[242],s162[244],s161[246],s160[248],s159[250],s158[252],s157[254],s156[256],s155[258],s154[260],s153[262],s152[264],s151[266],s150[268],s149[270],s148[272],s147[274],s146[276],s145[278],s144[280],s143[282],s142[284],s141[286],s140[288],s139[290],s138[292],s137[294],s136[296],s135[298],s134[300],s133[302],s132[304],s131[306],s130[308],s129[310],pp255[120],pp254[122],pp253[124],pp252[126],pp251[128],pp250[130],pp249[132],pp248[134],pp247[136],pp246[138],pp247[138],pp248[138],pp249[138],pp250[138],pp251[138]};
    CLA_268 KS_187(s187, c187, in187_1, in187_2);
    wire[265:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp118[5],pp118[6],pp118[7],pp118[8],pp118[9],pp120[8],pp122[7],pp124[6],pp126[5],pp128[4],pp130[3],pp132[2],pp134[1],pp136[0],s129[73],s130[73],s131[73],s132[73],s133[73],s134[73],s135[73],s136[73],s137[73],s138[73],s139[73],s140[73],s141[73],s142[73],s143[73],s144[73],s145[73],s146[73],s147[73],s148[73],s149[73],s150[73],s151[73],s152[73],s153[73],s154[73],s155[73],s156[73],s157[73],s158[73],s159[73],s160[73],s161[73],s162[73],s163[73],s164[73],s165[73],s166[73],s167[73],s168[73],s169[73],s170[73],s171[73],s172[73],s173[73],s174[73],s175[73],s176[73],s177[73],s178[73],s179[73],s180[73],s181[73],s182[73],s183[73],s184[73],s185[73],s186[73],s187[73],s187[74],s187[75],s187[76],s187[77],s187[78],s187[79],s187[80],s187[81],s187[82],s187[83],s187[84],s187[85],s187[86],s187[87],s187[88],s187[89],s187[90],s187[91],s187[92],s187[93],s187[94],s187[95],s187[96],s187[97],s187[98],s187[99],s187[100],s187[101],s187[102],s187[103],s187[104],s187[105],s187[106],s187[107],s187[108],s187[109],s187[110],s187[111],s187[112],s187[113],s187[114],s187[115],s187[116],s187[117],s187[118],s187[119],s187[120],s187[121],s187[122],s187[123],s187[124],s187[125],s187[126],s187[127],s187[128],s187[129],s187[130],s187[131],s187[132],s187[133],s187[134],s187[135],s187[136],s187[137],s187[138],s187[139],s187[140],s187[141],s187[142],s187[143],s187[144],s187[145],s187[146],s187[147],s187[148],s187[149],s187[150],s187[151],s187[152],s187[153],s187[154],s187[155],s187[156],s187[157],s187[158],s187[159],s187[160],s187[161],s187[162],s187[163],s187[164],s187[165],s187[166],s187[167],s187[168],s187[169],s187[170],s187[171],s187[172],s187[173],s187[174],s187[175],s187[176],s187[177],s187[178],s187[179],s187[180],s187[181],s187[182],s187[183],s187[184],s187[185],s187[186],s187[187],s187[188],s187[189],s187[190],s187[191],s187[192],s187[193],s187[194],s187[195],s186[197],s185[199],s184[201],s183[203],s182[205],s181[207],s180[209],s179[211],s178[213],s177[215],s176[217],s175[219],s174[221],s173[223],s172[225],s171[227],s170[229],s169[231],s168[233],s167[235],s166[237],s165[239],s164[241],s163[243],s162[245],s161[247],s160[249],s159[251],s158[253],s157[255],s156[257],s155[259],s154[261],s153[263],s152[265],s151[267],s150[269],s149[271],s148[273],s147[275],s146[277],s145[279],s144[281],s143[283],s142[285],s141[287],s140[289],s139[291],s138[293],s137[295],s136[297],s135[299],s134[301],s133[303],s132[305],s131[307],s130[309],s129[311],pp255[121],pp254[123],pp253[125],pp252[127],pp251[129],pp250[131],pp249[133],pp248[135],pp247[137],pp248[137],pp249[137],pp250[137],pp251[137]};
    assign in188_2 = {pp119[4],pp119[5],pp119[6],pp119[7],pp119[8],pp121[7],pp123[6],pp125[5],pp127[4],pp129[3],pp131[2],pp133[1],pp135[0],s129[72],s130[72],s131[72],s132[72],s133[72],s134[72],s135[72],s136[72],s137[72],s138[72],s139[72],s140[72],s141[72],s142[72],s143[72],s144[72],s145[72],s146[72],s147[72],s148[72],s149[72],s150[72],s151[72],s152[72],s153[72],s154[72],s155[72],s156[72],s157[72],s158[72],s159[72],s160[72],s161[72],s162[72],s163[72],s164[72],s165[72],s166[72],s167[72],s168[72],s169[72],s170[72],s171[72],s172[72],s173[72],s174[72],s175[72],s176[72],s177[72],s178[72],s179[72],s180[72],s181[72],s182[72],s183[72],s184[72],s185[72],s186[72],s187[72],s10[58],s11[58],s12[58],s13[58],s14[58],s15[58],s16[58],s17[58],s18[58],s19[58],s20[58],s21[58],s22[58],s23[58],s24[58],s25[58],s26[58],s27[58],s28[58],s29[58],s30[58],s31[58],s32[58],s33[58],s34[58],s35[58],s36[58],s37[58],s38[58],s39[58],s40[58],s41[58],s42[58],s42[59],s42[60],s42[61],s42[62],s42[63],s42[64],s42[65],s42[66],s42[67],s42[68],s42[69],s42[70],s42[71],s42[72],s42[73],s42[74],s42[75],s42[76],s42[77],s42[78],s42[79],s42[80],s42[81],s42[82],s42[83],s42[84],s42[85],s42[86],s42[87],s40[90],s38[93],s36[96],s34[99],s8[126],s7[128],s6[130],s5[132],s4[134],s3[136],s2[138],s1[140],s115[27],s113[30],s111[33],s109[36],s107[39],s105[42],s103[45],s101[48],s50[100],s49[102],s48[104],s47[106],s46[108],s45[110],s44[112],s43[114],s42[116],s41[118],s40[120],s39[122],s38[124],s37[126],s36[128],s35[130],s34[132],s33[134],s32[136],s31[138],s30[140],s29[142],s28[144],s27[146],s26[148],s25[150],s24[152],s23[154],s22[156],s21[158],s20[160],s19[162],s18[164],s17[166],s16[168],s15[170],s14[172],s13[174],s12[176],s11[178],s10[180],s187[196],s186[198],s185[200],s184[202],s183[204],s182[206],s181[208],s180[210],s179[212],s178[214],s177[216],s176[218],s175[220],s174[222],s173[224],s172[226],s171[228],s170[230],s169[232],s168[234],s167[236],s166[238],s165[240],s164[242],s163[244],s162[246],s161[248],s160[250],s159[252],s158[254],s157[256],s156[258],s155[260],s154[262],s153[264],s152[266],s151[268],s150[270],s149[272],s148[274],s147[276],s146[278],s145[280],s144[282],s143[284],s142[286],s141[288],s140[290],s139[292],s138[294],s137[296],s136[298],s135[300],s134[302],s133[304],s132[306],s131[308],s130[310],s129[312],pp255[122],pp254[124],pp253[126],pp252[128],pp251[130],pp250[132],pp249[134],pp248[136],pp249[136],pp250[136],pp251[136],pp252[136]};
    CLA_266 KS_188(s188, c188, in188_1, in188_2);
    wire[263:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp120[4],pp120[5],pp120[6],pp120[7],pp122[6],pp124[5],pp126[4],pp128[3],pp130[2],pp132[1],pp134[0],s129[71],s130[71],s131[71],s132[71],s133[71],s134[71],s135[71],s136[71],s137[71],s138[71],s139[71],s140[71],s141[71],s142[71],s143[71],s144[71],s145[71],s146[71],s147[71],s148[71],s149[71],s150[71],s151[71],s152[71],s153[71],s154[71],s155[71],s156[71],s157[71],s158[71],s159[71],s160[71],s161[71],s162[71],s163[71],s164[71],s165[71],s166[71],s167[71],s168[71],s169[71],s170[71],s171[71],s172[71],s173[71],s174[71],s175[71],s176[71],s177[71],s178[71],s179[71],s180[71],s181[71],s182[71],s183[71],s184[71],s185[71],s186[71],s187[71],s188[71],s188[72],s188[73],s188[74],s188[75],s188[76],s188[77],s188[78],s188[79],s188[80],s188[81],s188[82],s188[83],s188[84],s188[85],s188[86],s188[87],s188[88],s188[89],s188[90],s188[91],s188[92],s188[93],s188[94],s188[95],s188[96],s188[97],s188[98],s188[99],s188[100],s188[101],s188[102],s188[103],s188[104],s188[105],s188[106],s188[107],s188[108],s188[109],s188[110],s188[111],s188[112],s188[113],s188[114],s188[115],s188[116],s188[117],s188[118],s188[119],s188[120],s188[121],s188[122],s188[123],s188[124],s188[125],s188[126],s188[127],s188[128],s188[129],s188[130],s188[131],s188[132],s188[133],s188[134],s188[135],s188[136],s188[137],s188[138],s188[139],s188[140],s188[141],s188[142],s188[143],s188[144],s188[145],s188[146],s188[147],s188[148],s188[149],s188[150],s188[151],s188[152],s188[153],s188[154],s188[155],s188[156],s188[157],s188[158],s188[159],s188[160],s188[161],s188[162],s188[163],s188[164],s188[165],s188[166],s188[167],s188[168],s188[169],s188[170],s188[171],s188[172],s188[173],s188[174],s188[175],s188[176],s188[177],s188[178],s188[179],s188[180],s188[181],s188[182],s188[183],s188[184],s188[185],s188[186],s188[187],s188[188],s188[189],s188[190],s188[191],s188[192],s188[193],s188[194],s188[195],s187[197],s186[199],s185[201],s184[203],s183[205],s182[207],s181[209],s180[211],s179[213],s178[215],s177[217],s176[219],s175[221],s174[223],s173[225],s172[227],s171[229],s170[231],s169[233],s168[235],s167[237],s166[239],s165[241],s164[243],s163[245],s162[247],s161[249],s160[251],s159[253],s158[255],s157[257],s156[259],s155[261],s154[263],s153[265],s152[267],s151[269],s150[271],s149[273],s148[275],s147[277],s146[279],s145[281],s144[283],s143[285],s142[287],s141[289],s140[291],s139[293],s138[295],s137[297],s136[299],s135[301],s134[303],s133[305],s132[307],s131[309],s130[311],s129[313],pp255[123],pp254[125],pp253[127],pp252[129],pp251[131],pp250[133],pp249[135],pp250[135],pp251[135],pp252[135]};
    assign in189_2 = {pp121[3],pp121[4],pp121[5],pp121[6],pp123[5],pp125[4],pp127[3],pp129[2],pp131[1],pp133[0],s129[70],s130[70],s131[70],s132[70],s133[70],s134[70],s135[70],s136[70],s137[70],s138[70],s139[70],s140[70],s141[70],s142[70],s143[70],s144[70],s145[70],s146[70],s147[70],s148[70],s149[70],s150[70],s151[70],s152[70],s153[70],s154[70],s155[70],s156[70],s157[70],s158[70],s159[70],s160[70],s161[70],s162[70],s163[70],s164[70],s165[70],s166[70],s167[70],s168[70],s169[70],s170[70],s171[70],s172[70],s173[70],s174[70],s175[70],s176[70],s177[70],s178[70],s179[70],s180[70],s181[70],s182[70],s183[70],s184[70],s185[70],s186[70],s187[70],s188[70],s10[57],s11[57],s12[57],s13[57],s14[57],s15[57],s16[57],s17[57],s18[57],s19[57],s20[57],s21[57],s22[57],s23[57],s24[57],s25[57],s26[57],s27[57],s28[57],s29[57],s30[57],s31[57],s32[57],s33[57],s34[57],s35[57],s36[57],s37[57],s38[57],s39[57],s40[57],s41[57],s42[57],s43[57],s43[58],s43[59],s43[60],s43[61],s43[62],s43[63],s43[64],s43[65],s43[66],s43[67],s43[68],s43[69],s43[70],s43[71],s43[72],s43[73],s43[74],s43[75],s43[76],s43[77],s43[78],s43[79],s43[80],s43[81],s43[82],s43[83],s43[84],s43[85],s43[86],s41[89],s39[92],s37[95],s35[98],s9[125],s8[127],s7[129],s6[131],s5[133],s4[135],s3[137],s2[139],s1[141],s114[29],s112[32],s110[35],s108[38],s106[41],s104[44],s102[47],s100[50],s50[101],s49[103],s48[105],s47[107],s46[109],s45[111],s44[113],s43[115],s42[117],s41[119],s40[121],s39[123],s38[125],s37[127],s36[129],s35[131],s34[133],s33[135],s32[137],s31[139],s30[141],s29[143],s28[145],s27[147],s26[149],s25[151],s24[153],s23[155],s22[157],s21[159],s20[161],s19[163],s18[165],s17[167],s16[169],s15[171],s14[173],s13[175],s12[177],s11[179],s10[181],s188[196],s187[198],s186[200],s185[202],s184[204],s183[206],s182[208],s181[210],s180[212],s179[214],s178[216],s177[218],s176[220],s175[222],s174[224],s173[226],s172[228],s171[230],s170[232],s169[234],s168[236],s167[238],s166[240],s165[242],s164[244],s163[246],s162[248],s161[250],s160[252],s159[254],s158[256],s157[258],s156[260],s155[262],s154[264],s153[266],s152[268],s151[270],s150[272],s149[274],s148[276],s147[278],s146[280],s145[282],s144[284],s143[286],s142[288],s141[290],s140[292],s139[294],s138[296],s137[298],s136[300],s135[302],s134[304],s133[306],s132[308],s131[310],s130[312],s129[314],pp255[124],pp254[126],pp253[128],pp252[130],pp251[132],pp250[134],pp251[134],pp252[134],pp253[134]};
    CLA_264 KS_189(s189, c189, in189_1, in189_2);
    wire[261:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {pp122[3],pp122[4],pp122[5],pp124[4],pp126[3],pp128[2],pp130[1],pp132[0],s129[69],s130[69],s131[69],s132[69],s133[69],s134[69],s135[69],s136[69],s137[69],s138[69],s139[69],s140[69],s141[69],s142[69],s143[69],s144[69],s145[69],s146[69],s147[69],s148[69],s149[69],s150[69],s151[69],s152[69],s153[69],s154[69],s155[69],s156[69],s157[69],s158[69],s159[69],s160[69],s161[69],s162[69],s163[69],s164[69],s165[69],s166[69],s167[69],s168[69],s169[69],s170[69],s171[69],s172[69],s173[69],s174[69],s175[69],s176[69],s177[69],s178[69],s179[69],s180[69],s181[69],s182[69],s183[69],s184[69],s185[69],s186[69],s187[69],s188[69],s189[69],s189[70],s189[71],s189[72],s189[73],s189[74],s189[75],s189[76],s189[77],s189[78],s189[79],s189[80],s189[81],s189[82],s189[83],s189[84],s189[85],s189[86],s189[87],s189[88],s189[89],s189[90],s189[91],s189[92],s189[93],s189[94],s189[95],s189[96],s189[97],s189[98],s189[99],s189[100],s189[101],s189[102],s189[103],s189[104],s189[105],s189[106],s189[107],s189[108],s189[109],s189[110],s189[111],s189[112],s189[113],s189[114],s189[115],s189[116],s189[117],s189[118],s189[119],s189[120],s189[121],s189[122],s189[123],s189[124],s189[125],s189[126],s189[127],s189[128],s189[129],s189[130],s189[131],s189[132],s189[133],s189[134],s189[135],s189[136],s189[137],s189[138],s189[139],s189[140],s189[141],s189[142],s189[143],s189[144],s189[145],s189[146],s189[147],s189[148],s189[149],s189[150],s189[151],s189[152],s189[153],s189[154],s189[155],s189[156],s189[157],s189[158],s189[159],s189[160],s189[161],s189[162],s189[163],s189[164],s189[165],s189[166],s189[167],s189[168],s189[169],s189[170],s189[171],s189[172],s189[173],s189[174],s189[175],s189[176],s189[177],s189[178],s189[179],s189[180],s189[181],s189[182],s189[183],s189[184],s189[185],s189[186],s189[187],s189[188],s189[189],s189[190],s189[191],s189[192],s189[193],s189[194],s189[195],s188[197],s187[199],s186[201],s185[203],s184[205],s183[207],s182[209],s181[211],s180[213],s179[215],s178[217],s177[219],s176[221],s175[223],s174[225],s173[227],s172[229],s171[231],s170[233],s169[235],s168[237],s167[239],s166[241],s165[243],s164[245],s163[247],s162[249],s161[251],s160[253],s159[255],s158[257],s157[259],s156[261],s155[263],s154[265],s153[267],s152[269],s151[271],s150[273],s149[275],s148[277],s147[279],s146[281],s145[283],s144[285],s143[287],s142[289],s141[291],s140[293],s139[295],s138[297],s137[299],s136[301],s135[303],s134[305],s133[307],s132[309],s131[311],s130[313],s129[315],pp255[125],pp254[127],pp253[129],pp252[131],pp251[133],pp252[133],pp253[133]};
    assign in190_2 = {pp123[2],pp123[3],pp123[4],pp125[3],pp127[2],pp129[1],pp131[0],s129[68],s130[68],s131[68],s132[68],s133[68],s134[68],s135[68],s136[68],s137[68],s138[68],s139[68],s140[68],s141[68],s142[68],s143[68],s144[68],s145[68],s146[68],s147[68],s148[68],s149[68],s150[68],s151[68],s152[68],s153[68],s154[68],s155[68],s156[68],s157[68],s158[68],s159[68],s160[68],s161[68],s162[68],s163[68],s164[68],s165[68],s166[68],s167[68],s168[68],s169[68],s170[68],s171[68],s172[68],s173[68],s174[68],s175[68],s176[68],s177[68],s178[68],s179[68],s180[68],s181[68],s182[68],s183[68],s184[68],s185[68],s186[68],s187[68],s188[68],s189[68],s10[56],s11[56],s12[56],s13[56],s14[56],s15[56],s16[56],s17[56],s18[56],s19[56],s20[56],s21[56],s22[56],s23[56],s24[56],s25[56],s26[56],s27[56],s28[56],s29[56],s30[56],s31[56],s32[56],s33[56],s34[56],s35[56],s36[56],s37[56],s38[56],s39[56],s40[56],s41[56],s42[56],s43[56],s44[56],s44[57],s44[58],s44[59],s44[60],s44[61],s44[62],s44[63],s44[64],s44[65],s44[66],s44[67],s44[68],s44[69],s44[70],s44[71],s44[72],s44[73],s44[74],s44[75],s44[76],s44[77],s44[78],s44[79],s44[80],s44[81],s44[82],s44[83],s44[84],s44[85],s42[88],s40[91],s38[94],s36[97],s35[99],s9[126],s8[128],s7[130],s6[132],s5[134],s4[136],s3[138],s2[140],s1[142],s113[31],s111[34],s109[37],s107[40],s105[43],s103[46],s101[49],s51[100],s50[102],s49[104],s48[106],s47[108],s46[110],s45[112],s44[114],s43[116],s42[118],s41[120],s40[122],s39[124],s38[126],s37[128],s36[130],s35[132],s34[134],s33[136],s32[138],s31[140],s30[142],s29[144],s28[146],s27[148],s26[150],s25[152],s24[154],s23[156],s22[158],s21[160],s20[162],s19[164],s18[166],s17[168],s16[170],s15[172],s14[174],s13[176],s12[178],s11[180],s10[182],s189[196],s188[198],s187[200],s186[202],s185[204],s184[206],s183[208],s182[210],s181[212],s180[214],s179[216],s178[218],s177[220],s176[222],s175[224],s174[226],s173[228],s172[230],s171[232],s170[234],s169[236],s168[238],s167[240],s166[242],s165[244],s164[246],s163[248],s162[250],s161[252],s160[254],s159[256],s158[258],s157[260],s156[262],s155[264],s154[266],s153[268],s152[270],s151[272],s150[274],s149[276],s148[278],s147[280],s146[282],s145[284],s144[286],s143[288],s142[290],s141[292],s140[294],s139[296],s138[298],s137[300],s136[302],s135[304],s134[306],s133[308],s132[310],s131[312],s130[314],s129[316],pp255[126],pp254[128],pp253[130],pp252[132],pp253[132],pp254[132]};
    CLA_262 KS_190(s190, c190, in190_1, in190_2);
    wire[259:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {pp124[2],pp124[3],pp126[2],pp128[1],pp130[0],s129[67],s130[67],s131[67],s132[67],s133[67],s134[67],s135[67],s136[67],s137[67],s138[67],s139[67],s140[67],s141[67],s142[67],s143[67],s144[67],s145[67],s146[67],s147[67],s148[67],s149[67],s150[67],s151[67],s152[67],s153[67],s154[67],s155[67],s156[67],s157[67],s158[67],s159[67],s160[67],s161[67],s162[67],s163[67],s164[67],s165[67],s166[67],s167[67],s168[67],s169[67],s170[67],s171[67],s172[67],s173[67],s174[67],s175[67],s176[67],s177[67],s178[67],s179[67],s180[67],s181[67],s182[67],s183[67],s184[67],s185[67],s186[67],s187[67],s188[67],s189[67],s190[67],s190[68],s190[69],s190[70],s190[71],s190[72],s190[73],s190[74],s190[75],s190[76],s190[77],s190[78],s190[79],s190[80],s190[81],s190[82],s190[83],s190[84],s190[85],s190[86],s190[87],s190[88],s190[89],s190[90],s190[91],s190[92],s190[93],s190[94],s190[95],s190[96],s190[97],s190[98],s190[99],s190[100],s190[101],s190[102],s190[103],s190[104],s190[105],s190[106],s190[107],s190[108],s190[109],s190[110],s190[111],s190[112],s190[113],s190[114],s190[115],s190[116],s190[117],s190[118],s190[119],s190[120],s190[121],s190[122],s190[123],s190[124],s190[125],s190[126],s190[127],s190[128],s190[129],s190[130],s190[131],s190[132],s190[133],s190[134],s190[135],s190[136],s190[137],s190[138],s190[139],s190[140],s190[141],s190[142],s190[143],s190[144],s190[145],s190[146],s190[147],s190[148],s190[149],s190[150],s190[151],s190[152],s190[153],s190[154],s190[155],s190[156],s190[157],s190[158],s190[159],s190[160],s190[161],s190[162],s190[163],s190[164],s190[165],s190[166],s190[167],s190[168],s190[169],s190[170],s190[171],s190[172],s190[173],s190[174],s190[175],s190[176],s190[177],s190[178],s190[179],s190[180],s190[181],s190[182],s190[183],s190[184],s190[185],s190[186],s190[187],s190[188],s190[189],s190[190],s190[191],s190[192],s190[193],s190[194],s190[195],s189[197],s188[199],s187[201],s186[203],s185[205],s184[207],s183[209],s182[211],s181[213],s180[215],s179[217],s178[219],s177[221],s176[223],s175[225],s174[227],s173[229],s172[231],s171[233],s170[235],s169[237],s168[239],s167[241],s166[243],s165[245],s164[247],s163[249],s162[251],s161[253],s160[255],s159[257],s158[259],s157[261],s156[263],s155[265],s154[267],s153[269],s152[271],s151[273],s150[275],s149[277],s148[279],s147[281],s146[283],s145[285],s144[287],s143[289],s142[291],s141[293],s140[295],s139[297],s138[299],s137[301],s136[303],s135[305],s134[307],s133[309],s132[311],s131[313],s130[315],s129[317],pp255[127],pp254[129],pp253[131],pp254[131]};
    assign in191_2 = {pp125[1],pp125[2],pp127[1],pp129[0],s129[66],s130[66],s131[66],s132[66],s133[66],s134[66],s135[66],s136[66],s137[66],s138[66],s139[66],s140[66],s141[66],s142[66],s143[66],s144[66],s145[66],s146[66],s147[66],s148[66],s149[66],s150[66],s151[66],s152[66],s153[66],s154[66],s155[66],s156[66],s157[66],s158[66],s159[66],s160[66],s161[66],s162[66],s163[66],s164[66],s165[66],s166[66],s167[66],s168[66],s169[66],s170[66],s171[66],s172[66],s173[66],s174[66],s175[66],s176[66],s177[66],s178[66],s179[66],s180[66],s181[66],s182[66],s183[66],s184[66],s185[66],s186[66],s187[66],s188[66],s189[66],s190[66],s10[55],s11[55],s12[55],s13[55],s14[55],s15[55],s16[55],s17[55],s18[55],s19[55],s20[55],s21[55],s22[55],s23[55],s24[55],s25[55],s26[55],s27[55],s28[55],s29[55],s30[55],s31[55],s32[55],s33[55],s34[55],s35[55],s36[55],s37[55],s38[55],s39[55],s40[55],s41[55],s42[55],s43[55],s44[55],s45[55],s45[56],s45[57],s45[58],s45[59],s45[60],s45[61],s45[62],s45[63],s45[64],s45[65],s45[66],s45[67],s45[68],s45[69],s45[70],s45[71],s45[72],s45[73],s45[74],s45[75],s45[76],s45[77],s45[78],s45[79],s45[80],s45[81],s45[82],s45[83],s45[84],s43[87],s41[90],s39[93],s37[96],s36[98],s36[99],s9[127],s8[129],s7[131],s6[133],s5[135],s4[137],s3[139],s2[141],s1[143],s112[33],s110[36],s108[39],s106[42],s104[45],s102[48],s100[51],s51[101],s50[103],s49[105],s48[107],s47[109],s46[111],s45[113],s44[115],s43[117],s42[119],s41[121],s40[123],s39[125],s38[127],s37[129],s36[131],s35[133],s34[135],s33[137],s32[139],s31[141],s30[143],s29[145],s28[147],s27[149],s26[151],s25[153],s24[155],s23[157],s22[159],s21[161],s20[163],s19[165],s18[167],s17[169],s16[171],s15[173],s14[175],s13[177],s12[179],s11[181],s10[183],s190[196],s189[198],s188[200],s187[202],s186[204],s185[206],s184[208],s183[210],s182[212],s181[214],s180[216],s179[218],s178[220],s177[222],s176[224],s175[226],s174[228],s173[230],s172[232],s171[234],s170[236],s169[238],s168[240],s167[242],s166[244],s165[246],s164[248],s163[250],s162[252],s161[254],s160[256],s159[258],s158[260],s157[262],s156[264],s155[266],s154[268],s153[270],s152[272],s151[274],s150[276],s149[278],s148[280],s147[282],s146[284],s145[286],s144[288],s143[290],s142[292],s141[294],s140[296],s139[298],s138[300],s137[302],s136[304],s135[306],s134[308],s133[310],s132[312],s131[314],s130[316],s129[318],pp255[128],pp254[130],pp255[130]};
    CLA_260 KS_191(s191, c191, in191_1, in191_2);
    wire[257:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {pp126[1],pp128[0],s129[65],s130[65],s131[65],s132[65],s133[65],s134[65],s135[65],s136[65],s137[65],s138[65],s139[65],s140[65],s141[65],s142[65],s143[65],s144[65],s145[65],s146[65],s147[65],s148[65],s149[65],s150[65],s151[65],s152[65],s153[65],s154[65],s155[65],s156[65],s157[65],s158[65],s159[65],s160[65],s161[65],s162[65],s163[65],s164[65],s165[65],s166[65],s167[65],s168[65],s169[65],s170[65],s171[65],s172[65],s173[65],s174[65],s175[65],s176[65],s177[65],s178[65],s179[65],s180[65],s181[65],s182[65],s183[65],s184[65],s185[65],s186[65],s187[65],s188[65],s189[65],s190[65],s191[65],s191[66],s191[67],s191[68],s191[69],s191[70],s191[71],s191[72],s191[73],s191[74],s191[75],s191[76],s191[77],s191[78],s191[79],s191[80],s191[81],s191[82],s191[83],s191[84],s191[85],s191[86],s191[87],s191[88],s191[89],s191[90],s191[91],s191[92],s191[93],s191[94],s191[95],s191[96],s191[97],s191[98],s191[99],s191[100],s191[101],s191[102],s191[103],s191[104],s191[105],s191[106],s191[107],s191[108],s191[109],s191[110],s191[111],s191[112],s191[113],s191[114],s191[115],s191[116],s191[117],s191[118],s191[119],s191[120],s191[121],s191[122],s191[123],s191[124],s191[125],s191[126],s191[127],s191[128],s191[129],s191[130],s191[131],s191[132],s191[133],s191[134],s191[135],s191[136],s191[137],s191[138],s191[139],s191[140],s191[141],s191[142],s191[143],s191[144],s191[145],s191[146],s191[147],s191[148],s191[149],s191[150],s191[151],s191[152],s191[153],s191[154],s191[155],s191[156],s191[157],s191[158],s191[159],s191[160],s191[161],s191[162],s191[163],s191[164],s191[165],s191[166],s191[167],s191[168],s191[169],s191[170],s191[171],s191[172],s191[173],s191[174],s191[175],s191[176],s191[177],s191[178],s191[179],s191[180],s191[181],s191[182],s191[183],s191[184],s191[185],s191[186],s191[187],s191[188],s191[189],s191[190],s191[191],s191[192],s191[193],s191[194],s191[195],s190[197],s189[199],s188[201],s187[203],s186[205],s185[207],s184[209],s183[211],s182[213],s181[215],s180[217],s179[219],s178[221],s177[223],s176[225],s175[227],s174[229],s173[231],s172[233],s171[235],s170[237],s169[239],s168[241],s167[243],s166[245],s165[247],s164[249],s163[251],s162[253],s161[255],s160[257],s159[259],s158[261],s157[263],s156[265],s155[267],s154[269],s153[271],s152[273],s151[275],s150[277],s149[279],s148[281],s147[283],s146[285],s145[287],s144[289],s143[291],s142[293],s141[295],s140[297],s139[299],s138[301],s137[303],s136[305],s135[307],s134[309],s133[311],s132[313],s131[315],s130[317],s129[319],pp255[129]};
    assign in192_2 = {pp127[0],s129[64],s130[64],s131[64],s132[64],s133[64],s134[64],s135[64],s136[64],s137[64],s138[64],s139[64],s140[64],s141[64],s142[64],s143[64],s144[64],s145[64],s146[64],s147[64],s148[64],s149[64],s150[64],s151[64],s152[64],s153[64],s154[64],s155[64],s156[64],s157[64],s158[64],s159[64],s160[64],s161[64],s162[64],s163[64],s164[64],s165[64],s166[64],s167[64],s168[64],s169[64],s170[64],s171[64],s172[64],s173[64],s174[64],s175[64],s176[64],s177[64],s178[64],s179[64],s180[64],s181[64],s182[64],s183[64],s184[64],s185[64],s186[64],s187[64],s188[64],s189[64],s190[64],s191[64],s10[54],s11[54],s12[54],s13[54],s14[54],s15[54],s16[54],s17[54],s18[54],s19[54],s20[54],s21[54],s22[54],s23[54],s24[54],s25[54],s26[54],s27[54],s28[54],s29[54],s30[54],s31[54],s32[54],s33[54],s34[54],s35[54],s36[54],s37[54],s38[54],s39[54],s40[54],s41[54],s42[54],s43[54],s44[54],s45[54],s46[54],s46[55],s46[56],s46[57],s46[58],s46[59],s46[60],s46[61],s46[62],s46[63],s46[64],s46[65],s46[66],s46[67],s46[68],s46[69],s46[70],s46[71],s46[72],s46[73],s46[74],s46[75],s46[76],s46[77],s46[78],s46[79],s46[80],s46[81],s46[82],s46[83],s44[86],s42[89],s40[92],s38[95],s37[97],s37[98],s37[99],s9[128],s8[130],s7[132],s6[134],s5[136],s4[138],s3[140],s2[142],s1[144],s111[35],s109[38],s107[41],s105[44],s103[47],s101[50],s52[100],s51[102],s50[104],s49[106],s48[108],s47[110],s46[112],s45[114],s44[116],s43[118],s42[120],s41[122],s40[124],s39[126],s38[128],s37[130],s36[132],s35[134],s34[136],s33[138],s32[140],s31[142],s30[144],s29[146],s28[148],s27[150],s26[152],s25[154],s24[156],s23[158],s22[160],s21[162],s20[164],s19[166],s18[168],s17[170],s16[172],s15[174],s14[176],s13[178],s12[180],s11[182],s10[184],s191[196],s190[198],s189[200],s188[202],s187[204],s186[206],s185[208],s184[210],s183[212],s182[214],s181[216],s180[218],s179[220],s178[222],s177[224],s176[226],s175[228],s174[230],s173[232],s172[234],s171[236],s170[238],s169[240],s168[242],s167[244],s166[246],s165[248],s164[250],s163[252],s162[254],s161[256],s160[258],s159[260],s158[262],s157[264],s156[266],s155[268],s154[270],s153[272],s152[274],s151[276],s150[278],s149[280],s148[282],s147[284],s146[286],s145[288],s144[290],s143[292],s142[294],s141[296],s140[298],s139[300],s138[302],s137[304],s136[306],s135[308],s134[310],s133[312],s132[314],s131[316],s130[318],s129[320]};
    CLA_258 KS_192(s192, c192, in192_1, in192_2);

    /*Stage 3*/
    wire[447:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {pp10[22],pp10[23],pp10[24],pp10[25],pp10[26],pp10[27],pp10[28],pp10[29],pp10[30],pp10[31],pp10[32],pp10[33],pp10[34],pp10[35],pp10[36],pp10[37],pp10[38],pp10[39],pp10[40],pp10[41],pp10[42],pp10[43],pp10[44],pp10[45],pp10[46],pp10[47],pp10[48],pp10[49],pp10[50],pp10[51],pp10[52],pp10[53],pp12[52],pp14[51],pp16[50],pp18[49],pp20[48],pp22[47],pp24[46],pp26[45],pp28[44],pp30[43],pp32[42],pp34[41],pp36[40],pp38[39],pp40[38],pp42[37],pp44[36],pp46[35],pp48[34],pp50[33],pp52[32],pp54[31],pp56[30],pp58[29],pp60[28],pp62[27],pp64[26],pp66[25],pp68[24],pp70[23],pp72[22],pp74[21],pp76[20],pp78[19],pp80[18],pp82[17],pp83[17],pp84[17],pp85[17],pp86[17],pp87[17],pp88[17],pp89[17],pp90[17],pp91[17],pp92[17],pp93[17],pp94[17],pp95[17],pp96[17],pp97[17],pp98[17],pp99[17],pp108[9],pp110[8],pp112[7],pp114[6],pp116[5],pp118[4],pp120[3],pp122[2],pp124[1],pp126[0],s129[63],s130[63],s131[63],s132[63],s133[63],s134[63],s135[63],s136[63],s137[63],s138[63],s139[63],s140[63],s141[63],s142[63],s143[63],s144[63],s145[63],s146[63],s147[63],s148[63],s149[63],s150[63],s151[63],s152[63],s153[63],s154[63],s155[63],s156[63],s157[63],s158[63],s159[63],s160[63],s161[63],s162[63],s163[63],s164[63],s165[63],s166[63],s167[63],s168[63],s169[63],s170[63],s171[63],s172[63],s173[63],s174[63],s175[63],s176[63],s177[63],s178[63],s179[63],s180[63],s181[63],s182[63],s183[63],s184[63],s185[63],s186[63],s187[63],s188[63],s189[63],s190[63],s191[63],s192[63],s192[64],s192[65],s192[66],s192[67],s192[68],s192[69],s192[70],s192[71],s192[72],s192[73],s192[74],s192[75],s192[76],s192[77],s192[78],s192[79],s192[80],s192[81],s192[82],s192[83],s192[84],s192[85],s192[86],s192[87],s192[88],s192[89],s192[90],s192[91],s192[92],s192[93],s192[94],s192[95],s192[96],s192[97],s192[98],s192[99],s192[100],s192[101],s192[102],s192[103],s192[104],s192[105],s192[106],s192[107],s192[108],s192[109],s192[110],s192[111],s192[112],s192[113],s192[114],s192[115],s192[116],s192[117],s192[118],s192[119],s192[120],s192[121],s192[122],s192[123],s192[124],s192[125],s192[126],s192[127],s192[128],s192[129],s192[130],s192[131],s192[132],s192[133],s192[134],s192[135],s192[136],s192[137],s192[138],s192[139],s192[140],s192[141],s192[142],s192[143],s192[144],s192[145],s192[146],s192[147],s192[148],s192[149],s192[150],s192[151],s192[152],s192[153],s192[154],s192[155],s192[156],s192[157],s192[158],s192[159],s192[160],s192[161],s192[162],s192[163],s192[164],s192[165],s192[166],s192[167],s192[168],s192[169],s192[170],s192[171],s192[172],s192[173],s192[174],s192[175],s192[176],s192[177],s192[178],s192[179],s192[180],s192[181],s192[182],s192[183],s192[184],s192[185],s192[186],s192[187],s192[188],s192[189],s192[190],s192[191],s192[192],s192[193],s192[194],s192[195],s191[197],s190[199],s189[201],s188[203],s187[205],s186[207],s185[209],s184[211],s183[213],s182[215],s181[217],s180[219],s179[221],s178[223],s177[225],s176[227],s175[229],s174[231],s173[233],s172[235],s171[237],s170[239],s169[241],s168[243],s167[245],s166[247],s165[249],s164[251],s163[253],s162[255],s161[257],s160[259],s159[261],s158[263],s157[265],s156[267],s155[269],s154[271],s153[273],s152[275],s151[277],s150[279],s149[281],s148[283],s147[285],s146[287],s145[289],s144[291],s143[293],s142[295],s141[297],s140[299],s139[301],s138[303],s137[305],s136[307],s135[309],s134[311],s133[313],s132[315],s131[317],s130[319],s129[321],pp255[131],pp254[133],pp253[135],pp252[137],pp251[139],pp250[141],pp249[143],pp248[145],pp247[147],pp246[149],pp245[151],pp244[153],pp243[155],pp242[157],pp241[159],pp240[161],pp239[163],pp238[165],pp237[167],pp236[169],pp235[171],pp234[173],pp233[175],pp232[177],pp231[179],pp230[181],pp229[183],pp228[185],pp227[187],pp226[189],pp225[191],pp224[193],pp223[195],pp222[197],pp221[199],pp220[201],pp219[203],pp218[205],pp217[207],pp216[209],pp215[211],pp214[213],pp213[215],pp212[217],pp211[219],pp210[221],pp209[223],pp208[225],pp207[227],pp206[229],pp205[231],pp204[233],pp203[235],pp202[237],pp201[239],pp200[241],pp199[243],pp198[245],pp197[247],pp196[249],pp195[251],pp194[253],pp193[255],pp194[255],pp195[255],pp196[255],pp197[255],pp198[255],pp199[255],pp200[255],pp201[255],pp202[255],pp203[255],pp204[255],pp205[255],pp206[255],pp207[255],pp208[255],pp209[255],pp210[255],pp211[255],pp212[255],pp213[255],pp214[255],pp215[255],pp216[255],pp217[255],pp218[255],pp219[255],pp220[255],pp221[255],pp222[255],pp223[255],pp224[255]};
    assign in193_2 = {pp11[21],pp11[22],pp11[23],pp11[24],pp11[25],pp11[26],pp11[27],pp11[28],pp11[29],pp11[30],pp11[31],pp11[32],pp11[33],pp11[34],pp11[35],pp11[36],pp11[37],pp11[38],pp11[39],pp11[40],pp11[41],pp11[42],pp11[43],pp11[44],pp11[45],pp11[46],pp11[47],pp11[48],pp11[49],pp11[50],pp11[51],pp11[52],pp13[51],pp15[50],pp17[49],pp19[48],pp21[47],pp23[46],pp25[45],pp27[44],pp29[43],pp31[42],pp33[41],pp35[40],pp37[39],pp39[38],pp41[37],pp43[36],pp45[35],pp47[34],pp49[33],pp51[32],pp53[31],pp55[30],pp57[29],pp59[28],pp61[27],pp63[26],pp65[25],pp67[24],pp69[23],pp71[22],pp73[21],pp75[20],pp77[19],pp79[18],pp81[17],pp83[16],pp84[16],pp85[16],pp86[16],pp87[16],pp88[16],pp89[16],pp90[16],pp91[16],pp92[16],pp93[16],pp94[16],pp95[16],pp96[16],pp97[16],pp98[16],pp99[16],pp107[9],pp109[8],pp111[7],pp113[6],pp115[5],pp117[4],pp119[3],pp121[2],pp123[1],pp125[0],s129[62],s130[62],s131[62],s132[62],s133[62],s134[62],s135[62],s136[62],s137[62],s138[62],s139[62],s140[62],s141[62],s142[62],s143[62],s144[62],s145[62],s146[62],s147[62],s148[62],s149[62],s150[62],s151[62],s152[62],s153[62],s154[62],s155[62],s156[62],s157[62],s158[62],s159[62],s160[62],s161[62],s162[62],s163[62],s164[62],s165[62],s166[62],s167[62],s168[62],s169[62],s170[62],s171[62],s172[62],s173[62],s174[62],s175[62],s176[62],s177[62],s178[62],s179[62],s180[62],s181[62],s182[62],s183[62],s184[62],s185[62],s186[62],s187[62],s188[62],s189[62],s190[62],s191[62],s192[62],s10[53],s11[53],s12[53],s13[53],s14[53],s15[53],s16[53],s17[53],s18[53],s19[53],s20[53],s21[53],s22[53],s23[53],s24[53],s25[53],s26[53],s27[53],s28[53],s29[53],s30[53],s31[53],s32[53],s33[53],s34[53],s35[53],s36[53],s37[53],s38[53],s39[53],s40[53],s41[53],s42[53],s43[53],s44[53],s45[53],s46[53],s47[53],s47[54],s47[55],s47[56],s47[57],s47[58],s47[59],s47[60],s47[61],s47[62],s47[63],s47[64],s47[65],s47[66],s47[67],s47[68],s47[69],s47[70],s47[71],s47[72],s47[73],s47[74],s47[75],s47[76],s47[77],s47[78],s47[79],s47[80],s47[81],s47[82],s45[85],s43[88],s41[91],s39[94],s38[96],s38[97],s38[98],s38[99],s9[129],s8[131],s7[133],s6[135],s5[137],s4[139],s3[141],s2[143],s1[145],s110[37],s108[40],s106[43],s104[46],s102[49],s100[52],s52[101],s51[103],s50[105],s49[107],s48[109],s47[111],s46[113],s45[115],s44[117],s43[119],s42[121],s41[123],s40[125],s39[127],s38[129],s37[131],s36[133],s35[135],s34[137],s33[139],s32[141],s31[143],s30[145],s29[147],s28[149],s27[151],s26[153],s25[155],s24[157],s23[159],s22[161],s21[163],s20[165],s19[167],s18[169],s17[171],s16[173],s15[175],s14[177],s13[179],s12[181],s11[183],s10[185],s192[196],s191[198],s190[200],s189[202],s188[204],s187[206],s186[208],s185[210],s184[212],s183[214],s182[216],s181[218],s180[220],s179[222],s178[224],s177[226],s176[228],s175[230],s174[232],s173[234],s172[236],s171[238],s170[240],s169[242],s168[244],s167[246],s166[248],s165[250],s164[252],s163[254],s162[256],s161[258],s160[260],s159[262],s158[264],s157[266],s156[268],s155[270],s154[272],s153[274],s152[276],s151[278],s150[280],s149[282],s148[284],s147[286],s146[288],s145[290],s144[292],s143[294],s142[296],s141[298],s140[300],s139[302],s138[304],s137[306],s136[308],s135[310],s134[312],s133[314],s132[316],s131[318],s130[320],s129[322],pp255[132],pp254[134],pp253[136],pp252[138],pp251[140],pp250[142],pp249[144],pp248[146],pp247[148],pp246[150],pp245[152],pp244[154],pp243[156],pp242[158],pp241[160],pp240[162],pp239[164],pp238[166],pp237[168],pp236[170],pp235[172],pp234[174],pp233[176],pp232[178],pp231[180],pp230[182],pp229[184],pp228[186],pp227[188],pp226[190],pp225[192],pp224[194],pp223[196],pp222[198],pp221[200],pp220[202],pp219[204],pp218[206],pp217[208],pp216[210],pp215[212],pp214[214],pp213[216],pp212[218],pp211[220],pp210[222],pp209[224],pp208[226],pp207[228],pp206[230],pp205[232],pp204[234],pp203[236],pp202[238],pp201[240],pp200[242],pp199[244],pp198[246],pp197[248],pp196[250],pp195[252],pp194[254],pp195[254],pp196[254],pp197[254],pp198[254],pp199[254],pp200[254],pp201[254],pp202[254],pp203[254],pp204[254],pp205[254],pp206[254],pp207[254],pp208[254],pp209[254],pp210[254],pp211[254],pp212[254],pp213[254],pp214[254],pp215[254],pp216[254],pp217[254],pp218[254],pp219[254],pp220[254],pp221[254],pp222[254],pp223[254],pp224[254],pp225[254]};
    CLA_448 KS_193(s193, c193, in193_1, in193_2);
    wire[445:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {pp12[21],pp12[22],pp12[23],pp12[24],pp12[25],pp12[26],pp12[27],pp12[28],pp12[29],pp12[30],pp12[31],pp12[32],pp12[33],pp12[34],pp12[35],pp12[36],pp12[37],pp12[38],pp12[39],pp12[40],pp12[41],pp12[42],pp12[43],pp12[44],pp12[45],pp12[46],pp12[47],pp12[48],pp12[49],pp12[50],pp12[51],pp14[50],pp16[49],pp18[48],pp20[47],pp22[46],pp24[45],pp26[44],pp28[43],pp30[42],pp32[41],pp34[40],pp36[39],pp38[38],pp40[37],pp42[36],pp44[35],pp46[34],pp48[33],pp50[32],pp52[31],pp54[30],pp56[29],pp58[28],pp60[27],pp62[26],pp64[25],pp66[24],pp68[23],pp70[22],pp72[21],pp74[20],pp76[19],pp78[18],pp80[17],pp82[16],pp84[15],pp85[15],pp86[15],pp87[15],pp88[15],pp89[15],pp90[15],pp91[15],pp92[15],pp93[15],pp94[15],pp95[15],pp96[15],pp97[15],pp98[15],pp99[15],pp106[9],pp108[8],pp110[7],pp112[6],pp114[5],pp116[4],pp118[3],pp120[2],pp122[1],pp124[0],s129[61],s130[61],s131[61],s132[61],s133[61],s134[61],s135[61],s193[100],s193[101],s193[102],s193[103],s193[104],s193[105],s193[106],s193[107],s193[108],s193[109],s193[110],s193[111],s193[112],s193[113],s193[114],s193[115],s193[116],s193[117],s193[118],s193[119],s193[120],s193[121],s193[122],s193[123],s193[124],s193[125],s193[126],s193[127],s193[128],s193[129],s193[130],s193[131],s193[132],s193[133],s193[134],s193[135],s193[136],s193[137],s193[138],s193[139],s193[140],s193[141],s193[142],s193[143],s193[144],s193[145],s193[146],s193[147],s193[148],s193[149],s193[150],s193[151],s193[152],s193[153],s193[154],s193[155],s193[156],s193[157],s193[158],s193[159],s193[160],s193[161],s193[162],s193[163],s193[164],s193[165],s193[166],s193[167],s193[168],s193[169],s193[170],s193[171],s193[172],s193[173],s193[174],s193[175],s193[176],s193[177],s193[178],s193[179],s193[180],s193[181],s193[182],s193[183],s193[184],s193[185],s193[186],s193[187],s193[188],s193[189],s193[190],s193[191],s193[192],s193[193],s193[194],s193[195],s193[196],s193[197],s193[198],s193[199],s193[200],s193[201],s193[202],s193[203],s193[204],s193[205],s193[206],s193[207],s193[208],s193[209],s193[210],s193[211],s193[212],s193[213],s193[214],s193[215],s193[216],s193[217],s193[218],s193[219],s193[220],s193[221],s193[222],s193[223],s193[224],s193[225],s193[226],s193[227],s193[228],s193[229],s193[230],s193[231],s193[232],s193[233],s193[234],s193[235],s193[236],s193[237],s193[238],s193[239],s193[240],s193[241],s193[242],s193[243],s193[244],s193[245],s193[246],s193[247],s193[248],s193[249],s193[250],s193[251],s193[252],s193[253],s193[254],s193[255],s193[256],s193[257],s193[258],s193[259],s193[260],s193[261],s193[262],s193[263],s193[264],s193[265],s193[266],s193[267],s193[268],s193[269],s193[270],s193[271],s193[272],s193[273],s193[274],s193[275],s193[276],s193[277],s193[278],s193[279],s193[280],s193[281],s193[282],s193[283],s193[284],s193[285],s193[286],s193[287],s193[288],s193[289],s193[290],s193[291],s192[197],s191[199],s190[201],s189[203],s188[205],s187[207],s186[209],s185[211],s184[213],s183[215],s182[217],s181[219],s180[221],s179[223],s178[225],s177[227],s176[229],s175[231],s174[233],s173[235],s172[237],s171[239],s170[241],s169[243],s168[245],s167[247],s166[249],s165[251],s164[253],s163[255],s162[257],s161[259],s160[261],s159[263],s158[265],s157[267],s156[269],s155[271],s154[273],s153[275],s152[277],s151[279],s150[281],s149[283],s148[285],s147[287],s146[289],s145[291],s144[293],s143[295],s142[297],s141[299],s140[301],s139[303],s138[305],s137[307],s136[309],s135[311],s134[313],s133[315],s132[317],s131[319],s130[321],s129[323],pp255[133],pp254[135],pp253[137],pp252[139],pp251[141],pp250[143],pp249[145],pp248[147],pp247[149],pp246[151],pp245[153],pp244[155],pp243[157],pp242[159],pp241[161],pp240[163],pp239[165],pp238[167],pp237[169],pp236[171],pp235[173],pp234[175],pp233[177],pp232[179],pp231[181],pp230[183],pp229[185],pp228[187],pp227[189],pp226[191],pp225[193],pp224[195],pp223[197],pp222[199],pp221[201],pp220[203],pp219[205],pp218[207],pp217[209],pp216[211],pp215[213],pp214[215],pp213[217],pp212[219],pp211[221],pp210[223],pp209[225],pp208[227],pp207[229],pp206[231],pp205[233],pp204[235],pp203[237],pp202[239],pp201[241],pp200[243],pp199[245],pp198[247],pp197[249],pp196[251],pp195[253],pp196[253],pp197[253],pp198[253],pp199[253],pp200[253],pp201[253],pp202[253],pp203[253],pp204[253],pp205[253],pp206[253],pp207[253],pp208[253],pp209[253],pp210[253],pp211[253],pp212[253],pp213[253],pp214[253],pp215[253],pp216[253],pp217[253],pp218[253],pp219[253],pp220[253],pp221[253],pp222[253],pp223[253],pp224[253],pp225[253]};
    assign in194_2 = {pp13[20],pp13[21],pp13[22],pp13[23],pp13[24],pp13[25],pp13[26],pp13[27],pp13[28],pp13[29],pp13[30],pp13[31],pp13[32],pp13[33],pp13[34],pp13[35],pp13[36],pp13[37],pp13[38],pp13[39],pp13[40],pp13[41],pp13[42],pp13[43],pp13[44],pp13[45],pp13[46],pp13[47],pp13[48],pp13[49],pp13[50],pp15[49],pp17[48],pp19[47],pp21[46],pp23[45],pp25[44],pp27[43],pp29[42],pp31[41],pp33[40],pp35[39],pp37[38],pp39[37],pp41[36],pp43[35],pp45[34],pp47[33],pp49[32],pp51[31],pp53[30],pp55[29],pp57[28],pp59[27],pp61[26],pp63[25],pp65[24],pp67[23],pp69[22],pp71[21],pp73[20],pp75[19],pp77[18],pp79[17],pp81[16],pp83[15],pp85[14],pp86[14],pp87[14],pp88[14],pp89[14],pp90[14],pp91[14],pp92[14],pp93[14],pp94[14],pp95[14],pp96[14],pp97[14],pp98[14],pp99[14],pp105[9],pp107[8],pp109[7],pp111[6],pp113[5],pp115[4],pp117[3],pp119[2],pp121[1],pp123[0],s129[60],s130[60],s131[60],s132[60],s133[60],s134[60],s135[60],s136[60],s136[61],s137[61],s138[61],s139[61],s140[61],s141[61],s142[61],s143[61],s144[61],s145[61],s146[61],s147[61],s148[61],s149[61],s150[61],s151[61],s152[61],s153[61],s154[61],s155[61],s156[61],s157[61],s158[61],s159[61],s160[61],s161[61],s162[61],s163[61],s164[61],s165[61],s166[61],s167[61],s168[61],s169[61],s170[61],s171[61],s172[61],s173[61],s174[61],s175[61],s176[61],s177[61],s178[61],s179[61],s180[61],s181[61],s182[61],s183[61],s184[61],s185[61],s186[61],s187[61],s188[61],s189[61],s190[61],s191[61],s192[61],s10[52],s11[52],s12[52],s13[52],s14[52],s15[52],s16[52],s17[52],s18[52],s19[52],s20[52],s21[52],s22[52],s23[52],s24[52],s25[52],s26[52],s27[52],s28[52],s29[52],s30[52],s31[52],s32[52],s33[52],s34[52],s35[52],s36[52],s37[52],s38[52],s39[52],s40[52],s41[52],s42[52],s43[52],s44[52],s45[52],s46[52],s47[52],s48[52],s48[53],s48[54],s48[55],s48[56],s48[57],s48[58],s48[59],s48[60],s48[61],s48[62],s48[63],s48[64],s48[65],s48[66],s48[67],s48[68],s48[69],s48[70],s48[71],s48[72],s48[73],s48[74],s48[75],s48[76],s48[77],s48[78],s48[79],s48[80],s48[81],s46[84],s44[87],s42[90],s40[93],s39[95],s39[96],s39[97],s39[98],s39[99],s9[130],s8[132],s7[134],s6[136],s5[138],s4[140],s3[142],s2[144],s1[146],s109[39],s107[42],s105[45],s103[48],s101[51],s53[100],s52[102],s51[104],s50[106],s49[108],s48[110],s47[112],s46[114],s45[116],s44[118],s43[120],s42[122],s41[124],s40[126],s39[128],s38[130],s37[132],s36[134],s35[136],s34[138],s33[140],s32[142],s31[144],s30[146],s29[148],s28[150],s27[152],s26[154],s25[156],s24[158],s23[160],s22[162],s21[164],s20[166],s19[168],s18[170],s17[172],s16[174],s15[176],s14[178],s13[180],s12[182],s11[184],s10[186],s193[292],s192[198],s191[200],s190[202],s189[204],s188[206],s187[208],s186[210],s185[212],s184[214],s183[216],s182[218],s181[220],s180[222],s179[224],s178[226],s177[228],s176[230],s175[232],s174[234],s173[236],s172[238],s171[240],s170[242],s169[244],s168[246],s167[248],s166[250],s165[252],s164[254],s163[256],s162[258],s161[260],s160[262],s159[264],s158[266],s157[268],s156[270],s155[272],s154[274],s153[276],s152[278],s151[280],s150[282],s149[284],s148[286],s147[288],s146[290],s145[292],s144[294],s143[296],s142[298],s141[300],s140[302],s139[304],s138[306],s137[308],s136[310],s135[312],s134[314],s133[316],s132[318],s131[320],s130[322],s129[324],pp255[134],pp254[136],pp253[138],pp252[140],pp251[142],pp250[144],pp249[146],pp248[148],pp247[150],pp246[152],pp245[154],pp244[156],pp243[158],pp242[160],pp241[162],pp240[164],pp239[166],pp238[168],pp237[170],pp236[172],pp235[174],pp234[176],pp233[178],pp232[180],pp231[182],pp230[184],pp229[186],pp228[188],pp227[190],pp226[192],pp225[194],pp224[196],pp223[198],pp222[200],pp221[202],pp220[204],pp219[206],pp218[208],pp217[210],pp216[212],pp215[214],pp214[216],pp213[218],pp212[220],pp211[222],pp210[224],pp209[226],pp208[228],pp207[230],pp206[232],pp205[234],pp204[236],pp203[238],pp202[240],pp201[242],pp200[244],pp199[246],pp198[248],pp197[250],pp196[252],pp197[252],pp198[252],pp199[252],pp200[252],pp201[252],pp202[252],pp203[252],pp204[252],pp205[252],pp206[252],pp207[252],pp208[252],pp209[252],pp210[252],pp211[252],pp212[252],pp213[252],pp214[252],pp215[252],pp216[252],pp217[252],pp218[252],pp219[252],pp220[252],pp221[252],pp222[252],pp223[252],pp224[252],pp225[252],pp226[252]};
    CLA_446 KS_194(s194, c194, in194_1, in194_2);
    wire[443:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp14[20],pp14[21],pp14[22],pp14[23],pp14[24],pp14[25],pp14[26],pp14[27],pp14[28],pp14[29],pp14[30],pp14[31],pp14[32],pp14[33],pp14[34],pp14[35],pp14[36],pp14[37],pp14[38],pp14[39],pp14[40],pp14[41],pp14[42],pp14[43],pp14[44],pp14[45],pp14[46],pp14[47],pp14[48],pp14[49],pp16[48],pp18[47],pp20[46],pp22[45],pp24[44],pp26[43],pp28[42],pp30[41],pp32[40],pp34[39],pp36[38],pp38[37],pp40[36],pp42[35],pp44[34],pp46[33],pp48[32],pp50[31],pp52[30],pp54[29],pp56[28],pp58[27],pp60[26],pp62[25],pp64[24],pp66[23],pp68[22],pp70[21],pp72[20],pp74[19],pp76[18],pp78[17],pp80[16],pp82[15],pp84[14],pp86[13],pp87[13],pp88[13],pp89[13],pp90[13],pp91[13],pp92[13],pp93[13],pp94[13],pp95[13],pp96[13],pp97[13],pp98[13],pp99[13],pp104[9],pp106[8],pp108[7],pp110[6],pp112[5],pp114[4],pp116[3],pp118[2],pp120[1],pp122[0],s129[59],s130[59],s131[59],s132[59],s133[59],s134[59],s135[59],s136[59],s137[59],s137[60],s194[100],s194[101],s194[102],s194[103],s194[104],s194[105],s194[106],s194[107],s194[108],s194[109],s194[110],s194[111],s194[112],s194[113],s194[114],s194[115],s194[116],s194[117],s194[118],s194[119],s194[120],s194[121],s194[122],s194[123],s194[124],s194[125],s194[126],s194[127],s194[128],s194[129],s194[130],s194[131],s194[132],s194[133],s194[134],s194[135],s194[136],s194[137],s194[138],s194[139],s194[140],s194[141],s194[142],s194[143],s194[144],s194[145],s194[146],s194[147],s194[148],s194[149],s194[150],s194[151],s194[152],s194[153],s194[154],s194[155],s194[156],s194[157],s194[158],s194[159],s194[160],s194[161],s194[162],s194[163],s194[164],s194[165],s194[166],s194[167],s194[168],s194[169],s194[170],s194[171],s194[172],s194[173],s194[174],s194[175],s194[176],s194[177],s194[178],s194[179],s194[180],s194[181],s194[182],s194[183],s194[184],s194[185],s194[186],s194[187],s194[188],s194[189],s194[190],s194[191],s194[192],s194[193],s194[194],s194[195],s194[196],s194[197],s194[198],s194[199],s194[200],s194[201],s194[202],s194[203],s194[204],s194[205],s194[206],s194[207],s194[208],s194[209],s194[210],s194[211],s194[212],s194[213],s194[214],s194[215],s194[216],s194[217],s194[218],s194[219],s194[220],s194[221],s194[222],s194[223],s194[224],s194[225],s194[226],s194[227],s194[228],s194[229],s194[230],s194[231],s194[232],s194[233],s194[234],s194[235],s194[236],s194[237],s194[238],s194[239],s194[240],s194[241],s194[242],s194[243],s194[244],s194[245],s194[246],s194[247],s194[248],s194[249],s194[250],s194[251],s194[252],s194[253],s194[254],s194[255],s194[256],s194[257],s194[258],s194[259],s194[260],s194[261],s194[262],s194[263],s194[264],s194[265],s194[266],s194[267],s194[268],s194[269],s194[270],s194[271],s194[272],s194[273],s194[274],s194[275],s194[276],s194[277],s194[278],s194[279],s194[280],s194[281],s194[282],s194[283],s194[284],s194[285],s194[286],s194[287],s194[288],s194[289],s194[290],s194[291],s193[293],s192[199],s191[201],s190[203],s189[205],s188[207],s187[209],s186[211],s185[213],s184[215],s183[217],s182[219],s181[221],s180[223],s179[225],s178[227],s177[229],s176[231],s175[233],s174[235],s173[237],s172[239],s171[241],s170[243],s169[245],s168[247],s167[249],s166[251],s165[253],s164[255],s163[257],s162[259],s161[261],s160[263],s159[265],s158[267],s157[269],s156[271],s155[273],s154[275],s153[277],s152[279],s151[281],s150[283],s149[285],s148[287],s147[289],s146[291],s145[293],s144[295],s143[297],s142[299],s141[301],s140[303],s139[305],s138[307],s137[309],s136[311],s135[313],s134[315],s133[317],s132[319],s131[321],s130[323],s129[325],pp255[135],pp254[137],pp253[139],pp252[141],pp251[143],pp250[145],pp249[147],pp248[149],pp247[151],pp246[153],pp245[155],pp244[157],pp243[159],pp242[161],pp241[163],pp240[165],pp239[167],pp238[169],pp237[171],pp236[173],pp235[175],pp234[177],pp233[179],pp232[181],pp231[183],pp230[185],pp229[187],pp228[189],pp227[191],pp226[193],pp225[195],pp224[197],pp223[199],pp222[201],pp221[203],pp220[205],pp219[207],pp218[209],pp217[211],pp216[213],pp215[215],pp214[217],pp213[219],pp212[221],pp211[223],pp210[225],pp209[227],pp208[229],pp207[231],pp206[233],pp205[235],pp204[237],pp203[239],pp202[241],pp201[243],pp200[245],pp199[247],pp198[249],pp197[251],pp198[251],pp199[251],pp200[251],pp201[251],pp202[251],pp203[251],pp204[251],pp205[251],pp206[251],pp207[251],pp208[251],pp209[251],pp210[251],pp211[251],pp212[251],pp213[251],pp214[251],pp215[251],pp216[251],pp217[251],pp218[251],pp219[251],pp220[251],pp221[251],pp222[251],pp223[251],pp224[251],pp225[251],pp226[251]};
    assign in195_2 = {pp15[19],pp15[20],pp15[21],pp15[22],pp15[23],pp15[24],pp15[25],pp15[26],pp15[27],pp15[28],pp15[29],pp15[30],pp15[31],pp15[32],pp15[33],pp15[34],pp15[35],pp15[36],pp15[37],pp15[38],pp15[39],pp15[40],pp15[41],pp15[42],pp15[43],pp15[44],pp15[45],pp15[46],pp15[47],pp15[48],pp17[47],pp19[46],pp21[45],pp23[44],pp25[43],pp27[42],pp29[41],pp31[40],pp33[39],pp35[38],pp37[37],pp39[36],pp41[35],pp43[34],pp45[33],pp47[32],pp49[31],pp51[30],pp53[29],pp55[28],pp57[27],pp59[26],pp61[25],pp63[24],pp65[23],pp67[22],pp69[21],pp71[20],pp73[19],pp75[18],pp77[17],pp79[16],pp81[15],pp83[14],pp85[13],pp87[12],pp88[12],pp89[12],pp90[12],pp91[12],pp92[12],pp93[12],pp94[12],pp95[12],pp96[12],pp97[12],pp98[12],pp99[12],pp103[9],pp105[8],pp107[7],pp109[6],pp111[5],pp113[4],pp115[3],pp117[2],pp119[1],pp121[0],s129[58],s130[58],s131[58],s132[58],s133[58],s134[58],s135[58],s136[58],s137[58],s138[58],s138[59],s138[60],s139[60],s140[60],s141[60],s142[60],s143[60],s144[60],s145[60],s146[60],s147[60],s148[60],s149[60],s150[60],s151[60],s152[60],s153[60],s154[60],s155[60],s156[60],s157[60],s158[60],s159[60],s160[60],s161[60],s162[60],s163[60],s164[60],s165[60],s166[60],s167[60],s168[60],s169[60],s170[60],s171[60],s172[60],s173[60],s174[60],s175[60],s176[60],s177[60],s178[60],s179[60],s180[60],s181[60],s182[60],s183[60],s184[60],s185[60],s186[60],s187[60],s188[60],s189[60],s190[60],s191[60],s192[60],s10[51],s11[51],s12[51],s13[51],s14[51],s15[51],s16[51],s17[51],s18[51],s19[51],s20[51],s21[51],s22[51],s23[51],s24[51],s25[51],s26[51],s27[51],s28[51],s29[51],s30[51],s31[51],s32[51],s33[51],s34[51],s35[51],s36[51],s37[51],s38[51],s39[51],s40[51],s41[51],s42[51],s43[51],s44[51],s45[51],s46[51],s47[51],s48[51],s49[51],s49[52],s49[53],s49[54],s49[55],s49[56],s49[57],s49[58],s49[59],s49[60],s49[61],s49[62],s49[63],s49[64],s49[65],s49[66],s49[67],s49[68],s49[69],s49[70],s49[71],s49[72],s49[73],s49[74],s49[75],s49[76],s49[77],s49[78],s49[79],s49[80],s47[83],s45[86],s43[89],s41[92],s40[94],s40[95],s40[96],s40[97],s40[98],s40[99],s9[131],s8[133],s7[135],s6[137],s5[139],s4[141],s3[143],s2[145],s1[147],s108[41],s106[44],s104[47],s102[50],s100[53],s53[101],s52[103],s51[105],s50[107],s49[109],s48[111],s47[113],s46[115],s45[117],s44[119],s43[121],s42[123],s41[125],s40[127],s39[129],s38[131],s37[133],s36[135],s35[137],s34[139],s33[141],s32[143],s31[145],s30[147],s29[149],s28[151],s27[153],s26[155],s25[157],s24[159],s23[161],s22[163],s21[165],s20[167],s19[169],s18[171],s17[173],s16[175],s15[177],s14[179],s13[181],s12[183],s11[185],s10[187],s194[292],s193[294],s192[200],s191[202],s190[204],s189[206],s188[208],s187[210],s186[212],s185[214],s184[216],s183[218],s182[220],s181[222],s180[224],s179[226],s178[228],s177[230],s176[232],s175[234],s174[236],s173[238],s172[240],s171[242],s170[244],s169[246],s168[248],s167[250],s166[252],s165[254],s164[256],s163[258],s162[260],s161[262],s160[264],s159[266],s158[268],s157[270],s156[272],s155[274],s154[276],s153[278],s152[280],s151[282],s150[284],s149[286],s148[288],s147[290],s146[292],s145[294],s144[296],s143[298],s142[300],s141[302],s140[304],s139[306],s138[308],s137[310],s136[312],s135[314],s134[316],s133[318],s132[320],s131[322],s130[324],s129[326],pp255[136],pp254[138],pp253[140],pp252[142],pp251[144],pp250[146],pp249[148],pp248[150],pp247[152],pp246[154],pp245[156],pp244[158],pp243[160],pp242[162],pp241[164],pp240[166],pp239[168],pp238[170],pp237[172],pp236[174],pp235[176],pp234[178],pp233[180],pp232[182],pp231[184],pp230[186],pp229[188],pp228[190],pp227[192],pp226[194],pp225[196],pp224[198],pp223[200],pp222[202],pp221[204],pp220[206],pp219[208],pp218[210],pp217[212],pp216[214],pp215[216],pp214[218],pp213[220],pp212[222],pp211[224],pp210[226],pp209[228],pp208[230],pp207[232],pp206[234],pp205[236],pp204[238],pp203[240],pp202[242],pp201[244],pp200[246],pp199[248],pp198[250],pp199[250],pp200[250],pp201[250],pp202[250],pp203[250],pp204[250],pp205[250],pp206[250],pp207[250],pp208[250],pp209[250],pp210[250],pp211[250],pp212[250],pp213[250],pp214[250],pp215[250],pp216[250],pp217[250],pp218[250],pp219[250],pp220[250],pp221[250],pp222[250],pp223[250],pp224[250],pp225[250],pp226[250],pp227[250]};
    CLA_444 KS_195(s195, c195, in195_1, in195_2);
    wire[441:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp16[19],pp16[20],pp16[21],pp16[22],pp16[23],pp16[24],pp16[25],pp16[26],pp16[27],pp16[28],pp16[29],pp16[30],pp16[31],pp16[32],pp16[33],pp16[34],pp16[35],pp16[36],pp16[37],pp16[38],pp16[39],pp16[40],pp16[41],pp16[42],pp16[43],pp16[44],pp16[45],pp16[46],pp16[47],pp18[46],pp20[45],pp22[44],pp24[43],pp26[42],pp28[41],pp30[40],pp32[39],pp34[38],pp36[37],pp38[36],pp40[35],pp42[34],pp44[33],pp46[32],pp48[31],pp50[30],pp52[29],pp54[28],pp56[27],pp58[26],pp60[25],pp62[24],pp64[23],pp66[22],pp68[21],pp70[20],pp72[19],pp74[18],pp76[17],pp78[16],pp80[15],pp82[14],pp84[13],pp86[12],pp88[11],pp89[11],pp90[11],pp91[11],pp92[11],pp93[11],pp94[11],pp95[11],pp96[11],pp97[11],pp98[11],pp99[11],pp102[9],pp104[8],pp106[7],pp108[6],pp110[5],pp112[4],pp114[3],pp116[2],pp118[1],pp120[0],s129[57],s130[57],s131[57],s132[57],s133[57],s134[57],s135[57],s136[57],s137[57],s138[57],s139[57],s139[58],s139[59],s195[100],s195[101],s195[102],s195[103],s195[104],s195[105],s195[106],s195[107],s195[108],s195[109],s195[110],s195[111],s195[112],s195[113],s195[114],s195[115],s195[116],s195[117],s195[118],s195[119],s195[120],s195[121],s195[122],s195[123],s195[124],s195[125],s195[126],s195[127],s195[128],s195[129],s195[130],s195[131],s195[132],s195[133],s195[134],s195[135],s195[136],s195[137],s195[138],s195[139],s195[140],s195[141],s195[142],s195[143],s195[144],s195[145],s195[146],s195[147],s195[148],s195[149],s195[150],s195[151],s195[152],s195[153],s195[154],s195[155],s195[156],s195[157],s195[158],s195[159],s195[160],s195[161],s195[162],s195[163],s195[164],s195[165],s195[166],s195[167],s195[168],s195[169],s195[170],s195[171],s195[172],s195[173],s195[174],s195[175],s195[176],s195[177],s195[178],s195[179],s195[180],s195[181],s195[182],s195[183],s195[184],s195[185],s195[186],s195[187],s195[188],s195[189],s195[190],s195[191],s195[192],s195[193],s195[194],s195[195],s195[196],s195[197],s195[198],s195[199],s195[200],s195[201],s195[202],s195[203],s195[204],s195[205],s195[206],s195[207],s195[208],s195[209],s195[210],s195[211],s195[212],s195[213],s195[214],s195[215],s195[216],s195[217],s195[218],s195[219],s195[220],s195[221],s195[222],s195[223],s195[224],s195[225],s195[226],s195[227],s195[228],s195[229],s195[230],s195[231],s195[232],s195[233],s195[234],s195[235],s195[236],s195[237],s195[238],s195[239],s195[240],s195[241],s195[242],s195[243],s195[244],s195[245],s195[246],s195[247],s195[248],s195[249],s195[250],s195[251],s195[252],s195[253],s195[254],s195[255],s195[256],s195[257],s195[258],s195[259],s195[260],s195[261],s195[262],s195[263],s195[264],s195[265],s195[266],s195[267],s195[268],s195[269],s195[270],s195[271],s195[272],s195[273],s195[274],s195[275],s195[276],s195[277],s195[278],s195[279],s195[280],s195[281],s195[282],s195[283],s195[284],s195[285],s195[286],s195[287],s195[288],s195[289],s195[290],s195[291],s194[293],s193[295],s192[201],s191[203],s190[205],s189[207],s188[209],s187[211],s186[213],s185[215],s184[217],s183[219],s182[221],s181[223],s180[225],s179[227],s178[229],s177[231],s176[233],s175[235],s174[237],s173[239],s172[241],s171[243],s170[245],s169[247],s168[249],s167[251],s166[253],s165[255],s164[257],s163[259],s162[261],s161[263],s160[265],s159[267],s158[269],s157[271],s156[273],s155[275],s154[277],s153[279],s152[281],s151[283],s150[285],s149[287],s148[289],s147[291],s146[293],s145[295],s144[297],s143[299],s142[301],s141[303],s140[305],s139[307],s138[309],s137[311],s136[313],s135[315],s134[317],s133[319],s132[321],s131[323],s130[325],s129[327],pp255[137],pp254[139],pp253[141],pp252[143],pp251[145],pp250[147],pp249[149],pp248[151],pp247[153],pp246[155],pp245[157],pp244[159],pp243[161],pp242[163],pp241[165],pp240[167],pp239[169],pp238[171],pp237[173],pp236[175],pp235[177],pp234[179],pp233[181],pp232[183],pp231[185],pp230[187],pp229[189],pp228[191],pp227[193],pp226[195],pp225[197],pp224[199],pp223[201],pp222[203],pp221[205],pp220[207],pp219[209],pp218[211],pp217[213],pp216[215],pp215[217],pp214[219],pp213[221],pp212[223],pp211[225],pp210[227],pp209[229],pp208[231],pp207[233],pp206[235],pp205[237],pp204[239],pp203[241],pp202[243],pp201[245],pp200[247],pp199[249],pp200[249],pp201[249],pp202[249],pp203[249],pp204[249],pp205[249],pp206[249],pp207[249],pp208[249],pp209[249],pp210[249],pp211[249],pp212[249],pp213[249],pp214[249],pp215[249],pp216[249],pp217[249],pp218[249],pp219[249],pp220[249],pp221[249],pp222[249],pp223[249],pp224[249],pp225[249],pp226[249],pp227[249]};
    assign in196_2 = {pp17[18],pp17[19],pp17[20],pp17[21],pp17[22],pp17[23],pp17[24],pp17[25],pp17[26],pp17[27],pp17[28],pp17[29],pp17[30],pp17[31],pp17[32],pp17[33],pp17[34],pp17[35],pp17[36],pp17[37],pp17[38],pp17[39],pp17[40],pp17[41],pp17[42],pp17[43],pp17[44],pp17[45],pp17[46],pp19[45],pp21[44],pp23[43],pp25[42],pp27[41],pp29[40],pp31[39],pp33[38],pp35[37],pp37[36],pp39[35],pp41[34],pp43[33],pp45[32],pp47[31],pp49[30],pp51[29],pp53[28],pp55[27],pp57[26],pp59[25],pp61[24],pp63[23],pp65[22],pp67[21],pp69[20],pp71[19],pp73[18],pp75[17],pp77[16],pp79[15],pp81[14],pp83[13],pp85[12],pp87[11],pp89[10],pp90[10],pp91[10],pp92[10],pp93[10],pp94[10],pp95[10],pp96[10],pp97[10],pp98[10],pp99[10],pp101[9],pp103[8],pp105[7],pp107[6],pp109[5],pp111[4],pp113[3],pp115[2],pp117[1],pp119[0],s129[56],s130[56],s131[56],s132[56],s133[56],s134[56],s135[56],s136[56],s137[56],s138[56],s139[56],s140[56],s140[57],s140[58],s140[59],s141[59],s142[59],s143[59],s144[59],s145[59],s146[59],s147[59],s148[59],s149[59],s150[59],s151[59],s152[59],s153[59],s154[59],s155[59],s156[59],s157[59],s158[59],s159[59],s160[59],s161[59],s162[59],s163[59],s164[59],s165[59],s166[59],s167[59],s168[59],s169[59],s170[59],s171[59],s172[59],s173[59],s174[59],s175[59],s176[59],s177[59],s178[59],s179[59],s180[59],s181[59],s182[59],s183[59],s184[59],s185[59],s186[59],s187[59],s188[59],s189[59],s190[59],s191[59],s192[59],s10[50],s11[50],s12[50],s13[50],s14[50],s15[50],s16[50],s17[50],s18[50],s19[50],s20[50],s21[50],s22[50],s23[50],s24[50],s25[50],s26[50],s27[50],s28[50],s29[50],s30[50],s31[50],s32[50],s33[50],s34[50],s35[50],s36[50],s37[50],s38[50],s39[50],s40[50],s41[50],s42[50],s43[50],s44[50],s45[50],s46[50],s47[50],s48[50],s49[50],s50[50],s50[51],s50[52],s50[53],s50[54],s50[55],s50[56],s50[57],s50[58],s50[59],s50[60],s50[61],s50[62],s50[63],s50[64],s50[65],s50[66],s50[67],s50[68],s50[69],s50[70],s50[71],s50[72],s50[73],s50[74],s50[75],s50[76],s50[77],s50[78],s50[79],s48[82],s46[85],s44[88],s42[91],s41[93],s41[94],s41[95],s41[96],s41[97],s41[98],s41[99],s9[132],s8[134],s7[136],s6[138],s5[140],s4[142],s3[144],s2[146],s1[148],s107[43],s105[46],s103[49],s101[52],s54[100],s53[102],s52[104],s51[106],s50[108],s49[110],s48[112],s47[114],s46[116],s45[118],s44[120],s43[122],s42[124],s41[126],s40[128],s39[130],s38[132],s37[134],s36[136],s35[138],s34[140],s33[142],s32[144],s31[146],s30[148],s29[150],s28[152],s27[154],s26[156],s25[158],s24[160],s23[162],s22[164],s21[166],s20[168],s19[170],s18[172],s17[174],s16[176],s15[178],s14[180],s13[182],s12[184],s11[186],s10[188],s195[292],s194[294],s193[296],s192[202],s191[204],s190[206],s189[208],s188[210],s187[212],s186[214],s185[216],s184[218],s183[220],s182[222],s181[224],s180[226],s179[228],s178[230],s177[232],s176[234],s175[236],s174[238],s173[240],s172[242],s171[244],s170[246],s169[248],s168[250],s167[252],s166[254],s165[256],s164[258],s163[260],s162[262],s161[264],s160[266],s159[268],s158[270],s157[272],s156[274],s155[276],s154[278],s153[280],s152[282],s151[284],s150[286],s149[288],s148[290],s147[292],s146[294],s145[296],s144[298],s143[300],s142[302],s141[304],s140[306],s139[308],s138[310],s137[312],s136[314],s135[316],s134[318],s133[320],s132[322],s131[324],s130[326],s129[328],pp255[138],pp254[140],pp253[142],pp252[144],pp251[146],pp250[148],pp249[150],pp248[152],pp247[154],pp246[156],pp245[158],pp244[160],pp243[162],pp242[164],pp241[166],pp240[168],pp239[170],pp238[172],pp237[174],pp236[176],pp235[178],pp234[180],pp233[182],pp232[184],pp231[186],pp230[188],pp229[190],pp228[192],pp227[194],pp226[196],pp225[198],pp224[200],pp223[202],pp222[204],pp221[206],pp220[208],pp219[210],pp218[212],pp217[214],pp216[216],pp215[218],pp214[220],pp213[222],pp212[224],pp211[226],pp210[228],pp209[230],pp208[232],pp207[234],pp206[236],pp205[238],pp204[240],pp203[242],pp202[244],pp201[246],pp200[248],pp201[248],pp202[248],pp203[248],pp204[248],pp205[248],pp206[248],pp207[248],pp208[248],pp209[248],pp210[248],pp211[248],pp212[248],pp213[248],pp214[248],pp215[248],pp216[248],pp217[248],pp218[248],pp219[248],pp220[248],pp221[248],pp222[248],pp223[248],pp224[248],pp225[248],pp226[248],pp227[248],pp228[248]};
    CLA_442 KS_196(s196, c196, in196_1, in196_2);
    wire[439:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {pp18[18],pp18[19],pp18[20],pp18[21],pp18[22],pp18[23],pp18[24],pp18[25],pp18[26],pp18[27],pp18[28],pp18[29],pp18[30],pp18[31],pp18[32],pp18[33],pp18[34],pp18[35],pp18[36],pp18[37],pp18[38],pp18[39],pp18[40],pp18[41],pp18[42],pp18[43],pp18[44],pp18[45],pp20[44],pp22[43],pp24[42],pp26[41],pp28[40],pp30[39],pp32[38],pp34[37],pp36[36],pp38[35],pp40[34],pp42[33],pp44[32],pp46[31],pp48[30],pp50[29],pp52[28],pp54[27],pp56[26],pp58[25],pp60[24],pp62[23],pp64[22],pp66[21],pp68[20],pp70[19],pp72[18],pp74[17],pp76[16],pp78[15],pp80[14],pp82[13],pp84[12],pp86[11],pp88[10],s129[35],pp100[0],pp100[1],pp100[2],pp100[3],pp100[4],pp100[5],pp100[6],pp100[7],pp100[8],pp100[9],pp102[8],pp104[7],pp106[6],pp108[5],pp110[4],pp112[3],pp114[2],pp116[1],pp118[0],s129[55],s130[55],s131[55],s132[55],s133[55],s134[55],s135[55],s136[55],s137[55],s138[55],s139[55],s140[55],s141[55],s141[56],s141[57],s141[58],s196[100],s196[101],s196[102],s196[103],s196[104],s196[105],s196[106],s196[107],s196[108],s196[109],s196[110],s196[111],s196[112],s196[113],s196[114],s196[115],s196[116],s196[117],s196[118],s196[119],s196[120],s196[121],s196[122],s196[123],s196[124],s196[125],s196[126],s196[127],s196[128],s196[129],s196[130],s196[131],s196[132],s196[133],s196[134],s196[135],s196[136],s196[137],s196[138],s196[139],s196[140],s196[141],s196[142],s196[143],s196[144],s196[145],s196[146],s196[147],s196[148],s196[149],s196[150],s196[151],s196[152],s196[153],s196[154],s196[155],s196[156],s196[157],s196[158],s196[159],s196[160],s196[161],s196[162],s196[163],s196[164],s196[165],s196[166],s196[167],s196[168],s196[169],s196[170],s196[171],s196[172],s196[173],s196[174],s196[175],s196[176],s196[177],s196[178],s196[179],s196[180],s196[181],s196[182],s196[183],s196[184],s196[185],s196[186],s196[187],s196[188],s196[189],s196[190],s196[191],s196[192],s196[193],s196[194],s196[195],s196[196],s196[197],s196[198],s196[199],s196[200],s196[201],s196[202],s196[203],s196[204],s196[205],s196[206],s196[207],s196[208],s196[209],s196[210],s196[211],s196[212],s196[213],s196[214],s196[215],s196[216],s196[217],s196[218],s196[219],s196[220],s196[221],s196[222],s196[223],s196[224],s196[225],s196[226],s196[227],s196[228],s196[229],s196[230],s196[231],s196[232],s196[233],s196[234],s196[235],s196[236],s196[237],s196[238],s196[239],s196[240],s196[241],s196[242],s196[243],s196[244],s196[245],s196[246],s196[247],s196[248],s196[249],s196[250],s196[251],s196[252],s196[253],s196[254],s196[255],s196[256],s196[257],s196[258],s196[259],s196[260],s196[261],s196[262],s196[263],s196[264],s196[265],s196[266],s196[267],s196[268],s196[269],s196[270],s196[271],s196[272],s196[273],s196[274],s196[275],s196[276],s196[277],s196[278],s196[279],s196[280],s196[281],s196[282],s196[283],s196[284],s196[285],s196[286],s196[287],s196[288],s196[289],s196[290],s196[291],s195[293],s194[295],s193[297],s192[203],s191[205],s190[207],s189[209],s188[211],s187[213],s186[215],s185[217],s184[219],s183[221],s182[223],s181[225],s180[227],s179[229],s178[231],s177[233],s176[235],s175[237],s174[239],s173[241],s172[243],s171[245],s170[247],s169[249],s168[251],s167[253],s166[255],s165[257],s164[259],s163[261],s162[263],s161[265],s160[267],s159[269],s158[271],s157[273],s156[275],s155[277],s154[279],s153[281],s152[283],s151[285],s150[287],s149[289],s148[291],s147[293],s146[295],s145[297],s144[299],s143[301],s142[303],s141[305],s140[307],s139[309],s138[311],s137[313],s136[315],s135[317],s134[319],s133[321],s132[323],s131[325],s130[327],s129[329],pp255[139],pp254[141],pp253[143],pp252[145],pp251[147],pp250[149],pp249[151],pp248[153],pp247[155],pp246[157],pp245[159],pp244[161],pp243[163],pp242[165],pp241[167],pp240[169],pp239[171],pp238[173],pp237[175],pp236[177],pp235[179],pp234[181],pp233[183],pp232[185],pp231[187],pp230[189],pp229[191],pp228[193],pp227[195],pp226[197],pp225[199],pp224[201],pp223[203],pp222[205],pp221[207],pp220[209],pp219[211],pp218[213],pp217[215],pp216[217],pp215[219],pp214[221],pp213[223],pp212[225],pp211[227],pp210[229],pp209[231],pp208[233],pp207[235],pp206[237],pp205[239],pp204[241],pp203[243],pp202[245],pp201[247],pp202[247],pp203[247],pp204[247],pp205[247],pp206[247],pp207[247],pp208[247],pp209[247],pp210[247],pp211[247],pp212[247],pp213[247],pp214[247],pp215[247],pp216[247],pp217[247],pp218[247],pp219[247],pp220[247],pp221[247],pp222[247],pp223[247],pp224[247],pp225[247],pp226[247],pp227[247],pp228[247]};
    assign in197_2 = {pp19[17],pp19[18],pp19[19],pp19[20],pp19[21],pp19[22],pp19[23],pp19[24],pp19[25],pp19[26],pp19[27],pp19[28],pp19[29],pp19[30],pp19[31],pp19[32],pp19[33],pp19[34],pp19[35],pp19[36],pp19[37],pp19[38],pp19[39],pp19[40],pp19[41],pp19[42],pp19[43],pp19[44],pp21[43],pp23[42],pp25[41],pp27[40],pp29[39],pp31[38],pp33[37],pp35[36],pp37[35],pp39[34],pp41[33],pp43[32],pp45[31],pp47[30],pp49[29],pp51[28],pp53[27],pp55[26],pp57[25],pp59[24],pp61[23],pp63[22],pp65[21],pp67[20],pp69[19],pp71[18],pp73[17],pp75[16],pp77[15],pp79[14],pp81[13],pp83[12],pp85[11],pp87[10],s129[34],s130[34],s129[36],pp101[0],pp101[1],pp101[2],pp101[3],pp101[4],pp101[5],pp101[6],pp101[7],pp101[8],pp103[7],pp105[6],pp107[5],pp109[4],pp111[3],pp113[2],pp115[1],pp117[0],s129[54],s130[54],s131[54],s132[54],s133[54],s134[54],s135[54],s136[54],s137[54],s138[54],s139[54],s140[54],s141[54],s142[54],s142[55],s142[56],s142[57],s142[58],s143[58],s144[58],s145[58],s146[58],s147[58],s148[58],s149[58],s150[58],s151[58],s152[58],s153[58],s154[58],s155[58],s156[58],s157[58],s158[58],s159[58],s160[58],s161[58],s162[58],s163[58],s164[58],s165[58],s166[58],s167[58],s168[58],s169[58],s170[58],s171[58],s172[58],s173[58],s174[58],s175[58],s176[58],s177[58],s178[58],s179[58],s180[58],s181[58],s182[58],s183[58],s184[58],s185[58],s186[58],s187[58],s188[58],s189[58],s190[58],s191[58],s192[58],s10[49],s11[49],s12[49],s13[49],s14[49],s15[49],s16[49],s17[49],s18[49],s19[49],s20[49],s21[49],s22[49],s23[49],s24[49],s25[49],s26[49],s27[49],s28[49],s29[49],s30[49],s31[49],s32[49],s33[49],s34[49],s35[49],s36[49],s37[49],s38[49],s39[49],s40[49],s41[49],s42[49],s43[49],s44[49],s45[49],s46[49],s47[49],s48[49],s49[49],s50[49],s51[49],s51[50],s51[51],s51[52],s51[53],s51[54],s51[55],s51[56],s51[57],s51[58],s51[59],s51[60],s51[61],s51[62],s51[63],s51[64],s51[65],s51[66],s51[67],s51[68],s51[69],s51[70],s51[71],s51[72],s51[73],s51[74],s51[75],s51[76],s51[77],s51[78],s49[81],s47[84],s45[87],s43[90],s42[92],s42[93],s42[94],s42[95],s42[96],s42[97],s42[98],s42[99],s9[133],s8[135],s7[137],s6[139],s5[141],s4[143],s3[145],s2[147],s1[149],s106[45],s104[48],s102[51],s100[54],s54[101],s53[103],s52[105],s51[107],s50[109],s49[111],s48[113],s47[115],s46[117],s45[119],s44[121],s43[123],s42[125],s41[127],s40[129],s39[131],s38[133],s37[135],s36[137],s35[139],s34[141],s33[143],s32[145],s31[147],s30[149],s29[151],s28[153],s27[155],s26[157],s25[159],s24[161],s23[163],s22[165],s21[167],s20[169],s19[171],s18[173],s17[175],s16[177],s15[179],s14[181],s13[183],s12[185],s11[187],s10[189],s196[292],s195[294],s194[296],s193[298],s192[204],s191[206],s190[208],s189[210],s188[212],s187[214],s186[216],s185[218],s184[220],s183[222],s182[224],s181[226],s180[228],s179[230],s178[232],s177[234],s176[236],s175[238],s174[240],s173[242],s172[244],s171[246],s170[248],s169[250],s168[252],s167[254],s166[256],s165[258],s164[260],s163[262],s162[264],s161[266],s160[268],s159[270],s158[272],s157[274],s156[276],s155[278],s154[280],s153[282],s152[284],s151[286],s150[288],s149[290],s148[292],s147[294],s146[296],s145[298],s144[300],s143[302],s142[304],s141[306],s140[308],s139[310],s138[312],s137[314],s136[316],s135[318],s134[320],s133[322],s132[324],s131[326],s130[328],s129[330],pp255[140],pp254[142],pp253[144],pp252[146],pp251[148],pp250[150],pp249[152],pp248[154],pp247[156],pp246[158],pp245[160],pp244[162],pp243[164],pp242[166],pp241[168],pp240[170],pp239[172],pp238[174],pp237[176],pp236[178],pp235[180],pp234[182],pp233[184],pp232[186],pp231[188],pp230[190],pp229[192],pp228[194],pp227[196],pp226[198],pp225[200],pp224[202],pp223[204],pp222[206],pp221[208],pp220[210],pp219[212],pp218[214],pp217[216],pp216[218],pp215[220],pp214[222],pp213[224],pp212[226],pp211[228],pp210[230],pp209[232],pp208[234],pp207[236],pp206[238],pp205[240],pp204[242],pp203[244],pp202[246],pp203[246],pp204[246],pp205[246],pp206[246],pp207[246],pp208[246],pp209[246],pp210[246],pp211[246],pp212[246],pp213[246],pp214[246],pp215[246],pp216[246],pp217[246],pp218[246],pp219[246],pp220[246],pp221[246],pp222[246],pp223[246],pp224[246],pp225[246],pp226[246],pp227[246],pp228[246],pp229[246]};
    CLA_440 KS_197(s197, c197, in197_1, in197_2);
    wire[437:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {pp20[17],pp20[18],pp20[19],pp20[20],pp20[21],pp20[22],pp20[23],pp20[24],pp20[25],pp20[26],pp20[27],pp20[28],pp20[29],pp20[30],pp20[31],pp20[32],pp20[33],pp20[34],pp20[35],pp20[36],pp20[37],pp20[38],pp20[39],pp20[40],pp20[41],pp20[42],pp20[43],pp22[42],pp24[41],pp26[40],pp28[39],pp30[38],pp32[37],pp34[36],pp36[35],pp38[34],pp40[33],pp42[32],pp44[31],pp46[30],pp48[29],pp50[28],pp52[27],pp54[26],pp56[25],pp58[24],pp60[23],pp62[22],pp64[21],pp66[20],pp68[19],pp70[18],pp72[17],pp74[16],pp76[15],pp78[14],pp80[13],pp82[12],pp84[11],pp86[10],s129[33],s130[33],s131[33],s130[35],s129[37],pp102[0],pp102[1],pp102[2],pp102[3],pp102[4],pp102[5],pp102[6],pp102[7],pp104[6],pp106[5],pp108[4],pp110[3],pp112[2],pp114[1],pp116[0],s129[53],s130[53],s131[53],s132[53],s133[53],s134[53],s135[53],s136[53],s137[53],s138[53],s139[53],s140[53],s141[53],s142[53],s143[53],s143[54],s143[55],s143[56],s143[57],s197[100],s197[101],s197[102],s197[103],s197[104],s197[105],s197[106],s197[107],s197[108],s197[109],s197[110],s197[111],s197[112],s197[113],s197[114],s197[115],s197[116],s197[117],s197[118],s197[119],s197[120],s197[121],s197[122],s197[123],s197[124],s197[125],s197[126],s197[127],s197[128],s197[129],s197[130],s197[131],s197[132],s197[133],s197[134],s197[135],s197[136],s197[137],s197[138],s197[139],s197[140],s197[141],s197[142],s197[143],s197[144],s197[145],s197[146],s197[147],s197[148],s197[149],s197[150],s197[151],s197[152],s197[153],s197[154],s197[155],s197[156],s197[157],s197[158],s197[159],s197[160],s197[161],s197[162],s197[163],s197[164],s197[165],s197[166],s197[167],s197[168],s197[169],s197[170],s197[171],s197[172],s197[173],s197[174],s197[175],s197[176],s197[177],s197[178],s197[179],s197[180],s197[181],s197[182],s197[183],s197[184],s197[185],s197[186],s197[187],s197[188],s197[189],s197[190],s197[191],s197[192],s197[193],s197[194],s197[195],s197[196],s197[197],s197[198],s197[199],s197[200],s197[201],s197[202],s197[203],s197[204],s197[205],s197[206],s197[207],s197[208],s197[209],s197[210],s197[211],s197[212],s197[213],s197[214],s197[215],s197[216],s197[217],s197[218],s197[219],s197[220],s197[221],s197[222],s197[223],s197[224],s197[225],s197[226],s197[227],s197[228],s197[229],s197[230],s197[231],s197[232],s197[233],s197[234],s197[235],s197[236],s197[237],s197[238],s197[239],s197[240],s197[241],s197[242],s197[243],s197[244],s197[245],s197[246],s197[247],s197[248],s197[249],s197[250],s197[251],s197[252],s197[253],s197[254],s197[255],s197[256],s197[257],s197[258],s197[259],s197[260],s197[261],s197[262],s197[263],s197[264],s197[265],s197[266],s197[267],s197[268],s197[269],s197[270],s197[271],s197[272],s197[273],s197[274],s197[275],s197[276],s197[277],s197[278],s197[279],s197[280],s197[281],s197[282],s197[283],s197[284],s197[285],s197[286],s197[287],s197[288],s197[289],s197[290],s197[291],s196[293],s195[295],s194[297],s193[299],s192[205],s191[207],s190[209],s189[211],s188[213],s187[215],s186[217],s185[219],s184[221],s183[223],s182[225],s181[227],s180[229],s179[231],s178[233],s177[235],s176[237],s175[239],s174[241],s173[243],s172[245],s171[247],s170[249],s169[251],s168[253],s167[255],s166[257],s165[259],s164[261],s163[263],s162[265],s161[267],s160[269],s159[271],s158[273],s157[275],s156[277],s155[279],s154[281],s153[283],s152[285],s151[287],s150[289],s149[291],s148[293],s147[295],s146[297],s145[299],s144[301],s143[303],s142[305],s141[307],s140[309],s139[311],s138[313],s137[315],s136[317],s135[319],s134[321],s133[323],s132[325],s131[327],s130[329],s129[331],pp255[141],pp254[143],pp253[145],pp252[147],pp251[149],pp250[151],pp249[153],pp248[155],pp247[157],pp246[159],pp245[161],pp244[163],pp243[165],pp242[167],pp241[169],pp240[171],pp239[173],pp238[175],pp237[177],pp236[179],pp235[181],pp234[183],pp233[185],pp232[187],pp231[189],pp230[191],pp229[193],pp228[195],pp227[197],pp226[199],pp225[201],pp224[203],pp223[205],pp222[207],pp221[209],pp220[211],pp219[213],pp218[215],pp217[217],pp216[219],pp215[221],pp214[223],pp213[225],pp212[227],pp211[229],pp210[231],pp209[233],pp208[235],pp207[237],pp206[239],pp205[241],pp204[243],pp203[245],pp204[245],pp205[245],pp206[245],pp207[245],pp208[245],pp209[245],pp210[245],pp211[245],pp212[245],pp213[245],pp214[245],pp215[245],pp216[245],pp217[245],pp218[245],pp219[245],pp220[245],pp221[245],pp222[245],pp223[245],pp224[245],pp225[245],pp226[245],pp227[245],pp228[245],pp229[245]};
    assign in198_2 = {pp21[16],pp21[17],pp21[18],pp21[19],pp21[20],pp21[21],pp21[22],pp21[23],pp21[24],pp21[25],pp21[26],pp21[27],pp21[28],pp21[29],pp21[30],pp21[31],pp21[32],pp21[33],pp21[34],pp21[35],pp21[36],pp21[37],pp21[38],pp21[39],pp21[40],pp21[41],pp21[42],pp23[41],pp25[40],pp27[39],pp29[38],pp31[37],pp33[36],pp35[35],pp37[34],pp39[33],pp41[32],pp43[31],pp45[30],pp47[29],pp49[28],pp51[27],pp53[26],pp55[25],pp57[24],pp59[23],pp61[22],pp63[21],pp65[20],pp67[19],pp69[18],pp71[17],pp73[16],pp75[15],pp77[14],pp79[13],pp81[12],pp83[11],pp85[10],s129[32],s130[32],s131[32],s132[32],s131[34],s130[36],s129[38],pp103[0],pp103[1],pp103[2],pp103[3],pp103[4],pp103[5],pp103[6],pp105[5],pp107[4],pp109[3],pp111[2],pp113[1],pp115[0],s129[52],s130[52],s131[52],s132[52],s133[52],s134[52],s135[52],s136[52],s137[52],s138[52],s139[52],s140[52],s141[52],s142[52],s143[52],s144[52],s144[53],s144[54],s144[55],s144[56],s144[57],s145[57],s146[57],s147[57],s148[57],s149[57],s150[57],s151[57],s152[57],s153[57],s154[57],s155[57],s156[57],s157[57],s158[57],s159[57],s160[57],s161[57],s162[57],s163[57],s164[57],s165[57],s166[57],s167[57],s168[57],s169[57],s170[57],s171[57],s172[57],s173[57],s174[57],s175[57],s176[57],s177[57],s178[57],s179[57],s180[57],s181[57],s182[57],s183[57],s184[57],s185[57],s186[57],s187[57],s188[57],s189[57],s190[57],s191[57],s192[57],s10[48],s11[48],s12[48],s13[48],s14[48],s15[48],s16[48],s17[48],s18[48],s19[48],s20[48],s21[48],s22[48],s23[48],s24[48],s25[48],s26[48],s27[48],s28[48],s29[48],s30[48],s31[48],s32[48],s33[48],s34[48],s35[48],s36[48],s37[48],s38[48],s39[48],s40[48],s41[48],s42[48],s43[48],s44[48],s45[48],s46[48],s47[48],s48[48],s49[48],s50[48],s51[48],s52[48],s52[49],s52[50],s52[51],s52[52],s52[53],s52[54],s52[55],s52[56],s52[57],s52[58],s52[59],s52[60],s52[61],s52[62],s52[63],s52[64],s52[65],s52[66],s52[67],s52[68],s52[69],s52[70],s52[71],s52[72],s52[73],s52[74],s52[75],s52[76],s52[77],s50[80],s48[83],s46[86],s44[89],s43[91],s43[92],s43[93],s43[94],s43[95],s43[96],s43[97],s43[98],s43[99],s9[134],s8[136],s7[138],s6[140],s5[142],s4[144],s3[146],s2[148],s1[150],s105[47],s103[50],s101[53],s55[100],s54[102],s53[104],s52[106],s51[108],s50[110],s49[112],s48[114],s47[116],s46[118],s45[120],s44[122],s43[124],s42[126],s41[128],s40[130],s39[132],s38[134],s37[136],s36[138],s35[140],s34[142],s33[144],s32[146],s31[148],s30[150],s29[152],s28[154],s27[156],s26[158],s25[160],s24[162],s23[164],s22[166],s21[168],s20[170],s19[172],s18[174],s17[176],s16[178],s15[180],s14[182],s13[184],s12[186],s11[188],s10[190],s197[292],s196[294],s195[296],s194[298],s193[300],s192[206],s191[208],s190[210],s189[212],s188[214],s187[216],s186[218],s185[220],s184[222],s183[224],s182[226],s181[228],s180[230],s179[232],s178[234],s177[236],s176[238],s175[240],s174[242],s173[244],s172[246],s171[248],s170[250],s169[252],s168[254],s167[256],s166[258],s165[260],s164[262],s163[264],s162[266],s161[268],s160[270],s159[272],s158[274],s157[276],s156[278],s155[280],s154[282],s153[284],s152[286],s151[288],s150[290],s149[292],s148[294],s147[296],s146[298],s145[300],s144[302],s143[304],s142[306],s141[308],s140[310],s139[312],s138[314],s137[316],s136[318],s135[320],s134[322],s133[324],s132[326],s131[328],s130[330],s129[332],pp255[142],pp254[144],pp253[146],pp252[148],pp251[150],pp250[152],pp249[154],pp248[156],pp247[158],pp246[160],pp245[162],pp244[164],pp243[166],pp242[168],pp241[170],pp240[172],pp239[174],pp238[176],pp237[178],pp236[180],pp235[182],pp234[184],pp233[186],pp232[188],pp231[190],pp230[192],pp229[194],pp228[196],pp227[198],pp226[200],pp225[202],pp224[204],pp223[206],pp222[208],pp221[210],pp220[212],pp219[214],pp218[216],pp217[218],pp216[220],pp215[222],pp214[224],pp213[226],pp212[228],pp211[230],pp210[232],pp209[234],pp208[236],pp207[238],pp206[240],pp205[242],pp204[244],pp205[244],pp206[244],pp207[244],pp208[244],pp209[244],pp210[244],pp211[244],pp212[244],pp213[244],pp214[244],pp215[244],pp216[244],pp217[244],pp218[244],pp219[244],pp220[244],pp221[244],pp222[244],pp223[244],pp224[244],pp225[244],pp226[244],pp227[244],pp228[244],pp229[244],pp230[244]};
    CLA_438 KS_198(s198, c198, in198_1, in198_2);
    wire[435:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {pp22[16],pp22[17],pp22[18],pp22[19],pp22[20],pp22[21],pp22[22],pp22[23],pp22[24],pp22[25],pp22[26],pp22[27],pp22[28],pp22[29],pp22[30],pp22[31],pp22[32],pp22[33],pp22[34],pp22[35],pp22[36],pp22[37],pp22[38],pp22[39],pp22[40],pp22[41],pp24[40],pp26[39],pp28[38],pp30[37],pp32[36],pp34[35],pp36[34],pp38[33],pp40[32],pp42[31],pp44[30],pp46[29],pp48[28],pp50[27],pp52[26],pp54[25],pp56[24],pp58[23],pp60[22],pp62[21],pp64[20],pp66[19],pp68[18],pp70[17],pp72[16],pp74[15],pp76[14],pp78[13],pp80[12],pp82[11],pp84[10],s129[31],s130[31],s131[31],s132[31],s133[31],s132[33],s131[35],s130[37],s129[39],pp104[0],pp104[1],pp104[2],pp104[3],pp104[4],pp104[5],pp106[4],pp108[3],pp110[2],pp112[1],pp114[0],s129[51],s130[51],s131[51],s132[51],s133[51],s134[51],s135[51],s136[51],s137[51],s138[51],s139[51],s140[51],s141[51],s142[51],s143[51],s144[51],s145[51],s145[52],s145[53],s145[54],s145[55],s145[56],s198[100],s198[101],s198[102],s198[103],s198[104],s198[105],s198[106],s198[107],s198[108],s198[109],s198[110],s198[111],s198[112],s198[113],s198[114],s198[115],s198[116],s198[117],s198[118],s198[119],s198[120],s198[121],s198[122],s198[123],s198[124],s198[125],s198[126],s198[127],s198[128],s198[129],s198[130],s198[131],s198[132],s198[133],s198[134],s198[135],s198[136],s198[137],s198[138],s198[139],s198[140],s198[141],s198[142],s198[143],s198[144],s198[145],s198[146],s198[147],s198[148],s198[149],s198[150],s198[151],s198[152],s198[153],s198[154],s198[155],s198[156],s198[157],s198[158],s198[159],s198[160],s198[161],s198[162],s198[163],s198[164],s198[165],s198[166],s198[167],s198[168],s198[169],s198[170],s198[171],s198[172],s198[173],s198[174],s198[175],s198[176],s198[177],s198[178],s198[179],s198[180],s198[181],s198[182],s198[183],s198[184],s198[185],s198[186],s198[187],s198[188],s198[189],s198[190],s198[191],s198[192],s198[193],s198[194],s198[195],s198[196],s198[197],s198[198],s198[199],s198[200],s198[201],s198[202],s198[203],s198[204],s198[205],s198[206],s198[207],s198[208],s198[209],s198[210],s198[211],s198[212],s198[213],s198[214],s198[215],s198[216],s198[217],s198[218],s198[219],s198[220],s198[221],s198[222],s198[223],s198[224],s198[225],s198[226],s198[227],s198[228],s198[229],s198[230],s198[231],s198[232],s198[233],s198[234],s198[235],s198[236],s198[237],s198[238],s198[239],s198[240],s198[241],s198[242],s198[243],s198[244],s198[245],s198[246],s198[247],s198[248],s198[249],s198[250],s198[251],s198[252],s198[253],s198[254],s198[255],s198[256],s198[257],s198[258],s198[259],s198[260],s198[261],s198[262],s198[263],s198[264],s198[265],s198[266],s198[267],s198[268],s198[269],s198[270],s198[271],s198[272],s198[273],s198[274],s198[275],s198[276],s198[277],s198[278],s198[279],s198[280],s198[281],s198[282],s198[283],s198[284],s198[285],s198[286],s198[287],s198[288],s198[289],s198[290],s198[291],s197[293],s196[295],s195[297],s194[299],s193[301],s192[207],s191[209],s190[211],s189[213],s188[215],s187[217],s186[219],s185[221],s184[223],s183[225],s182[227],s181[229],s180[231],s179[233],s178[235],s177[237],s176[239],s175[241],s174[243],s173[245],s172[247],s171[249],s170[251],s169[253],s168[255],s167[257],s166[259],s165[261],s164[263],s163[265],s162[267],s161[269],s160[271],s159[273],s158[275],s157[277],s156[279],s155[281],s154[283],s153[285],s152[287],s151[289],s150[291],s149[293],s148[295],s147[297],s146[299],s145[301],s144[303],s143[305],s142[307],s141[309],s140[311],s139[313],s138[315],s137[317],s136[319],s135[321],s134[323],s133[325],s132[327],s131[329],s130[331],s129[333],pp255[143],pp254[145],pp253[147],pp252[149],pp251[151],pp250[153],pp249[155],pp248[157],pp247[159],pp246[161],pp245[163],pp244[165],pp243[167],pp242[169],pp241[171],pp240[173],pp239[175],pp238[177],pp237[179],pp236[181],pp235[183],pp234[185],pp233[187],pp232[189],pp231[191],pp230[193],pp229[195],pp228[197],pp227[199],pp226[201],pp225[203],pp224[205],pp223[207],pp222[209],pp221[211],pp220[213],pp219[215],pp218[217],pp217[219],pp216[221],pp215[223],pp214[225],pp213[227],pp212[229],pp211[231],pp210[233],pp209[235],pp208[237],pp207[239],pp206[241],pp205[243],pp206[243],pp207[243],pp208[243],pp209[243],pp210[243],pp211[243],pp212[243],pp213[243],pp214[243],pp215[243],pp216[243],pp217[243],pp218[243],pp219[243],pp220[243],pp221[243],pp222[243],pp223[243],pp224[243],pp225[243],pp226[243],pp227[243],pp228[243],pp229[243],pp230[243]};
    assign in199_2 = {pp23[15],pp23[16],pp23[17],pp23[18],pp23[19],pp23[20],pp23[21],pp23[22],pp23[23],pp23[24],pp23[25],pp23[26],pp23[27],pp23[28],pp23[29],pp23[30],pp23[31],pp23[32],pp23[33],pp23[34],pp23[35],pp23[36],pp23[37],pp23[38],pp23[39],pp23[40],pp25[39],pp27[38],pp29[37],pp31[36],pp33[35],pp35[34],pp37[33],pp39[32],pp41[31],pp43[30],pp45[29],pp47[28],pp49[27],pp51[26],pp53[25],pp55[24],pp57[23],pp59[22],pp61[21],pp63[20],pp65[19],pp67[18],pp69[17],pp71[16],pp73[15],pp75[14],pp77[13],pp79[12],pp81[11],pp83[10],s129[30],s130[30],s131[30],s132[30],s133[30],s134[30],s133[32],s132[34],s131[36],s130[38],s129[40],pp105[0],pp105[1],pp105[2],pp105[3],pp105[4],pp107[3],pp109[2],pp111[1],pp113[0],s129[50],s130[50],s131[50],s132[50],s133[50],s134[50],s135[50],s136[50],s137[50],s138[50],s139[50],s140[50],s141[50],s142[50],s143[50],s144[50],s145[50],s146[50],s146[51],s146[52],s146[53],s146[54],s146[55],s146[56],s147[56],s148[56],s149[56],s150[56],s151[56],s152[56],s153[56],s154[56],s155[56],s156[56],s157[56],s158[56],s159[56],s160[56],s161[56],s162[56],s163[56],s164[56],s165[56],s166[56],s167[56],s168[56],s169[56],s170[56],s171[56],s172[56],s173[56],s174[56],s175[56],s176[56],s177[56],s178[56],s179[56],s180[56],s181[56],s182[56],s183[56],s184[56],s185[56],s186[56],s187[56],s188[56],s189[56],s190[56],s191[56],s192[56],s10[47],s11[47],s12[47],s13[47],s14[47],s15[47],s16[47],s17[47],s18[47],s19[47],s20[47],s21[47],s22[47],s23[47],s24[47],s25[47],s26[47],s27[47],s28[47],s29[47],s30[47],s31[47],s32[47],s33[47],s34[47],s35[47],s36[47],s37[47],s38[47],s39[47],s40[47],s41[47],s42[47],s43[47],s44[47],s45[47],s46[47],s47[47],s48[47],s49[47],s50[47],s51[47],s52[47],s53[47],s53[48],s53[49],s53[50],s53[51],s53[52],s53[53],s53[54],s53[55],s53[56],s53[57],s53[58],s53[59],s53[60],s53[61],s53[62],s53[63],s53[64],s53[65],s53[66],s53[67],s53[68],s53[69],s53[70],s53[71],s53[72],s53[73],s53[74],s53[75],s53[76],s51[79],s49[82],s47[85],s45[88],s44[90],s44[91],s44[92],s44[93],s44[94],s44[95],s44[96],s44[97],s44[98],s44[99],s9[135],s8[137],s7[139],s6[141],s5[143],s4[145],s3[147],s2[149],s1[151],s104[49],s102[52],s100[55],s55[101],s54[103],s53[105],s52[107],s51[109],s50[111],s49[113],s48[115],s47[117],s46[119],s45[121],s44[123],s43[125],s42[127],s41[129],s40[131],s39[133],s38[135],s37[137],s36[139],s35[141],s34[143],s33[145],s32[147],s31[149],s30[151],s29[153],s28[155],s27[157],s26[159],s25[161],s24[163],s23[165],s22[167],s21[169],s20[171],s19[173],s18[175],s17[177],s16[179],s15[181],s14[183],s13[185],s12[187],s11[189],s10[191],s198[292],s197[294],s196[296],s195[298],s194[300],s193[302],s192[208],s191[210],s190[212],s189[214],s188[216],s187[218],s186[220],s185[222],s184[224],s183[226],s182[228],s181[230],s180[232],s179[234],s178[236],s177[238],s176[240],s175[242],s174[244],s173[246],s172[248],s171[250],s170[252],s169[254],s168[256],s167[258],s166[260],s165[262],s164[264],s163[266],s162[268],s161[270],s160[272],s159[274],s158[276],s157[278],s156[280],s155[282],s154[284],s153[286],s152[288],s151[290],s150[292],s149[294],s148[296],s147[298],s146[300],s145[302],s144[304],s143[306],s142[308],s141[310],s140[312],s139[314],s138[316],s137[318],s136[320],s135[322],s134[324],s133[326],s132[328],s131[330],s130[332],s129[334],pp255[144],pp254[146],pp253[148],pp252[150],pp251[152],pp250[154],pp249[156],pp248[158],pp247[160],pp246[162],pp245[164],pp244[166],pp243[168],pp242[170],pp241[172],pp240[174],pp239[176],pp238[178],pp237[180],pp236[182],pp235[184],pp234[186],pp233[188],pp232[190],pp231[192],pp230[194],pp229[196],pp228[198],pp227[200],pp226[202],pp225[204],pp224[206],pp223[208],pp222[210],pp221[212],pp220[214],pp219[216],pp218[218],pp217[220],pp216[222],pp215[224],pp214[226],pp213[228],pp212[230],pp211[232],pp210[234],pp209[236],pp208[238],pp207[240],pp206[242],pp207[242],pp208[242],pp209[242],pp210[242],pp211[242],pp212[242],pp213[242],pp214[242],pp215[242],pp216[242],pp217[242],pp218[242],pp219[242],pp220[242],pp221[242],pp222[242],pp223[242],pp224[242],pp225[242],pp226[242],pp227[242],pp228[242],pp229[242],pp230[242],pp231[242]};
    CLA_436 KS_199(s199, c199, in199_1, in199_2);
    wire[433:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {pp24[15],pp24[16],pp24[17],pp24[18],pp24[19],pp24[20],pp24[21],pp24[22],pp24[23],pp24[24],pp24[25],pp24[26],pp24[27],pp24[28],pp24[29],pp24[30],pp24[31],pp24[32],pp24[33],pp24[34],pp24[35],pp24[36],pp24[37],pp24[38],pp24[39],pp26[38],pp28[37],pp30[36],pp32[35],pp34[34],pp36[33],pp38[32],pp40[31],pp42[30],pp44[29],pp46[28],pp48[27],pp50[26],pp52[25],pp54[24],pp56[23],pp58[22],pp60[21],pp62[20],pp64[19],pp66[18],pp68[17],pp70[16],pp72[15],pp74[14],pp76[13],pp78[12],pp80[11],pp82[10],s129[29],s130[29],s131[29],s132[29],s133[29],s134[29],s135[29],s134[31],s133[33],s132[35],s131[37],s130[39],s129[41],pp106[0],pp106[1],pp106[2],pp106[3],pp108[2],pp110[1],pp112[0],s129[49],s130[49],s131[49],s132[49],s133[49],s134[49],s135[49],s136[49],s137[49],s138[49],s139[49],s140[49],s141[49],s142[49],s143[49],s144[49],s145[49],s146[49],s147[49],s147[50],s147[51],s147[52],s147[53],s147[54],s147[55],s199[100],s199[101],s199[102],s199[103],s199[104],s199[105],s199[106],s199[107],s199[108],s199[109],s199[110],s199[111],s199[112],s199[113],s199[114],s199[115],s199[116],s199[117],s199[118],s199[119],s199[120],s199[121],s199[122],s199[123],s199[124],s199[125],s199[126],s199[127],s199[128],s199[129],s199[130],s199[131],s199[132],s199[133],s199[134],s199[135],s199[136],s199[137],s199[138],s199[139],s199[140],s199[141],s199[142],s199[143],s199[144],s199[145],s199[146],s199[147],s199[148],s199[149],s199[150],s199[151],s199[152],s199[153],s199[154],s199[155],s199[156],s199[157],s199[158],s199[159],s199[160],s199[161],s199[162],s199[163],s199[164],s199[165],s199[166],s199[167],s199[168],s199[169],s199[170],s199[171],s199[172],s199[173],s199[174],s199[175],s199[176],s199[177],s199[178],s199[179],s199[180],s199[181],s199[182],s199[183],s199[184],s199[185],s199[186],s199[187],s199[188],s199[189],s199[190],s199[191],s199[192],s199[193],s199[194],s199[195],s199[196],s199[197],s199[198],s199[199],s199[200],s199[201],s199[202],s199[203],s199[204],s199[205],s199[206],s199[207],s199[208],s199[209],s199[210],s199[211],s199[212],s199[213],s199[214],s199[215],s199[216],s199[217],s199[218],s199[219],s199[220],s199[221],s199[222],s199[223],s199[224],s199[225],s199[226],s199[227],s199[228],s199[229],s199[230],s199[231],s199[232],s199[233],s199[234],s199[235],s199[236],s199[237],s199[238],s199[239],s199[240],s199[241],s199[242],s199[243],s199[244],s199[245],s199[246],s199[247],s199[248],s199[249],s199[250],s199[251],s199[252],s199[253],s199[254],s199[255],s199[256],s199[257],s199[258],s199[259],s199[260],s199[261],s199[262],s199[263],s199[264],s199[265],s199[266],s199[267],s199[268],s199[269],s199[270],s199[271],s199[272],s199[273],s199[274],s199[275],s199[276],s199[277],s199[278],s199[279],s199[280],s199[281],s199[282],s199[283],s199[284],s199[285],s199[286],s199[287],s199[288],s199[289],s199[290],s199[291],s198[293],s197[295],s196[297],s195[299],s194[301],s193[303],s192[209],s191[211],s190[213],s189[215],s188[217],s187[219],s186[221],s185[223],s184[225],s183[227],s182[229],s181[231],s180[233],s179[235],s178[237],s177[239],s176[241],s175[243],s174[245],s173[247],s172[249],s171[251],s170[253],s169[255],s168[257],s167[259],s166[261],s165[263],s164[265],s163[267],s162[269],s161[271],s160[273],s159[275],s158[277],s157[279],s156[281],s155[283],s154[285],s153[287],s152[289],s151[291],s150[293],s149[295],s148[297],s147[299],s146[301],s145[303],s144[305],s143[307],s142[309],s141[311],s140[313],s139[315],s138[317],s137[319],s136[321],s135[323],s134[325],s133[327],s132[329],s131[331],s130[333],s129[335],pp255[145],pp254[147],pp253[149],pp252[151],pp251[153],pp250[155],pp249[157],pp248[159],pp247[161],pp246[163],pp245[165],pp244[167],pp243[169],pp242[171],pp241[173],pp240[175],pp239[177],pp238[179],pp237[181],pp236[183],pp235[185],pp234[187],pp233[189],pp232[191],pp231[193],pp230[195],pp229[197],pp228[199],pp227[201],pp226[203],pp225[205],pp224[207],pp223[209],pp222[211],pp221[213],pp220[215],pp219[217],pp218[219],pp217[221],pp216[223],pp215[225],pp214[227],pp213[229],pp212[231],pp211[233],pp210[235],pp209[237],pp208[239],pp207[241],pp208[241],pp209[241],pp210[241],pp211[241],pp212[241],pp213[241],pp214[241],pp215[241],pp216[241],pp217[241],pp218[241],pp219[241],pp220[241],pp221[241],pp222[241],pp223[241],pp224[241],pp225[241],pp226[241],pp227[241],pp228[241],pp229[241],pp230[241],pp231[241]};
    assign in200_2 = {pp25[14],pp25[15],pp25[16],pp25[17],pp25[18],pp25[19],pp25[20],pp25[21],pp25[22],pp25[23],pp25[24],pp25[25],pp25[26],pp25[27],pp25[28],pp25[29],pp25[30],pp25[31],pp25[32],pp25[33],pp25[34],pp25[35],pp25[36],pp25[37],pp25[38],pp27[37],pp29[36],pp31[35],pp33[34],pp35[33],pp37[32],pp39[31],pp41[30],pp43[29],pp45[28],pp47[27],pp49[26],pp51[25],pp53[24],pp55[23],pp57[22],pp59[21],pp61[20],pp63[19],pp65[18],pp67[17],pp69[16],pp71[15],pp73[14],pp75[13],pp77[12],pp79[11],pp81[10],s129[28],s130[28],s131[28],s132[28],s133[28],s134[28],s135[28],s136[28],s135[30],s134[32],s133[34],s132[36],s131[38],s130[40],s129[42],pp107[0],pp107[1],pp107[2],pp109[1],pp111[0],s129[48],s130[48],s131[48],s132[48],s133[48],s134[48],s135[48],s136[48],s137[48],s138[48],s139[48],s140[48],s141[48],s142[48],s143[48],s144[48],s145[48],s146[48],s147[48],s148[48],s148[49],s148[50],s148[51],s148[52],s148[53],s148[54],s148[55],s149[55],s150[55],s151[55],s152[55],s153[55],s154[55],s155[55],s156[55],s157[55],s158[55],s159[55],s160[55],s161[55],s162[55],s163[55],s164[55],s165[55],s166[55],s167[55],s168[55],s169[55],s170[55],s171[55],s172[55],s173[55],s174[55],s175[55],s176[55],s177[55],s178[55],s179[55],s180[55],s181[55],s182[55],s183[55],s184[55],s185[55],s186[55],s187[55],s188[55],s189[55],s190[55],s191[55],s192[55],s10[46],s11[46],s12[46],s13[46],s14[46],s15[46],s16[46],s17[46],s18[46],s19[46],s20[46],s21[46],s22[46],s23[46],s24[46],s25[46],s26[46],s27[46],s28[46],s29[46],s30[46],s31[46],s32[46],s33[46],s34[46],s35[46],s36[46],s37[46],s38[46],s39[46],s40[46],s41[46],s42[46],s43[46],s44[46],s45[46],s46[46],s47[46],s48[46],s49[46],s50[46],s51[46],s52[46],s53[46],s54[46],s54[47],s54[48],s54[49],s54[50],s54[51],s54[52],s54[53],s54[54],s54[55],s54[56],s54[57],s54[58],s54[59],s54[60],s54[61],s54[62],s54[63],s54[64],s54[65],s54[66],s54[67],s54[68],s54[69],s54[70],s54[71],s54[72],s54[73],s54[74],s54[75],s52[78],s50[81],s48[84],s46[87],s45[89],s45[90],s45[91],s45[92],s45[93],s45[94],s45[95],s45[96],s45[97],s45[98],s45[99],s9[136],s8[138],s7[140],s6[142],s5[144],s4[146],s3[148],s2[150],s1[152],s103[51],s101[54],s56[100],s55[102],s54[104],s53[106],s52[108],s51[110],s50[112],s49[114],s48[116],s47[118],s46[120],s45[122],s44[124],s43[126],s42[128],s41[130],s40[132],s39[134],s38[136],s37[138],s36[140],s35[142],s34[144],s33[146],s32[148],s31[150],s30[152],s29[154],s28[156],s27[158],s26[160],s25[162],s24[164],s23[166],s22[168],s21[170],s20[172],s19[174],s18[176],s17[178],s16[180],s15[182],s14[184],s13[186],s12[188],s11[190],s10[192],s199[292],s198[294],s197[296],s196[298],s195[300],s194[302],s193[304],s192[210],s191[212],s190[214],s189[216],s188[218],s187[220],s186[222],s185[224],s184[226],s183[228],s182[230],s181[232],s180[234],s179[236],s178[238],s177[240],s176[242],s175[244],s174[246],s173[248],s172[250],s171[252],s170[254],s169[256],s168[258],s167[260],s166[262],s165[264],s164[266],s163[268],s162[270],s161[272],s160[274],s159[276],s158[278],s157[280],s156[282],s155[284],s154[286],s153[288],s152[290],s151[292],s150[294],s149[296],s148[298],s147[300],s146[302],s145[304],s144[306],s143[308],s142[310],s141[312],s140[314],s139[316],s138[318],s137[320],s136[322],s135[324],s134[326],s133[328],s132[330],s131[332],s130[334],s129[336],pp255[146],pp254[148],pp253[150],pp252[152],pp251[154],pp250[156],pp249[158],pp248[160],pp247[162],pp246[164],pp245[166],pp244[168],pp243[170],pp242[172],pp241[174],pp240[176],pp239[178],pp238[180],pp237[182],pp236[184],pp235[186],pp234[188],pp233[190],pp232[192],pp231[194],pp230[196],pp229[198],pp228[200],pp227[202],pp226[204],pp225[206],pp224[208],pp223[210],pp222[212],pp221[214],pp220[216],pp219[218],pp218[220],pp217[222],pp216[224],pp215[226],pp214[228],pp213[230],pp212[232],pp211[234],pp210[236],pp209[238],pp208[240],pp209[240],pp210[240],pp211[240],pp212[240],pp213[240],pp214[240],pp215[240],pp216[240],pp217[240],pp218[240],pp219[240],pp220[240],pp221[240],pp222[240],pp223[240],pp224[240],pp225[240],pp226[240],pp227[240],pp228[240],pp229[240],pp230[240],pp231[240],pp232[240]};
    CLA_434 KS_200(s200, c200, in200_1, in200_2);
    wire[431:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {pp26[14],pp26[15],pp26[16],pp26[17],pp26[18],pp26[19],pp26[20],pp26[21],pp26[22],pp26[23],pp26[24],pp26[25],pp26[26],pp26[27],pp26[28],pp26[29],pp26[30],pp26[31],pp26[32],pp26[33],pp26[34],pp26[35],pp26[36],pp26[37],pp28[36],pp30[35],pp32[34],pp34[33],pp36[32],pp38[31],pp40[30],pp42[29],pp44[28],pp46[27],pp48[26],pp50[25],pp52[24],pp54[23],pp56[22],pp58[21],pp60[20],pp62[19],pp64[18],pp66[17],pp68[16],pp70[15],pp72[14],pp74[13],pp76[12],pp78[11],pp80[10],s129[27],s130[27],s131[27],s132[27],s133[27],s134[27],s135[27],s136[27],s137[27],s136[29],s135[31],s134[33],s133[35],s132[37],s131[39],s130[41],s129[43],pp108[0],pp108[1],pp110[0],s129[47],s130[47],s131[47],s132[47],s133[47],s134[47],s135[47],s136[47],s137[47],s138[47],s139[47],s140[47],s141[47],s142[47],s143[47],s144[47],s145[47],s146[47],s147[47],s148[47],s149[47],s149[48],s149[49],s149[50],s149[51],s149[52],s149[53],s149[54],s200[100],s200[101],s200[102],s200[103],s200[104],s200[105],s200[106],s200[107],s200[108],s200[109],s200[110],s200[111],s200[112],s200[113],s200[114],s200[115],s200[116],s200[117],s200[118],s200[119],s200[120],s200[121],s200[122],s200[123],s200[124],s200[125],s200[126],s200[127],s200[128],s200[129],s200[130],s200[131],s200[132],s200[133],s200[134],s200[135],s200[136],s200[137],s200[138],s200[139],s200[140],s200[141],s200[142],s200[143],s200[144],s200[145],s200[146],s200[147],s200[148],s200[149],s200[150],s200[151],s200[152],s200[153],s200[154],s200[155],s200[156],s200[157],s200[158],s200[159],s200[160],s200[161],s200[162],s200[163],s200[164],s200[165],s200[166],s200[167],s200[168],s200[169],s200[170],s200[171],s200[172],s200[173],s200[174],s200[175],s200[176],s200[177],s200[178],s200[179],s200[180],s200[181],s200[182],s200[183],s200[184],s200[185],s200[186],s200[187],s200[188],s200[189],s200[190],s200[191],s200[192],s200[193],s200[194],s200[195],s200[196],s200[197],s200[198],s200[199],s200[200],s200[201],s200[202],s200[203],s200[204],s200[205],s200[206],s200[207],s200[208],s200[209],s200[210],s200[211],s200[212],s200[213],s200[214],s200[215],s200[216],s200[217],s200[218],s200[219],s200[220],s200[221],s200[222],s200[223],s200[224],s200[225],s200[226],s200[227],s200[228],s200[229],s200[230],s200[231],s200[232],s200[233],s200[234],s200[235],s200[236],s200[237],s200[238],s200[239],s200[240],s200[241],s200[242],s200[243],s200[244],s200[245],s200[246],s200[247],s200[248],s200[249],s200[250],s200[251],s200[252],s200[253],s200[254],s200[255],s200[256],s200[257],s200[258],s200[259],s200[260],s200[261],s200[262],s200[263],s200[264],s200[265],s200[266],s200[267],s200[268],s200[269],s200[270],s200[271],s200[272],s200[273],s200[274],s200[275],s200[276],s200[277],s200[278],s200[279],s200[280],s200[281],s200[282],s200[283],s200[284],s200[285],s200[286],s200[287],s200[288],s200[289],s200[290],s200[291],s199[293],s198[295],s197[297],s196[299],s195[301],s194[303],s193[305],s192[211],s191[213],s190[215],s189[217],s188[219],s187[221],s186[223],s185[225],s184[227],s183[229],s182[231],s181[233],s180[235],s179[237],s178[239],s177[241],s176[243],s175[245],s174[247],s173[249],s172[251],s171[253],s170[255],s169[257],s168[259],s167[261],s166[263],s165[265],s164[267],s163[269],s162[271],s161[273],s160[275],s159[277],s158[279],s157[281],s156[283],s155[285],s154[287],s153[289],s152[291],s151[293],s150[295],s149[297],s148[299],s147[301],s146[303],s145[305],s144[307],s143[309],s142[311],s141[313],s140[315],s139[317],s138[319],s137[321],s136[323],s135[325],s134[327],s133[329],s132[331],s131[333],s130[335],s129[337],pp255[147],pp254[149],pp253[151],pp252[153],pp251[155],pp250[157],pp249[159],pp248[161],pp247[163],pp246[165],pp245[167],pp244[169],pp243[171],pp242[173],pp241[175],pp240[177],pp239[179],pp238[181],pp237[183],pp236[185],pp235[187],pp234[189],pp233[191],pp232[193],pp231[195],pp230[197],pp229[199],pp228[201],pp227[203],pp226[205],pp225[207],pp224[209],pp223[211],pp222[213],pp221[215],pp220[217],pp219[219],pp218[221],pp217[223],pp216[225],pp215[227],pp214[229],pp213[231],pp212[233],pp211[235],pp210[237],pp209[239],pp210[239],pp211[239],pp212[239],pp213[239],pp214[239],pp215[239],pp216[239],pp217[239],pp218[239],pp219[239],pp220[239],pp221[239],pp222[239],pp223[239],pp224[239],pp225[239],pp226[239],pp227[239],pp228[239],pp229[239],pp230[239],pp231[239],pp232[239]};
    assign in201_2 = {pp27[13],pp27[14],pp27[15],pp27[16],pp27[17],pp27[18],pp27[19],pp27[20],pp27[21],pp27[22],pp27[23],pp27[24],pp27[25],pp27[26],pp27[27],pp27[28],pp27[29],pp27[30],pp27[31],pp27[32],pp27[33],pp27[34],pp27[35],pp27[36],pp29[35],pp31[34],pp33[33],pp35[32],pp37[31],pp39[30],pp41[29],pp43[28],pp45[27],pp47[26],pp49[25],pp51[24],pp53[23],pp55[22],pp57[21],pp59[20],pp61[19],pp63[18],pp65[17],pp67[16],pp69[15],pp71[14],pp73[13],pp75[12],pp77[11],pp79[10],s129[26],s130[26],s131[26],s132[26],s133[26],s134[26],s135[26],s136[26],s137[26],s138[26],s137[28],s136[30],s135[32],s134[34],s133[36],s132[38],s131[40],s130[42],s129[44],pp109[0],s129[46],s130[46],s131[46],s132[46],s133[46],s134[46],s135[46],s136[46],s137[46],s138[46],s139[46],s140[46],s141[46],s142[46],s143[46],s144[46],s145[46],s146[46],s147[46],s148[46],s149[46],s150[46],s150[47],s150[48],s150[49],s150[50],s150[51],s150[52],s150[53],s150[54],s151[54],s152[54],s153[54],s154[54],s155[54],s156[54],s157[54],s158[54],s159[54],s160[54],s161[54],s162[54],s163[54],s164[54],s165[54],s166[54],s167[54],s168[54],s169[54],s170[54],s171[54],s172[54],s173[54],s174[54],s175[54],s176[54],s177[54],s178[54],s179[54],s180[54],s181[54],s182[54],s183[54],s184[54],s185[54],s186[54],s187[54],s188[54],s189[54],s190[54],s191[54],s192[54],s10[45],s11[45],s12[45],s13[45],s14[45],s15[45],s16[45],s17[45],s18[45],s19[45],s20[45],s21[45],s22[45],s23[45],s24[45],s25[45],s26[45],s27[45],s28[45],s29[45],s30[45],s31[45],s32[45],s33[45],s34[45],s35[45],s36[45],s37[45],s38[45],s39[45],s40[45],s41[45],s42[45],s43[45],s44[45],s45[45],s46[45],s47[45],s48[45],s49[45],s50[45],s51[45],s52[45],s53[45],s54[45],s55[45],s55[46],s55[47],s55[48],s55[49],s55[50],s55[51],s55[52],s55[53],s55[54],s55[55],s55[56],s55[57],s55[58],s55[59],s55[60],s55[61],s55[62],s55[63],s55[64],s55[65],s55[66],s55[67],s55[68],s55[69],s55[70],s55[71],s55[72],s55[73],s55[74],s53[77],s51[80],s49[83],s47[86],s46[88],s46[89],s46[90],s46[91],s46[92],s46[93],s46[94],s46[95],s46[96],s46[97],s46[98],s46[99],s9[137],s8[139],s7[141],s6[143],s5[145],s4[147],s3[149],s2[151],s1[153],s102[53],s100[56],s56[101],s55[103],s54[105],s53[107],s52[109],s51[111],s50[113],s49[115],s48[117],s47[119],s46[121],s45[123],s44[125],s43[127],s42[129],s41[131],s40[133],s39[135],s38[137],s37[139],s36[141],s35[143],s34[145],s33[147],s32[149],s31[151],s30[153],s29[155],s28[157],s27[159],s26[161],s25[163],s24[165],s23[167],s22[169],s21[171],s20[173],s19[175],s18[177],s17[179],s16[181],s15[183],s14[185],s13[187],s12[189],s11[191],s10[193],s200[292],s199[294],s198[296],s197[298],s196[300],s195[302],s194[304],s193[306],s192[212],s191[214],s190[216],s189[218],s188[220],s187[222],s186[224],s185[226],s184[228],s183[230],s182[232],s181[234],s180[236],s179[238],s178[240],s177[242],s176[244],s175[246],s174[248],s173[250],s172[252],s171[254],s170[256],s169[258],s168[260],s167[262],s166[264],s165[266],s164[268],s163[270],s162[272],s161[274],s160[276],s159[278],s158[280],s157[282],s156[284],s155[286],s154[288],s153[290],s152[292],s151[294],s150[296],s149[298],s148[300],s147[302],s146[304],s145[306],s144[308],s143[310],s142[312],s141[314],s140[316],s139[318],s138[320],s137[322],s136[324],s135[326],s134[328],s133[330],s132[332],s131[334],s130[336],s129[338],pp255[148],pp254[150],pp253[152],pp252[154],pp251[156],pp250[158],pp249[160],pp248[162],pp247[164],pp246[166],pp245[168],pp244[170],pp243[172],pp242[174],pp241[176],pp240[178],pp239[180],pp238[182],pp237[184],pp236[186],pp235[188],pp234[190],pp233[192],pp232[194],pp231[196],pp230[198],pp229[200],pp228[202],pp227[204],pp226[206],pp225[208],pp224[210],pp223[212],pp222[214],pp221[216],pp220[218],pp219[220],pp218[222],pp217[224],pp216[226],pp215[228],pp214[230],pp213[232],pp212[234],pp211[236],pp210[238],pp211[238],pp212[238],pp213[238],pp214[238],pp215[238],pp216[238],pp217[238],pp218[238],pp219[238],pp220[238],pp221[238],pp222[238],pp223[238],pp224[238],pp225[238],pp226[238],pp227[238],pp228[238],pp229[238],pp230[238],pp231[238],pp232[238],pp233[238]};
    CLA_432 KS_201(s201, c201, in201_1, in201_2);
    wire[429:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp28[13],pp28[14],pp28[15],pp28[16],pp28[17],pp28[18],pp28[19],pp28[20],pp28[21],pp28[22],pp28[23],pp28[24],pp28[25],pp28[26],pp28[27],pp28[28],pp28[29],pp28[30],pp28[31],pp28[32],pp28[33],pp28[34],pp28[35],pp30[34],pp32[33],pp34[32],pp36[31],pp38[30],pp40[29],pp42[28],pp44[27],pp46[26],pp48[25],pp50[24],pp52[23],pp54[22],pp56[21],pp58[20],pp60[19],pp62[18],pp64[17],pp66[16],pp68[15],pp70[14],pp72[13],pp74[12],pp76[11],pp78[10],s129[25],s130[25],s131[25],s132[25],s133[25],s134[25],s135[25],s136[25],s137[25],s138[25],s139[25],s138[27],s137[29],s136[31],s135[33],s134[35],s133[37],s132[39],s131[41],s130[43],s129[45],s130[45],s131[45],s132[45],s133[45],s134[45],s135[45],s136[45],s137[45],s138[45],s139[45],s140[45],s141[45],s142[45],s143[45],s144[45],s145[45],s146[45],s147[45],s148[45],s149[45],s150[45],s151[45],s151[46],s151[47],s151[48],s151[49],s151[50],s151[51],s151[52],s151[53],s201[100],s201[101],s201[102],s201[103],s201[104],s201[105],s201[106],s201[107],s201[108],s201[109],s201[110],s201[111],s201[112],s201[113],s201[114],s201[115],s201[116],s201[117],s201[118],s201[119],s201[120],s201[121],s201[122],s201[123],s201[124],s201[125],s201[126],s201[127],s201[128],s201[129],s201[130],s201[131],s201[132],s201[133],s201[134],s201[135],s201[136],s201[137],s201[138],s201[139],s201[140],s201[141],s201[142],s201[143],s201[144],s201[145],s201[146],s201[147],s201[148],s201[149],s201[150],s201[151],s201[152],s201[153],s201[154],s201[155],s201[156],s201[157],s201[158],s201[159],s201[160],s201[161],s201[162],s201[163],s201[164],s201[165],s201[166],s201[167],s201[168],s201[169],s201[170],s201[171],s201[172],s201[173],s201[174],s201[175],s201[176],s201[177],s201[178],s201[179],s201[180],s201[181],s201[182],s201[183],s201[184],s201[185],s201[186],s201[187],s201[188],s201[189],s201[190],s201[191],s201[192],s201[193],s201[194],s201[195],s201[196],s201[197],s201[198],s201[199],s201[200],s201[201],s201[202],s201[203],s201[204],s201[205],s201[206],s201[207],s201[208],s201[209],s201[210],s201[211],s201[212],s201[213],s201[214],s201[215],s201[216],s201[217],s201[218],s201[219],s201[220],s201[221],s201[222],s201[223],s201[224],s201[225],s201[226],s201[227],s201[228],s201[229],s201[230],s201[231],s201[232],s201[233],s201[234],s201[235],s201[236],s201[237],s201[238],s201[239],s201[240],s201[241],s201[242],s201[243],s201[244],s201[245],s201[246],s201[247],s201[248],s201[249],s201[250],s201[251],s201[252],s201[253],s201[254],s201[255],s201[256],s201[257],s201[258],s201[259],s201[260],s201[261],s201[262],s201[263],s201[264],s201[265],s201[266],s201[267],s201[268],s201[269],s201[270],s201[271],s201[272],s201[273],s201[274],s201[275],s201[276],s201[277],s201[278],s201[279],s201[280],s201[281],s201[282],s201[283],s201[284],s201[285],s201[286],s201[287],s201[288],s201[289],s201[290],s201[291],s200[293],s199[295],s198[297],s197[299],s196[301],s195[303],s194[305],s193[307],s192[213],s191[215],s190[217],s189[219],s188[221],s187[223],s186[225],s185[227],s184[229],s183[231],s182[233],s181[235],s180[237],s179[239],s178[241],s177[243],s176[245],s175[247],s174[249],s173[251],s172[253],s171[255],s170[257],s169[259],s168[261],s167[263],s166[265],s165[267],s164[269],s163[271],s162[273],s161[275],s160[277],s159[279],s158[281],s157[283],s156[285],s155[287],s154[289],s153[291],s152[293],s151[295],s150[297],s149[299],s148[301],s147[303],s146[305],s145[307],s144[309],s143[311],s142[313],s141[315],s140[317],s139[319],s138[321],s137[323],s136[325],s135[327],s134[329],s133[331],s132[333],s131[335],s130[337],s129[339],pp255[149],pp254[151],pp253[153],pp252[155],pp251[157],pp250[159],pp249[161],pp248[163],pp247[165],pp246[167],pp245[169],pp244[171],pp243[173],pp242[175],pp241[177],pp240[179],pp239[181],pp238[183],pp237[185],pp236[187],pp235[189],pp234[191],pp233[193],pp232[195],pp231[197],pp230[199],pp229[201],pp228[203],pp227[205],pp226[207],pp225[209],pp224[211],pp223[213],pp222[215],pp221[217],pp220[219],pp219[221],pp218[223],pp217[225],pp216[227],pp215[229],pp214[231],pp213[233],pp212[235],pp211[237],pp212[237],pp213[237],pp214[237],pp215[237],pp216[237],pp217[237],pp218[237],pp219[237],pp220[237],pp221[237],pp222[237],pp223[237],pp224[237],pp225[237],pp226[237],pp227[237],pp228[237],pp229[237],pp230[237],pp231[237],pp232[237],pp233[237]};
    assign in202_2 = {pp29[12],pp29[13],pp29[14],pp29[15],pp29[16],pp29[17],pp29[18],pp29[19],pp29[20],pp29[21],pp29[22],pp29[23],pp29[24],pp29[25],pp29[26],pp29[27],pp29[28],pp29[29],pp29[30],pp29[31],pp29[32],pp29[33],pp29[34],pp31[33],pp33[32],pp35[31],pp37[30],pp39[29],pp41[28],pp43[27],pp45[26],pp47[25],pp49[24],pp51[23],pp53[22],pp55[21],pp57[20],pp59[19],pp61[18],pp63[17],pp65[16],pp67[15],pp69[14],pp71[13],pp73[12],pp75[11],pp77[10],s129[24],s130[24],s131[24],s132[24],s133[24],s134[24],s135[24],s136[24],s137[24],s138[24],s139[24],s140[24],s139[26],s138[28],s137[30],s136[32],s135[34],s134[36],s133[38],s132[40],s131[42],s130[44],s131[44],s132[44],s133[44],s134[44],s135[44],s136[44],s137[44],s138[44],s139[44],s140[44],s141[44],s142[44],s143[44],s144[44],s145[44],s146[44],s147[44],s148[44],s149[44],s150[44],s151[44],s152[44],s152[45],s152[46],s152[47],s152[48],s152[49],s152[50],s152[51],s152[52],s152[53],s153[53],s154[53],s155[53],s156[53],s157[53],s158[53],s159[53],s160[53],s161[53],s162[53],s163[53],s164[53],s165[53],s166[53],s167[53],s168[53],s169[53],s170[53],s171[53],s172[53],s173[53],s174[53],s175[53],s176[53],s177[53],s178[53],s179[53],s180[53],s181[53],s182[53],s183[53],s184[53],s185[53],s186[53],s187[53],s188[53],s189[53],s190[53],s191[53],s192[53],s10[44],s11[44],s12[44],s13[44],s14[44],s15[44],s16[44],s17[44],s18[44],s19[44],s20[44],s21[44],s22[44],s23[44],s24[44],s25[44],s26[44],s27[44],s28[44],s29[44],s30[44],s31[44],s32[44],s33[44],s34[44],s35[44],s36[44],s37[44],s38[44],s39[44],s40[44],s41[44],s42[44],s43[44],s44[44],s45[44],s46[44],s47[44],s48[44],s49[44],s50[44],s51[44],s52[44],s53[44],s54[44],s55[44],s56[44],s56[45],s56[46],s56[47],s56[48],s56[49],s56[50],s56[51],s56[52],s56[53],s56[54],s56[55],s56[56],s56[57],s56[58],s56[59],s56[60],s56[61],s56[62],s56[63],s56[64],s56[65],s56[66],s56[67],s56[68],s56[69],s56[70],s56[71],s56[72],s56[73],s54[76],s52[79],s50[82],s48[85],s47[87],s47[88],s47[89],s47[90],s47[91],s47[92],s47[93],s47[94],s47[95],s47[96],s47[97],s47[98],s47[99],s9[138],s8[140],s7[142],s6[144],s5[146],s4[148],s3[150],s2[152],s1[154],s101[55],s57[100],s56[102],s55[104],s54[106],s53[108],s52[110],s51[112],s50[114],s49[116],s48[118],s47[120],s46[122],s45[124],s44[126],s43[128],s42[130],s41[132],s40[134],s39[136],s38[138],s37[140],s36[142],s35[144],s34[146],s33[148],s32[150],s31[152],s30[154],s29[156],s28[158],s27[160],s26[162],s25[164],s24[166],s23[168],s22[170],s21[172],s20[174],s19[176],s18[178],s17[180],s16[182],s15[184],s14[186],s13[188],s12[190],s11[192],s10[194],s201[292],s200[294],s199[296],s198[298],s197[300],s196[302],s195[304],s194[306],s193[308],s192[214],s191[216],s190[218],s189[220],s188[222],s187[224],s186[226],s185[228],s184[230],s183[232],s182[234],s181[236],s180[238],s179[240],s178[242],s177[244],s176[246],s175[248],s174[250],s173[252],s172[254],s171[256],s170[258],s169[260],s168[262],s167[264],s166[266],s165[268],s164[270],s163[272],s162[274],s161[276],s160[278],s159[280],s158[282],s157[284],s156[286],s155[288],s154[290],s153[292],s152[294],s151[296],s150[298],s149[300],s148[302],s147[304],s146[306],s145[308],s144[310],s143[312],s142[314],s141[316],s140[318],s139[320],s138[322],s137[324],s136[326],s135[328],s134[330],s133[332],s132[334],s131[336],s130[338],s129[340],pp255[150],pp254[152],pp253[154],pp252[156],pp251[158],pp250[160],pp249[162],pp248[164],pp247[166],pp246[168],pp245[170],pp244[172],pp243[174],pp242[176],pp241[178],pp240[180],pp239[182],pp238[184],pp237[186],pp236[188],pp235[190],pp234[192],pp233[194],pp232[196],pp231[198],pp230[200],pp229[202],pp228[204],pp227[206],pp226[208],pp225[210],pp224[212],pp223[214],pp222[216],pp221[218],pp220[220],pp219[222],pp218[224],pp217[226],pp216[228],pp215[230],pp214[232],pp213[234],pp212[236],pp213[236],pp214[236],pp215[236],pp216[236],pp217[236],pp218[236],pp219[236],pp220[236],pp221[236],pp222[236],pp223[236],pp224[236],pp225[236],pp226[236],pp227[236],pp228[236],pp229[236],pp230[236],pp231[236],pp232[236],pp233[236],pp234[236]};
    CLA_430 KS_202(s202, c202, in202_1, in202_2);
    wire[427:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {pp30[12],pp30[13],pp30[14],pp30[15],pp30[16],pp30[17],pp30[18],pp30[19],pp30[20],pp30[21],pp30[22],pp30[23],pp30[24],pp30[25],pp30[26],pp30[27],pp30[28],pp30[29],pp30[30],pp30[31],pp30[32],pp30[33],pp32[32],pp34[31],pp36[30],pp38[29],pp40[28],pp42[27],pp44[26],pp46[25],pp48[24],pp50[23],pp52[22],pp54[21],pp56[20],pp58[19],pp60[18],pp62[17],pp64[16],pp66[15],pp68[14],pp70[13],pp72[12],pp74[11],pp76[10],s129[23],s130[23],s131[23],s132[23],s133[23],s134[23],s135[23],s136[23],s137[23],s138[23],s139[23],s140[23],s141[23],s140[25],s139[27],s138[29],s137[31],s136[33],s135[35],s134[37],s133[39],s132[41],s131[43],s132[43],s133[43],s134[43],s135[43],s136[43],s137[43],s138[43],s139[43],s140[43],s141[43],s142[43],s143[43],s144[43],s145[43],s146[43],s147[43],s148[43],s149[43],s150[43],s151[43],s152[43],s153[43],s153[44],s153[45],s153[46],s153[47],s153[48],s153[49],s153[50],s153[51],s153[52],s202[100],s202[101],s202[102],s202[103],s202[104],s202[105],s202[106],s202[107],s202[108],s202[109],s202[110],s202[111],s202[112],s202[113],s202[114],s202[115],s202[116],s202[117],s202[118],s202[119],s202[120],s202[121],s202[122],s202[123],s202[124],s202[125],s202[126],s202[127],s202[128],s202[129],s202[130],s202[131],s202[132],s202[133],s202[134],s202[135],s202[136],s202[137],s202[138],s202[139],s202[140],s202[141],s202[142],s202[143],s202[144],s202[145],s202[146],s202[147],s202[148],s202[149],s202[150],s202[151],s202[152],s202[153],s202[154],s202[155],s202[156],s202[157],s202[158],s202[159],s202[160],s202[161],s202[162],s202[163],s202[164],s202[165],s202[166],s202[167],s202[168],s202[169],s202[170],s202[171],s202[172],s202[173],s202[174],s202[175],s202[176],s202[177],s202[178],s202[179],s202[180],s202[181],s202[182],s202[183],s202[184],s202[185],s202[186],s202[187],s202[188],s202[189],s202[190],s202[191],s202[192],s202[193],s202[194],s202[195],s202[196],s202[197],s202[198],s202[199],s202[200],s202[201],s202[202],s202[203],s202[204],s202[205],s202[206],s202[207],s202[208],s202[209],s202[210],s202[211],s202[212],s202[213],s202[214],s202[215],s202[216],s202[217],s202[218],s202[219],s202[220],s202[221],s202[222],s202[223],s202[224],s202[225],s202[226],s202[227],s202[228],s202[229],s202[230],s202[231],s202[232],s202[233],s202[234],s202[235],s202[236],s202[237],s202[238],s202[239],s202[240],s202[241],s202[242],s202[243],s202[244],s202[245],s202[246],s202[247],s202[248],s202[249],s202[250],s202[251],s202[252],s202[253],s202[254],s202[255],s202[256],s202[257],s202[258],s202[259],s202[260],s202[261],s202[262],s202[263],s202[264],s202[265],s202[266],s202[267],s202[268],s202[269],s202[270],s202[271],s202[272],s202[273],s202[274],s202[275],s202[276],s202[277],s202[278],s202[279],s202[280],s202[281],s202[282],s202[283],s202[284],s202[285],s202[286],s202[287],s202[288],s202[289],s202[290],s202[291],s201[293],s200[295],s199[297],s198[299],s197[301],s196[303],s195[305],s194[307],s193[309],s192[215],s191[217],s190[219],s189[221],s188[223],s187[225],s186[227],s185[229],s184[231],s183[233],s182[235],s181[237],s180[239],s179[241],s178[243],s177[245],s176[247],s175[249],s174[251],s173[253],s172[255],s171[257],s170[259],s169[261],s168[263],s167[265],s166[267],s165[269],s164[271],s163[273],s162[275],s161[277],s160[279],s159[281],s158[283],s157[285],s156[287],s155[289],s154[291],s153[293],s152[295],s151[297],s150[299],s149[301],s148[303],s147[305],s146[307],s145[309],s144[311],s143[313],s142[315],s141[317],s140[319],s139[321],s138[323],s137[325],s136[327],s135[329],s134[331],s133[333],s132[335],s131[337],s130[339],s129[341],pp255[151],pp254[153],pp253[155],pp252[157],pp251[159],pp250[161],pp249[163],pp248[165],pp247[167],pp246[169],pp245[171],pp244[173],pp243[175],pp242[177],pp241[179],pp240[181],pp239[183],pp238[185],pp237[187],pp236[189],pp235[191],pp234[193],pp233[195],pp232[197],pp231[199],pp230[201],pp229[203],pp228[205],pp227[207],pp226[209],pp225[211],pp224[213],pp223[215],pp222[217],pp221[219],pp220[221],pp219[223],pp218[225],pp217[227],pp216[229],pp215[231],pp214[233],pp213[235],pp214[235],pp215[235],pp216[235],pp217[235],pp218[235],pp219[235],pp220[235],pp221[235],pp222[235],pp223[235],pp224[235],pp225[235],pp226[235],pp227[235],pp228[235],pp229[235],pp230[235],pp231[235],pp232[235],pp233[235],pp234[235]};
    assign in203_2 = {pp31[11],pp31[12],pp31[13],pp31[14],pp31[15],pp31[16],pp31[17],pp31[18],pp31[19],pp31[20],pp31[21],pp31[22],pp31[23],pp31[24],pp31[25],pp31[26],pp31[27],pp31[28],pp31[29],pp31[30],pp31[31],pp31[32],pp33[31],pp35[30],pp37[29],pp39[28],pp41[27],pp43[26],pp45[25],pp47[24],pp49[23],pp51[22],pp53[21],pp55[20],pp57[19],pp59[18],pp61[17],pp63[16],pp65[15],pp67[14],pp69[13],pp71[12],pp73[11],pp75[10],s129[22],s130[22],s131[22],s132[22],s133[22],s134[22],s135[22],s136[22],s137[22],s138[22],s139[22],s140[22],s141[22],s142[22],s141[24],s140[26],s139[28],s138[30],s137[32],s136[34],s135[36],s134[38],s133[40],s132[42],s133[42],s134[42],s135[42],s136[42],s137[42],s138[42],s139[42],s140[42],s141[42],s142[42],s143[42],s144[42],s145[42],s146[42],s147[42],s148[42],s149[42],s150[42],s151[42],s152[42],s153[42],s154[42],s154[43],s154[44],s154[45],s154[46],s154[47],s154[48],s154[49],s154[50],s154[51],s154[52],s155[52],s156[52],s157[52],s158[52],s159[52],s160[52],s161[52],s162[52],s163[52],s164[52],s165[52],s166[52],s167[52],s168[52],s169[52],s170[52],s171[52],s172[52],s173[52],s174[52],s175[52],s176[52],s177[52],s178[52],s179[52],s180[52],s181[52],s182[52],s183[52],s184[52],s185[52],s186[52],s187[52],s188[52],s189[52],s190[52],s191[52],s192[52],s10[43],s11[43],s12[43],s13[43],s14[43],s15[43],s16[43],s17[43],s18[43],s19[43],s20[43],s21[43],s22[43],s23[43],s24[43],s25[43],s26[43],s27[43],s28[43],s29[43],s30[43],s31[43],s32[43],s33[43],s34[43],s35[43],s36[43],s37[43],s38[43],s39[43],s40[43],s41[43],s42[43],s43[43],s44[43],s45[43],s46[43],s47[43],s48[43],s49[43],s50[43],s51[43],s52[43],s53[43],s54[43],s55[43],s56[43],s57[43],s57[44],s57[45],s57[46],s57[47],s57[48],s57[49],s57[50],s57[51],s57[52],s57[53],s57[54],s57[55],s57[56],s57[57],s57[58],s57[59],s57[60],s57[61],s57[62],s57[63],s57[64],s57[65],s57[66],s57[67],s57[68],s57[69],s57[70],s57[71],s57[72],s55[75],s53[78],s51[81],s49[84],s48[86],s48[87],s48[88],s48[89],s48[90],s48[91],s48[92],s48[93],s48[94],s48[95],s48[96],s48[97],s48[98],s48[99],s9[139],s8[141],s7[143],s6[145],s5[147],s4[149],s3[151],s2[153],s1[155],s100[57],s57[101],s56[103],s55[105],s54[107],s53[109],s52[111],s51[113],s50[115],s49[117],s48[119],s47[121],s46[123],s45[125],s44[127],s43[129],s42[131],s41[133],s40[135],s39[137],s38[139],s37[141],s36[143],s35[145],s34[147],s33[149],s32[151],s31[153],s30[155],s29[157],s28[159],s27[161],s26[163],s25[165],s24[167],s23[169],s22[171],s21[173],s20[175],s19[177],s18[179],s17[181],s16[183],s15[185],s14[187],s13[189],s12[191],s11[193],s10[195],s202[292],s201[294],s200[296],s199[298],s198[300],s197[302],s196[304],s195[306],s194[308],s193[310],s192[216],s191[218],s190[220],s189[222],s188[224],s187[226],s186[228],s185[230],s184[232],s183[234],s182[236],s181[238],s180[240],s179[242],s178[244],s177[246],s176[248],s175[250],s174[252],s173[254],s172[256],s171[258],s170[260],s169[262],s168[264],s167[266],s166[268],s165[270],s164[272],s163[274],s162[276],s161[278],s160[280],s159[282],s158[284],s157[286],s156[288],s155[290],s154[292],s153[294],s152[296],s151[298],s150[300],s149[302],s148[304],s147[306],s146[308],s145[310],s144[312],s143[314],s142[316],s141[318],s140[320],s139[322],s138[324],s137[326],s136[328],s135[330],s134[332],s133[334],s132[336],s131[338],s130[340],s129[342],pp255[152],pp254[154],pp253[156],pp252[158],pp251[160],pp250[162],pp249[164],pp248[166],pp247[168],pp246[170],pp245[172],pp244[174],pp243[176],pp242[178],pp241[180],pp240[182],pp239[184],pp238[186],pp237[188],pp236[190],pp235[192],pp234[194],pp233[196],pp232[198],pp231[200],pp230[202],pp229[204],pp228[206],pp227[208],pp226[210],pp225[212],pp224[214],pp223[216],pp222[218],pp221[220],pp220[222],pp219[224],pp218[226],pp217[228],pp216[230],pp215[232],pp214[234],pp215[234],pp216[234],pp217[234],pp218[234],pp219[234],pp220[234],pp221[234],pp222[234],pp223[234],pp224[234],pp225[234],pp226[234],pp227[234],pp228[234],pp229[234],pp230[234],pp231[234],pp232[234],pp233[234],pp234[234],pp235[234]};
    CLA_428 KS_203(s203, c203, in203_1, in203_2);
    wire[425:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {pp32[11],pp32[12],pp32[13],pp32[14],pp32[15],pp32[16],pp32[17],pp32[18],pp32[19],pp32[20],pp32[21],pp32[22],pp32[23],pp32[24],pp32[25],pp32[26],pp32[27],pp32[28],pp32[29],pp32[30],pp32[31],pp34[30],pp36[29],pp38[28],pp40[27],pp42[26],pp44[25],pp46[24],pp48[23],pp50[22],pp52[21],pp54[20],pp56[19],pp58[18],pp60[17],pp62[16],pp64[15],pp66[14],pp68[13],pp70[12],pp72[11],pp74[10],s129[21],s130[21],s131[21],s132[21],s133[21],s134[21],s135[21],s136[21],s137[21],s138[21],s139[21],s140[21],s141[21],s142[21],s143[21],s142[23],s141[25],s140[27],s139[29],s138[31],s137[33],s136[35],s135[37],s134[39],s133[41],s134[41],s135[41],s136[41],s137[41],s138[41],s139[41],s140[41],s141[41],s142[41],s143[41],s144[41],s145[41],s146[41],s147[41],s148[41],s149[41],s150[41],s151[41],s152[41],s153[41],s154[41],s155[41],s155[42],s155[43],s155[44],s155[45],s155[46],s155[47],s155[48],s155[49],s155[50],s155[51],s203[100],s203[101],s203[102],s203[103],s203[104],s203[105],s203[106],s203[107],s203[108],s203[109],s203[110],s203[111],s203[112],s203[113],s203[114],s203[115],s203[116],s203[117],s203[118],s203[119],s203[120],s203[121],s203[122],s203[123],s203[124],s203[125],s203[126],s203[127],s203[128],s203[129],s203[130],s203[131],s203[132],s203[133],s203[134],s203[135],s203[136],s203[137],s203[138],s203[139],s203[140],s203[141],s203[142],s203[143],s203[144],s203[145],s203[146],s203[147],s203[148],s203[149],s203[150],s203[151],s203[152],s203[153],s203[154],s203[155],s203[156],s203[157],s203[158],s203[159],s203[160],s203[161],s203[162],s203[163],s203[164],s203[165],s203[166],s203[167],s203[168],s203[169],s203[170],s203[171],s203[172],s203[173],s203[174],s203[175],s203[176],s203[177],s203[178],s203[179],s203[180],s203[181],s203[182],s203[183],s203[184],s203[185],s203[186],s203[187],s203[188],s203[189],s203[190],s203[191],s203[192],s203[193],s203[194],s203[195],s203[196],s203[197],s203[198],s203[199],s203[200],s203[201],s203[202],s203[203],s203[204],s203[205],s203[206],s203[207],s203[208],s203[209],s203[210],s203[211],s203[212],s203[213],s203[214],s203[215],s203[216],s203[217],s203[218],s203[219],s203[220],s203[221],s203[222],s203[223],s203[224],s203[225],s203[226],s203[227],s203[228],s203[229],s203[230],s203[231],s203[232],s203[233],s203[234],s203[235],s203[236],s203[237],s203[238],s203[239],s203[240],s203[241],s203[242],s203[243],s203[244],s203[245],s203[246],s203[247],s203[248],s203[249],s203[250],s203[251],s203[252],s203[253],s203[254],s203[255],s203[256],s203[257],s203[258],s203[259],s203[260],s203[261],s203[262],s203[263],s203[264],s203[265],s203[266],s203[267],s203[268],s203[269],s203[270],s203[271],s203[272],s203[273],s203[274],s203[275],s203[276],s203[277],s203[278],s203[279],s203[280],s203[281],s203[282],s203[283],s203[284],s203[285],s203[286],s203[287],s203[288],s203[289],s203[290],s203[291],s202[293],s201[295],s200[297],s199[299],s198[301],s197[303],s196[305],s195[307],s194[309],s193[311],s192[217],s191[219],s190[221],s189[223],s188[225],s187[227],s186[229],s185[231],s184[233],s183[235],s182[237],s181[239],s180[241],s179[243],s178[245],s177[247],s176[249],s175[251],s174[253],s173[255],s172[257],s171[259],s170[261],s169[263],s168[265],s167[267],s166[269],s165[271],s164[273],s163[275],s162[277],s161[279],s160[281],s159[283],s158[285],s157[287],s156[289],s155[291],s154[293],s153[295],s152[297],s151[299],s150[301],s149[303],s148[305],s147[307],s146[309],s145[311],s144[313],s143[315],s142[317],s141[319],s140[321],s139[323],s138[325],s137[327],s136[329],s135[331],s134[333],s133[335],s132[337],s131[339],s130[341],s129[343],pp255[153],pp254[155],pp253[157],pp252[159],pp251[161],pp250[163],pp249[165],pp248[167],pp247[169],pp246[171],pp245[173],pp244[175],pp243[177],pp242[179],pp241[181],pp240[183],pp239[185],pp238[187],pp237[189],pp236[191],pp235[193],pp234[195],pp233[197],pp232[199],pp231[201],pp230[203],pp229[205],pp228[207],pp227[209],pp226[211],pp225[213],pp224[215],pp223[217],pp222[219],pp221[221],pp220[223],pp219[225],pp218[227],pp217[229],pp216[231],pp215[233],pp216[233],pp217[233],pp218[233],pp219[233],pp220[233],pp221[233],pp222[233],pp223[233],pp224[233],pp225[233],pp226[233],pp227[233],pp228[233],pp229[233],pp230[233],pp231[233],pp232[233],pp233[233],pp234[233],pp235[233]};
    assign in204_2 = {pp33[10],pp33[11],pp33[12],pp33[13],pp33[14],pp33[15],pp33[16],pp33[17],pp33[18],pp33[19],pp33[20],pp33[21],pp33[22],pp33[23],pp33[24],pp33[25],pp33[26],pp33[27],pp33[28],pp33[29],pp33[30],pp35[29],pp37[28],pp39[27],pp41[26],pp43[25],pp45[24],pp47[23],pp49[22],pp51[21],pp53[20],pp55[19],pp57[18],pp59[17],pp61[16],pp63[15],pp65[14],pp67[13],pp69[12],pp71[11],pp73[10],s129[20],s130[20],s131[20],s132[20],s133[20],s134[20],s135[20],s136[20],s137[20],s138[20],s139[20],s140[20],s141[20],s142[20],s143[20],s144[20],s143[22],s142[24],s141[26],s140[28],s139[30],s138[32],s137[34],s136[36],s135[38],s134[40],s135[40],s136[40],s137[40],s138[40],s139[40],s140[40],s141[40],s142[40],s143[40],s144[40],s145[40],s146[40],s147[40],s148[40],s149[40],s150[40],s151[40],s152[40],s153[40],s154[40],s155[40],s156[40],s156[41],s156[42],s156[43],s156[44],s156[45],s156[46],s156[47],s156[48],s156[49],s156[50],s156[51],s157[51],s158[51],s159[51],s160[51],s161[51],s162[51],s163[51],s164[51],s165[51],s166[51],s167[51],s168[51],s169[51],s170[51],s171[51],s172[51],s173[51],s174[51],s175[51],s176[51],s177[51],s178[51],s179[51],s180[51],s181[51],s182[51],s183[51],s184[51],s185[51],s186[51],s187[51],s188[51],s189[51],s190[51],s191[51],s192[51],s10[42],s11[42],s12[42],s13[42],s14[42],s15[42],s16[42],s17[42],s18[42],s19[42],s20[42],s21[42],s22[42],s23[42],s24[42],s25[42],s26[42],s27[42],s28[42],s29[42],s30[42],s31[42],s32[42],s33[42],s34[42],s35[42],s36[42],s37[42],s38[42],s39[42],s40[42],s41[42],s42[42],s43[42],s44[42],s45[42],s46[42],s47[42],s48[42],s49[42],s50[42],s51[42],s52[42],s53[42],s54[42],s55[42],s56[42],s57[42],s58[42],s58[43],s58[44],s58[45],s58[46],s58[47],s58[48],s58[49],s58[50],s58[51],s58[52],s58[53],s58[54],s58[55],s58[56],s58[57],s58[58],s58[59],s58[60],s58[61],s58[62],s58[63],s58[64],s58[65],s58[66],s58[67],s58[68],s58[69],s58[70],s58[71],s56[74],s54[77],s52[80],s50[83],s49[85],s49[86],s49[87],s49[88],s49[89],s49[90],s49[91],s49[92],s49[93],s49[94],s49[95],s49[96],s49[97],s49[98],s49[99],s9[140],s8[142],s7[144],s6[146],s5[148],s4[150],s3[152],s2[154],s1[156],s58[100],s57[102],s56[104],s55[106],s54[108],s53[110],s52[112],s51[114],s50[116],s49[118],s48[120],s47[122],s46[124],s45[126],s44[128],s43[130],s42[132],s41[134],s40[136],s39[138],s38[140],s37[142],s36[144],s35[146],s34[148],s33[150],s32[152],s31[154],s30[156],s29[158],s28[160],s27[162],s26[164],s25[166],s24[168],s23[170],s22[172],s21[174],s20[176],s19[178],s18[180],s17[182],s16[184],s15[186],s14[188],s13[190],s12[192],s11[194],s10[196],s203[292],s202[294],s201[296],s200[298],s199[300],s198[302],s197[304],s196[306],s195[308],s194[310],s193[312],s192[218],s191[220],s190[222],s189[224],s188[226],s187[228],s186[230],s185[232],s184[234],s183[236],s182[238],s181[240],s180[242],s179[244],s178[246],s177[248],s176[250],s175[252],s174[254],s173[256],s172[258],s171[260],s170[262],s169[264],s168[266],s167[268],s166[270],s165[272],s164[274],s163[276],s162[278],s161[280],s160[282],s159[284],s158[286],s157[288],s156[290],s155[292],s154[294],s153[296],s152[298],s151[300],s150[302],s149[304],s148[306],s147[308],s146[310],s145[312],s144[314],s143[316],s142[318],s141[320],s140[322],s139[324],s138[326],s137[328],s136[330],s135[332],s134[334],s133[336],s132[338],s131[340],s130[342],s129[344],pp255[154],pp254[156],pp253[158],pp252[160],pp251[162],pp250[164],pp249[166],pp248[168],pp247[170],pp246[172],pp245[174],pp244[176],pp243[178],pp242[180],pp241[182],pp240[184],pp239[186],pp238[188],pp237[190],pp236[192],pp235[194],pp234[196],pp233[198],pp232[200],pp231[202],pp230[204],pp229[206],pp228[208],pp227[210],pp226[212],pp225[214],pp224[216],pp223[218],pp222[220],pp221[222],pp220[224],pp219[226],pp218[228],pp217[230],pp216[232],pp217[232],pp218[232],pp219[232],pp220[232],pp221[232],pp222[232],pp223[232],pp224[232],pp225[232],pp226[232],pp227[232],pp228[232],pp229[232],pp230[232],pp231[232],pp232[232],pp233[232],pp234[232],pp235[232],pp236[232]};
    CLA_426 KS_204(s204, c204, in204_1, in204_2);
    wire[423:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {pp34[10],pp34[11],pp34[12],pp34[13],pp34[14],pp34[15],pp34[16],pp34[17],pp34[18],pp34[19],pp34[20],pp34[21],pp34[22],pp34[23],pp34[24],pp34[25],pp34[26],pp34[27],pp34[28],pp34[29],pp36[28],pp38[27],pp40[26],pp42[25],pp44[24],pp46[23],pp48[22],pp50[21],pp52[20],pp54[19],pp56[18],pp58[17],pp60[16],pp62[15],pp64[14],pp66[13],pp68[12],pp70[11],pp72[10],s129[19],s130[19],s131[19],s132[19],s133[19],s134[19],s135[19],s136[19],s137[19],s138[19],s139[19],s140[19],s141[19],s142[19],s143[19],s144[19],s145[19],s144[21],s143[23],s142[25],s141[27],s140[29],s139[31],s138[33],s137[35],s136[37],s135[39],s136[39],s137[39],s138[39],s139[39],s140[39],s141[39],s142[39],s143[39],s144[39],s145[39],s146[39],s147[39],s148[39],s149[39],s150[39],s151[39],s152[39],s153[39],s154[39],s155[39],s156[39],s157[39],s157[40],s157[41],s157[42],s157[43],s157[44],s157[45],s157[46],s157[47],s157[48],s157[49],s157[50],s204[100],s204[101],s204[102],s204[103],s204[104],s204[105],s204[106],s204[107],s204[108],s204[109],s204[110],s204[111],s204[112],s204[113],s204[114],s204[115],s204[116],s204[117],s204[118],s204[119],s204[120],s204[121],s204[122],s204[123],s204[124],s204[125],s204[126],s204[127],s204[128],s204[129],s204[130],s204[131],s204[132],s204[133],s204[134],s204[135],s204[136],s204[137],s204[138],s204[139],s204[140],s204[141],s204[142],s204[143],s204[144],s204[145],s204[146],s204[147],s204[148],s204[149],s204[150],s204[151],s204[152],s204[153],s204[154],s204[155],s204[156],s204[157],s204[158],s204[159],s204[160],s204[161],s204[162],s204[163],s204[164],s204[165],s204[166],s204[167],s204[168],s204[169],s204[170],s204[171],s204[172],s204[173],s204[174],s204[175],s204[176],s204[177],s204[178],s204[179],s204[180],s204[181],s204[182],s204[183],s204[184],s204[185],s204[186],s204[187],s204[188],s204[189],s204[190],s204[191],s204[192],s204[193],s204[194],s204[195],s204[196],s204[197],s204[198],s204[199],s204[200],s204[201],s204[202],s204[203],s204[204],s204[205],s204[206],s204[207],s204[208],s204[209],s204[210],s204[211],s204[212],s204[213],s204[214],s204[215],s204[216],s204[217],s204[218],s204[219],s204[220],s204[221],s204[222],s204[223],s204[224],s204[225],s204[226],s204[227],s204[228],s204[229],s204[230],s204[231],s204[232],s204[233],s204[234],s204[235],s204[236],s204[237],s204[238],s204[239],s204[240],s204[241],s204[242],s204[243],s204[244],s204[245],s204[246],s204[247],s204[248],s204[249],s204[250],s204[251],s204[252],s204[253],s204[254],s204[255],s204[256],s204[257],s204[258],s204[259],s204[260],s204[261],s204[262],s204[263],s204[264],s204[265],s204[266],s204[267],s204[268],s204[269],s204[270],s204[271],s204[272],s204[273],s204[274],s204[275],s204[276],s204[277],s204[278],s204[279],s204[280],s204[281],s204[282],s204[283],s204[284],s204[285],s204[286],s204[287],s204[288],s204[289],s204[290],s204[291],s203[293],s202[295],s201[297],s200[299],s199[301],s198[303],s197[305],s196[307],s195[309],s194[311],s193[313],s192[219],s191[221],s190[223],s189[225],s188[227],s187[229],s186[231],s185[233],s184[235],s183[237],s182[239],s181[241],s180[243],s179[245],s178[247],s177[249],s176[251],s175[253],s174[255],s173[257],s172[259],s171[261],s170[263],s169[265],s168[267],s167[269],s166[271],s165[273],s164[275],s163[277],s162[279],s161[281],s160[283],s159[285],s158[287],s157[289],s156[291],s155[293],s154[295],s153[297],s152[299],s151[301],s150[303],s149[305],s148[307],s147[309],s146[311],s145[313],s144[315],s143[317],s142[319],s141[321],s140[323],s139[325],s138[327],s137[329],s136[331],s135[333],s134[335],s133[337],s132[339],s131[341],s130[343],s129[345],pp255[155],pp254[157],pp253[159],pp252[161],pp251[163],pp250[165],pp249[167],pp248[169],pp247[171],pp246[173],pp245[175],pp244[177],pp243[179],pp242[181],pp241[183],pp240[185],pp239[187],pp238[189],pp237[191],pp236[193],pp235[195],pp234[197],pp233[199],pp232[201],pp231[203],pp230[205],pp229[207],pp228[209],pp227[211],pp226[213],pp225[215],pp224[217],pp223[219],pp222[221],pp221[223],pp220[225],pp219[227],pp218[229],pp217[231],pp218[231],pp219[231],pp220[231],pp221[231],pp222[231],pp223[231],pp224[231],pp225[231],pp226[231],pp227[231],pp228[231],pp229[231],pp230[231],pp231[231],pp232[231],pp233[231],pp234[231],pp235[231],pp236[231]};
    assign in205_2 = {s193[12],pp35[10],pp35[11],pp35[12],pp35[13],pp35[14],pp35[15],pp35[16],pp35[17],pp35[18],pp35[19],pp35[20],pp35[21],pp35[22],pp35[23],pp35[24],pp35[25],pp35[26],pp35[27],pp35[28],pp37[27],pp39[26],pp41[25],pp43[24],pp45[23],pp47[22],pp49[21],pp51[20],pp53[19],pp55[18],pp57[17],pp59[16],pp61[15],pp63[14],pp65[13],pp67[12],pp69[11],pp71[10],s129[18],s130[18],s131[18],s132[18],s133[18],s134[18],s135[18],s136[18],s137[18],s138[18],s139[18],s140[18],s141[18],s142[18],s143[18],s144[18],s145[18],s146[18],s145[20],s144[22],s143[24],s142[26],s141[28],s140[30],s139[32],s138[34],s137[36],s136[38],s137[38],s138[38],s139[38],s140[38],s141[38],s142[38],s143[38],s144[38],s145[38],s146[38],s147[38],s148[38],s149[38],s150[38],s151[38],s152[38],s153[38],s154[38],s155[38],s156[38],s157[38],s158[38],s158[39],s158[40],s158[41],s158[42],s158[43],s158[44],s158[45],s158[46],s158[47],s158[48],s158[49],s158[50],s159[50],s160[50],s161[50],s162[50],s163[50],s164[50],s165[50],s166[50],s167[50],s168[50],s169[50],s170[50],s171[50],s172[50],s173[50],s174[50],s175[50],s176[50],s177[50],s178[50],s179[50],s180[50],s181[50],s182[50],s183[50],s184[50],s185[50],s186[50],s187[50],s188[50],s189[50],s190[50],s191[50],s192[50],s10[41],s11[41],s12[41],s13[41],s14[41],s15[41],s16[41],s17[41],s18[41],s19[41],s20[41],s21[41],s22[41],s23[41],s24[41],s25[41],s26[41],s27[41],s28[41],s29[41],s30[41],s31[41],s32[41],s33[41],s34[41],s35[41],s36[41],s37[41],s38[41],s39[41],s40[41],s41[41],s42[41],s43[41],s44[41],s45[41],s46[41],s47[41],s48[41],s49[41],s50[41],s51[41],s52[41],s53[41],s54[41],s55[41],s56[41],s57[41],s58[41],s59[41],s59[42],s59[43],s59[44],s59[45],s59[46],s59[47],s59[48],s59[49],s59[50],s59[51],s59[52],s59[53],s59[54],s59[55],s59[56],s59[57],s59[58],s59[59],s59[60],s59[61],s59[62],s59[63],s59[64],s59[65],s59[66],s59[67],s59[68],s59[69],s59[70],s57[73],s55[76],s53[79],s51[82],s50[84],s50[85],s50[86],s50[87],s50[88],s50[89],s50[90],s50[91],s50[92],s50[93],s50[94],s50[95],s50[96],s50[97],s50[98],s50[99],s9[141],s8[143],s7[145],s6[147],s5[149],s4[151],s3[153],s2[155],s1[157],s58[101],s57[103],s56[105],s55[107],s54[109],s53[111],s52[113],s51[115],s50[117],s49[119],s48[121],s47[123],s46[125],s45[127],s44[129],s43[131],s42[133],s41[135],s40[137],s39[139],s38[141],s37[143],s36[145],s35[147],s34[149],s33[151],s32[153],s31[155],s30[157],s29[159],s28[161],s27[163],s26[165],s25[167],s24[169],s23[171],s22[173],s21[175],s20[177],s19[179],s18[181],s17[183],s16[185],s15[187],s14[189],s13[191],s12[193],s11[195],s10[197],s204[292],s203[294],s202[296],s201[298],s200[300],s199[302],s198[304],s197[306],s196[308],s195[310],s194[312],s193[314],s192[220],s191[222],s190[224],s189[226],s188[228],s187[230],s186[232],s185[234],s184[236],s183[238],s182[240],s181[242],s180[244],s179[246],s178[248],s177[250],s176[252],s175[254],s174[256],s173[258],s172[260],s171[262],s170[264],s169[266],s168[268],s167[270],s166[272],s165[274],s164[276],s163[278],s162[280],s161[282],s160[284],s159[286],s158[288],s157[290],s156[292],s155[294],s154[296],s153[298],s152[300],s151[302],s150[304],s149[306],s148[308],s147[310],s146[312],s145[314],s144[316],s143[318],s142[320],s141[322],s140[324],s139[326],s138[328],s137[330],s136[332],s135[334],s134[336],s133[338],s132[340],s131[342],s130[344],s129[346],pp255[156],pp254[158],pp253[160],pp252[162],pp251[164],pp250[166],pp249[168],pp248[170],pp247[172],pp246[174],pp245[176],pp244[178],pp243[180],pp242[182],pp241[184],pp240[186],pp239[188],pp238[190],pp237[192],pp236[194],pp235[196],pp234[198],pp233[200],pp232[202],pp231[204],pp230[206],pp229[208],pp228[210],pp227[212],pp226[214],pp225[216],pp224[218],pp223[220],pp222[222],pp221[224],pp220[226],pp219[228],pp218[230],pp219[230],pp220[230],pp221[230],pp222[230],pp223[230],pp224[230],pp225[230],pp226[230],pp227[230],pp228[230],pp229[230],pp230[230],pp231[230],pp232[230],pp233[230],pp234[230],pp235[230],pp236[230],pp237[230]};
    CLA_424 KS_205(s205, c205, in205_1, in205_2);
    wire[421:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {s193[13],pp36[10],pp36[11],pp36[12],pp36[13],pp36[14],pp36[15],pp36[16],pp36[17],pp36[18],pp36[19],pp36[20],pp36[21],pp36[22],pp36[23],pp36[24],pp36[25],pp36[26],pp36[27],pp38[26],pp40[25],pp42[24],pp44[23],pp46[22],pp48[21],pp50[20],pp52[19],pp54[18],pp56[17],pp58[16],pp60[15],pp62[14],pp64[13],pp66[12],pp68[11],pp70[10],s129[17],s130[17],s131[17],s132[17],s133[17],s134[17],s135[17],s136[17],s137[17],s138[17],s139[17],s140[17],s141[17],s142[17],s143[17],s144[17],s145[17],s146[17],s147[17],s146[19],s145[21],s144[23],s143[25],s142[27],s141[29],s140[31],s139[33],s138[35],s137[37],s138[37],s139[37],s140[37],s141[37],s142[37],s143[37],s144[37],s145[37],s146[37],s147[37],s148[37],s149[37],s150[37],s151[37],s152[37],s153[37],s154[37],s155[37],s156[37],s157[37],s158[37],s159[37],s159[38],s159[39],s159[40],s159[41],s159[42],s159[43],s159[44],s159[45],s159[46],s159[47],s159[48],s159[49],s205[100],s205[101],s205[102],s205[103],s205[104],s205[105],s205[106],s205[107],s205[108],s205[109],s205[110],s205[111],s205[112],s205[113],s205[114],s205[115],s205[116],s205[117],s205[118],s205[119],s205[120],s205[121],s205[122],s205[123],s205[124],s205[125],s205[126],s205[127],s205[128],s205[129],s205[130],s205[131],s205[132],s205[133],s205[134],s205[135],s205[136],s205[137],s205[138],s205[139],s205[140],s205[141],s205[142],s205[143],s205[144],s205[145],s205[146],s205[147],s205[148],s205[149],s205[150],s205[151],s205[152],s205[153],s205[154],s205[155],s205[156],s205[157],s205[158],s205[159],s205[160],s205[161],s205[162],s205[163],s205[164],s205[165],s205[166],s205[167],s205[168],s205[169],s205[170],s205[171],s205[172],s205[173],s205[174],s205[175],s205[176],s205[177],s205[178],s205[179],s205[180],s205[181],s205[182],s205[183],s205[184],s205[185],s205[186],s205[187],s205[188],s205[189],s205[190],s205[191],s205[192],s205[193],s205[194],s205[195],s205[196],s205[197],s205[198],s205[199],s205[200],s205[201],s205[202],s205[203],s205[204],s205[205],s205[206],s205[207],s205[208],s205[209],s205[210],s205[211],s205[212],s205[213],s205[214],s205[215],s205[216],s205[217],s205[218],s205[219],s205[220],s205[221],s205[222],s205[223],s205[224],s205[225],s205[226],s205[227],s205[228],s205[229],s205[230],s205[231],s205[232],s205[233],s205[234],s205[235],s205[236],s205[237],s205[238],s205[239],s205[240],s205[241],s205[242],s205[243],s205[244],s205[245],s205[246],s205[247],s205[248],s205[249],s205[250],s205[251],s205[252],s205[253],s205[254],s205[255],s205[256],s205[257],s205[258],s205[259],s205[260],s205[261],s205[262],s205[263],s205[264],s205[265],s205[266],s205[267],s205[268],s205[269],s205[270],s205[271],s205[272],s205[273],s205[274],s205[275],s205[276],s205[277],s205[278],s205[279],s205[280],s205[281],s205[282],s205[283],s205[284],s205[285],s205[286],s205[287],s205[288],s205[289],s205[290],s205[291],s204[293],s203[295],s202[297],s201[299],s200[301],s199[303],s198[305],s197[307],s196[309],s195[311],s194[313],s193[315],s192[221],s191[223],s190[225],s189[227],s188[229],s187[231],s186[233],s185[235],s184[237],s183[239],s182[241],s181[243],s180[245],s179[247],s178[249],s177[251],s176[253],s175[255],s174[257],s173[259],s172[261],s171[263],s170[265],s169[267],s168[269],s167[271],s166[273],s165[275],s164[277],s163[279],s162[281],s161[283],s160[285],s159[287],s158[289],s157[291],s156[293],s155[295],s154[297],s153[299],s152[301],s151[303],s150[305],s149[307],s148[309],s147[311],s146[313],s145[315],s144[317],s143[319],s142[321],s141[323],s140[325],s139[327],s138[329],s137[331],s136[333],s135[335],s134[337],s133[339],s132[341],s131[343],s130[345],s129[347],pp255[157],pp254[159],pp253[161],pp252[163],pp251[165],pp250[167],pp249[169],pp248[171],pp247[173],pp246[175],pp245[177],pp244[179],pp243[181],pp242[183],pp241[185],pp240[187],pp239[189],pp238[191],pp237[193],pp236[195],pp235[197],pp234[199],pp233[201],pp232[203],pp231[205],pp230[207],pp229[209],pp228[211],pp227[213],pp226[215],pp225[217],pp224[219],pp223[221],pp222[223],pp221[225],pp220[227],pp219[229],pp220[229],pp221[229],pp222[229],pp223[229],pp224[229],pp225[229],pp226[229],pp227[229],pp228[229],pp229[229],pp230[229],pp231[229],pp232[229],pp233[229],pp234[229],pp235[229],pp236[229],pp237[229]};
    assign in206_2 = {s194[12],s193[14],pp37[10],pp37[11],pp37[12],pp37[13],pp37[14],pp37[15],pp37[16],pp37[17],pp37[18],pp37[19],pp37[20],pp37[21],pp37[22],pp37[23],pp37[24],pp37[25],pp37[26],pp39[25],pp41[24],pp43[23],pp45[22],pp47[21],pp49[20],pp51[19],pp53[18],pp55[17],pp57[16],pp59[15],pp61[14],pp63[13],pp65[12],pp67[11],pp69[10],s129[16],s130[16],s131[16],s132[16],s133[16],s134[16],s135[16],s136[16],s137[16],s138[16],s139[16],s140[16],s141[16],s142[16],s143[16],s144[16],s145[16],s146[16],s147[16],s148[16],s147[18],s146[20],s145[22],s144[24],s143[26],s142[28],s141[30],s140[32],s139[34],s138[36],s139[36],s140[36],s141[36],s142[36],s143[36],s144[36],s145[36],s146[36],s147[36],s148[36],s149[36],s150[36],s151[36],s152[36],s153[36],s154[36],s155[36],s156[36],s157[36],s158[36],s159[36],s160[36],s160[37],s160[38],s160[39],s160[40],s160[41],s160[42],s160[43],s160[44],s160[45],s160[46],s160[47],s160[48],s160[49],s161[49],s162[49],s163[49],s164[49],s165[49],s166[49],s167[49],s168[49],s169[49],s170[49],s171[49],s172[49],s173[49],s174[49],s175[49],s176[49],s177[49],s178[49],s179[49],s180[49],s181[49],s182[49],s183[49],s184[49],s185[49],s186[49],s187[49],s188[49],s189[49],s190[49],s191[49],s192[49],s10[40],s11[40],s12[40],s13[40],s14[40],s15[40],s16[40],s17[40],s18[40],s19[40],s20[40],s21[40],s22[40],s23[40],s24[40],s25[40],s26[40],s27[40],s28[40],s29[40],s30[40],s31[40],s32[40],s33[40],s34[40],s35[40],s36[40],s37[40],s38[40],s39[40],s40[40],s41[40],s42[40],s43[40],s44[40],s45[40],s46[40],s47[40],s48[40],s49[40],s50[40],s51[40],s52[40],s53[40],s54[40],s55[40],s56[40],s57[40],s58[40],s59[40],s60[40],s60[41],s60[42],s60[43],s60[44],s60[45],s60[46],s60[47],s60[48],s60[49],s60[50],s60[51],s60[52],s60[53],s60[54],s60[55],s60[56],s60[57],s60[58],s60[59],s60[60],s60[61],s60[62],s60[63],s60[64],s60[65],s60[66],s60[67],s60[68],s60[69],s58[72],s56[75],s54[78],s52[81],s51[83],s51[84],s51[85],s51[86],s51[87],s51[88],s51[89],s51[90],s51[91],s51[92],s51[93],s51[94],s51[95],s51[96],s51[97],s51[98],s51[99],s9[142],s8[144],s7[146],s6[148],s5[150],s4[152],s3[154],s2[156],s59[100],s58[102],s57[104],s56[106],s55[108],s54[110],s53[112],s52[114],s51[116],s50[118],s49[120],s48[122],s47[124],s46[126],s45[128],s44[130],s43[132],s42[134],s41[136],s40[138],s39[140],s38[142],s37[144],s36[146],s35[148],s34[150],s33[152],s32[154],s31[156],s30[158],s29[160],s28[162],s27[164],s26[166],s25[168],s24[170],s23[172],s22[174],s21[176],s20[178],s19[180],s18[182],s17[184],s16[186],s15[188],s14[190],s13[192],s12[194],s11[196],s10[198],s205[292],s204[294],s203[296],s202[298],s201[300],s200[302],s199[304],s198[306],s197[308],s196[310],s195[312],s194[314],s193[316],s192[222],s191[224],s190[226],s189[228],s188[230],s187[232],s186[234],s185[236],s184[238],s183[240],s182[242],s181[244],s180[246],s179[248],s178[250],s177[252],s176[254],s175[256],s174[258],s173[260],s172[262],s171[264],s170[266],s169[268],s168[270],s167[272],s166[274],s165[276],s164[278],s163[280],s162[282],s161[284],s160[286],s159[288],s158[290],s157[292],s156[294],s155[296],s154[298],s153[300],s152[302],s151[304],s150[306],s149[308],s148[310],s147[312],s146[314],s145[316],s144[318],s143[320],s142[322],s141[324],s140[326],s139[328],s138[330],s137[332],s136[334],s135[336],s134[338],s133[340],s132[342],s131[344],s130[346],s129[348],pp255[158],pp254[160],pp253[162],pp252[164],pp251[166],pp250[168],pp249[170],pp248[172],pp247[174],pp246[176],pp245[178],pp244[180],pp243[182],pp242[184],pp241[186],pp240[188],pp239[190],pp238[192],pp237[194],pp236[196],pp235[198],pp234[200],pp233[202],pp232[204],pp231[206],pp230[208],pp229[210],pp228[212],pp227[214],pp226[216],pp225[218],pp224[220],pp223[222],pp222[224],pp221[226],pp220[228],pp221[228],pp222[228],pp223[228],pp224[228],pp225[228],pp226[228],pp227[228],pp228[228],pp229[228],pp230[228],pp231[228],pp232[228],pp233[228],pp234[228],pp235[228],pp236[228],pp237[228],pp238[228]};
    CLA_422 KS_206(s206, c206, in206_1, in206_2);
    wire[419:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {s194[13],s193[15],pp38[10],pp38[11],pp38[12],pp38[13],pp38[14],pp38[15],pp38[16],pp38[17],pp38[18],pp38[19],pp38[20],pp38[21],pp38[22],pp38[23],pp38[24],pp38[25],pp40[24],pp42[23],pp44[22],pp46[21],pp48[20],pp50[19],pp52[18],pp54[17],pp56[16],pp58[15],pp60[14],pp62[13],pp64[12],pp66[11],pp68[10],s129[15],s130[15],s131[15],s132[15],s133[15],s134[15],s135[15],s136[15],s137[15],s138[15],s139[15],s140[15],s141[15],s142[15],s143[15],s144[15],s145[15],s146[15],s147[15],s148[15],s149[15],s148[17],s147[19],s146[21],s145[23],s144[25],s143[27],s142[29],s141[31],s140[33],s139[35],s140[35],s141[35],s142[35],s143[35],s144[35],s145[35],s146[35],s147[35],s148[35],s149[35],s150[35],s151[35],s152[35],s153[35],s154[35],s155[35],s156[35],s157[35],s158[35],s159[35],s160[35],s161[35],s161[36],s161[37],s161[38],s161[39],s161[40],s161[41],s161[42],s161[43],s161[44],s161[45],s161[46],s161[47],s161[48],s206[100],s206[101],s206[102],s206[103],s206[104],s206[105],s206[106],s206[107],s206[108],s206[109],s206[110],s206[111],s206[112],s206[113],s206[114],s206[115],s206[116],s206[117],s206[118],s206[119],s206[120],s206[121],s206[122],s206[123],s206[124],s206[125],s206[126],s206[127],s206[128],s206[129],s206[130],s206[131],s206[132],s206[133],s206[134],s206[135],s206[136],s206[137],s206[138],s206[139],s206[140],s206[141],s206[142],s206[143],s206[144],s206[145],s206[146],s206[147],s206[148],s206[149],s206[150],s206[151],s206[152],s206[153],s206[154],s206[155],s206[156],s206[157],s206[158],s206[159],s206[160],s206[161],s206[162],s206[163],s206[164],s206[165],s206[166],s206[167],s206[168],s206[169],s206[170],s206[171],s206[172],s206[173],s206[174],s206[175],s206[176],s206[177],s206[178],s206[179],s206[180],s206[181],s206[182],s206[183],s206[184],s206[185],s206[186],s206[187],s206[188],s206[189],s206[190],s206[191],s206[192],s206[193],s206[194],s206[195],s206[196],s206[197],s206[198],s206[199],s206[200],s206[201],s206[202],s206[203],s206[204],s206[205],s206[206],s206[207],s206[208],s206[209],s206[210],s206[211],s206[212],s206[213],s206[214],s206[215],s206[216],s206[217],s206[218],s206[219],s206[220],s206[221],s206[222],s206[223],s206[224],s206[225],s206[226],s206[227],s206[228],s206[229],s206[230],s206[231],s206[232],s206[233],s206[234],s206[235],s206[236],s206[237],s206[238],s206[239],s206[240],s206[241],s206[242],s206[243],s206[244],s206[245],s206[246],s206[247],s206[248],s206[249],s206[250],s206[251],s206[252],s206[253],s206[254],s206[255],s206[256],s206[257],s206[258],s206[259],s206[260],s206[261],s206[262],s206[263],s206[264],s206[265],s206[266],s206[267],s206[268],s206[269],s206[270],s206[271],s206[272],s206[273],s206[274],s206[275],s206[276],s206[277],s206[278],s206[279],s206[280],s206[281],s206[282],s206[283],s206[284],s206[285],s206[286],s206[287],s206[288],s206[289],s206[290],s206[291],s205[293],s204[295],s203[297],s202[299],s201[301],s200[303],s199[305],s198[307],s197[309],s196[311],s195[313],s194[315],s193[317],s192[223],s191[225],s190[227],s189[229],s188[231],s187[233],s186[235],s185[237],s184[239],s183[241],s182[243],s181[245],s180[247],s179[249],s178[251],s177[253],s176[255],s175[257],s174[259],s173[261],s172[263],s171[265],s170[267],s169[269],s168[271],s167[273],s166[275],s165[277],s164[279],s163[281],s162[283],s161[285],s160[287],s159[289],s158[291],s157[293],s156[295],s155[297],s154[299],s153[301],s152[303],s151[305],s150[307],s149[309],s148[311],s147[313],s146[315],s145[317],s144[319],s143[321],s142[323],s141[325],s140[327],s139[329],s138[331],s137[333],s136[335],s135[337],s134[339],s133[341],s132[343],s131[345],s130[347],s129[349],pp255[159],pp254[161],pp253[163],pp252[165],pp251[167],pp250[169],pp249[171],pp248[173],pp247[175],pp246[177],pp245[179],pp244[181],pp243[183],pp242[185],pp241[187],pp240[189],pp239[191],pp238[193],pp237[195],pp236[197],pp235[199],pp234[201],pp233[203],pp232[205],pp231[207],pp230[209],pp229[211],pp228[213],pp227[215],pp226[217],pp225[219],pp224[221],pp223[223],pp222[225],pp221[227],pp222[227],pp223[227],pp224[227],pp225[227],pp226[227],pp227[227],pp228[227],pp229[227],pp230[227],pp231[227],pp232[227],pp233[227],pp234[227],pp235[227],pp236[227],pp237[227],pp238[227]};
    assign in207_2 = {s195[12],s194[14],s193[16],pp39[10],pp39[11],pp39[12],pp39[13],pp39[14],pp39[15],pp39[16],pp39[17],pp39[18],pp39[19],pp39[20],pp39[21],pp39[22],pp39[23],pp39[24],pp41[23],pp43[22],pp45[21],pp47[20],pp49[19],pp51[18],pp53[17],pp55[16],pp57[15],pp59[14],pp61[13],pp63[12],pp65[11],pp67[10],s129[14],s130[14],s131[14],s132[14],s133[14],s134[14],s135[14],s136[14],s137[14],s138[14],s139[14],s140[14],s141[14],s142[14],s143[14],s144[14],s145[14],s146[14],s147[14],s148[14],s149[14],s150[14],s149[16],s148[18],s147[20],s146[22],s145[24],s144[26],s143[28],s142[30],s141[32],s140[34],s141[34],s142[34],s143[34],s144[34],s145[34],s146[34],s147[34],s148[34],s149[34],s150[34],s151[34],s152[34],s153[34],s154[34],s155[34],s156[34],s157[34],s158[34],s159[34],s160[34],s161[34],s162[34],s162[35],s162[36],s162[37],s162[38],s162[39],s162[40],s162[41],s162[42],s162[43],s162[44],s162[45],s162[46],s162[47],s162[48],s163[48],s164[48],s165[48],s166[48],s167[48],s168[48],s169[48],s170[48],s171[48],s172[48],s173[48],s174[48],s175[48],s176[48],s177[48],s178[48],s179[48],s180[48],s181[48],s182[48],s183[48],s184[48],s185[48],s186[48],s187[48],s188[48],s189[48],s190[48],s191[48],s192[48],s10[39],s11[39],s12[39],s13[39],s14[39],s15[39],s16[39],s17[39],s18[39],s19[39],s20[39],s21[39],s22[39],s23[39],s24[39],s25[39],s26[39],s27[39],s28[39],s29[39],s30[39],s31[39],s32[39],s33[39],s34[39],s35[39],s36[39],s37[39],s38[39],s39[39],s40[39],s41[39],s42[39],s43[39],s44[39],s45[39],s46[39],s47[39],s48[39],s49[39],s50[39],s51[39],s52[39],s53[39],s54[39],s55[39],s56[39],s57[39],s58[39],s59[39],s60[39],s61[39],s61[40],s61[41],s61[42],s61[43],s61[44],s61[45],s61[46],s61[47],s61[48],s61[49],s61[50],s61[51],s61[52],s61[53],s61[54],s61[55],s61[56],s61[57],s61[58],s61[59],s61[60],s61[61],s61[62],s61[63],s61[64],s61[65],s61[66],s61[67],s61[68],s59[71],s57[74],s55[77],s53[80],s52[82],s52[83],s52[84],s52[85],s52[86],s52[87],s52[88],s52[89],s52[90],s52[91],s52[92],s52[93],s52[94],s52[95],s52[96],s52[97],s52[98],s52[99],s9[143],s8[145],s7[147],s6[149],s5[151],s4[153],s3[155],s1[158],s59[101],s58[103],s57[105],s56[107],s55[109],s54[111],s53[113],s52[115],s51[117],s50[119],s49[121],s48[123],s47[125],s46[127],s45[129],s44[131],s43[133],s42[135],s41[137],s40[139],s39[141],s38[143],s37[145],s36[147],s35[149],s34[151],s33[153],s32[155],s31[157],s30[159],s29[161],s28[163],s27[165],s26[167],s25[169],s24[171],s23[173],s22[175],s21[177],s20[179],s19[181],s18[183],s17[185],s16[187],s15[189],s14[191],s13[193],s12[195],s11[197],s10[199],s206[292],s205[294],s204[296],s203[298],s202[300],s201[302],s200[304],s199[306],s198[308],s197[310],s196[312],s195[314],s194[316],s193[318],s192[224],s191[226],s190[228],s189[230],s188[232],s187[234],s186[236],s185[238],s184[240],s183[242],s182[244],s181[246],s180[248],s179[250],s178[252],s177[254],s176[256],s175[258],s174[260],s173[262],s172[264],s171[266],s170[268],s169[270],s168[272],s167[274],s166[276],s165[278],s164[280],s163[282],s162[284],s161[286],s160[288],s159[290],s158[292],s157[294],s156[296],s155[298],s154[300],s153[302],s152[304],s151[306],s150[308],s149[310],s148[312],s147[314],s146[316],s145[318],s144[320],s143[322],s142[324],s141[326],s140[328],s139[330],s138[332],s137[334],s136[336],s135[338],s134[340],s133[342],s132[344],s131[346],s130[348],s129[350],pp255[160],pp254[162],pp253[164],pp252[166],pp251[168],pp250[170],pp249[172],pp248[174],pp247[176],pp246[178],pp245[180],pp244[182],pp243[184],pp242[186],pp241[188],pp240[190],pp239[192],pp238[194],pp237[196],pp236[198],pp235[200],pp234[202],pp233[204],pp232[206],pp231[208],pp230[210],pp229[212],pp228[214],pp227[216],pp226[218],pp225[220],pp224[222],pp223[224],pp222[226],pp223[226],pp224[226],pp225[226],pp226[226],pp227[226],pp228[226],pp229[226],pp230[226],pp231[226],pp232[226],pp233[226],pp234[226],pp235[226],pp236[226],pp237[226],pp238[226],pp239[226]};
    CLA_420 KS_207(s207, c207, in207_1, in207_2);
    wire[417:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {s195[13],s194[15],s193[17],pp40[10],pp40[11],pp40[12],pp40[13],pp40[14],pp40[15],pp40[16],pp40[17],pp40[18],pp40[19],pp40[20],pp40[21],pp40[22],pp40[23],pp42[22],pp44[21],pp46[20],pp48[19],pp50[18],pp52[17],pp54[16],pp56[15],pp58[14],pp60[13],pp62[12],pp64[11],pp66[10],s129[13],s130[13],s131[13],s132[13],s133[13],s134[13],s135[13],s136[13],s137[13],s138[13],s139[13],s140[13],s141[13],s142[13],s143[13],s144[13],s145[13],s146[13],s147[13],s148[13],s149[13],s150[13],s151[13],s150[15],s149[17],s148[19],s147[21],s146[23],s145[25],s144[27],s143[29],s142[31],s141[33],s142[33],s143[33],s144[33],s145[33],s146[33],s147[33],s148[33],s149[33],s150[33],s151[33],s152[33],s153[33],s154[33],s155[33],s156[33],s157[33],s158[33],s159[33],s160[33],s161[33],s162[33],s163[33],s163[34],s163[35],s163[36],s163[37],s163[38],s163[39],s163[40],s163[41],s163[42],s163[43],s163[44],s163[45],s163[46],s163[47],s207[100],s207[101],s207[102],s207[103],s207[104],s207[105],s207[106],s207[107],s207[108],s207[109],s207[110],s207[111],s207[112],s207[113],s207[114],s207[115],s207[116],s207[117],s207[118],s207[119],s207[120],s207[121],s207[122],s207[123],s207[124],s207[125],s207[126],s207[127],s207[128],s207[129],s207[130],s207[131],s207[132],s207[133],s207[134],s207[135],s207[136],s207[137],s207[138],s207[139],s207[140],s207[141],s207[142],s207[143],s207[144],s207[145],s207[146],s207[147],s207[148],s207[149],s207[150],s207[151],s207[152],s207[153],s207[154],s207[155],s207[156],s207[157],s207[158],s207[159],s207[160],s207[161],s207[162],s207[163],s207[164],s207[165],s207[166],s207[167],s207[168],s207[169],s207[170],s207[171],s207[172],s207[173],s207[174],s207[175],s207[176],s207[177],s207[178],s207[179],s207[180],s207[181],s207[182],s207[183],s207[184],s207[185],s207[186],s207[187],s207[188],s207[189],s207[190],s207[191],s207[192],s207[193],s207[194],s207[195],s207[196],s207[197],s207[198],s207[199],s207[200],s207[201],s207[202],s207[203],s207[204],s207[205],s207[206],s207[207],s207[208],s207[209],s207[210],s207[211],s207[212],s207[213],s207[214],s207[215],s207[216],s207[217],s207[218],s207[219],s207[220],s207[221],s207[222],s207[223],s207[224],s207[225],s207[226],s207[227],s207[228],s207[229],s207[230],s207[231],s207[232],s207[233],s207[234],s207[235],s207[236],s207[237],s207[238],s207[239],s207[240],s207[241],s207[242],s207[243],s207[244],s207[245],s207[246],s207[247],s207[248],s207[249],s207[250],s207[251],s207[252],s207[253],s207[254],s207[255],s207[256],s207[257],s207[258],s207[259],s207[260],s207[261],s207[262],s207[263],s207[264],s207[265],s207[266],s207[267],s207[268],s207[269],s207[270],s207[271],s207[272],s207[273],s207[274],s207[275],s207[276],s207[277],s207[278],s207[279],s207[280],s207[281],s207[282],s207[283],s207[284],s207[285],s207[286],s207[287],s207[288],s207[289],s207[290],s207[291],s206[293],s205[295],s204[297],s203[299],s202[301],s201[303],s200[305],s199[307],s198[309],s197[311],s196[313],s195[315],s194[317],s193[319],s192[225],s191[227],s190[229],s189[231],s188[233],s187[235],s186[237],s185[239],s184[241],s183[243],s182[245],s181[247],s180[249],s179[251],s178[253],s177[255],s176[257],s175[259],s174[261],s173[263],s172[265],s171[267],s170[269],s169[271],s168[273],s167[275],s166[277],s165[279],s164[281],s163[283],s162[285],s161[287],s160[289],s159[291],s158[293],s157[295],s156[297],s155[299],s154[301],s153[303],s152[305],s151[307],s150[309],s149[311],s148[313],s147[315],s146[317],s145[319],s144[321],s143[323],s142[325],s141[327],s140[329],s139[331],s138[333],s137[335],s136[337],s135[339],s134[341],s133[343],s132[345],s131[347],s130[349],s129[351],pp255[161],pp254[163],pp253[165],pp252[167],pp251[169],pp250[171],pp249[173],pp248[175],pp247[177],pp246[179],pp245[181],pp244[183],pp243[185],pp242[187],pp241[189],pp240[191],pp239[193],pp238[195],pp237[197],pp236[199],pp235[201],pp234[203],pp233[205],pp232[207],pp231[209],pp230[211],pp229[213],pp228[215],pp227[217],pp226[219],pp225[221],pp224[223],pp223[225],pp224[225],pp225[225],pp226[225],pp227[225],pp228[225],pp229[225],pp230[225],pp231[225],pp232[225],pp233[225],pp234[225],pp235[225],pp236[225],pp237[225],pp238[225],pp239[225]};
    assign in208_2 = {s196[12],s195[14],s194[16],s193[18],pp41[10],pp41[11],pp41[12],pp41[13],pp41[14],pp41[15],pp41[16],pp41[17],pp41[18],pp41[19],pp41[20],pp41[21],pp41[22],pp43[21],pp45[20],pp47[19],pp49[18],pp51[17],pp53[16],pp55[15],pp57[14],pp59[13],pp61[12],pp63[11],pp65[10],s129[12],s130[12],s131[12],s132[12],s133[12],s134[12],s135[12],s136[12],s137[12],s138[12],s139[12],s140[12],s141[12],s142[12],s143[12],s144[12],s145[12],s146[12],s147[12],s148[12],s149[12],s150[12],s151[12],s152[12],s151[14],s150[16],s149[18],s148[20],s147[22],s146[24],s145[26],s144[28],s143[30],s142[32],s143[32],s144[32],s145[32],s146[32],s147[32],s148[32],s149[32],s150[32],s151[32],s152[32],s153[32],s154[32],s155[32],s156[32],s157[32],s158[32],s159[32],s160[32],s161[32],s162[32],s163[32],s164[32],s164[33],s164[34],s164[35],s164[36],s164[37],s164[38],s164[39],s164[40],s164[41],s164[42],s164[43],s164[44],s164[45],s164[46],s164[47],s165[47],s166[47],s167[47],s168[47],s169[47],s170[47],s171[47],s172[47],s173[47],s174[47],s175[47],s176[47],s177[47],s178[47],s179[47],s180[47],s181[47],s182[47],s183[47],s184[47],s185[47],s186[47],s187[47],s188[47],s189[47],s190[47],s191[47],s192[47],s10[38],s11[38],s12[38],s13[38],s14[38],s15[38],s16[38],s17[38],s18[38],s19[38],s20[38],s21[38],s22[38],s23[38],s24[38],s25[38],s26[38],s27[38],s28[38],s29[38],s30[38],s31[38],s32[38],s33[38],s34[38],s35[38],s36[38],s37[38],s38[38],s39[38],s40[38],s41[38],s42[38],s43[38],s44[38],s45[38],s46[38],s47[38],s48[38],s49[38],s50[38],s51[38],s52[38],s53[38],s54[38],s55[38],s56[38],s57[38],s58[38],s59[38],s60[38],s61[38],s62[38],s62[39],s62[40],s62[41],s62[42],s62[43],s62[44],s62[45],s62[46],s62[47],s62[48],s62[49],s62[50],s62[51],s62[52],s62[53],s62[54],s62[55],s62[56],s62[57],s62[58],s62[59],s62[60],s62[61],s62[62],s62[63],s62[64],s62[65],s62[66],s62[67],s60[70],s58[73],s56[76],s54[79],s53[81],s53[82],s53[83],s53[84],s53[85],s53[86],s53[87],s53[88],s53[89],s53[90],s53[91],s53[92],s53[93],s53[94],s53[95],s53[96],s53[97],s53[98],s53[99],s9[144],s8[146],s7[148],s6[150],s5[152],s4[154],s2[157],s60[100],s59[102],s58[104],s57[106],s56[108],s55[110],s54[112],s53[114],s52[116],s51[118],s50[120],s49[122],s48[124],s47[126],s46[128],s45[130],s44[132],s43[134],s42[136],s41[138],s40[140],s39[142],s38[144],s37[146],s36[148],s35[150],s34[152],s33[154],s32[156],s31[158],s30[160],s29[162],s28[164],s27[166],s26[168],s25[170],s24[172],s23[174],s22[176],s21[178],s20[180],s19[182],s18[184],s17[186],s16[188],s15[190],s14[192],s13[194],s12[196],s11[198],s10[200],s207[292],s206[294],s205[296],s204[298],s203[300],s202[302],s201[304],s200[306],s199[308],s198[310],s197[312],s196[314],s195[316],s194[318],s193[320],s192[226],s191[228],s190[230],s189[232],s188[234],s187[236],s186[238],s185[240],s184[242],s183[244],s182[246],s181[248],s180[250],s179[252],s178[254],s177[256],s176[258],s175[260],s174[262],s173[264],s172[266],s171[268],s170[270],s169[272],s168[274],s167[276],s166[278],s165[280],s164[282],s163[284],s162[286],s161[288],s160[290],s159[292],s158[294],s157[296],s156[298],s155[300],s154[302],s153[304],s152[306],s151[308],s150[310],s149[312],s148[314],s147[316],s146[318],s145[320],s144[322],s143[324],s142[326],s141[328],s140[330],s139[332],s138[334],s137[336],s136[338],s135[340],s134[342],s133[344],s132[346],s131[348],s130[350],s129[352],pp255[162],pp254[164],pp253[166],pp252[168],pp251[170],pp250[172],pp249[174],pp248[176],pp247[178],pp246[180],pp245[182],pp244[184],pp243[186],pp242[188],pp241[190],pp240[192],pp239[194],pp238[196],pp237[198],pp236[200],pp235[202],pp234[204],pp233[206],pp232[208],pp231[210],pp230[212],pp229[214],pp228[216],pp227[218],pp226[220],pp225[222],pp224[224],pp225[224],pp226[224],pp227[224],pp228[224],pp229[224],pp230[224],pp231[224],pp232[224],pp233[224],pp234[224],pp235[224],pp236[224],pp237[224],pp238[224],pp239[224],pp240[224]};
    CLA_418 KS_208(s208, c208, in208_1, in208_2);
    wire[415:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {s196[13],s195[15],s194[17],s193[19],pp42[10],pp42[11],pp42[12],pp42[13],pp42[14],pp42[15],pp42[16],pp42[17],pp42[18],pp42[19],pp42[20],pp42[21],pp44[20],pp46[19],pp48[18],pp50[17],pp52[16],pp54[15],pp56[14],pp58[13],pp60[12],pp62[11],pp64[10],s129[11],s130[11],s131[11],s132[11],s133[11],s134[11],s135[11],s136[11],s137[11],s138[11],s139[11],s140[11],s141[11],s142[11],s143[11],s144[11],s145[11],s146[11],s147[11],s148[11],s149[11],s150[11],s151[11],s152[11],s153[11],s152[13],s151[15],s150[17],s149[19],s148[21],s147[23],s146[25],s145[27],s144[29],s143[31],s144[31],s145[31],s146[31],s147[31],s148[31],s149[31],s150[31],s151[31],s152[31],s153[31],s154[31],s155[31],s156[31],s157[31],s158[31],s159[31],s160[31],s161[31],s162[31],s163[31],s164[31],s165[31],s165[32],s165[33],s165[34],s165[35],s165[36],s165[37],s165[38],s165[39],s165[40],s165[41],s165[42],s165[43],s165[44],s165[45],s165[46],s208[100],s208[101],s208[102],s208[103],s208[104],s208[105],s208[106],s208[107],s208[108],s208[109],s208[110],s208[111],s208[112],s208[113],s208[114],s208[115],s208[116],s208[117],s208[118],s208[119],s208[120],s208[121],s208[122],s208[123],s208[124],s208[125],s208[126],s208[127],s208[128],s208[129],s208[130],s208[131],s208[132],s208[133],s208[134],s208[135],s208[136],s208[137],s208[138],s208[139],s208[140],s208[141],s208[142],s208[143],s208[144],s208[145],s208[146],s208[147],s208[148],s208[149],s208[150],s208[151],s208[152],s208[153],s208[154],s208[155],s208[156],s208[157],s208[158],s208[159],s208[160],s208[161],s208[162],s208[163],s208[164],s208[165],s208[166],s208[167],s208[168],s208[169],s208[170],s208[171],s208[172],s208[173],s208[174],s208[175],s208[176],s208[177],s208[178],s208[179],s208[180],s208[181],s208[182],s208[183],s208[184],s208[185],s208[186],s208[187],s208[188],s208[189],s208[190],s208[191],s208[192],s208[193],s208[194],s208[195],s208[196],s208[197],s208[198],s208[199],s208[200],s208[201],s208[202],s208[203],s208[204],s208[205],s208[206],s208[207],s208[208],s208[209],s208[210],s208[211],s208[212],s208[213],s208[214],s208[215],s208[216],s208[217],s208[218],s208[219],s208[220],s208[221],s208[222],s208[223],s208[224],s208[225],s208[226],s208[227],s208[228],s208[229],s208[230],s208[231],s208[232],s208[233],s208[234],s208[235],s208[236],s208[237],s208[238],s208[239],s208[240],s208[241],s208[242],s208[243],s208[244],s208[245],s208[246],s208[247],s208[248],s208[249],s208[250],s208[251],s208[252],s208[253],s208[254],s208[255],s208[256],s208[257],s208[258],s208[259],s208[260],s208[261],s208[262],s208[263],s208[264],s208[265],s208[266],s208[267],s208[268],s208[269],s208[270],s208[271],s208[272],s208[273],s208[274],s208[275],s208[276],s208[277],s208[278],s208[279],s208[280],s208[281],s208[282],s208[283],s208[284],s208[285],s208[286],s208[287],s208[288],s208[289],s208[290],s208[291],s207[293],s206[295],s205[297],s204[299],s203[301],s202[303],s201[305],s200[307],s199[309],s198[311],s197[313],s196[315],s195[317],s194[319],s193[321],s192[227],s191[229],s190[231],s189[233],s188[235],s187[237],s186[239],s185[241],s184[243],s183[245],s182[247],s181[249],s180[251],s179[253],s178[255],s177[257],s176[259],s175[261],s174[263],s173[265],s172[267],s171[269],s170[271],s169[273],s168[275],s167[277],s166[279],s165[281],s164[283],s163[285],s162[287],s161[289],s160[291],s159[293],s158[295],s157[297],s156[299],s155[301],s154[303],s153[305],s152[307],s151[309],s150[311],s149[313],s148[315],s147[317],s146[319],s145[321],s144[323],s143[325],s142[327],s141[329],s140[331],s139[333],s138[335],s137[337],s136[339],s135[341],s134[343],s133[345],s132[347],s131[349],s130[351],s129[353],pp255[163],pp254[165],pp253[167],pp252[169],pp251[171],pp250[173],pp249[175],pp248[177],pp247[179],pp246[181],pp245[183],pp244[185],pp243[187],pp242[189],pp241[191],pp240[193],pp239[195],pp238[197],pp237[199],pp236[201],pp235[203],pp234[205],pp233[207],pp232[209],pp231[211],pp230[213],pp229[215],pp228[217],pp227[219],pp226[221],pp225[223],pp226[223],pp227[223],pp228[223],pp229[223],pp230[223],pp231[223],pp232[223],pp233[223],pp234[223],pp235[223],pp236[223],pp237[223],pp238[223],pp239[223],pp240[223]};
    assign in209_2 = {s197[12],s196[14],s195[16],s194[18],s193[20],pp43[10],pp43[11],pp43[12],pp43[13],pp43[14],pp43[15],pp43[16],pp43[17],pp43[18],pp43[19],pp43[20],pp45[19],pp47[18],pp49[17],pp51[16],pp53[15],pp55[14],pp57[13],pp59[12],pp61[11],pp63[10],s129[10],s130[10],s131[10],s132[10],s133[10],s134[10],s135[10],s136[10],s137[10],s138[10],s139[10],s140[10],s141[10],s142[10],s143[10],s144[10],s145[10],s146[10],s147[10],s148[10],s149[10],s150[10],s151[10],s152[10],s153[10],s154[10],s153[12],s152[14],s151[16],s150[18],s149[20],s148[22],s147[24],s146[26],s145[28],s144[30],s145[30],s146[30],s147[30],s148[30],s149[30],s150[30],s151[30],s152[30],s153[30],s154[30],s155[30],s156[30],s157[30],s158[30],s159[30],s160[30],s161[30],s162[30],s163[30],s164[30],s165[30],s166[30],s166[31],s166[32],s166[33],s166[34],s166[35],s166[36],s166[37],s166[38],s166[39],s166[40],s166[41],s166[42],s166[43],s166[44],s166[45],s166[46],s167[46],s168[46],s169[46],s170[46],s171[46],s172[46],s173[46],s174[46],s175[46],s176[46],s177[46],s178[46],s179[46],s180[46],s181[46],s182[46],s183[46],s184[46],s185[46],s186[46],s187[46],s188[46],s189[46],s190[46],s191[46],s192[46],s10[37],s11[37],s12[37],s13[37],s14[37],s15[37],s16[37],s17[37],s18[37],s19[37],s20[37],s21[37],s22[37],s23[37],s24[37],s25[37],s26[37],s27[37],s28[37],s29[37],s30[37],s31[37],s32[37],s33[37],s34[37],s35[37],s36[37],s37[37],s38[37],s39[37],s40[37],s41[37],s42[37],s43[37],s44[37],s45[37],s46[37],s47[37],s48[37],s49[37],s50[37],s51[37],s52[37],s53[37],s54[37],s55[37],s56[37],s57[37],s58[37],s59[37],s60[37],s61[37],s62[37],s63[37],s63[38],s63[39],s63[40],s63[41],s63[42],s63[43],s63[44],s63[45],s63[46],s63[47],s63[48],s63[49],s63[50],s63[51],s63[52],s63[53],s63[54],s63[55],s63[56],s63[57],s63[58],s63[59],s63[60],s63[61],s63[62],s63[63],s63[64],s63[65],s63[66],s61[69],s59[72],s57[75],s55[78],s54[80],s54[81],s54[82],s54[83],s54[84],s54[85],s54[86],s54[87],s54[88],s54[89],s54[90],s54[91],s54[92],s54[93],s54[94],s54[95],s54[96],s54[97],s54[98],s54[99],s9[145],s8[147],s7[149],s6[151],s5[153],s3[156],s1[159],s60[101],s59[103],s58[105],s57[107],s56[109],s55[111],s54[113],s53[115],s52[117],s51[119],s50[121],s49[123],s48[125],s47[127],s46[129],s45[131],s44[133],s43[135],s42[137],s41[139],s40[141],s39[143],s38[145],s37[147],s36[149],s35[151],s34[153],s33[155],s32[157],s31[159],s30[161],s29[163],s28[165],s27[167],s26[169],s25[171],s24[173],s23[175],s22[177],s21[179],s20[181],s19[183],s18[185],s17[187],s16[189],s15[191],s14[193],s13[195],s12[197],s11[199],s10[201],s208[292],s207[294],s206[296],s205[298],s204[300],s203[302],s202[304],s201[306],s200[308],s199[310],s198[312],s197[314],s196[316],s195[318],s194[320],s193[322],s192[228],s191[230],s190[232],s189[234],s188[236],s187[238],s186[240],s185[242],s184[244],s183[246],s182[248],s181[250],s180[252],s179[254],s178[256],s177[258],s176[260],s175[262],s174[264],s173[266],s172[268],s171[270],s170[272],s169[274],s168[276],s167[278],s166[280],s165[282],s164[284],s163[286],s162[288],s161[290],s160[292],s159[294],s158[296],s157[298],s156[300],s155[302],s154[304],s153[306],s152[308],s151[310],s150[312],s149[314],s148[316],s147[318],s146[320],s145[322],s144[324],s143[326],s142[328],s141[330],s140[332],s139[334],s138[336],s137[338],s136[340],s135[342],s134[344],s133[346],s132[348],s131[350],s130[352],s129[354],pp255[164],pp254[166],pp253[168],pp252[170],pp251[172],pp250[174],pp249[176],pp248[178],pp247[180],pp246[182],pp245[184],pp244[186],pp243[188],pp242[190],pp241[192],pp240[194],pp239[196],pp238[198],pp237[200],pp236[202],pp235[204],pp234[206],pp233[208],pp232[210],pp231[212],pp230[214],pp229[216],pp228[218],pp227[220],pp226[222],pp227[222],pp228[222],pp229[222],pp230[222],pp231[222],pp232[222],pp233[222],pp234[222],pp235[222],pp236[222],pp237[222],pp238[222],pp239[222],pp240[222],pp241[222]};
    CLA_416 KS_209(s209, c209, in209_1, in209_2);
    wire[413:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {s197[13],s196[15],s195[17],s194[19],s193[21],pp44[10],pp44[11],pp44[12],pp44[13],pp44[14],pp44[15],pp44[16],pp44[17],pp44[18],pp44[19],pp46[18],pp48[17],pp50[16],pp52[15],pp54[14],pp56[13],pp58[12],pp60[11],pp62[10],s193[41],s193[42],s193[43],s193[44],s193[45],s193[46],s193[47],s193[48],s193[49],s193[50],s193[51],s193[52],s193[53],s193[54],s193[55],s193[56],s193[57],s193[58],s193[59],s193[60],s193[61],s193[62],s193[63],s193[64],s193[65],s193[66],s193[67],s154[11],s153[13],s152[15],s151[17],s150[19],s149[21],s148[23],s147[25],s146[27],s145[29],s146[29],s147[29],s148[29],s149[29],s150[29],s151[29],s152[29],s153[29],s154[29],s155[29],s156[29],s157[29],s158[29],s159[29],s160[29],s161[29],s162[29],s163[29],s164[29],s165[29],s166[29],s167[29],s167[30],s167[31],s167[32],s167[33],s167[34],s167[35],s167[36],s167[37],s167[38],s167[39],s167[40],s167[41],s167[42],s167[43],s167[44],s167[45],s209[100],s209[101],s209[102],s209[103],s209[104],s209[105],s209[106],s209[107],s209[108],s209[109],s209[110],s209[111],s209[112],s209[113],s209[114],s209[115],s209[116],s209[117],s209[118],s209[119],s209[120],s209[121],s209[122],s209[123],s209[124],s209[125],s209[126],s209[127],s209[128],s209[129],s209[130],s209[131],s209[132],s209[133],s209[134],s209[135],s209[136],s209[137],s209[138],s209[139],s209[140],s209[141],s209[142],s209[143],s209[144],s209[145],s209[146],s209[147],s209[148],s209[149],s209[150],s209[151],s209[152],s209[153],s209[154],s209[155],s209[156],s209[157],s209[158],s209[159],s209[160],s209[161],s209[162],s209[163],s209[164],s209[165],s209[166],s209[167],s209[168],s209[169],s209[170],s209[171],s209[172],s209[173],s209[174],s209[175],s209[176],s209[177],s209[178],s209[179],s209[180],s209[181],s209[182],s209[183],s209[184],s209[185],s209[186],s209[187],s209[188],s209[189],s209[190],s209[191],s209[192],s209[193],s209[194],s209[195],s209[196],s209[197],s209[198],s209[199],s209[200],s209[201],s209[202],s209[203],s209[204],s209[205],s209[206],s209[207],s209[208],s209[209],s209[210],s209[211],s209[212],s209[213],s209[214],s209[215],s209[216],s209[217],s209[218],s209[219],s209[220],s209[221],s209[222],s209[223],s209[224],s209[225],s209[226],s209[227],s209[228],s209[229],s209[230],s209[231],s209[232],s209[233],s209[234],s209[235],s209[236],s209[237],s209[238],s209[239],s209[240],s209[241],s209[242],s209[243],s209[244],s209[245],s209[246],s209[247],s209[248],s209[249],s209[250],s209[251],s209[252],s209[253],s209[254],s209[255],s209[256],s209[257],s209[258],s209[259],s209[260],s209[261],s209[262],s209[263],s209[264],s209[265],s209[266],s209[267],s209[268],s209[269],s209[270],s209[271],s209[272],s209[273],s209[274],s209[275],s209[276],s209[277],s209[278],s209[279],s209[280],s209[281],s209[282],s209[283],s209[284],s209[285],s209[286],s209[287],s209[288],s209[289],s209[290],s209[291],s208[293],s207[295],s206[297],s205[299],s204[301],s203[303],s202[305],s201[307],s200[309],s199[311],s198[313],s197[315],s196[317],s195[319],s194[321],s193[323],s192[229],s191[231],s190[233],s189[235],s188[237],s187[239],s186[241],s185[243],s184[245],s183[247],s182[249],s181[251],s180[253],s179[255],s178[257],s177[259],s176[261],s175[263],s174[265],s173[267],s172[269],s171[271],s170[273],s169[275],s168[277],s167[279],s166[281],s165[283],s164[285],s163[287],s162[289],s161[291],s160[293],s159[295],s158[297],s157[299],s156[301],s155[303],s154[305],s153[307],s152[309],s151[311],s150[313],s149[315],s148[317],s147[319],s146[321],s145[323],s144[325],s143[327],s142[329],s141[331],s140[333],s139[335],s138[337],s137[339],s136[341],s135[343],s134[345],s133[347],s132[349],s131[351],s130[353],s129[355],pp255[165],pp254[167],pp253[169],pp252[171],pp251[173],pp250[175],pp249[177],pp248[179],pp247[181],pp246[183],pp245[185],pp244[187],pp243[189],pp242[191],pp241[193],pp240[195],pp239[197],pp238[199],pp237[201],pp236[203],pp235[205],pp234[207],pp233[209],pp232[211],pp231[213],pp230[215],pp229[217],pp228[219],pp227[221],pp228[221],pp229[221],pp230[221],pp231[221],pp232[221],pp233[221],pp234[221],pp235[221],pp236[221],pp237[221],pp238[221],pp239[221],pp240[221],pp241[221]};
    assign in210_2 = {s198[12],s197[14],s196[16],s195[18],s194[20],s193[22],pp45[10],pp45[11],pp45[12],pp45[13],pp45[14],pp45[15],pp45[16],pp45[17],pp45[18],pp47[17],pp49[16],pp51[15],pp53[14],pp55[13],pp57[12],pp59[11],pp61[10],s193[40],s194[40],s194[41],s194[42],s194[43],s194[44],s194[45],s194[46],s194[47],s194[48],s194[49],s194[50],s194[51],s194[52],s194[53],s194[54],s194[55],s194[56],s194[57],s194[58],s194[59],s194[60],s194[61],s194[62],s194[63],s194[64],s194[65],s194[66],s155[10],s154[12],s153[14],s152[16],s151[18],s150[20],s149[22],s148[24],s147[26],s146[28],s147[28],s148[28],s149[28],s150[28],s151[28],s152[28],s153[28],s154[28],s155[28],s156[28],s157[28],s158[28],s159[28],s160[28],s161[28],s162[28],s163[28],s164[28],s165[28],s166[28],s167[28],s168[28],s168[29],s168[30],s168[31],s168[32],s168[33],s168[34],s168[35],s168[36],s168[37],s168[38],s168[39],s168[40],s168[41],s168[42],s168[43],s168[44],s168[45],s169[45],s170[45],s171[45],s172[45],s173[45],s174[45],s175[45],s176[45],s177[45],s178[45],s179[45],s180[45],s181[45],s182[45],s183[45],s184[45],s185[45],s186[45],s187[45],s188[45],s189[45],s190[45],s191[45],s192[45],s10[36],s11[36],s12[36],s13[36],s14[36],s15[36],s16[36],s17[36],s18[36],s19[36],s20[36],s21[36],s22[36],s23[36],s24[36],s25[36],s26[36],s27[36],s28[36],s29[36],s30[36],s31[36],s32[36],s33[36],s34[36],s35[36],s36[36],s37[36],s38[36],s39[36],s40[36],s41[36],s42[36],s43[36],s44[36],s45[36],s46[36],s47[36],s48[36],s49[36],s50[36],s51[36],s52[36],s53[36],s54[36],s55[36],s56[36],s57[36],s58[36],s59[36],s60[36],s61[36],s62[36],s63[36],s64[36],s64[37],s64[38],s64[39],s64[40],s64[41],s64[42],s64[43],s64[44],s64[45],s64[46],s64[47],s64[48],s64[49],s64[50],s64[51],s64[52],s64[53],s64[54],s64[55],s64[56],s64[57],s64[58],s64[59],s64[60],s64[61],s64[62],s64[63],s64[64],s64[65],s62[68],s60[71],s58[74],s56[77],s55[79],s55[80],s55[81],s55[82],s55[83],s55[84],s55[85],s55[86],s55[87],s55[88],s55[89],s55[90],s55[91],s55[92],s55[93],s55[94],s55[95],s55[96],s55[97],s55[98],s55[99],s9[146],s8[148],s7[150],s6[152],s4[155],s2[158],s61[100],s60[102],s59[104],s58[106],s57[108],s56[110],s55[112],s54[114],s53[116],s52[118],s51[120],s50[122],s49[124],s48[126],s47[128],s46[130],s45[132],s44[134],s43[136],s42[138],s41[140],s40[142],s39[144],s38[146],s37[148],s36[150],s35[152],s34[154],s33[156],s32[158],s31[160],s30[162],s29[164],s28[166],s27[168],s26[170],s25[172],s24[174],s23[176],s22[178],s21[180],s20[182],s19[184],s18[186],s17[188],s16[190],s15[192],s14[194],s13[196],s12[198],s11[200],s10[202],s209[292],s208[294],s207[296],s206[298],s205[300],s204[302],s203[304],s202[306],s201[308],s200[310],s199[312],s198[314],s197[316],s196[318],s195[320],s194[322],s193[324],s192[230],s191[232],s190[234],s189[236],s188[238],s187[240],s186[242],s185[244],s184[246],s183[248],s182[250],s181[252],s180[254],s179[256],s178[258],s177[260],s176[262],s175[264],s174[266],s173[268],s172[270],s171[272],s170[274],s169[276],s168[278],s167[280],s166[282],s165[284],s164[286],s163[288],s162[290],s161[292],s160[294],s159[296],s158[298],s157[300],s156[302],s155[304],s154[306],s153[308],s152[310],s151[312],s150[314],s149[316],s148[318],s147[320],s146[322],s145[324],s144[326],s143[328],s142[330],s141[332],s140[334],s139[336],s138[338],s137[340],s136[342],s135[344],s134[346],s133[348],s132[350],s131[352],s130[354],s129[356],pp255[166],pp254[168],pp253[170],pp252[172],pp251[174],pp250[176],pp249[178],pp248[180],pp247[182],pp246[184],pp245[186],pp244[188],pp243[190],pp242[192],pp241[194],pp240[196],pp239[198],pp238[200],pp237[202],pp236[204],pp235[206],pp234[208],pp233[210],pp232[212],pp231[214],pp230[216],pp229[218],pp228[220],pp229[220],pp230[220],pp231[220],pp232[220],pp233[220],pp234[220],pp235[220],pp236[220],pp237[220],pp238[220],pp239[220],pp240[220],pp241[220],pp242[220]};
    CLA_414 KS_210(s210, c210, in210_1, in210_2);
    wire[411:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {s198[13],s197[15],s196[17],s195[19],s194[21],s193[23],pp46[10],pp46[11],pp46[12],pp46[13],pp46[14],pp46[15],pp46[16],pp46[17],pp48[16],pp50[15],pp52[14],pp54[13],pp56[12],pp58[11],pp60[10],s193[39],s194[39],s195[39],s195[40],s195[41],s195[42],s195[43],s195[44],s195[45],s195[46],s195[47],s195[48],s195[49],s195[50],s195[51],s195[52],s195[53],s195[54],s195[55],s195[56],s195[57],s195[58],s195[59],s195[60],s195[61],s195[62],s195[63],s195[64],s195[65],s193[68],s155[11],s154[13],s153[15],s152[17],s151[19],s150[21],s149[23],s148[25],s147[27],s148[27],s149[27],s150[27],s151[27],s152[27],s153[27],s154[27],s155[27],s156[27],s157[27],s158[27],s159[27],s160[27],s161[27],s162[27],s163[27],s164[27],s165[27],s166[27],s167[27],s168[27],s169[27],s169[28],s169[29],s169[30],s169[31],s169[32],s169[33],s169[34],s169[35],s169[36],s169[37],s169[38],s169[39],s169[40],s169[41],s169[42],s169[43],s169[44],s210[100],s210[101],s210[102],s210[103],s210[104],s210[105],s210[106],s210[107],s210[108],s210[109],s210[110],s210[111],s210[112],s210[113],s210[114],s210[115],s210[116],s210[117],s210[118],s210[119],s210[120],s210[121],s210[122],s210[123],s210[124],s210[125],s210[126],s210[127],s210[128],s210[129],s210[130],s210[131],s210[132],s210[133],s210[134],s210[135],s210[136],s210[137],s210[138],s210[139],s210[140],s210[141],s210[142],s210[143],s210[144],s210[145],s210[146],s210[147],s210[148],s210[149],s210[150],s210[151],s210[152],s210[153],s210[154],s210[155],s210[156],s210[157],s210[158],s210[159],s210[160],s210[161],s210[162],s210[163],s210[164],s210[165],s210[166],s210[167],s210[168],s210[169],s210[170],s210[171],s210[172],s210[173],s210[174],s210[175],s210[176],s210[177],s210[178],s210[179],s210[180],s210[181],s210[182],s210[183],s210[184],s210[185],s210[186],s210[187],s210[188],s210[189],s210[190],s210[191],s210[192],s210[193],s210[194],s210[195],s210[196],s210[197],s210[198],s210[199],s210[200],s210[201],s210[202],s210[203],s210[204],s210[205],s210[206],s210[207],s210[208],s210[209],s210[210],s210[211],s210[212],s210[213],s210[214],s210[215],s210[216],s210[217],s210[218],s210[219],s210[220],s210[221],s210[222],s210[223],s210[224],s210[225],s210[226],s210[227],s210[228],s210[229],s210[230],s210[231],s210[232],s210[233],s210[234],s210[235],s210[236],s210[237],s210[238],s210[239],s210[240],s210[241],s210[242],s210[243],s210[244],s210[245],s210[246],s210[247],s210[248],s210[249],s210[250],s210[251],s210[252],s210[253],s210[254],s210[255],s210[256],s210[257],s210[258],s210[259],s210[260],s210[261],s210[262],s210[263],s210[264],s210[265],s210[266],s210[267],s210[268],s210[269],s210[270],s210[271],s210[272],s210[273],s210[274],s210[275],s210[276],s210[277],s210[278],s210[279],s210[280],s210[281],s210[282],s210[283],s210[284],s210[285],s210[286],s210[287],s210[288],s210[289],s210[290],s210[291],s209[293],s208[295],s207[297],s206[299],s205[301],s204[303],s203[305],s202[307],s201[309],s200[311],s199[313],s198[315],s197[317],s196[319],s195[321],s194[323],s193[325],s192[231],s191[233],s190[235],s189[237],s188[239],s187[241],s186[243],s185[245],s184[247],s183[249],s182[251],s181[253],s180[255],s179[257],s178[259],s177[261],s176[263],s175[265],s174[267],s173[269],s172[271],s171[273],s170[275],s169[277],s168[279],s167[281],s166[283],s165[285],s164[287],s163[289],s162[291],s161[293],s160[295],s159[297],s158[299],s157[301],s156[303],s155[305],s154[307],s153[309],s152[311],s151[313],s150[315],s149[317],s148[319],s147[321],s146[323],s145[325],s144[327],s143[329],s142[331],s141[333],s140[335],s139[337],s138[339],s137[341],s136[343],s135[345],s134[347],s133[349],s132[351],s131[353],s130[355],s129[357],pp255[167],pp254[169],pp253[171],pp252[173],pp251[175],pp250[177],pp249[179],pp248[181],pp247[183],pp246[185],pp245[187],pp244[189],pp243[191],pp242[193],pp241[195],pp240[197],pp239[199],pp238[201],pp237[203],pp236[205],pp235[207],pp234[209],pp233[211],pp232[213],pp231[215],pp230[217],pp229[219],pp230[219],pp231[219],pp232[219],pp233[219],pp234[219],pp235[219],pp236[219],pp237[219],pp238[219],pp239[219],pp240[219],pp241[219],pp242[219]};
    assign in211_2 = {s199[12],s198[14],s197[16],s196[18],s195[20],s194[22],s193[24],pp47[10],pp47[11],pp47[12],pp47[13],pp47[14],pp47[15],pp47[16],pp49[15],pp51[14],pp53[13],pp55[12],pp57[11],pp59[10],s193[38],s194[38],s195[38],s196[38],s196[39],s196[40],s196[41],s196[42],s196[43],s196[44],s196[45],s196[46],s196[47],s196[48],s196[49],s196[50],s196[51],s196[52],s196[53],s196[54],s196[55],s196[56],s196[57],s196[58],s196[59],s196[60],s196[61],s196[62],s196[63],s196[64],s194[67],s156[10],s155[12],s154[14],s153[16],s152[18],s151[20],s150[22],s149[24],s148[26],s149[26],s150[26],s151[26],s152[26],s153[26],s154[26],s155[26],s156[26],s157[26],s158[26],s159[26],s160[26],s161[26],s162[26],s163[26],s164[26],s165[26],s166[26],s167[26],s168[26],s169[26],s170[26],s170[27],s170[28],s170[29],s170[30],s170[31],s170[32],s170[33],s170[34],s170[35],s170[36],s170[37],s170[38],s170[39],s170[40],s170[41],s170[42],s170[43],s170[44],s171[44],s172[44],s173[44],s174[44],s175[44],s176[44],s177[44],s178[44],s179[44],s180[44],s181[44],s182[44],s183[44],s184[44],s185[44],s186[44],s187[44],s188[44],s189[44],s190[44],s191[44],s192[44],s10[35],s11[35],s12[35],s13[35],s14[35],s15[35],s16[35],s17[35],s18[35],s19[35],s20[35],s21[35],s22[35],s23[35],s24[35],s25[35],s26[35],s27[35],s28[35],s29[35],s30[35],s31[35],s32[35],s33[35],s34[35],s35[35],s36[35],s37[35],s38[35],s39[35],s40[35],s41[35],s42[35],s43[35],s44[35],s45[35],s46[35],s47[35],s48[35],s49[35],s50[35],s51[35],s52[35],s53[35],s54[35],s55[35],s56[35],s57[35],s58[35],s59[35],s60[35],s61[35],s62[35],s63[35],s64[35],s65[35],s65[36],s65[37],s65[38],s65[39],s65[40],s65[41],s65[42],s65[43],s65[44],s65[45],s65[46],s65[47],s65[48],s65[49],s65[50],s65[51],s65[52],s65[53],s65[54],s65[55],s65[56],s65[57],s65[58],s65[59],s65[60],s65[61],s65[62],s65[63],s65[64],s63[67],s61[70],s59[73],s57[76],s56[78],s56[79],s56[80],s56[81],s56[82],s56[83],s56[84],s56[85],s56[86],s56[87],s56[88],s56[89],s56[90],s56[91],s56[92],s56[93],s56[94],s56[95],s56[96],s56[97],s56[98],s56[99],s9[147],s8[149],s7[151],s5[154],s3[157],s1[160],s61[101],s60[103],s59[105],s58[107],s57[109],s56[111],s55[113],s54[115],s53[117],s52[119],s51[121],s50[123],s49[125],s48[127],s47[129],s46[131],s45[133],s44[135],s43[137],s42[139],s41[141],s40[143],s39[145],s38[147],s37[149],s36[151],s35[153],s34[155],s33[157],s32[159],s31[161],s30[163],s29[165],s28[167],s27[169],s26[171],s25[173],s24[175],s23[177],s22[179],s21[181],s20[183],s19[185],s18[187],s17[189],s16[191],s15[193],s14[195],s13[197],s12[199],s11[201],s10[203],s210[292],s209[294],s208[296],s207[298],s206[300],s205[302],s204[304],s203[306],s202[308],s201[310],s200[312],s199[314],s198[316],s197[318],s196[320],s195[322],s194[324],s193[326],s192[232],s191[234],s190[236],s189[238],s188[240],s187[242],s186[244],s185[246],s184[248],s183[250],s182[252],s181[254],s180[256],s179[258],s178[260],s177[262],s176[264],s175[266],s174[268],s173[270],s172[272],s171[274],s170[276],s169[278],s168[280],s167[282],s166[284],s165[286],s164[288],s163[290],s162[292],s161[294],s160[296],s159[298],s158[300],s157[302],s156[304],s155[306],s154[308],s153[310],s152[312],s151[314],s150[316],s149[318],s148[320],s147[322],s146[324],s145[326],s144[328],s143[330],s142[332],s141[334],s140[336],s139[338],s138[340],s137[342],s136[344],s135[346],s134[348],s133[350],s132[352],s131[354],s130[356],s129[358],pp255[168],pp254[170],pp253[172],pp252[174],pp251[176],pp250[178],pp249[180],pp248[182],pp247[184],pp246[186],pp245[188],pp244[190],pp243[192],pp242[194],pp241[196],pp240[198],pp239[200],pp238[202],pp237[204],pp236[206],pp235[208],pp234[210],pp233[212],pp232[214],pp231[216],pp230[218],pp231[218],pp232[218],pp233[218],pp234[218],pp235[218],pp236[218],pp237[218],pp238[218],pp239[218],pp240[218],pp241[218],pp242[218],pp243[218]};
    CLA_412 KS_211(s211, c211, in211_1, in211_2);
    wire[409:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {s199[13],s198[15],s197[17],s196[19],s195[21],s194[23],s193[25],pp48[10],pp48[11],pp48[12],pp48[13],pp48[14],pp48[15],pp50[14],pp52[13],pp54[12],pp56[11],pp58[10],s193[37],s194[37],s195[37],s196[37],s197[37],s197[38],s197[39],s197[40],s197[41],s197[42],s197[43],s197[44],s197[45],s197[46],s197[47],s197[48],s197[49],s197[50],s197[51],s197[52],s197[53],s197[54],s197[55],s197[56],s197[57],s197[58],s197[59],s197[60],s197[61],s197[62],s197[63],s195[66],s193[69],s156[11],s155[13],s154[15],s153[17],s152[19],s151[21],s150[23],s149[25],s150[25],s151[25],s152[25],s153[25],s154[25],s155[25],s156[25],s157[25],s158[25],s159[25],s160[25],s161[25],s162[25],s163[25],s164[25],s165[25],s166[25],s167[25],s168[25],s169[25],s170[25],s171[25],s171[26],s171[27],s171[28],s171[29],s171[30],s171[31],s171[32],s171[33],s171[34],s171[35],s171[36],s171[37],s171[38],s171[39],s171[40],s171[41],s171[42],s171[43],s211[100],s211[101],s211[102],s211[103],s211[104],s211[105],s211[106],s211[107],s211[108],s211[109],s211[110],s211[111],s211[112],s211[113],s211[114],s211[115],s211[116],s211[117],s211[118],s211[119],s211[120],s211[121],s211[122],s211[123],s211[124],s211[125],s211[126],s211[127],s211[128],s211[129],s211[130],s211[131],s211[132],s211[133],s211[134],s211[135],s211[136],s211[137],s211[138],s211[139],s211[140],s211[141],s211[142],s211[143],s211[144],s211[145],s211[146],s211[147],s211[148],s211[149],s211[150],s211[151],s211[152],s211[153],s211[154],s211[155],s211[156],s211[157],s211[158],s211[159],s211[160],s211[161],s211[162],s211[163],s211[164],s211[165],s211[166],s211[167],s211[168],s211[169],s211[170],s211[171],s211[172],s211[173],s211[174],s211[175],s211[176],s211[177],s211[178],s211[179],s211[180],s211[181],s211[182],s211[183],s211[184],s211[185],s211[186],s211[187],s211[188],s211[189],s211[190],s211[191],s211[192],s211[193],s211[194],s211[195],s211[196],s211[197],s211[198],s211[199],s211[200],s211[201],s211[202],s211[203],s211[204],s211[205],s211[206],s211[207],s211[208],s211[209],s211[210],s211[211],s211[212],s211[213],s211[214],s211[215],s211[216],s211[217],s211[218],s211[219],s211[220],s211[221],s211[222],s211[223],s211[224],s211[225],s211[226],s211[227],s211[228],s211[229],s211[230],s211[231],s211[232],s211[233],s211[234],s211[235],s211[236],s211[237],s211[238],s211[239],s211[240],s211[241],s211[242],s211[243],s211[244],s211[245],s211[246],s211[247],s211[248],s211[249],s211[250],s211[251],s211[252],s211[253],s211[254],s211[255],s211[256],s211[257],s211[258],s211[259],s211[260],s211[261],s211[262],s211[263],s211[264],s211[265],s211[266],s211[267],s211[268],s211[269],s211[270],s211[271],s211[272],s211[273],s211[274],s211[275],s211[276],s211[277],s211[278],s211[279],s211[280],s211[281],s211[282],s211[283],s211[284],s211[285],s211[286],s211[287],s211[288],s211[289],s211[290],s211[291],s210[293],s209[295],s208[297],s207[299],s206[301],s205[303],s204[305],s203[307],s202[309],s201[311],s200[313],s199[315],s198[317],s197[319],s196[321],s195[323],s194[325],s193[327],s192[233],s191[235],s190[237],s189[239],s188[241],s187[243],s186[245],s185[247],s184[249],s183[251],s182[253],s181[255],s180[257],s179[259],s178[261],s177[263],s176[265],s175[267],s174[269],s173[271],s172[273],s171[275],s170[277],s169[279],s168[281],s167[283],s166[285],s165[287],s164[289],s163[291],s162[293],s161[295],s160[297],s159[299],s158[301],s157[303],s156[305],s155[307],s154[309],s153[311],s152[313],s151[315],s150[317],s149[319],s148[321],s147[323],s146[325],s145[327],s144[329],s143[331],s142[333],s141[335],s140[337],s139[339],s138[341],s137[343],s136[345],s135[347],s134[349],s133[351],s132[353],s131[355],s130[357],s129[359],pp255[169],pp254[171],pp253[173],pp252[175],pp251[177],pp250[179],pp249[181],pp248[183],pp247[185],pp246[187],pp245[189],pp244[191],pp243[193],pp242[195],pp241[197],pp240[199],pp239[201],pp238[203],pp237[205],pp236[207],pp235[209],pp234[211],pp233[213],pp232[215],pp231[217],pp232[217],pp233[217],pp234[217],pp235[217],pp236[217],pp237[217],pp238[217],pp239[217],pp240[217],pp241[217],pp242[217],pp243[217]};
    assign in212_2 = {s200[12],s199[14],s198[16],s197[18],s196[20],s195[22],s194[24],s193[26],pp49[10],pp49[11],pp49[12],pp49[13],pp49[14],pp51[13],pp53[12],pp55[11],pp57[10],s193[36],s194[36],s195[36],s196[36],s197[36],s198[36],s198[37],s198[38],s198[39],s198[40],s198[41],s198[42],s198[43],s198[44],s198[45],s198[46],s198[47],s198[48],s198[49],s198[50],s198[51],s198[52],s198[53],s198[54],s198[55],s198[56],s198[57],s198[58],s198[59],s198[60],s198[61],s198[62],s196[65],s194[68],s157[10],s156[12],s155[14],s154[16],s153[18],s152[20],s151[22],s150[24],s151[24],s152[24],s153[24],s154[24],s155[24],s156[24],s157[24],s158[24],s159[24],s160[24],s161[24],s162[24],s163[24],s164[24],s165[24],s166[24],s167[24],s168[24],s169[24],s170[24],s171[24],s172[24],s172[25],s172[26],s172[27],s172[28],s172[29],s172[30],s172[31],s172[32],s172[33],s172[34],s172[35],s172[36],s172[37],s172[38],s172[39],s172[40],s172[41],s172[42],s172[43],s173[43],s174[43],s175[43],s176[43],s177[43],s178[43],s179[43],s180[43],s181[43],s182[43],s183[43],s184[43],s185[43],s186[43],s187[43],s188[43],s189[43],s190[43],s191[43],s192[43],s10[34],s11[34],s12[34],s13[34],s14[34],s15[34],s16[34],s17[34],s18[34],s19[34],s20[34],s21[34],s22[34],s23[34],s24[34],s25[34],s26[34],s27[34],s28[34],s29[34],s30[34],s31[34],s32[34],s33[34],s34[34],s35[34],s36[34],s37[34],s38[34],s39[34],s40[34],s41[34],s42[34],s43[34],s44[34],s45[34],s46[34],s47[34],s48[34],s49[34],s50[34],s51[34],s52[34],s53[34],s54[34],s55[34],s56[34],s57[34],s58[34],s59[34],s60[34],s61[34],s62[34],s63[34],s64[34],s65[34],s66[34],s66[35],s66[36],s66[37],s66[38],s66[39],s66[40],s66[41],s66[42],s66[43],s66[44],s66[45],s66[46],s66[47],s66[48],s66[49],s66[50],s66[51],s66[52],s66[53],s66[54],s66[55],s66[56],s66[57],s66[58],s66[59],s66[60],s66[61],s66[62],s66[63],s64[66],s62[69],s60[72],s58[75],s57[77],s57[78],s57[79],s57[80],s57[81],s57[82],s57[83],s57[84],s57[85],s57[86],s57[87],s57[88],s57[89],s57[90],s57[91],s57[92],s57[93],s57[94],s57[95],s57[96],s57[97],s57[98],s57[99],s9[148],s8[150],s6[153],s4[156],s2[159],s62[100],s61[102],s60[104],s59[106],s58[108],s57[110],s56[112],s55[114],s54[116],s53[118],s52[120],s51[122],s50[124],s49[126],s48[128],s47[130],s46[132],s45[134],s44[136],s43[138],s42[140],s41[142],s40[144],s39[146],s38[148],s37[150],s36[152],s35[154],s34[156],s33[158],s32[160],s31[162],s30[164],s29[166],s28[168],s27[170],s26[172],s25[174],s24[176],s23[178],s22[180],s21[182],s20[184],s19[186],s18[188],s17[190],s16[192],s15[194],s14[196],s13[198],s12[200],s11[202],s10[204],s211[292],s210[294],s209[296],s208[298],s207[300],s206[302],s205[304],s204[306],s203[308],s202[310],s201[312],s200[314],s199[316],s198[318],s197[320],s196[322],s195[324],s194[326],s193[328],s192[234],s191[236],s190[238],s189[240],s188[242],s187[244],s186[246],s185[248],s184[250],s183[252],s182[254],s181[256],s180[258],s179[260],s178[262],s177[264],s176[266],s175[268],s174[270],s173[272],s172[274],s171[276],s170[278],s169[280],s168[282],s167[284],s166[286],s165[288],s164[290],s163[292],s162[294],s161[296],s160[298],s159[300],s158[302],s157[304],s156[306],s155[308],s154[310],s153[312],s152[314],s151[316],s150[318],s149[320],s148[322],s147[324],s146[326],s145[328],s144[330],s143[332],s142[334],s141[336],s140[338],s139[340],s138[342],s137[344],s136[346],s135[348],s134[350],s133[352],s132[354],s131[356],s130[358],s129[360],pp255[170],pp254[172],pp253[174],pp252[176],pp251[178],pp250[180],pp249[182],pp248[184],pp247[186],pp246[188],pp245[190],pp244[192],pp243[194],pp242[196],pp241[198],pp240[200],pp239[202],pp238[204],pp237[206],pp236[208],pp235[210],pp234[212],pp233[214],pp232[216],pp233[216],pp234[216],pp235[216],pp236[216],pp237[216],pp238[216],pp239[216],pp240[216],pp241[216],pp242[216],pp243[216],pp244[216]};
    CLA_410 KS_212(s212, c212, in212_1, in212_2);
    wire[407:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {s200[13],s199[15],s198[17],s197[19],s196[21],s195[23],s194[25],s193[27],pp50[10],pp50[11],pp50[12],pp50[13],pp52[12],pp54[11],pp56[10],s193[35],s194[35],s195[35],s196[35],s197[35],s198[35],s199[35],s199[36],s199[37],s199[38],s199[39],s199[40],s199[41],s199[42],s199[43],s199[44],s199[45],s199[46],s199[47],s199[48],s199[49],s199[50],s199[51],s199[52],s199[53],s199[54],s199[55],s199[56],s199[57],s199[58],s199[59],s199[60],s199[61],s197[64],s195[67],s193[70],s157[11],s156[13],s155[15],s154[17],s153[19],s152[21],s151[23],s152[23],s153[23],s154[23],s155[23],s156[23],s157[23],s158[23],s159[23],s160[23],s161[23],s162[23],s163[23],s164[23],s165[23],s166[23],s167[23],s168[23],s169[23],s170[23],s171[23],s172[23],s173[23],s173[24],s173[25],s173[26],s173[27],s173[28],s173[29],s173[30],s173[31],s173[32],s173[33],s173[34],s173[35],s173[36],s173[37],s173[38],s173[39],s173[40],s173[41],s173[42],s212[100],s212[101],s212[102],s212[103],s212[104],s212[105],s212[106],s212[107],s212[108],s212[109],s212[110],s212[111],s212[112],s212[113],s212[114],s212[115],s212[116],s212[117],s212[118],s212[119],s212[120],s212[121],s212[122],s212[123],s212[124],s212[125],s212[126],s212[127],s212[128],s212[129],s212[130],s212[131],s212[132],s212[133],s212[134],s212[135],s212[136],s212[137],s212[138],s212[139],s212[140],s212[141],s212[142],s212[143],s212[144],s212[145],s212[146],s212[147],s212[148],s212[149],s212[150],s212[151],s212[152],s212[153],s212[154],s212[155],s212[156],s212[157],s212[158],s212[159],s212[160],s212[161],s212[162],s212[163],s212[164],s212[165],s212[166],s212[167],s212[168],s212[169],s212[170],s212[171],s212[172],s212[173],s212[174],s212[175],s212[176],s212[177],s212[178],s212[179],s212[180],s212[181],s212[182],s212[183],s212[184],s212[185],s212[186],s212[187],s212[188],s212[189],s212[190],s212[191],s212[192],s212[193],s212[194],s212[195],s212[196],s212[197],s212[198],s212[199],s212[200],s212[201],s212[202],s212[203],s212[204],s212[205],s212[206],s212[207],s212[208],s212[209],s212[210],s212[211],s212[212],s212[213],s212[214],s212[215],s212[216],s212[217],s212[218],s212[219],s212[220],s212[221],s212[222],s212[223],s212[224],s212[225],s212[226],s212[227],s212[228],s212[229],s212[230],s212[231],s212[232],s212[233],s212[234],s212[235],s212[236],s212[237],s212[238],s212[239],s212[240],s212[241],s212[242],s212[243],s212[244],s212[245],s212[246],s212[247],s212[248],s212[249],s212[250],s212[251],s212[252],s212[253],s212[254],s212[255],s212[256],s212[257],s212[258],s212[259],s212[260],s212[261],s212[262],s212[263],s212[264],s212[265],s212[266],s212[267],s212[268],s212[269],s212[270],s212[271],s212[272],s212[273],s212[274],s212[275],s212[276],s212[277],s212[278],s212[279],s212[280],s212[281],s212[282],s212[283],s212[284],s212[285],s212[286],s212[287],s212[288],s212[289],s212[290],s212[291],s211[293],s210[295],s209[297],s208[299],s207[301],s206[303],s205[305],s204[307],s203[309],s202[311],s201[313],s200[315],s199[317],s198[319],s197[321],s196[323],s195[325],s194[327],s193[329],s192[235],s191[237],s190[239],s189[241],s188[243],s187[245],s186[247],s185[249],s184[251],s183[253],s182[255],s181[257],s180[259],s179[261],s178[263],s177[265],s176[267],s175[269],s174[271],s173[273],s172[275],s171[277],s170[279],s169[281],s168[283],s167[285],s166[287],s165[289],s164[291],s163[293],s162[295],s161[297],s160[299],s159[301],s158[303],s157[305],s156[307],s155[309],s154[311],s153[313],s152[315],s151[317],s150[319],s149[321],s148[323],s147[325],s146[327],s145[329],s144[331],s143[333],s142[335],s141[337],s140[339],s139[341],s138[343],s137[345],s136[347],s135[349],s134[351],s133[353],s132[355],s131[357],s130[359],s129[361],pp255[171],pp254[173],pp253[175],pp252[177],pp251[179],pp250[181],pp249[183],pp248[185],pp247[187],pp246[189],pp245[191],pp244[193],pp243[195],pp242[197],pp241[199],pp240[201],pp239[203],pp238[205],pp237[207],pp236[209],pp235[211],pp234[213],pp233[215],pp234[215],pp235[215],pp236[215],pp237[215],pp238[215],pp239[215],pp240[215],pp241[215],pp242[215],pp243[215],pp244[215]};
    assign in213_2 = {s201[12],s200[14],s199[16],s198[18],s197[20],s196[22],s195[24],s194[26],s193[28],pp51[10],pp51[11],pp51[12],pp53[11],pp55[10],s193[34],s194[34],s195[34],s196[34],s197[34],s198[34],s199[34],s200[34],s200[35],s200[36],s200[37],s200[38],s200[39],s200[40],s200[41],s200[42],s200[43],s200[44],s200[45],s200[46],s200[47],s200[48],s200[49],s200[50],s200[51],s200[52],s200[53],s200[54],s200[55],s200[56],s200[57],s200[58],s200[59],s200[60],s198[63],s196[66],s194[69],s158[10],s157[12],s156[14],s155[16],s154[18],s153[20],s152[22],s153[22],s154[22],s155[22],s156[22],s157[22],s158[22],s159[22],s160[22],s161[22],s162[22],s163[22],s164[22],s165[22],s166[22],s167[22],s168[22],s169[22],s170[22],s171[22],s172[22],s173[22],s174[22],s174[23],s174[24],s174[25],s174[26],s174[27],s174[28],s174[29],s174[30],s174[31],s174[32],s174[33],s174[34],s174[35],s174[36],s174[37],s174[38],s174[39],s174[40],s174[41],s174[42],s175[42],s176[42],s177[42],s178[42],s179[42],s180[42],s181[42],s182[42],s183[42],s184[42],s185[42],s186[42],s187[42],s188[42],s189[42],s190[42],s191[42],s192[42],s10[33],s11[33],s12[33],s13[33],s14[33],s15[33],s16[33],s17[33],s18[33],s19[33],s20[33],s21[33],s22[33],s23[33],s24[33],s25[33],s26[33],s27[33],s28[33],s29[33],s30[33],s31[33],s32[33],s33[33],s34[33],s35[33],s36[33],s37[33],s38[33],s39[33],s40[33],s41[33],s42[33],s43[33],s44[33],s45[33],s46[33],s47[33],s48[33],s49[33],s50[33],s51[33],s52[33],s53[33],s54[33],s55[33],s56[33],s57[33],s58[33],s59[33],s60[33],s61[33],s62[33],s63[33],s64[33],s65[33],s66[33],s67[33],s67[34],s67[35],s67[36],s67[37],s67[38],s67[39],s67[40],s67[41],s67[42],s67[43],s67[44],s67[45],s67[46],s67[47],s67[48],s67[49],s67[50],s67[51],s67[52],s67[53],s67[54],s67[55],s67[56],s67[57],s67[58],s67[59],s67[60],s67[61],s67[62],s65[65],s63[68],s61[71],s59[74],s58[76],s58[77],s58[78],s58[79],s58[80],s58[81],s58[82],s58[83],s58[84],s58[85],s58[86],s58[87],s58[88],s58[89],s58[90],s58[91],s58[92],s58[93],s58[94],s58[95],s58[96],s58[97],s58[98],s58[99],s9[149],s7[152],s5[155],s3[158],s1[161],s62[101],s61[103],s60[105],s59[107],s58[109],s57[111],s56[113],s55[115],s54[117],s53[119],s52[121],s51[123],s50[125],s49[127],s48[129],s47[131],s46[133],s45[135],s44[137],s43[139],s42[141],s41[143],s40[145],s39[147],s38[149],s37[151],s36[153],s35[155],s34[157],s33[159],s32[161],s31[163],s30[165],s29[167],s28[169],s27[171],s26[173],s25[175],s24[177],s23[179],s22[181],s21[183],s20[185],s19[187],s18[189],s17[191],s16[193],s15[195],s14[197],s13[199],s12[201],s11[203],s10[205],s212[292],s211[294],s210[296],s209[298],s208[300],s207[302],s206[304],s205[306],s204[308],s203[310],s202[312],s201[314],s200[316],s199[318],s198[320],s197[322],s196[324],s195[326],s194[328],s193[330],s192[236],s191[238],s190[240],s189[242],s188[244],s187[246],s186[248],s185[250],s184[252],s183[254],s182[256],s181[258],s180[260],s179[262],s178[264],s177[266],s176[268],s175[270],s174[272],s173[274],s172[276],s171[278],s170[280],s169[282],s168[284],s167[286],s166[288],s165[290],s164[292],s163[294],s162[296],s161[298],s160[300],s159[302],s158[304],s157[306],s156[308],s155[310],s154[312],s153[314],s152[316],s151[318],s150[320],s149[322],s148[324],s147[326],s146[328],s145[330],s144[332],s143[334],s142[336],s141[338],s140[340],s139[342],s138[344],s137[346],s136[348],s135[350],s134[352],s133[354],s132[356],s131[358],s130[360],s129[362],pp255[172],pp254[174],pp253[176],pp252[178],pp251[180],pp250[182],pp249[184],pp248[186],pp247[188],pp246[190],pp245[192],pp244[194],pp243[196],pp242[198],pp241[200],pp240[202],pp239[204],pp238[206],pp237[208],pp236[210],pp235[212],pp234[214],pp235[214],pp236[214],pp237[214],pp238[214],pp239[214],pp240[214],pp241[214],pp242[214],pp243[214],pp244[214],pp245[214]};
    CLA_408 KS_213(s213, c213, in213_1, in213_2);
    wire[405:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {s201[13],s200[15],s199[17],s198[19],s197[21],s196[23],s195[25],s194[27],s193[29],pp52[10],pp52[11],pp54[10],s193[33],s194[33],s195[33],s196[33],s197[33],s198[33],s199[33],s200[33],s201[33],s201[34],s201[35],s201[36],s201[37],s201[38],s201[39],s201[40],s201[41],s201[42],s201[43],s201[44],s201[45],s201[46],s201[47],s201[48],s201[49],s201[50],s201[51],s201[52],s201[53],s201[54],s201[55],s201[56],s201[57],s201[58],s201[59],s199[62],s197[65],s195[68],s193[71],s158[11],s157[13],s156[15],s155[17],s154[19],s153[21],s154[21],s155[21],s156[21],s157[21],s158[21],s159[21],s160[21],s161[21],s162[21],s163[21],s164[21],s165[21],s166[21],s167[21],s168[21],s169[21],s170[21],s171[21],s172[21],s173[21],s174[21],s175[21],s175[22],s175[23],s175[24],s175[25],s175[26],s175[27],s175[28],s175[29],s175[30],s175[31],s175[32],s175[33],s175[34],s175[35],s175[36],s175[37],s175[38],s175[39],s175[40],s175[41],s213[100],s213[101],s213[102],s213[103],s213[104],s213[105],s213[106],s213[107],s213[108],s213[109],s213[110],s213[111],s213[112],s213[113],s213[114],s213[115],s213[116],s213[117],s213[118],s213[119],s213[120],s213[121],s213[122],s213[123],s213[124],s213[125],s213[126],s213[127],s213[128],s213[129],s213[130],s213[131],s213[132],s213[133],s213[134],s213[135],s213[136],s213[137],s213[138],s213[139],s213[140],s213[141],s213[142],s213[143],s213[144],s213[145],s213[146],s213[147],s213[148],s213[149],s213[150],s213[151],s213[152],s213[153],s213[154],s213[155],s213[156],s213[157],s213[158],s213[159],s213[160],s213[161],s213[162],s213[163],s213[164],s213[165],s213[166],s213[167],s213[168],s213[169],s213[170],s213[171],s213[172],s213[173],s213[174],s213[175],s213[176],s213[177],s213[178],s213[179],s213[180],s213[181],s213[182],s213[183],s213[184],s213[185],s213[186],s213[187],s213[188],s213[189],s213[190],s213[191],s213[192],s213[193],s213[194],s213[195],s213[196],s213[197],s213[198],s213[199],s213[200],s213[201],s213[202],s213[203],s213[204],s213[205],s213[206],s213[207],s213[208],s213[209],s213[210],s213[211],s213[212],s213[213],s213[214],s213[215],s213[216],s213[217],s213[218],s213[219],s213[220],s213[221],s213[222],s213[223],s213[224],s213[225],s213[226],s213[227],s213[228],s213[229],s213[230],s213[231],s213[232],s213[233],s213[234],s213[235],s213[236],s213[237],s213[238],s213[239],s213[240],s213[241],s213[242],s213[243],s213[244],s213[245],s213[246],s213[247],s213[248],s213[249],s213[250],s213[251],s213[252],s213[253],s213[254],s213[255],s213[256],s213[257],s213[258],s213[259],s213[260],s213[261],s213[262],s213[263],s213[264],s213[265],s213[266],s213[267],s213[268],s213[269],s213[270],s213[271],s213[272],s213[273],s213[274],s213[275],s213[276],s213[277],s213[278],s213[279],s213[280],s213[281],s213[282],s213[283],s213[284],s213[285],s213[286],s213[287],s213[288],s213[289],s213[290],s213[291],s212[293],s211[295],s210[297],s209[299],s208[301],s207[303],s206[305],s205[307],s204[309],s203[311],s202[313],s201[315],s200[317],s199[319],s198[321],s197[323],s196[325],s195[327],s194[329],s193[331],s192[237],s191[239],s190[241],s189[243],s188[245],s187[247],s186[249],s185[251],s184[253],s183[255],s182[257],s181[259],s180[261],s179[263],s178[265],s177[267],s176[269],s175[271],s174[273],s173[275],s172[277],s171[279],s170[281],s169[283],s168[285],s167[287],s166[289],s165[291],s164[293],s163[295],s162[297],s161[299],s160[301],s159[303],s158[305],s157[307],s156[309],s155[311],s154[313],s153[315],s152[317],s151[319],s150[321],s149[323],s148[325],s147[327],s146[329],s145[331],s144[333],s143[335],s142[337],s141[339],s140[341],s139[343],s138[345],s137[347],s136[349],s135[351],s134[353],s133[355],s132[357],s131[359],s130[361],s129[363],pp255[173],pp254[175],pp253[177],pp252[179],pp251[181],pp250[183],pp249[185],pp248[187],pp247[189],pp246[191],pp245[193],pp244[195],pp243[197],pp242[199],pp241[201],pp240[203],pp239[205],pp238[207],pp237[209],pp236[211],pp235[213],pp236[213],pp237[213],pp238[213],pp239[213],pp240[213],pp241[213],pp242[213],pp243[213],pp244[213],pp245[213]};
    assign in214_2 = {s202[12],s201[14],s200[16],s199[18],s198[20],s197[22],s196[24],s195[26],s194[28],s193[30],pp53[10],s193[32],s194[32],s195[32],s196[32],s197[32],s198[32],s199[32],s200[32],s201[32],s202[32],s202[33],s202[34],s202[35],s202[36],s202[37],s202[38],s202[39],s202[40],s202[41],s202[42],s202[43],s202[44],s202[45],s202[46],s202[47],s202[48],s202[49],s202[50],s202[51],s202[52],s202[53],s202[54],s202[55],s202[56],s202[57],s202[58],s200[61],s198[64],s196[67],s194[70],s159[10],s158[12],s157[14],s156[16],s155[18],s154[20],s155[20],s156[20],s157[20],s158[20],s159[20],s160[20],s161[20],s162[20],s163[20],s164[20],s165[20],s166[20],s167[20],s168[20],s169[20],s170[20],s171[20],s172[20],s173[20],s174[20],s175[20],s176[20],s176[21],s176[22],s176[23],s176[24],s176[25],s176[26],s176[27],s176[28],s176[29],s176[30],s176[31],s176[32],s176[33],s176[34],s176[35],s176[36],s176[37],s176[38],s176[39],s176[40],s176[41],s177[41],s178[41],s179[41],s180[41],s181[41],s182[41],s183[41],s184[41],s185[41],s186[41],s187[41],s188[41],s189[41],s190[41],s191[41],s192[41],s10[32],s11[32],s12[32],s13[32],s14[32],s15[32],s16[32],s17[32],s18[32],s19[32],s20[32],s21[32],s22[32],s23[32],s24[32],s25[32],s26[32],s27[32],s28[32],s29[32],s30[32],s31[32],s32[32],s33[32],s34[32],s35[32],s36[32],s37[32],s38[32],s39[32],s40[32],s41[32],s42[32],s43[32],s44[32],s45[32],s46[32],s47[32],s48[32],s49[32],s50[32],s51[32],s52[32],s53[32],s54[32],s55[32],s56[32],s57[32],s58[32],s59[32],s60[32],s61[32],s62[32],s63[32],s64[32],s65[32],s66[32],s67[32],s68[32],s68[33],s68[34],s68[35],s68[36],s68[37],s68[38],s68[39],s68[40],s68[41],s68[42],s68[43],s68[44],s68[45],s68[46],s68[47],s68[48],s68[49],s68[50],s68[51],s68[52],s68[53],s68[54],s68[55],s68[56],s68[57],s68[58],s68[59],s68[60],s68[61],s66[64],s64[67],s62[70],s60[73],s59[75],s59[76],s59[77],s59[78],s59[79],s59[80],s59[81],s59[82],s59[83],s59[84],s59[85],s59[86],s59[87],s59[88],s59[89],s59[90],s59[91],s59[92],s59[93],s59[94],s59[95],s59[96],s59[97],s59[98],s59[99],s8[151],s6[154],s4[157],s2[160],s63[100],s62[102],s61[104],s60[106],s59[108],s58[110],s57[112],s56[114],s55[116],s54[118],s53[120],s52[122],s51[124],s50[126],s49[128],s48[130],s47[132],s46[134],s45[136],s44[138],s43[140],s42[142],s41[144],s40[146],s39[148],s38[150],s37[152],s36[154],s35[156],s34[158],s33[160],s32[162],s31[164],s30[166],s29[168],s28[170],s27[172],s26[174],s25[176],s24[178],s23[180],s22[182],s21[184],s20[186],s19[188],s18[190],s17[192],s16[194],s15[196],s14[198],s13[200],s12[202],s11[204],s10[206],s213[292],s212[294],s211[296],s210[298],s209[300],s208[302],s207[304],s206[306],s205[308],s204[310],s203[312],s202[314],s201[316],s200[318],s199[320],s198[322],s197[324],s196[326],s195[328],s194[330],s193[332],s192[238],s191[240],s190[242],s189[244],s188[246],s187[248],s186[250],s185[252],s184[254],s183[256],s182[258],s181[260],s180[262],s179[264],s178[266],s177[268],s176[270],s175[272],s174[274],s173[276],s172[278],s171[280],s170[282],s169[284],s168[286],s167[288],s166[290],s165[292],s164[294],s163[296],s162[298],s161[300],s160[302],s159[304],s158[306],s157[308],s156[310],s155[312],s154[314],s153[316],s152[318],s151[320],s150[322],s149[324],s148[326],s147[328],s146[330],s145[332],s144[334],s143[336],s142[338],s141[340],s140[342],s139[344],s138[346],s137[348],s136[350],s135[352],s134[354],s133[356],s132[358],s131[360],s130[362],s129[364],pp255[174],pp254[176],pp253[178],pp252[180],pp251[182],pp250[184],pp249[186],pp248[188],pp247[190],pp246[192],pp245[194],pp244[196],pp243[198],pp242[200],pp241[202],pp240[204],pp239[206],pp238[208],pp237[210],pp236[212],pp237[212],pp238[212],pp239[212],pp240[212],pp241[212],pp242[212],pp243[212],pp244[212],pp245[212],pp246[212]};
    CLA_406 KS_214(s214, c214, in214_1, in214_2);
    wire[403:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {s202[13],s201[15],s200[17],s199[19],s198[21],s197[23],s196[25],s195[27],s194[29],s193[31],s194[31],s195[31],s196[31],s197[31],s198[31],s199[31],s200[31],s201[31],s202[31],s203[31],s203[32],s203[33],s203[34],s203[35],s203[36],s203[37],s203[38],s203[39],s203[40],s203[41],s203[42],s203[43],s203[44],s203[45],s203[46],s203[47],s203[48],s203[49],s203[50],s203[51],s203[52],s203[53],s203[54],s203[55],s203[56],s203[57],s201[60],s199[63],s197[66],s195[69],s193[72],s159[11],s158[13],s157[15],s156[17],s155[19],s156[19],s157[19],s158[19],s159[19],s160[19],s161[19],s162[19],s163[19],s164[19],s165[19],s166[19],s167[19],s168[19],s169[19],s170[19],s171[19],s172[19],s173[19],s174[19],s175[19],s176[19],s177[19],s177[20],s177[21],s177[22],s177[23],s177[24],s177[25],s177[26],s177[27],s177[28],s177[29],s177[30],s177[31],s177[32],s177[33],s177[34],s177[35],s177[36],s177[37],s177[38],s177[39],s177[40],s214[100],s214[101],s214[102],s214[103],s214[104],s214[105],s214[106],s214[107],s214[108],s214[109],s214[110],s214[111],s214[112],s214[113],s214[114],s214[115],s214[116],s214[117],s214[118],s214[119],s214[120],s214[121],s214[122],s214[123],s214[124],s214[125],s214[126],s214[127],s214[128],s214[129],s214[130],s214[131],s214[132],s214[133],s214[134],s214[135],s214[136],s214[137],s214[138],s214[139],s214[140],s214[141],s214[142],s214[143],s214[144],s214[145],s214[146],s214[147],s214[148],s214[149],s214[150],s214[151],s214[152],s214[153],s214[154],s214[155],s214[156],s214[157],s214[158],s214[159],s214[160],s214[161],s214[162],s214[163],s214[164],s214[165],s214[166],s214[167],s214[168],s214[169],s214[170],s214[171],s214[172],s214[173],s214[174],s214[175],s214[176],s214[177],s214[178],s214[179],s214[180],s214[181],s214[182],s214[183],s214[184],s214[185],s214[186],s214[187],s214[188],s214[189],s214[190],s214[191],s214[192],s214[193],s214[194],s214[195],s214[196],s214[197],s214[198],s214[199],s214[200],s214[201],s214[202],s214[203],s214[204],s214[205],s214[206],s214[207],s214[208],s214[209],s214[210],s214[211],s214[212],s214[213],s214[214],s214[215],s214[216],s214[217],s214[218],s214[219],s214[220],s214[221],s214[222],s214[223],s214[224],s214[225],s214[226],s214[227],s214[228],s214[229],s214[230],s214[231],s214[232],s214[233],s214[234],s214[235],s214[236],s214[237],s214[238],s214[239],s214[240],s214[241],s214[242],s214[243],s214[244],s214[245],s214[246],s214[247],s214[248],s214[249],s214[250],s214[251],s214[252],s214[253],s214[254],s214[255],s214[256],s214[257],s214[258],s214[259],s214[260],s214[261],s214[262],s214[263],s214[264],s214[265],s214[266],s214[267],s214[268],s214[269],s214[270],s214[271],s214[272],s214[273],s214[274],s214[275],s214[276],s214[277],s214[278],s214[279],s214[280],s214[281],s214[282],s214[283],s214[284],s214[285],s214[286],s214[287],s214[288],s214[289],s214[290],s214[291],s213[293],s212[295],s211[297],s210[299],s209[301],s208[303],s207[305],s206[307],s205[309],s204[311],s203[313],s202[315],s201[317],s200[319],s199[321],s198[323],s197[325],s196[327],s195[329],s194[331],s193[333],s192[239],s191[241],s190[243],s189[245],s188[247],s187[249],s186[251],s185[253],s184[255],s183[257],s182[259],s181[261],s180[263],s179[265],s178[267],s177[269],s176[271],s175[273],s174[275],s173[277],s172[279],s171[281],s170[283],s169[285],s168[287],s167[289],s166[291],s165[293],s164[295],s163[297],s162[299],s161[301],s160[303],s159[305],s158[307],s157[309],s156[311],s155[313],s154[315],s153[317],s152[319],s151[321],s150[323],s149[325],s148[327],s147[329],s146[331],s145[333],s144[335],s143[337],s142[339],s141[341],s140[343],s139[345],s138[347],s137[349],s136[351],s135[353],s134[355],s133[357],s132[359],s131[361],s130[363],s129[365],pp255[175],pp254[177],pp253[179],pp252[181],pp251[183],pp250[185],pp249[187],pp248[189],pp247[191],pp246[193],pp245[195],pp244[197],pp243[199],pp242[201],pp241[203],pp240[205],pp239[207],pp238[209],pp237[211],pp238[211],pp239[211],pp240[211],pp241[211],pp242[211],pp243[211],pp244[211],pp245[211],pp246[211]};
    assign in215_2 = {s203[12],s202[14],s201[16],s200[18],s199[20],s198[22],s197[24],s196[26],s195[28],s194[30],s195[30],s196[30],s197[30],s198[30],s199[30],s200[30],s201[30],s202[30],s203[30],s204[30],s204[31],s204[32],s204[33],s204[34],s204[35],s204[36],s204[37],s204[38],s204[39],s204[40],s204[41],s204[42],s204[43],s204[44],s204[45],s204[46],s204[47],s204[48],s204[49],s204[50],s204[51],s204[52],s204[53],s204[54],s204[55],s204[56],s202[59],s200[62],s198[65],s196[68],s194[71],s160[10],s159[12],s158[14],s157[16],s156[18],s157[18],s158[18],s159[18],s160[18],s161[18],s162[18],s163[18],s164[18],s165[18],s166[18],s167[18],s168[18],s169[18],s170[18],s171[18],s172[18],s173[18],s174[18],s175[18],s176[18],s177[18],s178[18],s178[19],s178[20],s178[21],s178[22],s178[23],s178[24],s178[25],s178[26],s178[27],s178[28],s178[29],s178[30],s178[31],s178[32],s178[33],s178[34],s178[35],s178[36],s178[37],s178[38],s178[39],s178[40],s179[40],s180[40],s181[40],s182[40],s183[40],s184[40],s185[40],s186[40],s187[40],s188[40],s189[40],s190[40],s191[40],s192[40],s10[31],s11[31],s12[31],s13[31],s14[31],s15[31],s16[31],s17[31],s18[31],s19[31],s20[31],s21[31],s22[31],s23[31],s24[31],s25[31],s26[31],s27[31],s28[31],s29[31],s30[31],s31[31],s32[31],s33[31],s34[31],s35[31],s36[31],s37[31],s38[31],s39[31],s40[31],s41[31],s42[31],s43[31],s44[31],s45[31],s46[31],s47[31],s48[31],s49[31],s50[31],s51[31],s52[31],s53[31],s54[31],s55[31],s56[31],s57[31],s58[31],s59[31],s60[31],s61[31],s62[31],s63[31],s64[31],s65[31],s66[31],s67[31],s68[31],s69[31],s69[32],s69[33],s69[34],s69[35],s69[36],s69[37],s69[38],s69[39],s69[40],s69[41],s69[42],s69[43],s69[44],s69[45],s69[46],s69[47],s69[48],s69[49],s69[50],s69[51],s69[52],s69[53],s69[54],s69[55],s69[56],s69[57],s69[58],s69[59],s69[60],s67[63],s65[66],s63[69],s61[72],s60[74],s60[75],s60[76],s60[77],s60[78],s60[79],s60[80],s60[81],s60[82],s60[83],s60[84],s60[85],s60[86],s60[87],s60[88],s60[89],s60[90],s60[91],s60[92],s60[93],s60[94],s60[95],s60[96],s60[97],s60[98],s9[150],s7[153],s5[156],s3[159],s1[162],s63[101],s62[103],s61[105],s60[107],s59[109],s58[111],s57[113],s56[115],s55[117],s54[119],s53[121],s52[123],s51[125],s50[127],s49[129],s48[131],s47[133],s46[135],s45[137],s44[139],s43[141],s42[143],s41[145],s40[147],s39[149],s38[151],s37[153],s36[155],s35[157],s34[159],s33[161],s32[163],s31[165],s30[167],s29[169],s28[171],s27[173],s26[175],s25[177],s24[179],s23[181],s22[183],s21[185],s20[187],s19[189],s18[191],s17[193],s16[195],s15[197],s14[199],s13[201],s12[203],s11[205],s10[207],s214[292],s213[294],s212[296],s211[298],s210[300],s209[302],s208[304],s207[306],s206[308],s205[310],s204[312],s203[314],s202[316],s201[318],s200[320],s199[322],s198[324],s197[326],s196[328],s195[330],s194[332],s193[334],s192[240],s191[242],s190[244],s189[246],s188[248],s187[250],s186[252],s185[254],s184[256],s183[258],s182[260],s181[262],s180[264],s179[266],s178[268],s177[270],s176[272],s175[274],s174[276],s173[278],s172[280],s171[282],s170[284],s169[286],s168[288],s167[290],s166[292],s165[294],s164[296],s163[298],s162[300],s161[302],s160[304],s159[306],s158[308],s157[310],s156[312],s155[314],s154[316],s153[318],s152[320],s151[322],s150[324],s149[326],s148[328],s147[330],s146[332],s145[334],s144[336],s143[338],s142[340],s141[342],s140[344],s139[346],s138[348],s137[350],s136[352],s135[354],s134[356],s133[358],s132[360],s131[362],s130[364],s129[366],pp255[176],pp254[178],pp253[180],pp252[182],pp251[184],pp250[186],pp249[188],pp248[190],pp247[192],pp246[194],pp245[196],pp244[198],pp243[200],pp242[202],pp241[204],pp240[206],pp239[208],pp238[210],pp239[210],pp240[210],pp241[210],pp242[210],pp243[210],pp244[210],pp245[210],pp246[210],pp247[210]};
    CLA_404 KS_215(s215, c215, in215_1, in215_2);
    wire[401:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {s203[13],s202[15],s201[17],s200[19],s199[21],s198[23],s197[25],s196[27],s195[29],s196[29],s197[29],s198[29],s199[29],s200[29],s201[29],s202[29],s203[29],s204[29],s205[29],s205[30],s205[31],s205[32],s205[33],s205[34],s205[35],s205[36],s205[37],s205[38],s205[39],s205[40],s205[41],s205[42],s205[43],s205[44],s205[45],s205[46],s205[47],s205[48],s205[49],s205[50],s205[51],s205[52],s205[53],s205[54],s205[55],s203[58],s201[61],s199[64],s197[67],s195[70],s193[73],s160[11],s159[13],s158[15],s157[17],s158[17],s159[17],s160[17],s161[17],s162[17],s163[17],s164[17],s165[17],s166[17],s167[17],s168[17],s169[17],s170[17],s171[17],s172[17],s173[17],s174[17],s175[17],s176[17],s177[17],s178[17],s179[17],s179[18],s179[19],s179[20],s179[21],s179[22],s179[23],s179[24],s179[25],s179[26],s179[27],s179[28],s179[29],s179[30],s179[31],s179[32],s179[33],s179[34],s179[35],s179[36],s179[37],s179[38],s179[39],s215[100],s215[101],s215[102],s215[103],s215[104],s215[105],s215[106],s215[107],s215[108],s215[109],s215[110],s215[111],s215[112],s215[113],s215[114],s215[115],s215[116],s215[117],s215[118],s215[119],s215[120],s215[121],s215[122],s215[123],s215[124],s215[125],s215[126],s215[127],s215[128],s215[129],s215[130],s215[131],s215[132],s215[133],s215[134],s215[135],s215[136],s215[137],s215[138],s215[139],s215[140],s215[141],s215[142],s215[143],s215[144],s215[145],s215[146],s215[147],s215[148],s215[149],s215[150],s215[151],s215[152],s215[153],s215[154],s215[155],s215[156],s215[157],s215[158],s215[159],s215[160],s215[161],s215[162],s215[163],s215[164],s215[165],s215[166],s215[167],s215[168],s215[169],s215[170],s215[171],s215[172],s215[173],s215[174],s215[175],s215[176],s215[177],s215[178],s215[179],s215[180],s215[181],s215[182],s215[183],s215[184],s215[185],s215[186],s215[187],s215[188],s215[189],s215[190],s215[191],s215[192],s215[193],s215[194],s215[195],s215[196],s215[197],s215[198],s215[199],s215[200],s215[201],s215[202],s215[203],s215[204],s215[205],s215[206],s215[207],s215[208],s215[209],s215[210],s215[211],s215[212],s215[213],s215[214],s215[215],s215[216],s215[217],s215[218],s215[219],s215[220],s215[221],s215[222],s215[223],s215[224],s215[225],s215[226],s215[227],s215[228],s215[229],s215[230],s215[231],s215[232],s215[233],s215[234],s215[235],s215[236],s215[237],s215[238],s215[239],s215[240],s215[241],s215[242],s215[243],s215[244],s215[245],s215[246],s215[247],s215[248],s215[249],s215[250],s215[251],s215[252],s215[253],s215[254],s215[255],s215[256],s215[257],s215[258],s215[259],s215[260],s215[261],s215[262],s215[263],s215[264],s215[265],s215[266],s215[267],s215[268],s215[269],s215[270],s215[271],s215[272],s215[273],s215[274],s215[275],s215[276],s215[277],s215[278],s215[279],s215[280],s215[281],s215[282],s215[283],s215[284],s215[285],s215[286],s215[287],s215[288],s215[289],s215[290],s215[291],s214[293],s213[295],s212[297],s211[299],s210[301],s209[303],s208[305],s207[307],s206[309],s205[311],s204[313],s203[315],s202[317],s201[319],s200[321],s199[323],s198[325],s197[327],s196[329],s195[331],s194[333],s193[335],s192[241],s191[243],s190[245],s189[247],s188[249],s187[251],s186[253],s185[255],s184[257],s183[259],s182[261],s181[263],s180[265],s179[267],s178[269],s177[271],s176[273],s175[275],s174[277],s173[279],s172[281],s171[283],s170[285],s169[287],s168[289],s167[291],s166[293],s165[295],s164[297],s163[299],s162[301],s161[303],s160[305],s159[307],s158[309],s157[311],s156[313],s155[315],s154[317],s153[319],s152[321],s151[323],s150[325],s149[327],s148[329],s147[331],s146[333],s145[335],s144[337],s143[339],s142[341],s141[343],s140[345],s139[347],s138[349],s137[351],s136[353],s135[355],s134[357],s133[359],s132[361],s131[363],s130[365],s129[367],pp255[177],pp254[179],pp253[181],pp252[183],pp251[185],pp250[187],pp249[189],pp248[191],pp247[193],pp246[195],pp245[197],pp244[199],pp243[201],pp242[203],pp241[205],pp240[207],pp239[209],pp240[209],pp241[209],pp242[209],pp243[209],pp244[209],pp245[209],pp246[209],pp247[209]};
    assign in216_2 = {s204[12],s203[14],s202[16],s201[18],s200[20],s199[22],s198[24],s197[26],s196[28],s197[28],s198[28],s199[28],s200[28],s201[28],s202[28],s203[28],s204[28],s205[28],s206[28],s206[29],s206[30],s206[31],s206[32],s206[33],s206[34],s206[35],s206[36],s206[37],s206[38],s206[39],s206[40],s206[41],s206[42],s206[43],s206[44],s206[45],s206[46],s206[47],s206[48],s206[49],s206[50],s206[51],s206[52],s206[53],s206[54],s204[57],s202[60],s200[63],s198[66],s196[69],s194[72],s161[10],s160[12],s159[14],s158[16],s159[16],s160[16],s161[16],s162[16],s163[16],s164[16],s165[16],s166[16],s167[16],s168[16],s169[16],s170[16],s171[16],s172[16],s173[16],s174[16],s175[16],s176[16],s177[16],s178[16],s179[16],s180[16],s180[17],s180[18],s180[19],s180[20],s180[21],s180[22],s180[23],s180[24],s180[25],s180[26],s180[27],s180[28],s180[29],s180[30],s180[31],s180[32],s180[33],s180[34],s180[35],s180[36],s180[37],s180[38],s180[39],s181[39],s182[39],s183[39],s184[39],s185[39],s186[39],s187[39],s188[39],s189[39],s190[39],s191[39],s192[39],s10[30],s11[30],s12[30],s13[30],s14[30],s15[30],s16[30],s17[30],s18[30],s19[30],s20[30],s21[30],s22[30],s23[30],s24[30],s25[30],s26[30],s27[30],s28[30],s29[30],s30[30],s31[30],s32[30],s33[30],s34[30],s35[30],s36[30],s37[30],s38[30],s39[30],s40[30],s41[30],s42[30],s43[30],s44[30],s45[30],s46[30],s47[30],s48[30],s49[30],s50[30],s51[30],s52[30],s53[30],s54[30],s55[30],s56[30],s57[30],s58[30],s59[30],s60[30],s61[30],s62[30],s63[30],s64[30],s65[30],s66[30],s67[30],s68[30],s69[30],s70[30],s70[31],s70[32],s70[33],s70[34],s70[35],s70[36],s70[37],s70[38],s70[39],s70[40],s70[41],s70[42],s70[43],s70[44],s70[45],s70[46],s70[47],s70[48],s70[49],s70[50],s70[51],s70[52],s70[53],s70[54],s70[55],s70[56],s70[57],s70[58],s70[59],s68[62],s66[65],s64[68],s62[71],s61[73],s61[74],s61[75],s61[76],s61[77],s61[78],s61[79],s61[80],s61[81],s61[82],s61[83],s61[84],s61[85],s61[86],s61[87],s61[88],s61[89],s61[90],s61[91],s61[92],s61[93],s61[94],s61[95],s61[96],s61[97],s60[99],s8[152],s6[155],s4[158],s2[161],s64[100],s63[102],s62[104],s61[106],s60[108],s59[110],s58[112],s57[114],s56[116],s55[118],s54[120],s53[122],s52[124],s51[126],s50[128],s49[130],s48[132],s47[134],s46[136],s45[138],s44[140],s43[142],s42[144],s41[146],s40[148],s39[150],s38[152],s37[154],s36[156],s35[158],s34[160],s33[162],s32[164],s31[166],s30[168],s29[170],s28[172],s27[174],s26[176],s25[178],s24[180],s23[182],s22[184],s21[186],s20[188],s19[190],s18[192],s17[194],s16[196],s15[198],s14[200],s13[202],s12[204],s11[206],s10[208],s215[292],s214[294],s213[296],s212[298],s211[300],s210[302],s209[304],s208[306],s207[308],s206[310],s205[312],s204[314],s203[316],s202[318],s201[320],s200[322],s199[324],s198[326],s197[328],s196[330],s195[332],s194[334],s193[336],s192[242],s191[244],s190[246],s189[248],s188[250],s187[252],s186[254],s185[256],s184[258],s183[260],s182[262],s181[264],s180[266],s179[268],s178[270],s177[272],s176[274],s175[276],s174[278],s173[280],s172[282],s171[284],s170[286],s169[288],s168[290],s167[292],s166[294],s165[296],s164[298],s163[300],s162[302],s161[304],s160[306],s159[308],s158[310],s157[312],s156[314],s155[316],s154[318],s153[320],s152[322],s151[324],s150[326],s149[328],s148[330],s147[332],s146[334],s145[336],s144[338],s143[340],s142[342],s141[344],s140[346],s139[348],s138[350],s137[352],s136[354],s135[356],s134[358],s133[360],s132[362],s131[364],s130[366],s129[368],pp255[178],pp254[180],pp253[182],pp252[184],pp251[186],pp250[188],pp249[190],pp248[192],pp247[194],pp246[196],pp245[198],pp244[200],pp243[202],pp242[204],pp241[206],pp240[208],pp241[208],pp242[208],pp243[208],pp244[208],pp245[208],pp246[208],pp247[208],pp248[208]};
    CLA_402 KS_216(s216, c216, in216_1, in216_2);
    wire[399:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {s204[13],s203[15],s202[17],s201[19],s200[21],s199[23],s198[25],s197[27],s198[27],s199[27],s200[27],s201[27],s202[27],s203[27],s204[27],s205[27],s206[27],s207[27],s207[28],s207[29],s207[30],s207[31],s207[32],s207[33],s207[34],s207[35],s207[36],s207[37],s207[38],s207[39],s207[40],s207[41],s207[42],s207[43],s207[44],s207[45],s207[46],s207[47],s207[48],s207[49],s207[50],s207[51],s207[52],s207[53],s205[56],s203[59],s201[62],s199[65],s197[68],s195[71],s193[74],s161[11],s160[13],s159[15],s160[15],s161[15],s162[15],s163[15],s164[15],s165[15],s166[15],s167[15],s168[15],s169[15],s170[15],s171[15],s172[15],s173[15],s174[15],s175[15],s176[15],s177[15],s178[15],s179[15],s180[15],s181[15],s181[16],s181[17],s181[18],s181[19],s181[20],s181[21],s181[22],s181[23],s181[24],s181[25],s181[26],s181[27],s181[28],s181[29],s181[30],s181[31],s181[32],s181[33],s181[34],s181[35],s181[36],s181[37],s181[38],s216[100],s216[101],s216[102],s216[103],s216[104],s216[105],s216[106],s216[107],s216[108],s216[109],s216[110],s216[111],s216[112],s216[113],s216[114],s216[115],s216[116],s216[117],s216[118],s216[119],s216[120],s216[121],s216[122],s216[123],s216[124],s216[125],s216[126],s216[127],s216[128],s216[129],s216[130],s216[131],s216[132],s216[133],s216[134],s216[135],s216[136],s216[137],s216[138],s216[139],s216[140],s216[141],s216[142],s216[143],s216[144],s216[145],s216[146],s216[147],s216[148],s216[149],s216[150],s216[151],s216[152],s216[153],s216[154],s216[155],s216[156],s216[157],s216[158],s216[159],s216[160],s216[161],s216[162],s216[163],s216[164],s216[165],s216[166],s216[167],s216[168],s216[169],s216[170],s216[171],s216[172],s216[173],s216[174],s216[175],s216[176],s216[177],s216[178],s216[179],s216[180],s216[181],s216[182],s216[183],s216[184],s216[185],s216[186],s216[187],s216[188],s216[189],s216[190],s216[191],s216[192],s216[193],s216[194],s216[195],s216[196],s216[197],s216[198],s216[199],s216[200],s216[201],s216[202],s216[203],s216[204],s216[205],s216[206],s216[207],s216[208],s216[209],s216[210],s216[211],s216[212],s216[213],s216[214],s216[215],s216[216],s216[217],s216[218],s216[219],s216[220],s216[221],s216[222],s216[223],s216[224],s216[225],s216[226],s216[227],s216[228],s216[229],s216[230],s216[231],s216[232],s216[233],s216[234],s216[235],s216[236],s216[237],s216[238],s216[239],s216[240],s216[241],s216[242],s216[243],s216[244],s216[245],s216[246],s216[247],s216[248],s216[249],s216[250],s216[251],s216[252],s216[253],s216[254],s216[255],s216[256],s216[257],s216[258],s216[259],s216[260],s216[261],s216[262],s216[263],s216[264],s216[265],s216[266],s216[267],s216[268],s216[269],s216[270],s216[271],s216[272],s216[273],s216[274],s216[275],s216[276],s216[277],s216[278],s216[279],s216[280],s216[281],s216[282],s216[283],s216[284],s216[285],s216[286],s216[287],s216[288],s216[289],s216[290],s216[291],s215[293],s214[295],s213[297],s212[299],s211[301],s210[303],s209[305],s208[307],s207[309],s206[311],s205[313],s204[315],s203[317],s202[319],s201[321],s200[323],s199[325],s198[327],s197[329],s196[331],s195[333],s194[335],s193[337],s192[243],s191[245],s190[247],s189[249],s188[251],s187[253],s186[255],s185[257],s184[259],s183[261],s182[263],s181[265],s180[267],s179[269],s178[271],s177[273],s176[275],s175[277],s174[279],s173[281],s172[283],s171[285],s170[287],s169[289],s168[291],s167[293],s166[295],s165[297],s164[299],s163[301],s162[303],s161[305],s160[307],s159[309],s158[311],s157[313],s156[315],s155[317],s154[319],s153[321],s152[323],s151[325],s150[327],s149[329],s148[331],s147[333],s146[335],s145[337],s144[339],s143[341],s142[343],s141[345],s140[347],s139[349],s138[351],s137[353],s136[355],s135[357],s134[359],s133[361],s132[363],s131[365],s130[367],s129[369],pp255[179],pp254[181],pp253[183],pp252[185],pp251[187],pp250[189],pp249[191],pp248[193],pp247[195],pp246[197],pp245[199],pp244[201],pp243[203],pp242[205],pp241[207],pp242[207],pp243[207],pp244[207],pp245[207],pp246[207],pp247[207],pp248[207]};
    assign in217_2 = {s205[12],s204[14],s203[16],s202[18],s201[20],s200[22],s199[24],s198[26],s199[26],s200[26],s201[26],s202[26],s203[26],s204[26],s205[26],s206[26],s207[26],s208[26],s208[27],s208[28],s208[29],s208[30],s208[31],s208[32],s208[33],s208[34],s208[35],s208[36],s208[37],s208[38],s208[39],s208[40],s208[41],s208[42],s208[43],s208[44],s208[45],s208[46],s208[47],s208[48],s208[49],s208[50],s208[51],s208[52],s206[55],s204[58],s202[61],s200[64],s198[67],s196[70],s194[73],s162[10],s161[12],s160[14],s161[14],s162[14],s163[14],s164[14],s165[14],s166[14],s167[14],s168[14],s169[14],s170[14],s171[14],s172[14],s173[14],s174[14],s175[14],s176[14],s177[14],s178[14],s179[14],s180[14],s181[14],s182[14],s182[15],s182[16],s182[17],s182[18],s182[19],s182[20],s182[21],s182[22],s182[23],s182[24],s182[25],s182[26],s182[27],s182[28],s182[29],s182[30],s182[31],s182[32],s182[33],s182[34],s182[35],s182[36],s182[37],s182[38],s183[38],s184[38],s185[38],s186[38],s187[38],s188[38],s189[38],s190[38],s191[38],s192[38],s10[29],s11[29],s12[29],s13[29],s14[29],s15[29],s16[29],s17[29],s18[29],s19[29],s20[29],s21[29],s22[29],s23[29],s24[29],s25[29],s26[29],s27[29],s28[29],s29[29],s30[29],s31[29],s32[29],s33[29],s34[29],s35[29],s36[29],s37[29],s38[29],s39[29],s40[29],s41[29],s42[29],s43[29],s44[29],s45[29],s46[29],s47[29],s48[29],s49[29],s50[29],s51[29],s52[29],s53[29],s54[29],s55[29],s56[29],s57[29],s58[29],s59[29],s60[29],s61[29],s62[29],s63[29],s64[29],s65[29],s66[29],s67[29],s68[29],s69[29],s70[29],s71[29],s71[30],s71[31],s71[32],s71[33],s71[34],s71[35],s71[36],s71[37],s71[38],s71[39],s71[40],s71[41],s71[42],s71[43],s71[44],s71[45],s71[46],s71[47],s71[48],s71[49],s71[50],s71[51],s71[52],s71[53],s71[54],s71[55],s71[56],s71[57],s71[58],s69[61],s67[64],s65[67],s63[70],s62[72],s62[73],s62[74],s62[75],s62[76],s62[77],s62[78],s62[79],s62[80],s62[81],s62[82],s62[83],s62[84],s62[85],s62[86],s62[87],s62[88],s62[89],s62[90],s62[91],s62[92],s62[93],s62[94],s62[95],s62[96],s61[98],s9[151],s7[154],s5[157],s3[160],s1[163],s64[101],s63[103],s62[105],s61[107],s60[109],s59[111],s58[113],s57[115],s56[117],s55[119],s54[121],s53[123],s52[125],s51[127],s50[129],s49[131],s48[133],s47[135],s46[137],s45[139],s44[141],s43[143],s42[145],s41[147],s40[149],s39[151],s38[153],s37[155],s36[157],s35[159],s34[161],s33[163],s32[165],s31[167],s30[169],s29[171],s28[173],s27[175],s26[177],s25[179],s24[181],s23[183],s22[185],s21[187],s20[189],s19[191],s18[193],s17[195],s16[197],s15[199],s14[201],s13[203],s12[205],s11[207],s10[209],s216[292],s215[294],s214[296],s213[298],s212[300],s211[302],s210[304],s209[306],s208[308],s207[310],s206[312],s205[314],s204[316],s203[318],s202[320],s201[322],s200[324],s199[326],s198[328],s197[330],s196[332],s195[334],s194[336],s193[338],s192[244],s191[246],s190[248],s189[250],s188[252],s187[254],s186[256],s185[258],s184[260],s183[262],s182[264],s181[266],s180[268],s179[270],s178[272],s177[274],s176[276],s175[278],s174[280],s173[282],s172[284],s171[286],s170[288],s169[290],s168[292],s167[294],s166[296],s165[298],s164[300],s163[302],s162[304],s161[306],s160[308],s159[310],s158[312],s157[314],s156[316],s155[318],s154[320],s153[322],s152[324],s151[326],s150[328],s149[330],s148[332],s147[334],s146[336],s145[338],s144[340],s143[342],s142[344],s141[346],s140[348],s139[350],s138[352],s137[354],s136[356],s135[358],s134[360],s133[362],s132[364],s131[366],s130[368],s129[370],pp255[180],pp254[182],pp253[184],pp252[186],pp251[188],pp250[190],pp249[192],pp248[194],pp247[196],pp246[198],pp245[200],pp244[202],pp243[204],pp242[206],pp243[206],pp244[206],pp245[206],pp246[206],pp247[206],pp248[206],pp249[206]};
    CLA_400 KS_217(s217, c217, in217_1, in217_2);
    wire[397:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {s205[13],s204[15],s203[17],s202[19],s201[21],s200[23],s199[25],s200[25],s201[25],s202[25],s203[25],s204[25],s205[25],s206[25],s207[25],s208[25],s209[25],s209[26],s209[27],s209[28],s209[29],s209[30],s209[31],s209[32],s209[33],s209[34],s209[35],s209[36],s209[37],s209[38],s209[39],s209[40],s209[41],s209[42],s209[43],s209[44],s209[45],s209[46],s209[47],s209[48],s209[49],s209[50],s209[51],s207[54],s205[57],s203[60],s201[63],s199[66],s197[69],s195[72],s193[75],s162[11],s161[13],s162[13],s163[13],s164[13],s165[13],s166[13],s167[13],s168[13],s169[13],s170[13],s171[13],s172[13],s173[13],s174[13],s175[13],s176[13],s177[13],s178[13],s179[13],s180[13],s181[13],s182[13],s183[13],s183[14],s183[15],s183[16],s183[17],s183[18],s183[19],s183[20],s183[21],s183[22],s183[23],s183[24],s183[25],s183[26],s183[27],s183[28],s183[29],s183[30],s183[31],s183[32],s183[33],s183[34],s183[35],s183[36],s183[37],s217[100],s217[101],s217[102],s217[103],s217[104],s217[105],s217[106],s217[107],s217[108],s217[109],s217[110],s217[111],s217[112],s217[113],s217[114],s217[115],s217[116],s217[117],s217[118],s217[119],s217[120],s217[121],s217[122],s217[123],s217[124],s217[125],s217[126],s217[127],s217[128],s217[129],s217[130],s217[131],s217[132],s217[133],s217[134],s217[135],s217[136],s217[137],s217[138],s217[139],s217[140],s217[141],s217[142],s217[143],s217[144],s217[145],s217[146],s217[147],s217[148],s217[149],s217[150],s217[151],s217[152],s217[153],s217[154],s217[155],s217[156],s217[157],s217[158],s217[159],s217[160],s217[161],s217[162],s217[163],s217[164],s217[165],s217[166],s217[167],s217[168],s217[169],s217[170],s217[171],s217[172],s217[173],s217[174],s217[175],s217[176],s217[177],s217[178],s217[179],s217[180],s217[181],s217[182],s217[183],s217[184],s217[185],s217[186],s217[187],s217[188],s217[189],s217[190],s217[191],s217[192],s217[193],s217[194],s217[195],s217[196],s217[197],s217[198],s217[199],s217[200],s217[201],s217[202],s217[203],s217[204],s217[205],s217[206],s217[207],s217[208],s217[209],s217[210],s217[211],s217[212],s217[213],s217[214],s217[215],s217[216],s217[217],s217[218],s217[219],s217[220],s217[221],s217[222],s217[223],s217[224],s217[225],s217[226],s217[227],s217[228],s217[229],s217[230],s217[231],s217[232],s217[233],s217[234],s217[235],s217[236],s217[237],s217[238],s217[239],s217[240],s217[241],s217[242],s217[243],s217[244],s217[245],s217[246],s217[247],s217[248],s217[249],s217[250],s217[251],s217[252],s217[253],s217[254],s217[255],s217[256],s217[257],s217[258],s217[259],s217[260],s217[261],s217[262],s217[263],s217[264],s217[265],s217[266],s217[267],s217[268],s217[269],s217[270],s217[271],s217[272],s217[273],s217[274],s217[275],s217[276],s217[277],s217[278],s217[279],s217[280],s217[281],s217[282],s217[283],s217[284],s217[285],s217[286],s217[287],s217[288],s217[289],s217[290],s217[291],s216[293],s215[295],s214[297],s213[299],s212[301],s211[303],s210[305],s209[307],s208[309],s207[311],s206[313],s205[315],s204[317],s203[319],s202[321],s201[323],s200[325],s199[327],s198[329],s197[331],s196[333],s195[335],s194[337],s193[339],s192[245],s191[247],s190[249],s189[251],s188[253],s187[255],s186[257],s185[259],s184[261],s183[263],s182[265],s181[267],s180[269],s179[271],s178[273],s177[275],s176[277],s175[279],s174[281],s173[283],s172[285],s171[287],s170[289],s169[291],s168[293],s167[295],s166[297],s165[299],s164[301],s163[303],s162[305],s161[307],s160[309],s159[311],s158[313],s157[315],s156[317],s155[319],s154[321],s153[323],s152[325],s151[327],s150[329],s149[331],s148[333],s147[335],s146[337],s145[339],s144[341],s143[343],s142[345],s141[347],s140[349],s139[351],s138[353],s137[355],s136[357],s135[359],s134[361],s133[363],s132[365],s131[367],s130[369],s129[371],pp255[181],pp254[183],pp253[185],pp252[187],pp251[189],pp250[191],pp249[193],pp248[195],pp247[197],pp246[199],pp245[201],pp244[203],pp243[205],pp244[205],pp245[205],pp246[205],pp247[205],pp248[205],pp249[205]};
    assign in218_2 = {s206[12],s205[14],s204[16],s203[18],s202[20],s201[22],s200[24],s201[24],s202[24],s203[24],s204[24],s205[24],s206[24],s207[24],s208[24],s209[24],s210[24],s210[25],s210[26],s210[27],s210[28],s210[29],s210[30],s210[31],s210[32],s210[33],s210[34],s210[35],s210[36],s210[37],s210[38],s210[39],s210[40],s210[41],s210[42],s210[43],s210[44],s210[45],s210[46],s210[47],s210[48],s210[49],s210[50],s208[53],s206[56],s204[59],s202[62],s200[65],s198[68],s196[71],s194[74],s163[10],s162[12],s163[12],s164[12],s165[12],s166[12],s167[12],s168[12],s169[12],s170[12],s171[12],s172[12],s173[12],s174[12],s175[12],s176[12],s177[12],s178[12],s179[12],s180[12],s181[12],s182[12],s183[12],s184[12],s184[13],s184[14],s184[15],s184[16],s184[17],s184[18],s184[19],s184[20],s184[21],s184[22],s184[23],s184[24],s184[25],s184[26],s184[27],s184[28],s184[29],s184[30],s184[31],s184[32],s184[33],s184[34],s184[35],s184[36],s184[37],s185[37],s186[37],s187[37],s188[37],s189[37],s190[37],s191[37],s192[37],s10[28],s11[28],s12[28],s13[28],s14[28],s15[28],s16[28],s17[28],s18[28],s19[28],s20[28],s21[28],s22[28],s23[28],s24[28],s25[28],s26[28],s27[28],s28[28],s29[28],s30[28],s31[28],s32[28],s33[28],s34[28],s35[28],s36[28],s37[28],s38[28],s39[28],s40[28],s41[28],s42[28],s43[28],s44[28],s45[28],s46[28],s47[28],s48[28],s49[28],s50[28],s51[28],s52[28],s53[28],s54[28],s55[28],s56[28],s57[28],s58[28],s59[28],s60[28],s61[28],s62[28],s63[28],s64[28],s65[28],s66[28],s67[28],s68[28],s69[28],s70[28],s71[28],s72[28],s72[29],s72[30],s72[31],s72[32],s72[33],s72[34],s72[35],s72[36],s72[37],s72[38],s72[39],s72[40],s72[41],s72[42],s72[43],s72[44],s72[45],s72[46],s72[47],s72[48],s72[49],s72[50],s72[51],s72[52],s72[53],s72[54],s72[55],s72[56],s72[57],s70[60],s68[63],s66[66],s64[69],s63[71],s63[72],s63[73],s63[74],s63[75],s63[76],s63[77],s63[78],s63[79],s63[80],s63[81],s63[82],s63[83],s63[84],s63[85],s63[86],s63[87],s63[88],s63[89],s63[90],s63[91],s63[92],s63[93],s63[94],s63[95],s62[97],s61[99],s8[153],s6[156],s4[159],s2[162],s65[100],s64[102],s63[104],s62[106],s61[108],s60[110],s59[112],s58[114],s57[116],s56[118],s55[120],s54[122],s53[124],s52[126],s51[128],s50[130],s49[132],s48[134],s47[136],s46[138],s45[140],s44[142],s43[144],s42[146],s41[148],s40[150],s39[152],s38[154],s37[156],s36[158],s35[160],s34[162],s33[164],s32[166],s31[168],s30[170],s29[172],s28[174],s27[176],s26[178],s25[180],s24[182],s23[184],s22[186],s21[188],s20[190],s19[192],s18[194],s17[196],s16[198],s15[200],s14[202],s13[204],s12[206],s11[208],s10[210],s217[292],s216[294],s215[296],s214[298],s213[300],s212[302],s211[304],s210[306],s209[308],s208[310],s207[312],s206[314],s205[316],s204[318],s203[320],s202[322],s201[324],s200[326],s199[328],s198[330],s197[332],s196[334],s195[336],s194[338],s193[340],s192[246],s191[248],s190[250],s189[252],s188[254],s187[256],s186[258],s185[260],s184[262],s183[264],s182[266],s181[268],s180[270],s179[272],s178[274],s177[276],s176[278],s175[280],s174[282],s173[284],s172[286],s171[288],s170[290],s169[292],s168[294],s167[296],s166[298],s165[300],s164[302],s163[304],s162[306],s161[308],s160[310],s159[312],s158[314],s157[316],s156[318],s155[320],s154[322],s153[324],s152[326],s151[328],s150[330],s149[332],s148[334],s147[336],s146[338],s145[340],s144[342],s143[344],s142[346],s141[348],s140[350],s139[352],s138[354],s137[356],s136[358],s135[360],s134[362],s133[364],s132[366],s131[368],s130[370],s129[372],pp255[182],pp254[184],pp253[186],pp252[188],pp251[190],pp250[192],pp249[194],pp248[196],pp247[198],pp246[200],pp245[202],pp244[204],pp245[204],pp246[204],pp247[204],pp248[204],pp249[204],pp250[204]};
    CLA_398 KS_218(s218, c218, in218_1, in218_2);
    wire[395:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {s206[13],s205[15],s204[17],s203[19],s202[21],s201[23],s202[23],s203[23],s204[23],s205[23],s206[23],s207[23],s208[23],s209[23],s210[23],s211[23],s211[24],s211[25],s211[26],s211[27],s211[28],s211[29],s211[30],s211[31],s211[32],s211[33],s211[34],s211[35],s211[36],s211[37],s211[38],s211[39],s211[40],s211[41],s211[42],s211[43],s211[44],s211[45],s211[46],s211[47],s211[48],s211[49],s209[52],s207[55],s205[58],s203[61],s201[64],s199[67],s197[70],s195[73],s193[76],s163[11],s164[11],s165[11],s166[11],s167[11],s168[11],s169[11],s170[11],s171[11],s172[11],s173[11],s174[11],s175[11],s176[11],s177[11],s178[11],s179[11],s180[11],s181[11],s182[11],s183[11],s184[11],s185[11],s185[12],s185[13],s185[14],s185[15],s185[16],s185[17],s185[18],s185[19],s185[20],s185[21],s185[22],s185[23],s185[24],s185[25],s185[26],s185[27],s185[28],s185[29],s185[30],s185[31],s185[32],s185[33],s185[34],s185[35],s185[36],s218[100],s218[101],s218[102],s218[103],s218[104],s218[105],s218[106],s218[107],s218[108],s218[109],s218[110],s218[111],s218[112],s218[113],s218[114],s218[115],s218[116],s218[117],s218[118],s218[119],s218[120],s218[121],s218[122],s218[123],s218[124],s218[125],s218[126],s218[127],s218[128],s218[129],s218[130],s218[131],s218[132],s218[133],s218[134],s218[135],s218[136],s218[137],s218[138],s218[139],s218[140],s218[141],s218[142],s218[143],s218[144],s218[145],s218[146],s218[147],s218[148],s218[149],s218[150],s218[151],s218[152],s218[153],s218[154],s218[155],s218[156],s218[157],s218[158],s218[159],s218[160],s218[161],s218[162],s218[163],s218[164],s218[165],s218[166],s218[167],s218[168],s218[169],s218[170],s218[171],s218[172],s218[173],s218[174],s218[175],s218[176],s218[177],s218[178],s218[179],s218[180],s218[181],s218[182],s218[183],s218[184],s218[185],s218[186],s218[187],s218[188],s218[189],s218[190],s218[191],s218[192],s218[193],s218[194],s218[195],s218[196],s218[197],s218[198],s218[199],s218[200],s218[201],s218[202],s218[203],s218[204],s218[205],s218[206],s218[207],s218[208],s218[209],s218[210],s218[211],s218[212],s218[213],s218[214],s218[215],s218[216],s218[217],s218[218],s218[219],s218[220],s218[221],s218[222],s218[223],s218[224],s218[225],s218[226],s218[227],s218[228],s218[229],s218[230],s218[231],s218[232],s218[233],s218[234],s218[235],s218[236],s218[237],s218[238],s218[239],s218[240],s218[241],s218[242],s218[243],s218[244],s218[245],s218[246],s218[247],s218[248],s218[249],s218[250],s218[251],s218[252],s218[253],s218[254],s218[255],s218[256],s218[257],s218[258],s218[259],s218[260],s218[261],s218[262],s218[263],s218[264],s218[265],s218[266],s218[267],s218[268],s218[269],s218[270],s218[271],s218[272],s218[273],s218[274],s218[275],s218[276],s218[277],s218[278],s218[279],s218[280],s218[281],s218[282],s218[283],s218[284],s218[285],s218[286],s218[287],s218[288],s218[289],s218[290],s218[291],s217[293],s216[295],s215[297],s214[299],s213[301],s212[303],s211[305],s210[307],s209[309],s208[311],s207[313],s206[315],s205[317],s204[319],s203[321],s202[323],s201[325],s200[327],s199[329],s198[331],s197[333],s196[335],s195[337],s194[339],s193[341],s192[247],s191[249],s190[251],s189[253],s188[255],s187[257],s186[259],s185[261],s184[263],s183[265],s182[267],s181[269],s180[271],s179[273],s178[275],s177[277],s176[279],s175[281],s174[283],s173[285],s172[287],s171[289],s170[291],s169[293],s168[295],s167[297],s166[299],s165[301],s164[303],s163[305],s162[307],s161[309],s160[311],s159[313],s158[315],s157[317],s156[319],s155[321],s154[323],s153[325],s152[327],s151[329],s150[331],s149[333],s148[335],s147[337],s146[339],s145[341],s144[343],s143[345],s142[347],s141[349],s140[351],s139[353],s138[355],s137[357],s136[359],s135[361],s134[363],s133[365],s132[367],s131[369],s130[371],s129[373],pp255[183],pp254[185],pp253[187],pp252[189],pp251[191],pp250[193],pp249[195],pp248[197],pp247[199],pp246[201],pp245[203],pp246[203],pp247[203],pp248[203],pp249[203],pp250[203]};
    assign in219_2 = {s207[12],s206[14],s205[16],s204[18],s203[20],s202[22],s203[22],s204[22],s205[22],s206[22],s207[22],s208[22],s209[22],s210[22],s211[22],s212[22],s212[23],s212[24],s212[25],s212[26],s212[27],s212[28],s212[29],s212[30],s212[31],s212[32],s212[33],s212[34],s212[35],s212[36],s212[37],s212[38],s212[39],s212[40],s212[41],s212[42],s212[43],s212[44],s212[45],s212[46],s212[47],s212[48],s210[51],s208[54],s206[57],s204[60],s202[63],s200[66],s198[69],s196[72],s194[75],s164[10],s165[10],s166[10],s167[10],s168[10],s169[10],s170[10],s171[10],s172[10],s173[10],s174[10],s175[10],s176[10],s177[10],s178[10],s179[10],s180[10],s181[10],s182[10],s183[10],s184[10],s185[10],s186[10],s186[11],s186[12],s186[13],s186[14],s186[15],s186[16],s186[17],s186[18],s186[19],s186[20],s186[21],s186[22],s186[23],s186[24],s186[25],s186[26],s186[27],s186[28],s186[29],s186[30],s186[31],s186[32],s186[33],s186[34],s186[35],s186[36],s187[36],s188[36],s189[36],s190[36],s191[36],s192[36],s10[27],s11[27],s12[27],s13[27],s14[27],s15[27],s16[27],s17[27],s18[27],s19[27],s20[27],s21[27],s22[27],s23[27],s24[27],s25[27],s26[27],s27[27],s28[27],s29[27],s30[27],s31[27],s32[27],s33[27],s34[27],s35[27],s36[27],s37[27],s38[27],s39[27],s40[27],s41[27],s42[27],s43[27],s44[27],s45[27],s46[27],s47[27],s48[27],s49[27],s50[27],s51[27],s52[27],s53[27],s54[27],s55[27],s56[27],s57[27],s58[27],s59[27],s60[27],s61[27],s62[27],s63[27],s64[27],s65[27],s66[27],s67[27],s68[27],s69[27],s70[27],s71[27],s72[27],s73[27],s73[28],s73[29],s73[30],s73[31],s73[32],s73[33],s73[34],s73[35],s73[36],s73[37],s73[38],s73[39],s73[40],s73[41],s73[42],s73[43],s73[44],s73[45],s73[46],s73[47],s73[48],s73[49],s73[50],s73[51],s73[52],s73[53],s73[54],s73[55],s73[56],s71[59],s69[62],s67[65],s65[68],s64[70],s64[71],s64[72],s64[73],s64[74],s64[75],s64[76],s64[77],s64[78],s64[79],s64[80],s64[81],s64[82],s64[83],s64[84],s64[85],s64[86],s64[87],s64[88],s64[89],s64[90],s64[91],s64[92],s64[93],s64[94],s63[96],s62[98],s9[152],s7[155],s5[158],s3[161],s1[164],s65[101],s64[103],s63[105],s62[107],s61[109],s60[111],s59[113],s58[115],s57[117],s56[119],s55[121],s54[123],s53[125],s52[127],s51[129],s50[131],s49[133],s48[135],s47[137],s46[139],s45[141],s44[143],s43[145],s42[147],s41[149],s40[151],s39[153],s38[155],s37[157],s36[159],s35[161],s34[163],s33[165],s32[167],s31[169],s30[171],s29[173],s28[175],s27[177],s26[179],s25[181],s24[183],s23[185],s22[187],s21[189],s20[191],s19[193],s18[195],s17[197],s16[199],s15[201],s14[203],s13[205],s12[207],s11[209],s10[211],s218[292],s217[294],s216[296],s215[298],s214[300],s213[302],s212[304],s211[306],s210[308],s209[310],s208[312],s207[314],s206[316],s205[318],s204[320],s203[322],s202[324],s201[326],s200[328],s199[330],s198[332],s197[334],s196[336],s195[338],s194[340],s193[342],s192[248],s191[250],s190[252],s189[254],s188[256],s187[258],s186[260],s185[262],s184[264],s183[266],s182[268],s181[270],s180[272],s179[274],s178[276],s177[278],s176[280],s175[282],s174[284],s173[286],s172[288],s171[290],s170[292],s169[294],s168[296],s167[298],s166[300],s165[302],s164[304],s163[306],s162[308],s161[310],s160[312],s159[314],s158[316],s157[318],s156[320],s155[322],s154[324],s153[326],s152[328],s151[330],s150[332],s149[334],s148[336],s147[338],s146[340],s145[342],s144[344],s143[346],s142[348],s141[350],s140[352],s139[354],s138[356],s137[358],s136[360],s135[362],s134[364],s133[366],s132[368],s131[370],s130[372],s129[374],pp255[184],pp254[186],pp253[188],pp252[190],pp251[192],pp250[194],pp249[196],pp248[198],pp247[200],pp246[202],pp247[202],pp248[202],pp249[202],pp250[202],pp251[202]};
    CLA_396 KS_219(s219, c219, in219_1, in219_2);
    wire[393:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {s207[13],s206[15],s205[17],s204[19],s203[21],s204[21],s205[21],s206[21],s207[21],s208[21],s209[21],s210[21],s211[21],s212[21],s213[21],s213[22],s213[23],s213[24],s213[25],s213[26],s213[27],s213[28],s213[29],s213[30],s213[31],s213[32],s213[33],s213[34],s213[35],s213[36],s213[37],s213[38],s213[39],s213[40],s213[41],s213[42],s213[43],s213[44],s213[45],s213[46],s213[47],s211[50],s209[53],s207[56],s205[59],s203[62],s201[65],s199[68],s197[71],s195[74],s193[77],s193[78],s193[79],s193[80],s193[81],s193[82],s193[83],s193[84],s193[85],s193[86],s193[87],s193[88],s193[89],s193[90],s193[91],s193[92],s193[93],s193[94],s193[95],s193[96],s193[97],s193[98],s193[99],s187[10],s187[11],s187[12],s187[13],s187[14],s187[15],s187[16],s187[17],s187[18],s187[19],s187[20],s187[21],s187[22],s187[23],s187[24],s187[25],s187[26],s187[27],s187[28],s187[29],s187[30],s187[31],s187[32],s187[33],s187[34],s187[35],s219[100],s219[101],s219[102],s219[103],s219[104],s219[105],s219[106],s219[107],s219[108],s219[109],s219[110],s219[111],s219[112],s219[113],s219[114],s219[115],s219[116],s219[117],s219[118],s219[119],s219[120],s219[121],s219[122],s219[123],s219[124],s219[125],s219[126],s219[127],s219[128],s219[129],s219[130],s219[131],s219[132],s219[133],s219[134],s219[135],s219[136],s219[137],s219[138],s219[139],s219[140],s219[141],s219[142],s219[143],s219[144],s219[145],s219[146],s219[147],s219[148],s219[149],s219[150],s219[151],s219[152],s219[153],s219[154],s219[155],s219[156],s219[157],s219[158],s219[159],s219[160],s219[161],s219[162],s219[163],s219[164],s219[165],s219[166],s219[167],s219[168],s219[169],s219[170],s219[171],s219[172],s219[173],s219[174],s219[175],s219[176],s219[177],s219[178],s219[179],s219[180],s219[181],s219[182],s219[183],s219[184],s219[185],s219[186],s219[187],s219[188],s219[189],s219[190],s219[191],s219[192],s219[193],s219[194],s219[195],s219[196],s219[197],s219[198],s219[199],s219[200],s219[201],s219[202],s219[203],s219[204],s219[205],s219[206],s219[207],s219[208],s219[209],s219[210],s219[211],s219[212],s219[213],s219[214],s219[215],s219[216],s219[217],s219[218],s219[219],s219[220],s219[221],s219[222],s219[223],s219[224],s219[225],s219[226],s219[227],s219[228],s219[229],s219[230],s219[231],s219[232],s219[233],s219[234],s219[235],s219[236],s219[237],s219[238],s219[239],s219[240],s219[241],s219[242],s219[243],s219[244],s219[245],s219[246],s219[247],s219[248],s219[249],s219[250],s219[251],s219[252],s219[253],s219[254],s219[255],s219[256],s219[257],s219[258],s219[259],s219[260],s219[261],s219[262],s219[263],s219[264],s219[265],s219[266],s219[267],s219[268],s219[269],s219[270],s219[271],s219[272],s219[273],s219[274],s219[275],s219[276],s219[277],s219[278],s219[279],s219[280],s219[281],s219[282],s219[283],s219[284],s219[285],s219[286],s219[287],s219[288],s219[289],s219[290],s219[291],s218[293],s217[295],s216[297],s215[299],s214[301],s213[303],s212[305],s211[307],s210[309],s209[311],s208[313],s207[315],s206[317],s205[319],s204[321],s203[323],s202[325],s201[327],s200[329],s199[331],s198[333],s197[335],s196[337],s195[339],s194[341],s193[343],s192[249],s191[251],s190[253],s189[255],s188[257],s187[259],s186[261],s185[263],s184[265],s183[267],s182[269],s181[271],s180[273],s179[275],s178[277],s177[279],s176[281],s175[283],s174[285],s173[287],s172[289],s171[291],s170[293],s169[295],s168[297],s167[299],s166[301],s165[303],s164[305],s163[307],s162[309],s161[311],s160[313],s159[315],s158[317],s157[319],s156[321],s155[323],s154[325],s153[327],s152[329],s151[331],s150[333],s149[335],s148[337],s147[339],s146[341],s145[343],s144[345],s143[347],s142[349],s141[351],s140[353],s139[355],s138[357],s137[359],s136[361],s135[363],s134[365],s133[367],s132[369],s131[371],s130[373],s129[375],pp255[185],pp254[187],pp253[189],pp252[191],pp251[193],pp250[195],pp249[197],pp248[199],pp247[201],pp248[201],pp249[201],pp250[201],pp251[201]};
    assign in220_2 = {s208[12],s207[14],s206[16],s205[18],s204[20],s205[20],s206[20],s207[20],s208[20],s209[20],s210[20],s211[20],s212[20],s213[20],s214[20],s214[21],s214[22],s214[23],s214[24],s214[25],s214[26],s214[27],s214[28],s214[29],s214[30],s214[31],s214[32],s214[33],s214[34],s214[35],s214[36],s214[37],s214[38],s214[39],s214[40],s214[41],s214[42],s214[43],s214[44],s214[45],s214[46],s212[49],s210[52],s208[55],s206[58],s204[61],s202[64],s200[67],s198[70],s196[73],s194[76],s194[77],s194[78],s194[79],s194[80],s194[81],s194[82],s194[83],s194[84],s194[85],s194[86],s194[87],s194[88],s194[89],s194[90],s194[91],s194[92],s194[93],s194[94],s194[95],s194[96],s194[97],s194[98],s194[99],s188[10],s188[11],s188[12],s188[13],s188[14],s188[15],s188[16],s188[17],s188[18],s188[19],s188[20],s188[21],s188[22],s188[23],s188[24],s188[25],s188[26],s188[27],s188[28],s188[29],s188[30],s188[31],s188[32],s188[33],s188[34],s188[35],s189[35],s190[35],s191[35],s192[35],s10[26],s11[26],s12[26],s13[26],s14[26],s15[26],s16[26],s17[26],s18[26],s19[26],s20[26],s21[26],s22[26],s23[26],s24[26],s25[26],s26[26],s27[26],s28[26],s29[26],s30[26],s31[26],s32[26],s33[26],s34[26],s35[26],s36[26],s37[26],s38[26],s39[26],s40[26],s41[26],s42[26],s43[26],s44[26],s45[26],s46[26],s47[26],s48[26],s49[26],s50[26],s51[26],s52[26],s53[26],s54[26],s55[26],s56[26],s57[26],s58[26],s59[26],s60[26],s61[26],s62[26],s63[26],s64[26],s65[26],s66[26],s67[26],s68[26],s69[26],s70[26],s71[26],s72[26],s73[26],s74[26],s74[27],s74[28],s74[29],s74[30],s74[31],s74[32],s74[33],s74[34],s74[35],s74[36],s74[37],s74[38],s74[39],s74[40],s74[41],s74[42],s74[43],s74[44],s74[45],s74[46],s74[47],s74[48],s74[49],s74[50],s74[51],s74[52],s74[53],s74[54],s74[55],s72[58],s70[61],s68[64],s66[67],s65[69],s65[70],s65[71],s65[72],s65[73],s65[74],s65[75],s65[76],s65[77],s65[78],s65[79],s65[80],s65[81],s65[82],s65[83],s65[84],s65[85],s65[86],s65[87],s65[88],s65[89],s65[90],s65[91],s65[92],s65[93],s64[95],s63[97],s62[99],s8[154],s6[157],s4[160],s2[163],s66[100],s65[102],s64[104],s63[106],s62[108],s61[110],s60[112],s59[114],s58[116],s57[118],s56[120],s55[122],s54[124],s53[126],s52[128],s51[130],s50[132],s49[134],s48[136],s47[138],s46[140],s45[142],s44[144],s43[146],s42[148],s41[150],s40[152],s39[154],s38[156],s37[158],s36[160],s35[162],s34[164],s33[166],s32[168],s31[170],s30[172],s29[174],s28[176],s27[178],s26[180],s25[182],s24[184],s23[186],s22[188],s21[190],s20[192],s19[194],s18[196],s17[198],s16[200],s15[202],s14[204],s13[206],s12[208],s11[210],s10[212],s219[292],s218[294],s217[296],s216[298],s215[300],s214[302],s213[304],s212[306],s211[308],s210[310],s209[312],s208[314],s207[316],s206[318],s205[320],s204[322],s203[324],s202[326],s201[328],s200[330],s199[332],s198[334],s197[336],s196[338],s195[340],s194[342],s193[344],s192[250],s191[252],s190[254],s189[256],s188[258],s187[260],s186[262],s185[264],s184[266],s183[268],s182[270],s181[272],s180[274],s179[276],s178[278],s177[280],s176[282],s175[284],s174[286],s173[288],s172[290],s171[292],s170[294],s169[296],s168[298],s167[300],s166[302],s165[304],s164[306],s163[308],s162[310],s161[312],s160[314],s159[316],s158[318],s157[320],s156[322],s155[324],s154[326],s153[328],s152[330],s151[332],s150[334],s149[336],s148[338],s147[340],s146[342],s145[344],s144[346],s143[348],s142[350],s141[352],s140[354],s139[356],s138[358],s137[360],s136[362],s135[364],s134[366],s133[368],s132[370],s131[372],s130[374],s129[376],pp255[186],pp254[188],pp253[190],pp252[192],pp251[194],pp250[196],pp249[198],pp248[200],pp249[200],pp250[200],pp251[200],pp252[200]};
    CLA_394 KS_220(s220, c220, in220_1, in220_2);
    wire[391:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {s208[13],s207[15],s206[17],s205[19],s206[19],s207[19],s208[19],s209[19],s210[19],s211[19],s212[19],s213[19],s214[19],s215[19],s215[20],s215[21],s215[22],s215[23],s215[24],s215[25],s215[26],s215[27],s215[28],s215[29],s215[30],s215[31],s215[32],s215[33],s215[34],s215[35],s215[36],s215[37],s215[38],s215[39],s215[40],s215[41],s215[42],s215[43],s215[44],s215[45],s213[48],s211[51],s209[54],s207[57],s205[60],s203[63],s201[66],s199[69],s197[72],s195[75],s195[76],s195[77],s195[78],s195[79],s195[80],s195[81],s195[82],s195[83],s195[84],s195[85],s195[86],s195[87],s195[88],s195[89],s195[90],s195[91],s195[92],s195[93],s195[94],s195[95],s195[96],s195[97],s195[98],s195[99],s189[10],s189[11],s189[12],s189[13],s189[14],s189[15],s189[16],s189[17],s189[18],s189[19],s189[20],s189[21],s189[22],s189[23],s189[24],s189[25],s189[26],s189[27],s189[28],s189[29],s189[30],s189[31],s189[32],s189[33],s189[34],s220[100],s220[101],s220[102],s220[103],s220[104],s220[105],s220[106],s220[107],s220[108],s220[109],s220[110],s220[111],s220[112],s220[113],s220[114],s220[115],s220[116],s220[117],s220[118],s220[119],s220[120],s220[121],s220[122],s220[123],s220[124],s220[125],s220[126],s220[127],s220[128],s220[129],s220[130],s220[131],s220[132],s220[133],s220[134],s220[135],s220[136],s220[137],s220[138],s220[139],s220[140],s220[141],s220[142],s220[143],s220[144],s220[145],s220[146],s220[147],s220[148],s220[149],s220[150],s220[151],s220[152],s220[153],s220[154],s220[155],s220[156],s220[157],s220[158],s220[159],s220[160],s220[161],s220[162],s220[163],s220[164],s220[165],s220[166],s220[167],s220[168],s220[169],s220[170],s220[171],s220[172],s220[173],s220[174],s220[175],s220[176],s220[177],s220[178],s220[179],s220[180],s220[181],s220[182],s220[183],s220[184],s220[185],s220[186],s220[187],s220[188],s220[189],s220[190],s220[191],s220[192],s220[193],s220[194],s220[195],s220[196],s220[197],s220[198],s220[199],s220[200],s220[201],s220[202],s220[203],s220[204],s220[205],s220[206],s220[207],s220[208],s220[209],s220[210],s220[211],s220[212],s220[213],s220[214],s220[215],s220[216],s220[217],s220[218],s220[219],s220[220],s220[221],s220[222],s220[223],s220[224],s220[225],s220[226],s220[227],s220[228],s220[229],s220[230],s220[231],s220[232],s220[233],s220[234],s220[235],s220[236],s220[237],s220[238],s220[239],s220[240],s220[241],s220[242],s220[243],s220[244],s220[245],s220[246],s220[247],s220[248],s220[249],s220[250],s220[251],s220[252],s220[253],s220[254],s220[255],s220[256],s220[257],s220[258],s220[259],s220[260],s220[261],s220[262],s220[263],s220[264],s220[265],s220[266],s220[267],s220[268],s220[269],s220[270],s220[271],s220[272],s220[273],s220[274],s220[275],s220[276],s220[277],s220[278],s220[279],s220[280],s220[281],s220[282],s220[283],s220[284],s220[285],s220[286],s220[287],s220[288],s220[289],s220[290],s220[291],s219[293],s218[295],s217[297],s216[299],s215[301],s214[303],s213[305],s212[307],s211[309],s210[311],s209[313],s208[315],s207[317],s206[319],s205[321],s204[323],s203[325],s202[327],s201[329],s200[331],s199[333],s198[335],s197[337],s196[339],s195[341],s194[343],s193[345],s192[251],s191[253],s190[255],s189[257],s188[259],s187[261],s186[263],s185[265],s184[267],s183[269],s182[271],s181[273],s180[275],s179[277],s178[279],s177[281],s176[283],s175[285],s174[287],s173[289],s172[291],s171[293],s170[295],s169[297],s168[299],s167[301],s166[303],s165[305],s164[307],s163[309],s162[311],s161[313],s160[315],s159[317],s158[319],s157[321],s156[323],s155[325],s154[327],s153[329],s152[331],s151[333],s150[335],s149[337],s148[339],s147[341],s146[343],s145[345],s144[347],s143[349],s142[351],s141[353],s140[355],s139[357],s138[359],s137[361],s136[363],s135[365],s134[367],s133[369],s132[371],s131[373],s130[375],s129[377],pp255[187],pp254[189],pp253[191],pp252[193],pp251[195],pp250[197],pp249[199],pp250[199],pp251[199],pp252[199]};
    assign in221_2 = {s209[12],s208[14],s207[16],s206[18],s207[18],s208[18],s209[18],s210[18],s211[18],s212[18],s213[18],s214[18],s215[18],s216[18],s216[19],s216[20],s216[21],s216[22],s216[23],s216[24],s216[25],s216[26],s216[27],s216[28],s216[29],s216[30],s216[31],s216[32],s216[33],s216[34],s216[35],s216[36],s216[37],s216[38],s216[39],s216[40],s216[41],s216[42],s216[43],s216[44],s214[47],s212[50],s210[53],s208[56],s206[59],s204[62],s202[65],s200[68],s198[71],s196[74],s196[75],s196[76],s196[77],s196[78],s196[79],s196[80],s196[81],s196[82],s196[83],s196[84],s196[85],s196[86],s196[87],s196[88],s196[89],s196[90],s196[91],s196[92],s196[93],s196[94],s196[95],s196[96],s196[97],s196[98],s196[99],s190[10],s190[11],s190[12],s190[13],s190[14],s190[15],s190[16],s190[17],s190[18],s190[19],s190[20],s190[21],s190[22],s190[23],s190[24],s190[25],s190[26],s190[27],s190[28],s190[29],s190[30],s190[31],s190[32],s190[33],s190[34],s191[34],s192[34],s10[25],s11[25],s12[25],s13[25],s14[25],s15[25],s16[25],s17[25],s18[25],s19[25],s20[25],s21[25],s22[25],s23[25],s24[25],s25[25],s26[25],s27[25],s28[25],s29[25],s30[25],s31[25],s32[25],s33[25],s34[25],s35[25],s36[25],s37[25],s38[25],s39[25],s40[25],s41[25],s42[25],s43[25],s44[25],s45[25],s46[25],s47[25],s48[25],s49[25],s50[25],s51[25],s52[25],s53[25],s54[25],s55[25],s56[25],s57[25],s58[25],s59[25],s60[25],s61[25],s62[25],s63[25],s64[25],s65[25],s66[25],s67[25],s68[25],s69[25],s70[25],s71[25],s72[25],s73[25],s74[25],s75[25],s75[26],s75[27],s75[28],s75[29],s75[30],s75[31],s75[32],s75[33],s75[34],s75[35],s75[36],s75[37],s75[38],s75[39],s75[40],s75[41],s75[42],s75[43],s75[44],s75[45],s75[46],s75[47],s75[48],s75[49],s75[50],s75[51],s75[52],s75[53],s75[54],s73[57],s71[60],s69[63],s67[66],s66[68],s66[69],s66[70],s66[71],s66[72],s66[73],s66[74],s66[75],s66[76],s66[77],s66[78],s66[79],s66[80],s66[81],s66[82],s66[83],s66[84],s66[85],s66[86],s66[87],s66[88],s66[89],s66[90],s66[91],s66[92],s65[94],s64[96],s63[98],s9[153],s7[156],s5[159],s3[162],s1[165],s66[101],s65[103],s64[105],s63[107],s62[109],s61[111],s60[113],s59[115],s58[117],s57[119],s56[121],s55[123],s54[125],s53[127],s52[129],s51[131],s50[133],s49[135],s48[137],s47[139],s46[141],s45[143],s44[145],s43[147],s42[149],s41[151],s40[153],s39[155],s38[157],s37[159],s36[161],s35[163],s34[165],s33[167],s32[169],s31[171],s30[173],s29[175],s28[177],s27[179],s26[181],s25[183],s24[185],s23[187],s22[189],s21[191],s20[193],s19[195],s18[197],s17[199],s16[201],s15[203],s14[205],s13[207],s12[209],s11[211],s10[213],s220[292],s219[294],s218[296],s217[298],s216[300],s215[302],s214[304],s213[306],s212[308],s211[310],s210[312],s209[314],s208[316],s207[318],s206[320],s205[322],s204[324],s203[326],s202[328],s201[330],s200[332],s199[334],s198[336],s197[338],s196[340],s195[342],s194[344],s193[346],s192[252],s191[254],s190[256],s189[258],s188[260],s187[262],s186[264],s185[266],s184[268],s183[270],s182[272],s181[274],s180[276],s179[278],s178[280],s177[282],s176[284],s175[286],s174[288],s173[290],s172[292],s171[294],s170[296],s169[298],s168[300],s167[302],s166[304],s165[306],s164[308],s163[310],s162[312],s161[314],s160[316],s159[318],s158[320],s157[322],s156[324],s155[326],s154[328],s153[330],s152[332],s151[334],s150[336],s149[338],s148[340],s147[342],s146[344],s145[346],s144[348],s143[350],s142[352],s141[354],s140[356],s139[358],s138[360],s137[362],s136[364],s135[366],s134[368],s133[370],s132[372],s131[374],s130[376],s129[378],pp255[188],pp254[190],pp253[192],pp252[194],pp251[196],pp250[198],pp251[198],pp252[198],pp253[198]};
    CLA_392 KS_221(s221, c221, in221_1, in221_2);
    wire[389:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {s209[13],s208[15],s207[17],s208[17],s209[17],s210[17],s211[17],s212[17],s213[17],s214[17],s215[17],s216[17],s217[17],s217[18],s217[19],s217[20],s217[21],s217[22],s217[23],s217[24],s217[25],s217[26],s217[27],s217[28],s217[29],s217[30],s217[31],s217[32],s217[33],s217[34],s217[35],s217[36],s217[37],s217[38],s217[39],s217[40],s217[41],s217[42],s217[43],s215[46],s213[49],s211[52],s209[55],s207[58],s205[61],s203[64],s201[67],s199[70],s197[73],s197[74],s197[75],s197[76],s197[77],s197[78],s197[79],s197[80],s197[81],s197[82],s197[83],s197[84],s197[85],s197[86],s197[87],s197[88],s197[89],s197[90],s197[91],s197[92],s197[93],s197[94],s197[95],s197[96],s197[97],s197[98],s197[99],s191[10],s191[11],s191[12],s191[13],s191[14],s191[15],s191[16],s191[17],s191[18],s191[19],s191[20],s191[21],s191[22],s191[23],s191[24],s191[25],s191[26],s191[27],s191[28],s191[29],s191[30],s191[31],s191[32],s191[33],s221[100],s221[101],s221[102],s221[103],s221[104],s221[105],s221[106],s221[107],s221[108],s221[109],s221[110],s221[111],s221[112],s221[113],s221[114],s221[115],s221[116],s221[117],s221[118],s221[119],s221[120],s221[121],s221[122],s221[123],s221[124],s221[125],s221[126],s221[127],s221[128],s221[129],s221[130],s221[131],s221[132],s221[133],s221[134],s221[135],s221[136],s221[137],s221[138],s221[139],s221[140],s221[141],s221[142],s221[143],s221[144],s221[145],s221[146],s221[147],s221[148],s221[149],s221[150],s221[151],s221[152],s221[153],s221[154],s221[155],s221[156],s221[157],s221[158],s221[159],s221[160],s221[161],s221[162],s221[163],s221[164],s221[165],s221[166],s221[167],s221[168],s221[169],s221[170],s221[171],s221[172],s221[173],s221[174],s221[175],s221[176],s221[177],s221[178],s221[179],s221[180],s221[181],s221[182],s221[183],s221[184],s221[185],s221[186],s221[187],s221[188],s221[189],s221[190],s221[191],s221[192],s221[193],s221[194],s221[195],s221[196],s221[197],s221[198],s221[199],s221[200],s221[201],s221[202],s221[203],s221[204],s221[205],s221[206],s221[207],s221[208],s221[209],s221[210],s221[211],s221[212],s221[213],s221[214],s221[215],s221[216],s221[217],s221[218],s221[219],s221[220],s221[221],s221[222],s221[223],s221[224],s221[225],s221[226],s221[227],s221[228],s221[229],s221[230],s221[231],s221[232],s221[233],s221[234],s221[235],s221[236],s221[237],s221[238],s221[239],s221[240],s221[241],s221[242],s221[243],s221[244],s221[245],s221[246],s221[247],s221[248],s221[249],s221[250],s221[251],s221[252],s221[253],s221[254],s221[255],s221[256],s221[257],s221[258],s221[259],s221[260],s221[261],s221[262],s221[263],s221[264],s221[265],s221[266],s221[267],s221[268],s221[269],s221[270],s221[271],s221[272],s221[273],s221[274],s221[275],s221[276],s221[277],s221[278],s221[279],s221[280],s221[281],s221[282],s221[283],s221[284],s221[285],s221[286],s221[287],s221[288],s221[289],s221[290],s221[291],s220[293],s219[295],s218[297],s217[299],s216[301],s215[303],s214[305],s213[307],s212[309],s211[311],s210[313],s209[315],s208[317],s207[319],s206[321],s205[323],s204[325],s203[327],s202[329],s201[331],s200[333],s199[335],s198[337],s197[339],s196[341],s195[343],s194[345],s193[347],s192[253],s191[255],s190[257],s189[259],s188[261],s187[263],s186[265],s185[267],s184[269],s183[271],s182[273],s181[275],s180[277],s179[279],s178[281],s177[283],s176[285],s175[287],s174[289],s173[291],s172[293],s171[295],s170[297],s169[299],s168[301],s167[303],s166[305],s165[307],s164[309],s163[311],s162[313],s161[315],s160[317],s159[319],s158[321],s157[323],s156[325],s155[327],s154[329],s153[331],s152[333],s151[335],s150[337],s149[339],s148[341],s147[343],s146[345],s145[347],s144[349],s143[351],s142[353],s141[355],s140[357],s139[359],s138[361],s137[363],s136[365],s135[367],s134[369],s133[371],s132[373],s131[375],s130[377],s129[379],pp255[189],pp254[191],pp253[193],pp252[195],pp251[197],pp252[197],pp253[197]};
    assign in222_2 = {s210[12],s209[14],s208[16],s209[16],s210[16],s211[16],s212[16],s213[16],s214[16],s215[16],s216[16],s217[16],s218[16],s218[17],s218[18],s218[19],s218[20],s218[21],s218[22],s218[23],s218[24],s218[25],s218[26],s218[27],s218[28],s218[29],s218[30],s218[31],s218[32],s218[33],s218[34],s218[35],s218[36],s218[37],s218[38],s218[39],s218[40],s218[41],s218[42],s216[45],s214[48],s212[51],s210[54],s208[57],s206[60],s204[63],s202[66],s200[69],s198[72],s198[73],s198[74],s198[75],s198[76],s198[77],s198[78],s198[79],s198[80],s198[81],s198[82],s198[83],s198[84],s198[85],s198[86],s198[87],s198[88],s198[89],s198[90],s198[91],s198[92],s198[93],s198[94],s198[95],s198[96],s198[97],s198[98],s198[99],s192[10],s192[11],s192[12],s192[13],s192[14],s192[15],s192[16],s192[17],s192[18],s192[19],s192[20],s192[21],s192[22],s192[23],s192[24],s192[25],s192[26],s192[27],s192[28],s192[29],s192[30],s192[31],s192[32],s192[33],s10[24],s11[24],s12[24],s13[24],s14[24],s15[24],s16[24],s17[24],s18[24],s19[24],s20[24],s21[24],s22[24],s23[24],s24[24],s25[24],s26[24],s27[24],s28[24],s29[24],s30[24],s31[24],s32[24],s33[24],s34[24],s35[24],s36[24],s37[24],s38[24],s39[24],s40[24],s41[24],s42[24],s43[24],s44[24],s45[24],s46[24],s47[24],s48[24],s49[24],s50[24],s51[24],s52[24],s53[24],s54[24],s55[24],s56[24],s57[24],s58[24],s59[24],s60[24],s61[24],s62[24],s63[24],s64[24],s65[24],s66[24],s67[24],s68[24],s69[24],s70[24],s71[24],s72[24],s73[24],s74[24],s75[24],s76[24],s76[25],s76[26],s76[27],s76[28],s76[29],s76[30],s76[31],s76[32],s76[33],s76[34],s76[35],s76[36],s76[37],s76[38],s76[39],s76[40],s76[41],s76[42],s76[43],s76[44],s76[45],s76[46],s76[47],s76[48],s76[49],s76[50],s76[51],s76[52],s76[53],s74[56],s72[59],s70[62],s68[65],s67[67],s67[68],s67[69],s67[70],s67[71],s67[72],s67[73],s67[74],s67[75],s67[76],s67[77],s67[78],s67[79],s67[80],s67[81],s67[82],s67[83],s67[84],s67[85],s67[86],s67[87],s67[88],s67[89],s67[90],s67[91],s66[93],s65[95],s64[97],s63[99],s8[155],s6[158],s4[161],s2[164],s67[100],s66[102],s65[104],s64[106],s63[108],s62[110],s61[112],s60[114],s59[116],s58[118],s57[120],s56[122],s55[124],s54[126],s53[128],s52[130],s51[132],s50[134],s49[136],s48[138],s47[140],s46[142],s45[144],s44[146],s43[148],s42[150],s41[152],s40[154],s39[156],s38[158],s37[160],s36[162],s35[164],s34[166],s33[168],s32[170],s31[172],s30[174],s29[176],s28[178],s27[180],s26[182],s25[184],s24[186],s23[188],s22[190],s21[192],s20[194],s19[196],s18[198],s17[200],s16[202],s15[204],s14[206],s13[208],s12[210],s11[212],s10[214],s221[292],s220[294],s219[296],s218[298],s217[300],s216[302],s215[304],s214[306],s213[308],s212[310],s211[312],s210[314],s209[316],s208[318],s207[320],s206[322],s205[324],s204[326],s203[328],s202[330],s201[332],s200[334],s199[336],s198[338],s197[340],s196[342],s195[344],s194[346],s193[348],s192[254],s191[256],s190[258],s189[260],s188[262],s187[264],s186[266],s185[268],s184[270],s183[272],s182[274],s181[276],s180[278],s179[280],s178[282],s177[284],s176[286],s175[288],s174[290],s173[292],s172[294],s171[296],s170[298],s169[300],s168[302],s167[304],s166[306],s165[308],s164[310],s163[312],s162[314],s161[316],s160[318],s159[320],s158[322],s157[324],s156[326],s155[328],s154[330],s153[332],s152[334],s151[336],s150[338],s149[340],s148[342],s147[344],s146[346],s145[348],s144[350],s143[352],s142[354],s141[356],s140[358],s139[360],s138[362],s137[364],s136[366],s135[368],s134[370],s133[372],s132[374],s131[376],s130[378],s129[380],pp255[190],pp254[192],pp253[194],pp252[196],pp253[196],pp254[196]};
    CLA_390 KS_222(s222, c222, in222_1, in222_2);
    wire[387:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {s210[13],s209[15],s210[15],s211[15],s212[15],s213[15],s214[15],s215[15],s216[15],s217[15],s218[15],s219[15],s219[16],s219[17],s219[18],s219[19],s219[20],s219[21],s219[22],s219[23],s219[24],s219[25],s219[26],s219[27],s219[28],s219[29],s219[30],s219[31],s219[32],s219[33],s219[34],s219[35],s219[36],s219[37],s219[38],s219[39],s219[40],s219[41],s217[44],s215[47],s213[50],s211[53],s209[56],s207[59],s205[62],s203[65],s201[68],s199[71],s199[72],s199[73],s199[74],s199[75],s199[76],s199[77],s199[78],s199[79],s199[80],s199[81],s199[82],s199[83],s199[84],s199[85],s199[86],s199[87],s199[88],s199[89],s199[90],s199[91],s199[92],s199[93],s199[94],s199[95],s199[96],s199[97],s199[98],s199[99],s200[99],s201[99],s202[99],s203[99],s204[99],s205[99],s206[99],s207[99],s208[99],s209[99],s210[99],s211[99],s212[99],s213[99],s214[99],s215[99],s216[99],s217[99],s218[99],s219[99],s220[99],s221[99],s222[99],s222[100],s222[101],s222[102],s222[103],s222[104],s222[105],s222[106],s222[107],s222[108],s222[109],s222[110],s222[111],s222[112],s222[113],s222[114],s222[115],s222[116],s222[117],s222[118],s222[119],s222[120],s222[121],s222[122],s222[123],s222[124],s222[125],s222[126],s222[127],s222[128],s222[129],s222[130],s222[131],s222[132],s222[133],s222[134],s222[135],s222[136],s222[137],s222[138],s222[139],s222[140],s222[141],s222[142],s222[143],s222[144],s222[145],s222[146],s222[147],s222[148],s222[149],s222[150],s222[151],s222[152],s222[153],s222[154],s222[155],s222[156],s222[157],s222[158],s222[159],s222[160],s222[161],s222[162],s222[163],s222[164],s222[165],s222[166],s222[167],s222[168],s222[169],s222[170],s222[171],s222[172],s222[173],s222[174],s222[175],s222[176],s222[177],s222[178],s222[179],s222[180],s222[181],s222[182],s222[183],s222[184],s222[185],s222[186],s222[187],s222[188],s222[189],s222[190],s222[191],s222[192],s222[193],s222[194],s222[195],s222[196],s222[197],s222[198],s222[199],s222[200],s222[201],s222[202],s222[203],s222[204],s222[205],s222[206],s222[207],s222[208],s222[209],s222[210],s222[211],s222[212],s222[213],s222[214],s222[215],s222[216],s222[217],s222[218],s222[219],s222[220],s222[221],s222[222],s222[223],s222[224],s222[225],s222[226],s222[227],s222[228],s222[229],s222[230],s222[231],s222[232],s222[233],s222[234],s222[235],s222[236],s222[237],s222[238],s222[239],s222[240],s222[241],s222[242],s222[243],s222[244],s222[245],s222[246],s222[247],s222[248],s222[249],s222[250],s222[251],s222[252],s222[253],s222[254],s222[255],s222[256],s222[257],s222[258],s222[259],s222[260],s222[261],s222[262],s222[263],s222[264],s222[265],s222[266],s222[267],s222[268],s222[269],s222[270],s222[271],s222[272],s222[273],s222[274],s222[275],s222[276],s222[277],s222[278],s222[279],s222[280],s222[281],s222[282],s222[283],s222[284],s222[285],s222[286],s222[287],s222[288],s222[289],s222[290],s222[291],s221[293],s220[295],s219[297],s218[299],s217[301],s216[303],s215[305],s214[307],s213[309],s212[311],s211[313],s210[315],s209[317],s208[319],s207[321],s206[323],s205[325],s204[327],s203[329],s202[331],s201[333],s200[335],s199[337],s198[339],s197[341],s196[343],s195[345],s194[347],s193[349],s192[255],s191[257],s190[259],s189[261],s188[263],s187[265],s186[267],s185[269],s184[271],s183[273],s182[275],s181[277],s180[279],s179[281],s178[283],s177[285],s176[287],s175[289],s174[291],s173[293],s172[295],s171[297],s170[299],s169[301],s168[303],s167[305],s166[307],s165[309],s164[311],s163[313],s162[315],s161[317],s160[319],s159[321],s158[323],s157[325],s156[327],s155[329],s154[331],s153[333],s152[335],s151[337],s150[339],s149[341],s148[343],s147[345],s146[347],s145[349],s144[351],s143[353],s142[355],s141[357],s140[359],s139[361],s138[363],s137[365],s136[367],s135[369],s134[371],s133[373],s132[375],s131[377],s130[379],s129[381],pp255[191],pp254[193],pp253[195],pp254[195]};
    assign in223_2 = {s211[12],s210[14],s211[14],s212[14],s213[14],s214[14],s215[14],s216[14],s217[14],s218[14],s219[14],s220[14],s220[15],s220[16],s220[17],s220[18],s220[19],s220[20],s220[21],s220[22],s220[23],s220[24],s220[25],s220[26],s220[27],s220[28],s220[29],s220[30],s220[31],s220[32],s220[33],s220[34],s220[35],s220[36],s220[37],s220[38],s220[39],s220[40],s218[43],s216[46],s214[49],s212[52],s210[55],s208[58],s206[61],s204[64],s202[67],s200[70],s200[71],s200[72],s200[73],s200[74],s200[75],s200[76],s200[77],s200[78],s200[79],s200[80],s200[81],s200[82],s200[83],s200[84],s200[85],s200[86],s200[87],s200[88],s200[89],s200[90],s200[91],s200[92],s200[93],s200[94],s200[95],s200[96],s200[97],s200[98],s201[98],s202[98],s203[98],s204[98],s205[98],s206[98],s207[98],s208[98],s209[98],s210[98],s211[98],s212[98],s213[98],s214[98],s215[98],s216[98],s217[98],s218[98],s219[98],s220[98],s221[98],s222[98],s10[23],s11[23],s12[23],s13[23],s14[23],s15[23],s16[23],s17[23],s18[23],s19[23],s20[23],s21[23],s22[23],s23[23],s24[23],s25[23],s26[23],s27[23],s28[23],s29[23],s30[23],s31[23],s32[23],s33[23],s34[23],s35[23],s36[23],s37[23],s38[23],s39[23],s40[23],s41[23],s42[23],s43[23],s44[23],s45[23],s46[23],s47[23],s48[23],s49[23],s50[23],s51[23],s52[23],s53[23],s54[23],s55[23],s56[23],s57[23],s58[23],s59[23],s60[23],s61[23],s62[23],s63[23],s64[23],s65[23],s66[23],s67[23],s68[23],s69[23],s70[23],s71[23],s72[23],s73[23],s74[23],s75[23],s76[23],s77[23],s77[24],s77[25],s77[26],s77[27],s77[28],s77[29],s77[30],s77[31],s77[32],s77[33],s77[34],s77[35],s77[36],s77[37],s77[38],s77[39],s77[40],s77[41],s77[42],s77[43],s77[44],s77[45],s77[46],s77[47],s77[48],s77[49],s77[50],s77[51],s77[52],s75[55],s73[58],s71[61],s69[64],s68[66],s68[67],s68[68],s68[69],s68[70],s68[71],s68[72],s68[73],s68[74],s68[75],s68[76],s68[77],s68[78],s68[79],s68[80],s68[81],s68[82],s68[83],s68[84],s68[85],s68[86],s68[87],s68[88],s68[89],s68[90],s67[92],s66[94],s65[96],s64[98],s9[154],s7[157],s5[160],s3[163],s1[166],s67[101],s66[103],s65[105],s64[107],s63[109],s62[111],s61[113],s60[115],s59[117],s58[119],s57[121],s56[123],s55[125],s54[127],s53[129],s52[131],s51[133],s50[135],s49[137],s48[139],s47[141],s46[143],s45[145],s44[147],s43[149],s42[151],s41[153],s40[155],s39[157],s38[159],s37[161],s36[163],s35[165],s34[167],s33[169],s32[171],s31[173],s30[175],s29[177],s28[179],s27[181],s26[183],s25[185],s24[187],s23[189],s22[191],s21[193],s20[195],s19[197],s18[199],s17[201],s16[203],s15[205],s14[207],s13[209],s12[211],s11[213],s10[215],s222[292],s221[294],s220[296],s219[298],s218[300],s217[302],s216[304],s215[306],s214[308],s213[310],s212[312],s211[314],s210[316],s209[318],s208[320],s207[322],s206[324],s205[326],s204[328],s203[330],s202[332],s201[334],s200[336],s199[338],s198[340],s197[342],s196[344],s195[346],s194[348],s193[350],s192[256],s191[258],s190[260],s189[262],s188[264],s187[266],s186[268],s185[270],s184[272],s183[274],s182[276],s181[278],s180[280],s179[282],s178[284],s177[286],s176[288],s175[290],s174[292],s173[294],s172[296],s171[298],s170[300],s169[302],s168[304],s167[306],s166[308],s165[310],s164[312],s163[314],s162[316],s161[318],s160[320],s159[322],s158[324],s157[326],s156[328],s155[330],s154[332],s153[334],s152[336],s151[338],s150[340],s149[342],s148[344],s147[346],s146[348],s145[350],s144[352],s143[354],s142[356],s141[358],s140[360],s139[362],s138[364],s137[366],s136[368],s135[370],s134[372],s133[374],s132[376],s131[378],s130[380],s129[382],pp255[192],pp254[194],pp255[194]};
    CLA_388 KS_223(s223, c223, in223_1, in223_2);
    wire[385:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {s211[13],s212[13],s213[13],s214[13],s215[13],s216[13],s217[13],s218[13],s219[13],s220[13],s221[13],s221[14],s221[15],s221[16],s221[17],s221[18],s221[19],s221[20],s221[21],s221[22],s221[23],s221[24],s221[25],s221[26],s221[27],s221[28],s221[29],s221[30],s221[31],s221[32],s221[33],s221[34],s221[35],s221[36],s221[37],s221[38],s221[39],s219[42],s217[45],s215[48],s213[51],s211[54],s209[57],s207[60],s205[63],s203[66],s201[69],s201[70],s201[71],s201[72],s201[73],s201[74],s201[75],s201[76],s201[77],s201[78],s201[79],s201[80],s201[81],s201[82],s201[83],s201[84],s201[85],s201[86],s201[87],s201[88],s201[89],s201[90],s201[91],s201[92],s201[93],s201[94],s201[95],s201[96],s201[97],s202[97],s203[97],s204[97],s205[97],s206[97],s207[97],s208[97],s209[97],s210[97],s211[97],s212[97],s213[97],s214[97],s215[97],s216[97],s217[97],s218[97],s219[97],s220[97],s221[97],s222[97],s223[97],s223[98],s223[99],s223[100],s223[101],s223[102],s223[103],s223[104],s223[105],s223[106],s223[107],s223[108],s223[109],s223[110],s223[111],s223[112],s223[113],s223[114],s223[115],s223[116],s223[117],s223[118],s223[119],s223[120],s223[121],s223[122],s223[123],s223[124],s223[125],s223[126],s223[127],s223[128],s223[129],s223[130],s223[131],s223[132],s223[133],s223[134],s223[135],s223[136],s223[137],s223[138],s223[139],s223[140],s223[141],s223[142],s223[143],s223[144],s223[145],s223[146],s223[147],s223[148],s223[149],s223[150],s223[151],s223[152],s223[153],s223[154],s223[155],s223[156],s223[157],s223[158],s223[159],s223[160],s223[161],s223[162],s223[163],s223[164],s223[165],s223[166],s223[167],s223[168],s223[169],s223[170],s223[171],s223[172],s223[173],s223[174],s223[175],s223[176],s223[177],s223[178],s223[179],s223[180],s223[181],s223[182],s223[183],s223[184],s223[185],s223[186],s223[187],s223[188],s223[189],s223[190],s223[191],s223[192],s223[193],s223[194],s223[195],s223[196],s223[197],s223[198],s223[199],s223[200],s223[201],s223[202],s223[203],s223[204],s223[205],s223[206],s223[207],s223[208],s223[209],s223[210],s223[211],s223[212],s223[213],s223[214],s223[215],s223[216],s223[217],s223[218],s223[219],s223[220],s223[221],s223[222],s223[223],s223[224],s223[225],s223[226],s223[227],s223[228],s223[229],s223[230],s223[231],s223[232],s223[233],s223[234],s223[235],s223[236],s223[237],s223[238],s223[239],s223[240],s223[241],s223[242],s223[243],s223[244],s223[245],s223[246],s223[247],s223[248],s223[249],s223[250],s223[251],s223[252],s223[253],s223[254],s223[255],s223[256],s223[257],s223[258],s223[259],s223[260],s223[261],s223[262],s223[263],s223[264],s223[265],s223[266],s223[267],s223[268],s223[269],s223[270],s223[271],s223[272],s223[273],s223[274],s223[275],s223[276],s223[277],s223[278],s223[279],s223[280],s223[281],s223[282],s223[283],s223[284],s223[285],s223[286],s223[287],s223[288],s223[289],s223[290],s223[291],s222[293],s221[295],s220[297],s219[299],s218[301],s217[303],s216[305],s215[307],s214[309],s213[311],s212[313],s211[315],s210[317],s209[319],s208[321],s207[323],s206[325],s205[327],s204[329],s203[331],s202[333],s201[335],s200[337],s199[339],s198[341],s197[343],s196[345],s195[347],s194[349],s193[351],s192[257],s191[259],s190[261],s189[263],s188[265],s187[267],s186[269],s185[271],s184[273],s183[275],s182[277],s181[279],s180[281],s179[283],s178[285],s177[287],s176[289],s175[291],s174[293],s173[295],s172[297],s171[299],s170[301],s169[303],s168[305],s167[307],s166[309],s165[311],s164[313],s163[315],s162[317],s161[319],s160[321],s159[323],s158[325],s157[327],s156[329],s155[331],s154[333],s153[335],s152[337],s151[339],s150[341],s149[343],s148[345],s147[347],s146[349],s145[351],s144[353],s143[355],s142[357],s141[359],s140[361],s139[363],s138[365],s137[367],s136[369],s135[371],s134[373],s133[375],s132[377],s131[379],s130[381],s129[383],pp255[193]};
    assign in224_2 = {s212[12],s213[12],s214[12],s215[12],s216[12],s217[12],s218[12],s219[12],s220[12],s221[12],s222[12],s222[13],s222[14],s222[15],s222[16],s222[17],s222[18],s222[19],s222[20],s222[21],s222[22],s222[23],s222[24],s222[25],s222[26],s222[27],s222[28],s222[29],s222[30],s222[31],s222[32],s222[33],s222[34],s222[35],s222[36],s222[37],s222[38],s220[41],s218[44],s216[47],s214[50],s212[53],s210[56],s208[59],s206[62],s204[65],s202[68],s202[69],s202[70],s202[71],s202[72],s202[73],s202[74],s202[75],s202[76],s202[77],s202[78],s202[79],s202[80],s202[81],s202[82],s202[83],s202[84],s202[85],s202[86],s202[87],s202[88],s202[89],s202[90],s202[91],s202[92],s202[93],s202[94],s202[95],s202[96],s203[96],s204[96],s205[96],s206[96],s207[96],s208[96],s209[96],s210[96],s211[96],s212[96],s213[96],s214[96],s215[96],s216[96],s217[96],s218[96],s219[96],s220[96],s221[96],s222[96],s223[96],s10[22],s11[22],s12[22],s13[22],s14[22],s15[22],s16[22],s17[22],s18[22],s19[22],s20[22],s21[22],s22[22],s23[22],s24[22],s25[22],s26[22],s27[22],s28[22],s29[22],s30[22],s31[22],s32[22],s33[22],s34[22],s35[22],s36[22],s37[22],s38[22],s39[22],s40[22],s41[22],s42[22],s43[22],s44[22],s45[22],s46[22],s47[22],s48[22],s49[22],s50[22],s51[22],s52[22],s53[22],s54[22],s55[22],s56[22],s57[22],s58[22],s59[22],s60[22],s61[22],s62[22],s63[22],s64[22],s65[22],s66[22],s67[22],s68[22],s69[22],s70[22],s71[22],s72[22],s73[22],s74[22],s75[22],s76[22],s77[22],s78[22],s78[23],s78[24],s78[25],s78[26],s78[27],s78[28],s78[29],s78[30],s78[31],s78[32],s78[33],s78[34],s78[35],s78[36],s78[37],s78[38],s78[39],s78[40],s78[41],s78[42],s78[43],s78[44],s78[45],s78[46],s78[47],s78[48],s78[49],s78[50],s78[51],s76[54],s74[57],s72[60],s70[63],s69[65],s69[66],s69[67],s69[68],s69[69],s69[70],s69[71],s69[72],s69[73],s69[74],s69[75],s69[76],s69[77],s69[78],s69[79],s69[80],s69[81],s69[82],s69[83],s69[84],s69[85],s69[86],s69[87],s69[88],s69[89],s68[91],s67[93],s66[95],s65[97],s64[99],s8[156],s6[159],s4[162],s2[165],s68[100],s67[102],s66[104],s65[106],s64[108],s63[110],s62[112],s61[114],s60[116],s59[118],s58[120],s57[122],s56[124],s55[126],s54[128],s53[130],s52[132],s51[134],s50[136],s49[138],s48[140],s47[142],s46[144],s45[146],s44[148],s43[150],s42[152],s41[154],s40[156],s39[158],s38[160],s37[162],s36[164],s35[166],s34[168],s33[170],s32[172],s31[174],s30[176],s29[178],s28[180],s27[182],s26[184],s25[186],s24[188],s23[190],s22[192],s21[194],s20[196],s19[198],s18[200],s17[202],s16[204],s15[206],s14[208],s13[210],s12[212],s11[214],s10[216],s223[292],s222[294],s221[296],s220[298],s219[300],s218[302],s217[304],s216[306],s215[308],s214[310],s213[312],s212[314],s211[316],s210[318],s209[320],s208[322],s207[324],s206[326],s205[328],s204[330],s203[332],s202[334],s201[336],s200[338],s199[340],s198[342],s197[344],s196[346],s195[348],s194[350],s193[352],s193[353],s193[354],s193[355],s193[356],s193[357],s193[358],s193[359],s193[360],s193[361],s193[362],s193[363],s193[364],s193[365],s193[366],s193[367],s193[368],s193[369],s193[370],s193[371],s193[372],s193[373],s193[374],s193[375],s193[376],s193[377],s193[378],s193[379],s193[380],s193[381],s193[382],s193[383],s193[384],s193[385],s193[386],s193[387],s193[388],s193[389],s193[390],s193[391],s193[392],s193[393],s193[394],s193[395],s193[396],s193[397],s193[398],s193[399],s193[400],s193[401],s193[402],s193[403],s193[404],s193[405],s193[406],s193[407],s193[408],s193[409],s193[410],s193[411],s193[412],s193[413],s193[414],s193[415],s193[416]};
    CLA_386 KS_224(s224, c224, in224_1, in224_2);

    /*Stage 4*/
    wire[479:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {pp0[16],pp0[17],pp0[18],pp0[19],pp10[10],pp10[11],pp10[12],pp10[13],pp10[14],pp10[15],pp10[16],pp10[17],pp10[18],pp10[19],pp10[20],pp10[21],pp12[20],pp14[19],pp16[18],pp18[17],pp20[16],pp22[15],pp24[14],pp26[13],pp28[12],pp30[11],pp32[10],s193[11],s194[11],s195[11],s196[11],s197[11],s198[11],s199[11],s200[11],s201[11],s202[11],s203[11],s204[11],s205[11],s206[11],s207[11],s208[11],s209[11],s210[11],s211[11],s212[11],s213[11],s214[11],s215[11],s216[11],s217[11],s218[11],s219[11],s220[11],s221[11],s222[11],s223[11],s223[12],s223[13],s223[14],s223[15],s223[16],s223[17],s223[18],s223[19],s223[20],s223[21],s223[22],s223[23],s223[24],s223[25],s223[26],s223[27],s223[28],s223[29],s223[30],s223[31],s223[32],s223[33],s223[34],s223[35],s223[36],s223[37],s221[40],s219[43],s217[46],s215[49],s213[52],s211[55],s209[58],s207[61],s205[64],s203[67],s203[68],s203[69],s203[70],s203[71],s203[72],s203[73],s203[74],s203[75],s203[76],s203[77],s203[78],s203[79],s203[80],s203[81],s203[82],s203[83],s203[84],s203[85],s203[86],s203[87],s203[88],s203[89],s203[90],s203[91],s203[92],s203[93],s203[94],s203[95],s204[95],s205[95],s206[95],s207[95],s208[95],s209[95],s210[95],s211[95],s212[95],s213[95],s214[95],s215[95],s216[95],s217[95],s218[95],s219[95],s220[95],s221[95],s222[95],s223[95],s224[95],s224[96],s224[97],s224[98],s224[99],s224[100],s224[101],s224[102],s224[103],s224[104],s224[105],s224[106],s224[107],s224[108],s224[109],s224[110],s224[111],s224[112],s224[113],s224[114],s224[115],s224[116],s224[117],s224[118],s224[119],s224[120],s224[121],s224[122],s224[123],s224[124],s224[125],s224[126],s224[127],s224[128],s224[129],s224[130],s224[131],s224[132],s224[133],s224[134],s224[135],s224[136],s224[137],s224[138],s224[139],s224[140],s224[141],s224[142],s224[143],s224[144],s224[145],s224[146],s224[147],s224[148],s224[149],s224[150],s224[151],s224[152],s224[153],s224[154],s224[155],s224[156],s224[157],s224[158],s224[159],s224[160],s224[161],s224[162],s224[163],s224[164],s224[165],s224[166],s224[167],s224[168],s224[169],s224[170],s224[171],s224[172],s224[173],s224[174],s224[175],s224[176],s224[177],s224[178],s224[179],s224[180],s224[181],s224[182],s224[183],s224[184],s224[185],s224[186],s224[187],s224[188],s224[189],s224[190],s224[191],s224[192],s224[193],s224[194],s224[195],s224[196],s224[197],s224[198],s224[199],s224[200],s224[201],s224[202],s224[203],s224[204],s224[205],s224[206],s224[207],s224[208],s224[209],s224[210],s224[211],s224[212],s224[213],s224[214],s224[215],s224[216],s224[217],s224[218],s224[219],s224[220],s224[221],s224[222],s224[223],s224[224],s224[225],s224[226],s224[227],s224[228],s224[229],s224[230],s224[231],s224[232],s224[233],s224[234],s224[235],s224[236],s224[237],s224[238],s224[239],s224[240],s224[241],s224[242],s224[243],s224[244],s224[245],s224[246],s224[247],s224[248],s224[249],s224[250],s224[251],s224[252],s224[253],s224[254],s224[255],s224[256],s224[257],s224[258],s224[259],s224[260],s224[261],s224[262],s224[263],s224[264],s224[265],s224[266],s224[267],s224[268],s224[269],s224[270],s224[271],s224[272],s224[273],s224[274],s224[275],s224[276],s224[277],s224[278],s224[279],s224[280],s224[281],s224[282],s224[283],s224[284],s224[285],s224[286],s224[287],s224[288],s224[289],s224[290],s224[291],s223[293],s222[295],s221[297],s220[299],s219[301],s218[303],s217[305],s216[307],s215[309],s214[311],s213[313],s212[315],s211[317],s210[319],s209[321],s208[323],s207[325],s206[327],s205[329],s204[331],s203[333],s202[335],s201[337],s200[339],s199[341],s198[343],s197[345],s196[347],s195[349],s194[351],s194[352],s194[353],s194[354],s194[355],s194[356],s194[357],s194[358],s194[359],s194[360],s194[361],s194[362],s194[363],s194[364],s194[365],s194[366],s194[367],s194[368],s194[369],s194[370],s194[371],s194[372],s194[373],s194[374],s194[375],s194[376],s194[377],s194[378],s194[379],s194[380],s194[381],s194[382],s194[383],s194[384],s194[385],s194[386],s194[387],s194[388],s194[389],s194[390],s194[391],s194[392],s194[393],s194[394],s194[395],s194[396],s194[397],s194[398],s194[399],s194[400],s194[401],s194[402],s194[403],s194[404],s194[405],s194[406],s194[407],s194[408],s194[409],s194[410],s194[411],s194[412],s194[413],s194[414],s194[415],s193[417],pp255[195],pp254[197],pp253[199],pp252[201],pp251[203],pp250[205],pp249[207],pp248[209],pp247[211],pp246[213],pp245[215],pp244[217],pp243[219],pp242[221],pp241[223],pp240[225],pp239[227],pp238[229],pp237[231],pp236[233],pp235[235],pp234[237],pp233[239],pp232[241],pp231[243],pp230[245],pp229[247],pp228[249],pp227[251],pp226[253],pp225[255],pp226[255],pp227[255],pp228[255],pp229[255],pp230[255],pp231[255],pp232[255],pp233[255],pp234[255],pp235[255],pp236[255],pp237[255],pp238[255],pp239[255],pp240[255]};
    assign in225_2 = {pp1[15],pp1[16],pp1[17],pp1[18],pp0[20],pp11[10],pp11[11],pp11[12],pp11[13],pp11[14],pp11[15],pp11[16],pp11[17],pp11[18],pp11[19],pp11[20],pp13[19],pp15[18],pp17[17],pp19[16],pp21[15],pp23[14],pp25[13],pp27[12],pp29[11],pp31[10],s193[10],s194[10],s195[10],s196[10],s197[10],s198[10],s199[10],s200[10],s201[10],s202[10],s203[10],s204[10],s205[10],s206[10],s207[10],s208[10],s209[10],s210[10],s211[10],s212[10],s213[10],s214[10],s215[10],s216[10],s217[10],s218[10],s219[10],s220[10],s221[10],s222[10],s223[10],s224[10],s224[11],s224[12],s224[13],s224[14],s224[15],s224[16],s224[17],s224[18],s224[19],s224[20],s224[21],s224[22],s224[23],s224[24],s224[25],s224[26],s224[27],s224[28],s224[29],s224[30],s224[31],s224[32],s224[33],s224[34],s224[35],s224[36],s222[39],s220[42],s218[45],s216[48],s214[51],s212[54],s210[57],s208[60],s206[63],s204[66],s204[67],s204[68],s204[69],s204[70],s204[71],s204[72],s204[73],s204[74],s204[75],s204[76],s204[77],s204[78],s204[79],s204[80],s204[81],s204[82],s204[83],s204[84],s204[85],s204[86],s204[87],s204[88],s204[89],s204[90],s204[91],s204[92],s204[93],s204[94],s205[94],s206[94],s207[94],s208[94],s209[94],s210[94],s211[94],s212[94],s213[94],s214[94],s215[94],s216[94],s217[94],s218[94],s219[94],s220[94],s221[94],s222[94],s223[94],s224[94],s10[21],s11[21],s12[21],s13[21],s14[21],s15[21],s16[21],s17[21],s18[21],s19[21],s20[21],s21[21],s22[21],s23[21],s24[21],s25[21],s26[21],s27[21],s28[21],s29[21],s30[21],s31[21],s32[21],s33[21],s34[21],s35[21],s36[21],s37[21],s38[21],s39[21],s40[21],s41[21],s42[21],s43[21],s44[21],s45[21],s46[21],s47[21],s48[21],s49[21],s50[21],s51[21],s52[21],s53[21],s54[21],s55[21],s56[21],s57[21],s58[21],s59[21],s60[21],s61[21],s62[21],s63[21],s64[21],s65[21],s66[21],s67[21],s68[21],s69[21],s70[21],s71[21],s72[21],s73[21],s74[21],s75[21],s76[21],s77[21],s78[21],s79[21],s79[22],s79[23],s79[24],s79[25],s79[26],s79[27],s79[28],s79[29],s79[30],s79[31],s79[32],s79[33],s79[34],s79[35],s79[36],s79[37],s79[38],s79[39],s79[40],s79[41],s79[42],s79[43],s79[44],s79[45],s79[46],s79[47],s79[48],s79[49],s79[50],s77[53],s75[56],s73[59],s71[62],s70[64],s70[65],s70[66],s70[67],s70[68],s70[69],s70[70],s70[71],s70[72],s70[73],s70[74],s70[75],s70[76],s70[77],s70[78],s70[79],s70[80],s70[81],s70[82],s70[83],s70[84],s70[85],s70[86],s70[87],s70[88],s69[90],s68[92],s67[94],s66[96],s65[98],s9[155],s7[158],s5[161],s3[164],s1[167],s68[101],s67[103],s66[105],s65[107],s64[109],s63[111],s62[113],s61[115],s60[117],s59[119],s58[121],s57[123],s56[125],s55[127],s54[129],s53[131],s52[133],s51[135],s50[137],s49[139],s48[141],s47[143],s46[145],s45[147],s44[149],s43[151],s42[153],s41[155],s40[157],s39[159],s38[161],s37[163],s36[165],s35[167],s34[169],s33[171],s32[173],s31[175],s30[177],s29[179],s28[181],s27[183],s26[185],s25[187],s24[189],s23[191],s22[193],s21[195],s20[197],s19[199],s18[201],s17[203],s16[205],s15[207],s14[209],s13[211],s12[213],s11[215],s10[217],s224[292],s223[294],s222[296],s221[298],s220[300],s219[302],s218[304],s217[306],s216[308],s215[310],s214[312],s213[314],s212[316],s211[318],s210[320],s209[322],s208[324],s207[326],s206[328],s205[330],s204[332],s203[334],s202[336],s201[338],s200[340],s199[342],s198[344],s197[346],s196[348],s195[350],s195[351],s195[352],s195[353],s195[354],s195[355],s195[356],s195[357],s195[358],s195[359],s195[360],s195[361],s195[362],s195[363],s195[364],s195[365],s195[366],s195[367],s195[368],s195[369],s195[370],s195[371],s195[372],s195[373],s195[374],s195[375],s195[376],s195[377],s195[378],s195[379],s195[380],s195[381],s195[382],s195[383],s195[384],s195[385],s195[386],s195[387],s195[388],s195[389],s195[390],s195[391],s195[392],s195[393],s195[394],s195[395],s195[396],s195[397],s195[398],s195[399],s195[400],s195[401],s195[402],s195[403],s195[404],s195[405],s195[406],s195[407],s195[408],s195[409],s195[410],s195[411],s195[412],s195[413],s195[414],s194[416],s193[418],pp255[196],pp254[198],pp253[200],pp252[202],pp251[204],pp250[206],pp249[208],pp248[210],pp247[212],pp246[214],pp245[216],pp244[218],pp243[220],pp242[222],pp241[224],pp240[226],pp239[228],pp238[230],pp237[232],pp236[234],pp235[236],pp234[238],pp233[240],pp232[242],pp231[244],pp230[246],pp229[248],pp228[250],pp227[252],pp226[254],pp227[254],pp228[254],pp229[254],pp230[254],pp231[254],pp232[254],pp233[254],pp234[254],pp235[254],pp236[254],pp237[254],pp238[254],pp239[254],pp240[254],pp241[254]};
    CLA_480 KS_225(s225, c225, in225_1, in225_2);
    wire[477:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {pp2[15],pp2[16],pp2[17],pp1[19],pp0[21],pp12[10],pp12[11],pp12[12],pp12[13],pp12[14],pp12[15],pp12[16],pp12[17],pp12[18],pp12[19],pp14[18],pp16[17],pp18[16],pp20[15],pp22[14],pp24[13],pp26[12],pp28[11],pp30[10],s225[25],s225[26],s225[27],s225[28],s225[29],s225[30],s225[31],s225[32],s225[33],s225[34],s225[35],s225[36],s225[37],s225[38],s225[39],s225[40],s225[41],s225[42],s225[43],s225[44],s225[45],s225[46],s225[47],s225[48],s225[49],s225[50],s225[51],s225[52],s225[53],s225[54],s225[55],s225[56],s225[57],s225[58],s225[59],s225[60],s225[61],s225[62],s225[63],s225[64],s225[65],s225[66],s225[67],s225[68],s225[69],s225[70],s225[71],s225[72],s225[73],s225[74],s225[75],s225[76],s225[77],s225[78],s225[79],s225[80],s225[81],s225[82],s225[83],s223[38],s221[41],s219[44],s217[47],s215[50],s213[53],s211[56],s209[59],s207[62],s205[65],s205[66],s205[67],s205[68],s205[69],s205[70],s205[71],s225[100],s225[101],s225[102],s225[103],s225[104],s225[105],s225[106],s225[107],s225[108],s225[109],s225[110],s225[111],s225[112],s225[113],s225[114],s225[115],s225[116],s225[117],s225[118],s225[119],s225[120],s225[121],s225[122],s225[123],s225[124],s225[125],s225[126],s225[127],s225[128],s225[129],s225[130],s225[131],s225[132],s225[133],s225[134],s225[135],s225[136],s225[137],s225[138],s225[139],s225[140],s225[141],s225[142],s225[143],s225[144],s225[145],s225[146],s225[147],s225[148],s225[149],s225[150],s225[151],s225[152],s225[153],s225[154],s225[155],s225[156],s225[157],s225[158],s225[159],s225[160],s225[161],s225[162],s225[163],s225[164],s225[165],s225[166],s225[167],s225[168],s225[169],s225[170],s225[171],s225[172],s225[173],s225[174],s225[175],s225[176],s225[177],s225[178],s225[179],s225[180],s225[181],s225[182],s225[183],s225[184],s225[185],s225[186],s225[187],s225[188],s225[189],s225[190],s225[191],s225[192],s225[193],s225[194],s225[195],s225[196],s225[197],s225[198],s225[199],s225[200],s225[201],s225[202],s225[203],s225[204],s225[205],s225[206],s225[207],s225[208],s225[209],s225[210],s225[211],s225[212],s225[213],s225[214],s225[215],s225[216],s225[217],s225[218],s225[219],s225[220],s225[221],s225[222],s225[223],s225[224],s225[225],s225[226],s225[227],s225[228],s225[229],s225[230],s225[231],s225[232],s225[233],s225[234],s225[235],s225[236],s225[237],s225[238],s225[239],s225[240],s225[241],s225[242],s225[243],s225[244],s225[245],s225[246],s225[247],s225[248],s225[249],s225[250],s225[251],s225[252],s225[253],s225[254],s225[255],s225[256],s225[257],s225[258],s225[259],s225[260],s225[261],s225[262],s225[263],s225[264],s225[265],s225[266],s225[267],s225[268],s225[269],s225[270],s225[271],s225[272],s225[273],s225[274],s225[275],s225[276],s225[277],s225[278],s225[279],s225[280],s225[281],s225[282],s225[283],s225[284],s225[285],s225[286],s225[287],s225[288],s225[289],s225[290],s225[291],s225[292],s225[293],s225[294],s225[295],s225[296],s225[297],s225[298],s225[299],s225[300],s225[301],s225[302],s225[303],s225[304],s225[305],s225[306],s225[307],s225[308],s225[309],s225[310],s225[311],s225[312],s225[313],s225[314],s225[315],s225[316],s225[317],s225[318],s225[319],s225[320],s225[321],s225[322],s225[323],s225[324],s225[325],s225[326],s225[327],s225[328],s225[329],s225[330],s225[331],s225[332],s225[333],s225[334],s225[335],s225[336],s225[337],s225[338],s225[339],s224[293],s223[295],s222[297],s221[299],s220[301],s219[303],s218[305],s217[307],s216[309],s215[311],s214[313],s213[315],s212[317],s211[319],s210[321],s209[323],s208[325],s207[327],s206[329],s205[331],s204[333],s203[335],s202[337],s201[339],s200[341],s199[343],s198[345],s197[347],s196[349],s196[350],s196[351],s196[352],s196[353],s196[354],s196[355],s196[356],s196[357],s196[358],s196[359],s196[360],s196[361],s196[362],s196[363],s196[364],s196[365],s196[366],s196[367],s196[368],s196[369],s196[370],s196[371],s196[372],s196[373],s196[374],s196[375],s196[376],s196[377],s196[378],s196[379],s196[380],s196[381],s196[382],s196[383],s196[384],s196[385],s196[386],s196[387],s196[388],s196[389],s196[390],s196[391],s196[392],s196[393],s196[394],s196[395],s196[396],s196[397],s196[398],s196[399],s196[400],s196[401],s196[402],s196[403],s196[404],s196[405],s196[406],s196[407],s196[408],s196[409],s196[410],s196[411],s196[412],s196[413],s195[415],s194[417],s193[419],pp255[197],pp254[199],pp253[201],pp252[203],pp251[205],pp250[207],pp249[209],pp248[211],pp247[213],pp246[215],pp245[217],pp244[219],pp243[221],pp242[223],pp241[225],pp240[227],pp239[229],pp238[231],pp237[233],pp236[235],pp235[237],pp234[239],pp233[241],pp232[243],pp231[245],pp230[247],pp229[249],pp228[251],pp227[253],pp228[253],pp229[253],pp230[253],pp231[253],pp232[253],pp233[253],pp234[253],pp235[253],pp236[253],pp237[253],pp238[253],pp239[253],pp240[253],pp241[253]};
    assign in226_2 = {pp3[14],pp3[15],pp3[16],pp2[18],pp1[20],pp0[22],pp13[10],pp13[11],pp13[12],pp13[13],pp13[14],pp13[15],pp13[16],pp13[17],pp13[18],pp15[17],pp17[16],pp19[15],pp21[14],pp23[13],pp25[12],pp27[11],pp29[10],s225[24],pp0[41],pp0[42],pp0[43],pp0[44],pp0[45],pp0[46],pp0[47],pp0[48],pp0[49],pp0[50],pp0[51],pp0[52],pp0[53],pp0[54],pp0[55],pp0[56],pp0[57],pp0[58],pp0[59],pp0[60],pp0[61],pp0[62],pp0[63],pp0[64],pp0[65],pp0[66],pp0[67],pp0[68],pp0[69],pp0[70],pp0[71],pp0[72],pp0[73],pp0[74],pp0[75],pp0[76],pp0[77],pp0[78],pp0[79],pp0[80],pp0[81],pp0[82],pp0[83],pp0[84],pp0[85],pp0[86],pp0[87],pp0[88],pp0[89],pp0[90],pp0[91],pp0[92],pp0[93],pp0[94],pp0[95],pp0[96],pp0[97],pp0[98],pp0[99],s224[37],s222[40],s220[43],s218[46],s216[49],s214[52],s212[55],s210[58],s208[61],s206[64],s206[65],s206[66],s206[67],s206[68],s206[69],s206[70],s205[72],s205[73],s205[74],s205[75],s205[76],s205[77],s205[78],s205[79],s205[80],s205[81],s205[82],s205[83],s205[84],s205[85],s205[86],s205[87],s205[88],s205[89],s205[90],s205[91],s205[92],s205[93],s206[93],s207[93],s208[93],s209[93],s210[93],s211[93],s212[93],s213[93],s214[93],s215[93],s216[93],s217[93],s218[93],s219[93],s220[93],s221[93],s222[93],s223[93],s224[93],s10[20],s11[20],s12[20],s13[20],s14[20],s15[20],s16[20],s17[20],s18[20],s19[20],s20[20],s21[20],s22[20],s23[20],s24[20],s25[20],s26[20],s27[20],s28[20],s29[20],s30[20],s31[20],s32[20],s33[20],s34[20],s35[20],s36[20],s37[20],s38[20],s39[20],s40[20],s41[20],s42[20],s43[20],s44[20],s45[20],s46[20],s47[20],s48[20],s49[20],s50[20],s51[20],s52[20],s53[20],s54[20],s55[20],s56[20],s57[20],s58[20],s59[20],s60[20],s61[20],s62[20],s63[20],s64[20],s65[20],s66[20],s67[20],s68[20],s69[20],s70[20],s71[20],s72[20],s73[20],s74[20],s75[20],s76[20],s77[20],s78[20],s79[20],s80[20],s80[21],s80[22],s80[23],s80[24],s80[25],s80[26],s80[27],s80[28],s80[29],s80[30],s80[31],s80[32],s80[33],s80[34],s80[35],s80[36],s80[37],s80[38],s80[39],s80[40],s80[41],s80[42],s80[43],s80[44],s80[45],s80[46],s80[47],s80[48],s80[49],s78[52],s76[55],s74[58],s72[61],s71[63],s71[64],s71[65],s71[66],s71[67],s71[68],s71[69],s71[70],s71[71],s71[72],s71[73],s71[74],s71[75],s71[76],s71[77],s71[78],s71[79],s71[80],s71[81],s71[82],s71[83],s71[84],s71[85],s71[86],s71[87],s70[89],s69[91],s68[93],s67[95],s66[97],s65[99],s8[157],s6[160],s4[163],s2[166],s69[100],s68[102],s67[104],s66[106],s65[108],s64[110],s63[112],s62[114],s61[116],s60[118],s59[120],s58[122],s57[124],s56[126],s55[128],s54[130],s53[132],s52[134],s51[136],s50[138],s49[140],s48[142],s47[144],s46[146],s45[148],s44[150],s43[152],s42[154],s41[156],s40[158],s39[160],s38[162],s37[164],s36[166],s35[168],s34[170],s33[172],s32[174],s31[176],s30[178],s29[180],s28[182],s27[184],s26[186],s25[188],s24[190],s23[192],s22[194],s21[196],s20[198],s19[200],s18[202],s17[204],s16[206],s15[208],s14[210],s13[212],s12[214],s11[216],s10[218],s225[340],s224[294],s223[296],s222[298],s221[300],s220[302],s219[304],s218[306],s217[308],s216[310],s215[312],s214[314],s213[316],s212[318],s211[320],s210[322],s209[324],s208[326],s207[328],s206[330],s205[332],s204[334],s203[336],s202[338],s201[340],s200[342],s199[344],s198[346],s197[348],s197[349],s197[350],s197[351],s197[352],s197[353],s197[354],s197[355],s197[356],s197[357],s197[358],s197[359],s197[360],s197[361],s197[362],s197[363],s197[364],s197[365],s197[366],s197[367],s197[368],s197[369],s197[370],s197[371],s197[372],s197[373],s197[374],s197[375],s197[376],s197[377],s197[378],s197[379],s197[380],s197[381],s197[382],s197[383],s197[384],s197[385],s197[386],s197[387],s197[388],s197[389],s197[390],s197[391],s197[392],s197[393],s197[394],s197[395],s197[396],s197[397],s197[398],s197[399],s197[400],s197[401],s197[402],s197[403],s197[404],s197[405],s197[406],s197[407],s197[408],s197[409],s197[410],s197[411],s197[412],s196[414],s195[416],s194[418],s193[420],pp255[198],pp254[200],pp253[202],pp252[204],pp251[206],pp250[208],pp249[210],pp248[212],pp247[214],pp246[216],pp245[218],pp244[220],pp243[222],pp242[224],pp241[226],pp240[228],pp239[230],pp238[232],pp237[234],pp236[236],pp235[238],pp234[240],pp233[242],pp232[244],pp231[246],pp230[248],pp229[250],pp228[252],pp229[252],pp230[252],pp231[252],pp232[252],pp233[252],pp234[252],pp235[252],pp236[252],pp237[252],pp238[252],pp239[252],pp240[252],pp241[252],pp242[252]};
    CLA_478 KS_226(s226, c226, in226_1, in226_2);
    wire[475:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {pp4[14],pp4[15],pp3[17],pp2[19],pp1[21],pp0[23],pp14[10],pp14[11],pp14[12],pp14[13],pp14[14],pp14[15],pp14[16],pp14[17],pp16[16],pp18[15],pp20[14],pp22[13],pp24[12],pp26[11],pp28[10],s225[23],s226[23],s226[24],s226[25],s226[26],s226[27],s226[28],s226[29],s226[30],s226[31],s226[32],s226[33],s226[34],s226[35],s226[36],s226[37],s226[38],s226[39],s226[40],s226[41],s226[42],s226[43],s226[44],s226[45],s226[46],s226[47],s226[48],s226[49],s226[50],s226[51],s226[52],s226[53],s226[54],s226[55],s226[56],s226[57],s226[58],s226[59],s226[60],s226[61],s226[62],s226[63],s226[64],s226[65],s226[66],s226[67],s226[68],s226[69],s226[70],s226[71],s226[72],s226[73],s226[74],s226[75],s226[76],s226[77],s226[78],s226[79],s226[80],s226[81],s226[82],s225[84],s223[39],s221[42],s219[45],s217[48],s215[51],s213[54],s211[57],s209[60],s207[63],s207[64],s207[65],s207[66],s207[67],s207[68],s207[69],s206[71],s226[100],s226[101],s226[102],s226[103],s226[104],s226[105],s226[106],s226[107],s226[108],s226[109],s226[110],s226[111],s226[112],s226[113],s226[114],s226[115],s226[116],s226[117],s226[118],s226[119],s226[120],s226[121],s226[122],s226[123],s226[124],s226[125],s226[126],s226[127],s226[128],s226[129],s226[130],s226[131],s226[132],s226[133],s226[134],s226[135],s226[136],s226[137],s226[138],s226[139],s226[140],s226[141],s226[142],s226[143],s226[144],s226[145],s226[146],s226[147],s226[148],s226[149],s226[150],s226[151],s226[152],s226[153],s226[154],s226[155],s226[156],s226[157],s226[158],s226[159],s226[160],s226[161],s226[162],s226[163],s226[164],s226[165],s226[166],s226[167],s226[168],s226[169],s226[170],s226[171],s226[172],s226[173],s226[174],s226[175],s226[176],s226[177],s226[178],s226[179],s226[180],s226[181],s226[182],s226[183],s226[184],s226[185],s226[186],s226[187],s226[188],s226[189],s226[190],s226[191],s226[192],s226[193],s226[194],s226[195],s226[196],s226[197],s226[198],s226[199],s226[200],s226[201],s226[202],s226[203],s226[204],s226[205],s226[206],s226[207],s226[208],s226[209],s226[210],s226[211],s226[212],s226[213],s226[214],s226[215],s226[216],s226[217],s226[218],s226[219],s226[220],s226[221],s226[222],s226[223],s226[224],s226[225],s226[226],s226[227],s226[228],s226[229],s226[230],s226[231],s226[232],s226[233],s226[234],s226[235],s226[236],s226[237],s226[238],s226[239],s226[240],s226[241],s226[242],s226[243],s226[244],s226[245],s226[246],s226[247],s226[248],s226[249],s226[250],s226[251],s226[252],s226[253],s226[254],s226[255],s226[256],s226[257],s226[258],s226[259],s226[260],s226[261],s226[262],s226[263],s226[264],s226[265],s226[266],s226[267],s226[268],s226[269],s226[270],s226[271],s226[272],s226[273],s226[274],s226[275],s226[276],s226[277],s226[278],s226[279],s226[280],s226[281],s226[282],s226[283],s226[284],s226[285],s226[286],s226[287],s226[288],s226[289],s226[290],s226[291],s226[292],s226[293],s226[294],s226[295],s226[296],s226[297],s226[298],s226[299],s226[300],s226[301],s226[302],s226[303],s226[304],s226[305],s226[306],s226[307],s226[308],s226[309],s226[310],s226[311],s226[312],s226[313],s226[314],s226[315],s226[316],s226[317],s226[318],s226[319],s226[320],s226[321],s226[322],s226[323],s226[324],s226[325],s226[326],s226[327],s226[328],s226[329],s226[330],s226[331],s226[332],s226[333],s226[334],s226[335],s226[336],s226[337],s226[338],s226[339],s225[341],s224[295],s223[297],s222[299],s221[301],s220[303],s219[305],s218[307],s217[309],s216[311],s215[313],s214[315],s213[317],s212[319],s211[321],s210[323],s209[325],s208[327],s207[329],s206[331],s205[333],s204[335],s203[337],s202[339],s201[341],s200[343],s199[345],s198[347],s198[348],s198[349],s198[350],s198[351],s198[352],s198[353],s198[354],s198[355],s198[356],s198[357],s198[358],s198[359],s198[360],s198[361],s198[362],s198[363],s198[364],s198[365],s198[366],s198[367],s198[368],s198[369],s198[370],s198[371],s198[372],s198[373],s198[374],s198[375],s198[376],s198[377],s198[378],s198[379],s198[380],s198[381],s198[382],s198[383],s198[384],s198[385],s198[386],s198[387],s198[388],s198[389],s198[390],s198[391],s198[392],s198[393],s198[394],s198[395],s198[396],s198[397],s198[398],s198[399],s198[400],s198[401],s198[402],s198[403],s198[404],s198[405],s198[406],s198[407],s198[408],s198[409],s198[410],s198[411],s197[413],s196[415],s195[417],s194[419],s193[421],pp255[199],pp254[201],pp253[203],pp252[205],pp251[207],pp250[209],pp249[211],pp248[213],pp247[215],pp246[217],pp245[219],pp244[221],pp243[223],pp242[225],pp241[227],pp240[229],pp239[231],pp238[233],pp237[235],pp236[237],pp235[239],pp234[241],pp233[243],pp232[245],pp231[247],pp230[249],pp229[251],pp230[251],pp231[251],pp232[251],pp233[251],pp234[251],pp235[251],pp236[251],pp237[251],pp238[251],pp239[251],pp240[251],pp241[251],pp242[251]};
    assign in227_2 = {pp5[13],pp5[14],pp4[16],pp3[18],pp2[20],pp1[22],pp0[24],pp15[10],pp15[11],pp15[12],pp15[13],pp15[14],pp15[15],pp15[16],pp17[15],pp19[14],pp21[13],pp23[12],pp25[11],pp27[10],s225[22],s226[22],pp0[40],pp1[40],pp1[41],pp1[42],pp1[43],pp1[44],pp1[45],pp1[46],pp1[47],pp1[48],pp1[49],pp1[50],pp1[51],pp1[52],pp1[53],pp1[54],pp1[55],pp1[56],pp1[57],pp1[58],pp1[59],pp1[60],pp1[61],pp1[62],pp1[63],pp1[64],pp1[65],pp1[66],pp1[67],pp1[68],pp1[69],pp1[70],pp1[71],pp1[72],pp1[73],pp1[74],pp1[75],pp1[76],pp1[77],pp1[78],pp1[79],pp1[80],pp1[81],pp1[82],pp1[83],pp1[84],pp1[85],pp1[86],pp1[87],pp1[88],pp1[89],pp1[90],pp1[91],pp1[92],pp1[93],pp1[94],pp1[95],pp1[96],pp1[97],pp1[98],s226[83],s224[38],s222[41],s220[44],s218[47],s216[50],s214[53],s212[56],s210[59],s208[62],s208[63],s208[64],s208[65],s208[66],s208[67],s208[68],s207[70],s206[72],s206[73],s206[74],s206[75],s206[76],s206[77],s206[78],s206[79],s206[80],s206[81],s206[82],s206[83],s206[84],s206[85],s206[86],s206[87],s206[88],s206[89],s206[90],s206[91],s206[92],s207[92],s208[92],s209[92],s210[92],s211[92],s212[92],s213[92],s214[92],s215[92],s216[92],s217[92],s218[92],s219[92],s220[92],s221[92],s222[92],s223[92],s224[92],s10[19],s11[19],s12[19],s13[19],s14[19],s15[19],s16[19],s17[19],s18[19],s19[19],s20[19],s21[19],s22[19],s23[19],s24[19],s25[19],s26[19],s27[19],s28[19],s29[19],s30[19],s31[19],s32[19],s33[19],s34[19],s35[19],s36[19],s37[19],s38[19],s39[19],s40[19],s41[19],s42[19],s43[19],s44[19],s45[19],s46[19],s47[19],s48[19],s49[19],s50[19],s51[19],s52[19],s53[19],s54[19],s55[19],s56[19],s57[19],s58[19],s59[19],s60[19],s61[19],s62[19],s63[19],s64[19],s65[19],s66[19],s67[19],s68[19],s69[19],s70[19],s71[19],s72[19],s73[19],s74[19],s75[19],s76[19],s77[19],s78[19],s79[19],s80[19],s81[19],s81[20],s81[21],s81[22],s81[23],s81[24],s81[25],s81[26],s81[27],s81[28],s81[29],s81[30],s81[31],s81[32],s81[33],s81[34],s81[35],s81[36],s81[37],s81[38],s81[39],s81[40],s81[41],s81[42],s81[43],s81[44],s81[45],s81[46],s81[47],s81[48],s79[51],s77[54],s75[57],s73[60],s72[62],s72[63],s72[64],s72[65],s72[66],s72[67],s72[68],s72[69],s72[70],s72[71],s72[72],s72[73],s72[74],s72[75],s72[76],s72[77],s72[78],s72[79],s72[80],s72[81],s72[82],s72[83],s72[84],s72[85],s72[86],s71[88],s70[90],s69[92],s68[94],s67[96],s66[98],s9[156],s7[159],s5[162],s3[165],s1[168],s69[101],s68[103],s67[105],s66[107],s65[109],s64[111],s63[113],s62[115],s61[117],s60[119],s59[121],s58[123],s57[125],s56[127],s55[129],s54[131],s53[133],s52[135],s51[137],s50[139],s49[141],s48[143],s47[145],s46[147],s45[149],s44[151],s43[153],s42[155],s41[157],s40[159],s39[161],s38[163],s37[165],s36[167],s35[169],s34[171],s33[173],s32[175],s31[177],s30[179],s29[181],s28[183],s27[185],s26[187],s25[189],s24[191],s23[193],s22[195],s21[197],s20[199],s19[201],s18[203],s17[205],s16[207],s15[209],s14[211],s13[213],s12[215],s11[217],s10[219],s226[340],s225[342],s224[296],s223[298],s222[300],s221[302],s220[304],s219[306],s218[308],s217[310],s216[312],s215[314],s214[316],s213[318],s212[320],s211[322],s210[324],s209[326],s208[328],s207[330],s206[332],s205[334],s204[336],s203[338],s202[340],s201[342],s200[344],s199[346],s199[347],s199[348],s199[349],s199[350],s199[351],s199[352],s199[353],s199[354],s199[355],s199[356],s199[357],s199[358],s199[359],s199[360],s199[361],s199[362],s199[363],s199[364],s199[365],s199[366],s199[367],s199[368],s199[369],s199[370],s199[371],s199[372],s199[373],s199[374],s199[375],s199[376],s199[377],s199[378],s199[379],s199[380],s199[381],s199[382],s199[383],s199[384],s199[385],s199[386],s199[387],s199[388],s199[389],s199[390],s199[391],s199[392],s199[393],s199[394],s199[395],s199[396],s199[397],s199[398],s199[399],s199[400],s199[401],s199[402],s199[403],s199[404],s199[405],s199[406],s199[407],s199[408],s199[409],s199[410],s198[412],s197[414],s196[416],s195[418],s194[420],s193[422],pp255[200],pp254[202],pp253[204],pp252[206],pp251[208],pp250[210],pp249[212],pp248[214],pp247[216],pp246[218],pp245[220],pp244[222],pp243[224],pp242[226],pp241[228],pp240[230],pp239[232],pp238[234],pp237[236],pp236[238],pp235[240],pp234[242],pp233[244],pp232[246],pp231[248],pp230[250],pp231[250],pp232[250],pp233[250],pp234[250],pp235[250],pp236[250],pp237[250],pp238[250],pp239[250],pp240[250],pp241[250],pp242[250],pp243[250]};
    CLA_476 KS_227(s227, c227, in227_1, in227_2);
    wire[473:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {pp6[13],pp5[15],pp4[17],pp3[19],pp2[21],pp1[23],pp0[25],pp16[10],pp16[11],pp16[12],pp16[13],pp16[14],pp16[15],pp18[14],pp20[13],pp22[12],pp24[11],pp26[10],s225[21],s226[21],s227[21],s227[22],s227[23],s227[24],s227[25],s227[26],s227[27],s227[28],s227[29],s227[30],s227[31],s227[32],s227[33],s227[34],s227[35],s227[36],s227[37],s227[38],s227[39],s227[40],s227[41],s227[42],s227[43],s227[44],s227[45],s227[46],s227[47],s227[48],s227[49],s227[50],s227[51],s227[52],s227[53],s227[54],s227[55],s227[56],s227[57],s227[58],s227[59],s227[60],s227[61],s227[62],s227[63],s227[64],s227[65],s227[66],s227[67],s227[68],s227[69],s227[70],s227[71],s227[72],s227[73],s227[74],s227[75],s227[76],s227[77],s227[78],s227[79],s227[80],s227[81],s227[82],s225[85],s223[40],s221[43],s219[46],s217[49],s215[52],s213[55],s211[58],s209[61],s209[62],s209[63],s209[64],s209[65],s209[66],s209[67],s208[69],s207[71],s227[100],s227[101],s227[102],s227[103],s227[104],s227[105],s227[106],s227[107],s227[108],s227[109],s227[110],s227[111],s227[112],s227[113],s227[114],s227[115],s227[116],s227[117],s227[118],s227[119],s227[120],s227[121],s227[122],s227[123],s227[124],s227[125],s227[126],s227[127],s227[128],s227[129],s227[130],s227[131],s227[132],s227[133],s227[134],s227[135],s227[136],s227[137],s227[138],s227[139],s227[140],s227[141],s227[142],s227[143],s227[144],s227[145],s227[146],s227[147],s227[148],s227[149],s227[150],s227[151],s227[152],s227[153],s227[154],s227[155],s227[156],s227[157],s227[158],s227[159],s227[160],s227[161],s227[162],s227[163],s227[164],s227[165],s227[166],s227[167],s227[168],s227[169],s227[170],s227[171],s227[172],s227[173],s227[174],s227[175],s227[176],s227[177],s227[178],s227[179],s227[180],s227[181],s227[182],s227[183],s227[184],s227[185],s227[186],s227[187],s227[188],s227[189],s227[190],s227[191],s227[192],s227[193],s227[194],s227[195],s227[196],s227[197],s227[198],s227[199],s227[200],s227[201],s227[202],s227[203],s227[204],s227[205],s227[206],s227[207],s227[208],s227[209],s227[210],s227[211],s227[212],s227[213],s227[214],s227[215],s227[216],s227[217],s227[218],s227[219],s227[220],s227[221],s227[222],s227[223],s227[224],s227[225],s227[226],s227[227],s227[228],s227[229],s227[230],s227[231],s227[232],s227[233],s227[234],s227[235],s227[236],s227[237],s227[238],s227[239],s227[240],s227[241],s227[242],s227[243],s227[244],s227[245],s227[246],s227[247],s227[248],s227[249],s227[250],s227[251],s227[252],s227[253],s227[254],s227[255],s227[256],s227[257],s227[258],s227[259],s227[260],s227[261],s227[262],s227[263],s227[264],s227[265],s227[266],s227[267],s227[268],s227[269],s227[270],s227[271],s227[272],s227[273],s227[274],s227[275],s227[276],s227[277],s227[278],s227[279],s227[280],s227[281],s227[282],s227[283],s227[284],s227[285],s227[286],s227[287],s227[288],s227[289],s227[290],s227[291],s227[292],s227[293],s227[294],s227[295],s227[296],s227[297],s227[298],s227[299],s227[300],s227[301],s227[302],s227[303],s227[304],s227[305],s227[306],s227[307],s227[308],s227[309],s227[310],s227[311],s227[312],s227[313],s227[314],s227[315],s227[316],s227[317],s227[318],s227[319],s227[320],s227[321],s227[322],s227[323],s227[324],s227[325],s227[326],s227[327],s227[328],s227[329],s227[330],s227[331],s227[332],s227[333],s227[334],s227[335],s227[336],s227[337],s227[338],s227[339],s226[341],s225[343],s224[297],s223[299],s222[301],s221[303],s220[305],s219[307],s218[309],s217[311],s216[313],s215[315],s214[317],s213[319],s212[321],s211[323],s210[325],s209[327],s208[329],s207[331],s206[333],s205[335],s204[337],s203[339],s202[341],s201[343],s200[345],s200[346],s200[347],s200[348],s200[349],s200[350],s200[351],s200[352],s200[353],s200[354],s200[355],s200[356],s200[357],s200[358],s200[359],s200[360],s200[361],s200[362],s200[363],s200[364],s200[365],s200[366],s200[367],s200[368],s200[369],s200[370],s200[371],s200[372],s200[373],s200[374],s200[375],s200[376],s200[377],s200[378],s200[379],s200[380],s200[381],s200[382],s200[383],s200[384],s200[385],s200[386],s200[387],s200[388],s200[389],s200[390],s200[391],s200[392],s200[393],s200[394],s200[395],s200[396],s200[397],s200[398],s200[399],s200[400],s200[401],s200[402],s200[403],s200[404],s200[405],s200[406],s200[407],s200[408],s200[409],s199[411],s198[413],s197[415],s196[417],s195[419],s194[421],s193[423],pp255[201],pp254[203],pp253[205],pp252[207],pp251[209],pp250[211],pp249[213],pp248[215],pp247[217],pp246[219],pp245[221],pp244[223],pp243[225],pp242[227],pp241[229],pp240[231],pp239[233],pp238[235],pp237[237],pp236[239],pp235[241],pp234[243],pp233[245],pp232[247],pp231[249],pp232[249],pp233[249],pp234[249],pp235[249],pp236[249],pp237[249],pp238[249],pp239[249],pp240[249],pp241[249],pp242[249],pp243[249]};
    assign in228_2 = {pp7[12],pp6[14],pp5[16],pp4[18],pp3[20],pp2[22],pp1[24],s225[10],pp17[10],pp17[11],pp17[12],pp17[13],pp17[14],pp19[13],pp21[12],pp23[11],pp25[10],s225[20],s226[20],s227[20],pp0[39],pp1[39],pp2[39],pp2[40],pp2[41],pp2[42],pp2[43],pp2[44],pp2[45],pp2[46],pp2[47],pp2[48],pp2[49],pp2[50],pp2[51],pp2[52],pp2[53],pp2[54],pp2[55],pp2[56],pp2[57],pp2[58],pp2[59],pp2[60],pp2[61],pp2[62],pp2[63],pp2[64],pp2[65],pp2[66],pp2[67],pp2[68],pp2[69],pp2[70],pp2[71],pp2[72],pp2[73],pp2[74],pp2[75],pp2[76],pp2[77],pp2[78],pp2[79],pp2[80],pp2[81],pp2[82],pp2[83],pp2[84],pp2[85],pp2[86],pp2[87],pp2[88],pp2[89],pp2[90],pp2[91],pp2[92],pp2[93],pp2[94],pp2[95],pp2[96],pp2[97],pp1[99],s226[84],s224[39],s222[42],s220[45],s218[48],s216[51],s214[54],s212[57],s210[60],s210[61],s210[62],s210[63],s210[64],s210[65],s210[66],s209[68],s208[70],s207[72],s207[73],s207[74],s207[75],s207[76],s207[77],s207[78],s207[79],s207[80],s207[81],s207[82],s207[83],s207[84],s207[85],s207[86],s207[87],s207[88],s207[89],s207[90],s207[91],s208[91],s209[91],s210[91],s211[91],s212[91],s213[91],s214[91],s215[91],s216[91],s217[91],s218[91],s219[91],s220[91],s221[91],s222[91],s223[91],s224[91],s10[18],s11[18],s12[18],s13[18],s14[18],s15[18],s16[18],s17[18],s18[18],s19[18],s20[18],s21[18],s22[18],s23[18],s24[18],s25[18],s26[18],s27[18],s28[18],s29[18],s30[18],s31[18],s32[18],s33[18],s34[18],s35[18],s36[18],s37[18],s38[18],s39[18],s40[18],s41[18],s42[18],s43[18],s44[18],s45[18],s46[18],s47[18],s48[18],s49[18],s50[18],s51[18],s52[18],s53[18],s54[18],s55[18],s56[18],s57[18],s58[18],s59[18],s60[18],s61[18],s62[18],s63[18],s64[18],s65[18],s66[18],s67[18],s68[18],s69[18],s70[18],s71[18],s72[18],s73[18],s74[18],s75[18],s76[18],s77[18],s78[18],s79[18],s80[18],s81[18],s82[18],s82[19],s82[20],s82[21],s82[22],s82[23],s82[24],s82[25],s82[26],s82[27],s82[28],s82[29],s82[30],s82[31],s82[32],s82[33],s82[34],s82[35],s82[36],s82[37],s82[38],s82[39],s82[40],s82[41],s82[42],s82[43],s82[44],s82[45],s82[46],s82[47],s80[50],s78[53],s76[56],s74[59],s73[61],s73[62],s73[63],s73[64],s73[65],s73[66],s73[67],s73[68],s73[69],s73[70],s73[71],s73[72],s73[73],s73[74],s73[75],s73[76],s73[77],s73[78],s73[79],s73[80],s73[81],s73[82],s73[83],s73[84],s73[85],s72[87],s71[89],s70[91],s69[93],s68[95],s67[97],s66[99],s8[158],s6[161],s4[164],s2[167],s70[100],s69[102],s68[104],s67[106],s66[108],s65[110],s64[112],s63[114],s62[116],s61[118],s60[120],s59[122],s58[124],s57[126],s56[128],s55[130],s54[132],s53[134],s52[136],s51[138],s50[140],s49[142],s48[144],s47[146],s46[148],s45[150],s44[152],s43[154],s42[156],s41[158],s40[160],s39[162],s38[164],s37[166],s36[168],s35[170],s34[172],s33[174],s32[176],s31[178],s30[180],s29[182],s28[184],s27[186],s26[188],s25[190],s24[192],s23[194],s22[196],s21[198],s20[200],s19[202],s18[204],s17[206],s16[208],s15[210],s14[212],s13[214],s12[216],s11[218],s10[220],s227[340],s226[342],s225[344],s224[298],s223[300],s222[302],s221[304],s220[306],s219[308],s218[310],s217[312],s216[314],s215[316],s214[318],s213[320],s212[322],s211[324],s210[326],s209[328],s208[330],s207[332],s206[334],s205[336],s204[338],s203[340],s202[342],s201[344],s201[345],s201[346],s201[347],s201[348],s201[349],s201[350],s201[351],s201[352],s201[353],s201[354],s201[355],s201[356],s201[357],s201[358],s201[359],s201[360],s201[361],s201[362],s201[363],s201[364],s201[365],s201[366],s201[367],s201[368],s201[369],s201[370],s201[371],s201[372],s201[373],s201[374],s201[375],s201[376],s201[377],s201[378],s201[379],s201[380],s201[381],s201[382],s201[383],s201[384],s201[385],s201[386],s201[387],s201[388],s201[389],s201[390],s201[391],s201[392],s201[393],s201[394],s201[395],s201[396],s201[397],s201[398],s201[399],s201[400],s201[401],s201[402],s201[403],s201[404],s201[405],s201[406],s201[407],s201[408],s200[410],s199[412],s198[414],s197[416],s196[418],s195[420],s194[422],s193[424],pp255[202],pp254[204],pp253[206],pp252[208],pp251[210],pp250[212],pp249[214],pp248[216],pp247[218],pp246[220],pp245[222],pp244[224],pp243[226],pp242[228],pp241[230],pp240[232],pp239[234],pp238[236],pp237[238],pp236[240],pp235[242],pp234[244],pp233[246],pp232[248],pp233[248],pp234[248],pp235[248],pp236[248],pp237[248],pp238[248],pp239[248],pp240[248],pp241[248],pp242[248],pp243[248],pp244[248]};
    CLA_474 KS_228(s228, c228, in228_1, in228_2);
    wire[471:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {pp7[13],pp6[15],pp5[17],pp4[19],pp3[21],pp2[23],pp0[26],s225[11],pp18[10],pp18[11],pp18[12],pp18[13],pp20[12],pp22[11],pp24[10],s225[19],s226[19],s227[19],s228[19],s228[20],s228[21],s228[22],s228[23],s228[24],s228[25],s228[26],s228[27],s228[28],s228[29],s228[30],s228[31],s228[32],s228[33],s228[34],s228[35],s228[36],s228[37],s228[38],s228[39],s228[40],s228[41],s228[42],s228[43],s228[44],s228[45],s228[46],s228[47],s228[48],s228[49],s228[50],s228[51],s228[52],s228[53],s228[54],s228[55],s228[56],s228[57],s228[58],s228[59],s228[60],s228[61],s228[62],s228[63],s228[64],s228[65],s228[66],s228[67],s228[68],s228[69],s228[70],s228[71],s228[72],s228[73],s228[74],s228[75],s228[76],s228[77],s228[78],s228[79],s228[80],s228[81],s227[83],s225[86],s223[41],s221[44],s219[47],s217[50],s215[53],s213[56],s211[59],s211[60],s211[61],s211[62],s211[63],s211[64],s211[65],s210[67],s209[69],s208[71],s228[100],s228[101],s228[102],s228[103],s228[104],s228[105],s228[106],s228[107],s228[108],s228[109],s228[110],s228[111],s228[112],s228[113],s228[114],s228[115],s228[116],s228[117],s228[118],s228[119],s228[120],s228[121],s228[122],s228[123],s228[124],s228[125],s228[126],s228[127],s228[128],s228[129],s228[130],s228[131],s228[132],s228[133],s228[134],s228[135],s228[136],s228[137],s228[138],s228[139],s228[140],s228[141],s228[142],s228[143],s228[144],s228[145],s228[146],s228[147],s228[148],s228[149],s228[150],s228[151],s228[152],s228[153],s228[154],s228[155],s228[156],s228[157],s228[158],s228[159],s228[160],s228[161],s228[162],s228[163],s228[164],s228[165],s228[166],s228[167],s228[168],s228[169],s228[170],s228[171],s228[172],s228[173],s228[174],s228[175],s228[176],s228[177],s228[178],s228[179],s228[180],s228[181],s228[182],s228[183],s228[184],s228[185],s228[186],s228[187],s228[188],s228[189],s228[190],s228[191],s228[192],s228[193],s228[194],s228[195],s228[196],s228[197],s228[198],s228[199],s228[200],s228[201],s228[202],s228[203],s228[204],s228[205],s228[206],s228[207],s228[208],s228[209],s228[210],s228[211],s228[212],s228[213],s228[214],s228[215],s228[216],s228[217],s228[218],s228[219],s228[220],s228[221],s228[222],s228[223],s228[224],s228[225],s228[226],s228[227],s228[228],s228[229],s228[230],s228[231],s228[232],s228[233],s228[234],s228[235],s228[236],s228[237],s228[238],s228[239],s228[240],s228[241],s228[242],s228[243],s228[244],s228[245],s228[246],s228[247],s228[248],s228[249],s228[250],s228[251],s228[252],s228[253],s228[254],s228[255],s228[256],s228[257],s228[258],s228[259],s228[260],s228[261],s228[262],s228[263],s228[264],s228[265],s228[266],s228[267],s228[268],s228[269],s228[270],s228[271],s228[272],s228[273],s228[274],s228[275],s228[276],s228[277],s228[278],s228[279],s228[280],s228[281],s228[282],s228[283],s228[284],s228[285],s228[286],s228[287],s228[288],s228[289],s228[290],s228[291],s228[292],s228[293],s228[294],s228[295],s228[296],s228[297],s228[298],s228[299],s228[300],s228[301],s228[302],s228[303],s228[304],s228[305],s228[306],s228[307],s228[308],s228[309],s228[310],s228[311],s228[312],s228[313],s228[314],s228[315],s228[316],s228[317],s228[318],s228[319],s228[320],s228[321],s228[322],s228[323],s228[324],s228[325],s228[326],s228[327],s228[328],s228[329],s228[330],s228[331],s228[332],s228[333],s228[334],s228[335],s228[336],s228[337],s228[338],s228[339],s227[341],s226[343],s225[345],s224[299],s223[301],s222[303],s221[305],s220[307],s219[309],s218[311],s217[313],s216[315],s215[317],s214[319],s213[321],s212[323],s211[325],s210[327],s209[329],s208[331],s207[333],s206[335],s205[337],s204[339],s203[341],s202[343],s202[344],s202[345],s202[346],s202[347],s202[348],s202[349],s202[350],s202[351],s202[352],s202[353],s202[354],s202[355],s202[356],s202[357],s202[358],s202[359],s202[360],s202[361],s202[362],s202[363],s202[364],s202[365],s202[366],s202[367],s202[368],s202[369],s202[370],s202[371],s202[372],s202[373],s202[374],s202[375],s202[376],s202[377],s202[378],s202[379],s202[380],s202[381],s202[382],s202[383],s202[384],s202[385],s202[386],s202[387],s202[388],s202[389],s202[390],s202[391],s202[392],s202[393],s202[394],s202[395],s202[396],s202[397],s202[398],s202[399],s202[400],s202[401],s202[402],s202[403],s202[404],s202[405],s202[406],s202[407],s201[409],s200[411],s199[413],s198[415],s197[417],s196[419],s195[421],s194[423],s193[425],pp255[203],pp254[205],pp253[207],pp252[209],pp251[211],pp250[213],pp249[215],pp248[217],pp247[219],pp246[221],pp245[223],pp244[225],pp243[227],pp242[229],pp241[231],pp240[233],pp239[235],pp238[237],pp237[239],pp236[241],pp235[243],pp234[245],pp233[247],pp234[247],pp235[247],pp236[247],pp237[247],pp238[247],pp239[247],pp240[247],pp241[247],pp242[247],pp243[247],pp244[247]};
    assign in229_2 = {pp8[12],pp7[14],pp6[16],pp5[18],pp4[20],pp3[22],pp1[25],s226[10],s225[12],pp19[10],pp19[11],pp19[12],pp21[11],pp23[10],s225[18],s226[18],s227[18],s228[18],pp0[38],pp1[38],pp2[38],pp3[38],pp3[39],pp3[40],pp3[41],pp3[42],pp3[43],pp3[44],pp3[45],pp3[46],pp3[47],pp3[48],pp3[49],pp3[50],pp3[51],pp3[52],pp3[53],pp3[54],pp3[55],pp3[56],pp3[57],pp3[58],pp3[59],pp3[60],pp3[61],pp3[62],pp3[63],pp3[64],pp3[65],pp3[66],pp3[67],pp3[68],pp3[69],pp3[70],pp3[71],pp3[72],pp3[73],pp3[74],pp3[75],pp3[76],pp3[77],pp3[78],pp3[79],pp3[80],pp3[81],pp3[82],pp3[83],pp3[84],pp3[85],pp3[86],pp3[87],pp3[88],pp3[89],pp3[90],pp3[91],pp3[92],pp3[93],pp3[94],pp3[95],pp3[96],pp2[98],s228[82],s226[85],s224[40],s222[43],s220[46],s218[49],s216[52],s214[55],s212[58],s212[59],s212[60],s212[61],s212[62],s212[63],s212[64],s211[66],s210[68],s209[70],s208[72],s208[73],s208[74],s208[75],s208[76],s208[77],s208[78],s208[79],s208[80],s208[81],s208[82],s208[83],s208[84],s208[85],s208[86],s208[87],s208[88],s208[89],s208[90],s209[90],s210[90],s211[90],s212[90],s213[90],s214[90],s215[90],s216[90],s217[90],s218[90],s219[90],s220[90],s221[90],s222[90],s223[90],s224[90],s10[17],s11[17],s12[17],s13[17],s14[17],s15[17],s16[17],s17[17],s18[17],s19[17],s20[17],s21[17],s22[17],s23[17],s24[17],s25[17],s26[17],s27[17],s28[17],s29[17],s30[17],s31[17],s32[17],s33[17],s34[17],s35[17],s36[17],s37[17],s38[17],s39[17],s40[17],s41[17],s42[17],s43[17],s44[17],s45[17],s46[17],s47[17],s48[17],s49[17],s50[17],s51[17],s52[17],s53[17],s54[17],s55[17],s56[17],s57[17],s58[17],s59[17],s60[17],s61[17],s62[17],s63[17],s64[17],s65[17],s66[17],s67[17],s68[17],s69[17],s70[17],s71[17],s72[17],s73[17],s74[17],s75[17],s76[17],s77[17],s78[17],s79[17],s80[17],s81[17],s82[17],s83[17],s83[18],s83[19],s83[20],s83[21],s83[22],s83[23],s83[24],s83[25],s83[26],s83[27],s83[28],s83[29],s83[30],s83[31],s83[32],s83[33],s83[34],s83[35],s83[36],s83[37],s83[38],s83[39],s83[40],s83[41],s83[42],s83[43],s83[44],s83[45],s83[46],s81[49],s79[52],s77[55],s75[58],s74[60],s74[61],s74[62],s74[63],s74[64],s74[65],s74[66],s74[67],s74[68],s74[69],s74[70],s74[71],s74[72],s74[73],s74[74],s74[75],s74[76],s74[77],s74[78],s74[79],s74[80],s74[81],s74[82],s74[83],s74[84],s73[86],s72[88],s71[90],s70[92],s69[94],s68[96],s67[98],s9[157],s7[160],s5[163],s3[166],s1[169],s70[101],s69[103],s68[105],s67[107],s66[109],s65[111],s64[113],s63[115],s62[117],s61[119],s60[121],s59[123],s58[125],s57[127],s56[129],s55[131],s54[133],s53[135],s52[137],s51[139],s50[141],s49[143],s48[145],s47[147],s46[149],s45[151],s44[153],s43[155],s42[157],s41[159],s40[161],s39[163],s38[165],s37[167],s36[169],s35[171],s34[173],s33[175],s32[177],s31[179],s30[181],s29[183],s28[185],s27[187],s26[189],s25[191],s24[193],s23[195],s22[197],s21[199],s20[201],s19[203],s18[205],s17[207],s16[209],s15[211],s14[213],s13[215],s12[217],s11[219],s10[221],s228[340],s227[342],s226[344],s225[346],s224[300],s223[302],s222[304],s221[306],s220[308],s219[310],s218[312],s217[314],s216[316],s215[318],s214[320],s213[322],s212[324],s211[326],s210[328],s209[330],s208[332],s207[334],s206[336],s205[338],s204[340],s203[342],s203[343],s203[344],s203[345],s203[346],s203[347],s203[348],s203[349],s203[350],s203[351],s203[352],s203[353],s203[354],s203[355],s203[356],s203[357],s203[358],s203[359],s203[360],s203[361],s203[362],s203[363],s203[364],s203[365],s203[366],s203[367],s203[368],s203[369],s203[370],s203[371],s203[372],s203[373],s203[374],s203[375],s203[376],s203[377],s203[378],s203[379],s203[380],s203[381],s203[382],s203[383],s203[384],s203[385],s203[386],s203[387],s203[388],s203[389],s203[390],s203[391],s203[392],s203[393],s203[394],s203[395],s203[396],s203[397],s203[398],s203[399],s203[400],s203[401],s203[402],s203[403],s203[404],s203[405],s203[406],s202[408],s201[410],s200[412],s199[414],s198[416],s197[418],s196[420],s195[422],s194[424],s193[426],pp255[204],pp254[206],pp253[208],pp252[210],pp251[212],pp250[214],pp249[216],pp248[218],pp247[220],pp246[222],pp245[224],pp244[226],pp243[228],pp242[230],pp241[232],pp240[234],pp239[236],pp238[238],pp237[240],pp236[242],pp235[244],pp234[246],pp235[246],pp236[246],pp237[246],pp238[246],pp239[246],pp240[246],pp241[246],pp242[246],pp243[246],pp244[246],pp245[246]};
    CLA_472 KS_229(s229, c229, in229_1, in229_2);
    wire[469:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp8[13],pp7[15],pp6[17],pp5[19],pp4[21],pp2[24],pp0[27],s226[11],s225[13],pp20[10],pp20[11],pp22[10],s225[17],s226[17],s227[17],s228[17],s229[17],s229[18],s229[19],s229[20],s229[21],s229[22],s229[23],s229[24],s229[25],s229[26],s229[27],s229[28],s229[29],s229[30],s229[31],s229[32],s229[33],s229[34],s229[35],s229[36],s229[37],s229[38],s229[39],s229[40],s229[41],s229[42],s229[43],s229[44],s229[45],s229[46],s229[47],s229[48],s229[49],s229[50],s229[51],s229[52],s229[53],s229[54],s229[55],s229[56],s229[57],s229[58],s229[59],s229[60],s229[61],s229[62],s229[63],s229[64],s229[65],s229[66],s229[67],s229[68],s229[69],s229[70],s229[71],s229[72],s229[73],s229[74],s229[75],s229[76],s229[77],s229[78],s229[79],s229[80],s229[81],s227[84],s225[87],s223[42],s221[45],s219[48],s217[51],s215[54],s213[57],s213[58],s213[59],s213[60],s213[61],s213[62],s213[63],s212[65],s211[67],s210[69],s209[71],s229[100],s229[101],s229[102],s229[103],s229[104],s229[105],s229[106],s229[107],s229[108],s229[109],s229[110],s229[111],s229[112],s229[113],s229[114],s229[115],s229[116],s229[117],s229[118],s229[119],s229[120],s229[121],s229[122],s229[123],s229[124],s229[125],s229[126],s229[127],s229[128],s229[129],s229[130],s229[131],s229[132],s229[133],s229[134],s229[135],s229[136],s229[137],s229[138],s229[139],s229[140],s229[141],s229[142],s229[143],s229[144],s229[145],s229[146],s229[147],s229[148],s229[149],s229[150],s229[151],s229[152],s229[153],s229[154],s229[155],s229[156],s229[157],s229[158],s229[159],s229[160],s229[161],s229[162],s229[163],s229[164],s229[165],s229[166],s229[167],s229[168],s229[169],s229[170],s229[171],s229[172],s229[173],s229[174],s229[175],s229[176],s229[177],s229[178],s229[179],s229[180],s229[181],s229[182],s229[183],s229[184],s229[185],s229[186],s229[187],s229[188],s229[189],s229[190],s229[191],s229[192],s229[193],s229[194],s229[195],s229[196],s229[197],s229[198],s229[199],s229[200],s229[201],s229[202],s229[203],s229[204],s229[205],s229[206],s229[207],s229[208],s229[209],s229[210],s229[211],s229[212],s229[213],s229[214],s229[215],s229[216],s229[217],s229[218],s229[219],s229[220],s229[221],s229[222],s229[223],s229[224],s229[225],s229[226],s229[227],s229[228],s229[229],s229[230],s229[231],s229[232],s229[233],s229[234],s229[235],s229[236],s229[237],s229[238],s229[239],s229[240],s229[241],s229[242],s229[243],s229[244],s229[245],s229[246],s229[247],s229[248],s229[249],s229[250],s229[251],s229[252],s229[253],s229[254],s229[255],s229[256],s229[257],s229[258],s229[259],s229[260],s229[261],s229[262],s229[263],s229[264],s229[265],s229[266],s229[267],s229[268],s229[269],s229[270],s229[271],s229[272],s229[273],s229[274],s229[275],s229[276],s229[277],s229[278],s229[279],s229[280],s229[281],s229[282],s229[283],s229[284],s229[285],s229[286],s229[287],s229[288],s229[289],s229[290],s229[291],s229[292],s229[293],s229[294],s229[295],s229[296],s229[297],s229[298],s229[299],s229[300],s229[301],s229[302],s229[303],s229[304],s229[305],s229[306],s229[307],s229[308],s229[309],s229[310],s229[311],s229[312],s229[313],s229[314],s229[315],s229[316],s229[317],s229[318],s229[319],s229[320],s229[321],s229[322],s229[323],s229[324],s229[325],s229[326],s229[327],s229[328],s229[329],s229[330],s229[331],s229[332],s229[333],s229[334],s229[335],s229[336],s229[337],s229[338],s229[339],s228[341],s227[343],s226[345],s225[347],s224[301],s223[303],s222[305],s221[307],s220[309],s219[311],s218[313],s217[315],s216[317],s215[319],s214[321],s213[323],s212[325],s211[327],s210[329],s209[331],s208[333],s207[335],s206[337],s205[339],s204[341],s204[342],s204[343],s204[344],s204[345],s204[346],s204[347],s204[348],s204[349],s204[350],s204[351],s204[352],s204[353],s204[354],s204[355],s204[356],s204[357],s204[358],s204[359],s204[360],s204[361],s204[362],s204[363],s204[364],s204[365],s204[366],s204[367],s204[368],s204[369],s204[370],s204[371],s204[372],s204[373],s204[374],s204[375],s204[376],s204[377],s204[378],s204[379],s204[380],s204[381],s204[382],s204[383],s204[384],s204[385],s204[386],s204[387],s204[388],s204[389],s204[390],s204[391],s204[392],s204[393],s204[394],s204[395],s204[396],s204[397],s204[398],s204[399],s204[400],s204[401],s204[402],s204[403],s204[404],s204[405],s203[407],s202[409],s201[411],s200[413],s199[415],s198[417],s197[419],s196[421],s195[423],s194[425],s193[427],pp255[205],pp254[207],pp253[209],pp252[211],pp251[213],pp250[215],pp249[217],pp248[219],pp247[221],pp246[223],pp245[225],pp244[227],pp243[229],pp242[231],pp241[233],pp240[235],pp239[237],pp238[239],pp237[241],pp236[243],pp235[245],pp236[245],pp237[245],pp238[245],pp239[245],pp240[245],pp241[245],pp242[245],pp243[245],pp244[245],pp245[245]};
    assign in230_2 = {pp9[12],pp8[14],pp7[16],pp6[18],pp5[20],pp3[23],pp1[26],s227[10],s226[12],s225[14],pp21[10],s225[16],s226[16],s227[16],s228[16],s229[16],pp0[37],pp1[37],pp2[37],pp3[37],pp4[37],pp4[38],pp4[39],pp4[40],pp4[41],pp4[42],pp4[43],pp4[44],pp4[45],pp4[46],pp4[47],pp4[48],pp4[49],pp4[50],pp4[51],pp4[52],pp4[53],pp4[54],pp4[55],pp4[56],pp4[57],pp4[58],pp4[59],pp4[60],pp4[61],pp4[62],pp4[63],pp4[64],pp4[65],pp4[66],pp4[67],pp4[68],pp4[69],pp4[70],pp4[71],pp4[72],pp4[73],pp4[74],pp4[75],pp4[76],pp4[77],pp4[78],pp4[79],pp4[80],pp4[81],pp4[82],pp4[83],pp4[84],pp4[85],pp4[86],pp4[87],pp4[88],pp4[89],pp4[90],pp4[91],pp4[92],pp4[93],pp4[94],pp4[95],pp3[97],pp2[99],s228[83],s226[86],s224[41],s222[44],s220[47],s218[50],s216[53],s214[56],s214[57],s214[58],s214[59],s214[60],s214[61],s214[62],s213[64],s212[66],s211[68],s210[70],s209[72],s209[73],s209[74],s209[75],s209[76],s209[77],s209[78],s209[79],s209[80],s209[81],s209[82],s209[83],s209[84],s209[85],s209[86],s209[87],s209[88],s209[89],s210[89],s211[89],s212[89],s213[89],s214[89],s215[89],s216[89],s217[89],s218[89],s219[89],s220[89],s221[89],s222[89],s223[89],s224[89],s10[16],s11[16],s12[16],s13[16],s14[16],s15[16],s16[16],s17[16],s18[16],s19[16],s20[16],s21[16],s22[16],s23[16],s24[16],s25[16],s26[16],s27[16],s28[16],s29[16],s30[16],s31[16],s32[16],s33[16],s34[16],s35[16],s36[16],s37[16],s38[16],s39[16],s40[16],s41[16],s42[16],s43[16],s44[16],s45[16],s46[16],s47[16],s48[16],s49[16],s50[16],s51[16],s52[16],s53[16],s54[16],s55[16],s56[16],s57[16],s58[16],s59[16],s60[16],s61[16],s62[16],s63[16],s64[16],s65[16],s66[16],s67[16],s68[16],s69[16],s70[16],s71[16],s72[16],s73[16],s74[16],s75[16],s76[16],s77[16],s78[16],s79[16],s80[16],s81[16],s82[16],s83[16],s84[16],s84[17],s84[18],s84[19],s84[20],s84[21],s84[22],s84[23],s84[24],s84[25],s84[26],s84[27],s84[28],s84[29],s84[30],s84[31],s84[32],s84[33],s84[34],s84[35],s84[36],s84[37],s84[38],s84[39],s84[40],s84[41],s84[42],s84[43],s84[44],s84[45],s82[48],s80[51],s78[54],s76[57],s75[59],s75[60],s75[61],s75[62],s75[63],s75[64],s75[65],s75[66],s75[67],s75[68],s75[69],s75[70],s75[71],s75[72],s75[73],s75[74],s75[75],s75[76],s75[77],s75[78],s75[79],s75[80],s75[81],s75[82],s75[83],s74[85],s73[87],s72[89],s71[91],s70[93],s69[95],s68[97],s67[99],s8[159],s6[162],s4[165],s2[168],s71[100],s70[102],s69[104],s68[106],s67[108],s66[110],s65[112],s64[114],s63[116],s62[118],s61[120],s60[122],s59[124],s58[126],s57[128],s56[130],s55[132],s54[134],s53[136],s52[138],s51[140],s50[142],s49[144],s48[146],s47[148],s46[150],s45[152],s44[154],s43[156],s42[158],s41[160],s40[162],s39[164],s38[166],s37[168],s36[170],s35[172],s34[174],s33[176],s32[178],s31[180],s30[182],s29[184],s28[186],s27[188],s26[190],s25[192],s24[194],s23[196],s22[198],s21[200],s20[202],s19[204],s18[206],s17[208],s16[210],s15[212],s14[214],s13[216],s12[218],s11[220],s10[222],s229[340],s228[342],s227[344],s226[346],s225[348],s224[302],s223[304],s222[306],s221[308],s220[310],s219[312],s218[314],s217[316],s216[318],s215[320],s214[322],s213[324],s212[326],s211[328],s210[330],s209[332],s208[334],s207[336],s206[338],s205[340],s205[341],s205[342],s205[343],s205[344],s205[345],s205[346],s205[347],s205[348],s205[349],s205[350],s205[351],s205[352],s205[353],s205[354],s205[355],s205[356],s205[357],s205[358],s205[359],s205[360],s205[361],s205[362],s205[363],s205[364],s205[365],s205[366],s205[367],s205[368],s205[369],s205[370],s205[371],s205[372],s205[373],s205[374],s205[375],s205[376],s205[377],s205[378],s205[379],s205[380],s205[381],s205[382],s205[383],s205[384],s205[385],s205[386],s205[387],s205[388],s205[389],s205[390],s205[391],s205[392],s205[393],s205[394],s205[395],s205[396],s205[397],s205[398],s205[399],s205[400],s205[401],s205[402],s205[403],s205[404],s204[406],s203[408],s202[410],s201[412],s200[414],s199[416],s198[418],s197[420],s196[422],s195[424],s194[426],s193[428],pp255[206],pp254[208],pp253[210],pp252[212],pp251[214],pp250[216],pp249[218],pp248[220],pp247[222],pp246[224],pp245[226],pp244[228],pp243[230],pp242[232],pp241[234],pp240[236],pp239[238],pp238[240],pp237[242],pp236[244],pp237[244],pp238[244],pp239[244],pp240[244],pp241[244],pp242[244],pp243[244],pp244[244],pp245[244],pp246[244]};
    CLA_470 KS_230(s230, c230, in230_1, in230_2);
    wire[467:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp9[13],pp8[15],pp7[17],pp6[19],pp4[22],pp2[25],pp0[28],s227[11],s226[13],s225[15],s226[15],s227[15],s228[15],s229[15],s230[15],s230[16],s230[17],s230[18],s230[19],s230[20],s230[21],s230[22],s230[23],s230[24],s230[25],s230[26],s230[27],s230[28],s230[29],s230[30],s230[31],s230[32],s230[33],s230[34],s230[35],s230[36],s230[37],s230[38],s230[39],s230[40],s230[41],s230[42],s230[43],s230[44],s230[45],s230[46],s230[47],s230[48],s230[49],s230[50],s230[51],s230[52],s230[53],s230[54],s230[55],s230[56],s230[57],s230[58],s230[59],s230[60],s230[61],s230[62],s230[63],s230[64],s230[65],s230[66],s230[67],s230[68],s230[69],s230[70],s230[71],s230[72],s230[73],s230[74],s230[75],s230[76],s230[77],s230[78],s230[79],s230[80],s229[82],s227[85],s225[88],s223[43],s221[46],s219[49],s217[52],s215[55],s215[56],s215[57],s215[58],s215[59],s215[60],s215[61],s214[63],s213[65],s212[67],s211[69],s210[71],s230[100],s230[101],s230[102],s230[103],s230[104],s230[105],s230[106],s230[107],s230[108],s230[109],s230[110],s230[111],s230[112],s230[113],s230[114],s230[115],s230[116],s230[117],s230[118],s230[119],s230[120],s230[121],s230[122],s230[123],s230[124],s230[125],s230[126],s230[127],s230[128],s230[129],s230[130],s230[131],s230[132],s230[133],s230[134],s230[135],s230[136],s230[137],s230[138],s230[139],s230[140],s230[141],s230[142],s230[143],s230[144],s230[145],s230[146],s230[147],s230[148],s230[149],s230[150],s230[151],s230[152],s230[153],s230[154],s230[155],s230[156],s230[157],s230[158],s230[159],s230[160],s230[161],s230[162],s230[163],s230[164],s230[165],s230[166],s230[167],s230[168],s230[169],s230[170],s230[171],s230[172],s230[173],s230[174],s230[175],s230[176],s230[177],s230[178],s230[179],s230[180],s230[181],s230[182],s230[183],s230[184],s230[185],s230[186],s230[187],s230[188],s230[189],s230[190],s230[191],s230[192],s230[193],s230[194],s230[195],s230[196],s230[197],s230[198],s230[199],s230[200],s230[201],s230[202],s230[203],s230[204],s230[205],s230[206],s230[207],s230[208],s230[209],s230[210],s230[211],s230[212],s230[213],s230[214],s230[215],s230[216],s230[217],s230[218],s230[219],s230[220],s230[221],s230[222],s230[223],s230[224],s230[225],s230[226],s230[227],s230[228],s230[229],s230[230],s230[231],s230[232],s230[233],s230[234],s230[235],s230[236],s230[237],s230[238],s230[239],s230[240],s230[241],s230[242],s230[243],s230[244],s230[245],s230[246],s230[247],s230[248],s230[249],s230[250],s230[251],s230[252],s230[253],s230[254],s230[255],s230[256],s230[257],s230[258],s230[259],s230[260],s230[261],s230[262],s230[263],s230[264],s230[265],s230[266],s230[267],s230[268],s230[269],s230[270],s230[271],s230[272],s230[273],s230[274],s230[275],s230[276],s230[277],s230[278],s230[279],s230[280],s230[281],s230[282],s230[283],s230[284],s230[285],s230[286],s230[287],s230[288],s230[289],s230[290],s230[291],s230[292],s230[293],s230[294],s230[295],s230[296],s230[297],s230[298],s230[299],s230[300],s230[301],s230[302],s230[303],s230[304],s230[305],s230[306],s230[307],s230[308],s230[309],s230[310],s230[311],s230[312],s230[313],s230[314],s230[315],s230[316],s230[317],s230[318],s230[319],s230[320],s230[321],s230[322],s230[323],s230[324],s230[325],s230[326],s230[327],s230[328],s230[329],s230[330],s230[331],s230[332],s230[333],s230[334],s230[335],s230[336],s230[337],s230[338],s230[339],s229[341],s228[343],s227[345],s226[347],s225[349],s224[303],s223[305],s222[307],s221[309],s220[311],s219[313],s218[315],s217[317],s216[319],s215[321],s214[323],s213[325],s212[327],s211[329],s210[331],s209[333],s208[335],s207[337],s206[339],s206[340],s206[341],s206[342],s206[343],s206[344],s206[345],s206[346],s206[347],s206[348],s206[349],s206[350],s206[351],s206[352],s206[353],s206[354],s206[355],s206[356],s206[357],s206[358],s206[359],s206[360],s206[361],s206[362],s206[363],s206[364],s206[365],s206[366],s206[367],s206[368],s206[369],s206[370],s206[371],s206[372],s206[373],s206[374],s206[375],s206[376],s206[377],s206[378],s206[379],s206[380],s206[381],s206[382],s206[383],s206[384],s206[385],s206[386],s206[387],s206[388],s206[389],s206[390],s206[391],s206[392],s206[393],s206[394],s206[395],s206[396],s206[397],s206[398],s206[399],s206[400],s206[401],s206[402],s206[403],s205[405],s204[407],s203[409],s202[411],s201[413],s200[415],s199[417],s198[419],s197[421],s196[423],s195[425],s194[427],s193[429],pp255[207],pp254[209],pp253[211],pp252[213],pp251[215],pp250[217],pp249[219],pp248[221],pp247[223],pp246[225],pp245[227],pp244[229],pp243[231],pp242[233],pp241[235],pp240[237],pp239[239],pp238[241],pp237[243],pp238[243],pp239[243],pp240[243],pp241[243],pp242[243],pp243[243],pp244[243],pp245[243],pp246[243]};
    assign in231_2 = {pp13[9],pp9[14],pp8[16],pp7[18],pp5[21],pp3[24],pp1[27],s228[10],s227[12],s226[14],s227[14],s228[14],s229[14],s230[14],pp0[36],pp1[36],pp2[36],pp3[36],pp4[36],pp5[36],pp5[37],pp5[38],pp5[39],pp5[40],pp5[41],pp5[42],pp5[43],pp5[44],pp5[45],pp5[46],pp5[47],pp5[48],pp5[49],pp5[50],pp5[51],pp5[52],pp5[53],pp5[54],pp5[55],pp5[56],pp5[57],pp5[58],pp5[59],pp5[60],pp5[61],pp5[62],pp5[63],pp5[64],pp5[65],pp5[66],pp5[67],pp5[68],pp5[69],pp5[70],pp5[71],pp5[72],pp5[73],pp5[74],pp5[75],pp5[76],pp5[77],pp5[78],pp5[79],pp5[80],pp5[81],pp5[82],pp5[83],pp5[84],pp5[85],pp5[86],pp5[87],pp5[88],pp5[89],pp5[90],pp5[91],pp5[92],pp5[93],pp5[94],pp4[96],pp3[98],s230[81],s228[84],s226[87],s224[42],s222[45],s220[48],s218[51],s216[54],s216[55],s216[56],s216[57],s216[58],s216[59],s216[60],s215[62],s214[64],s213[66],s212[68],s211[70],s210[72],s210[73],s210[74],s210[75],s210[76],s210[77],s210[78],s210[79],s210[80],s210[81],s210[82],s210[83],s210[84],s210[85],s210[86],s210[87],s210[88],s211[88],s212[88],s213[88],s214[88],s215[88],s216[88],s217[88],s218[88],s219[88],s220[88],s221[88],s222[88],s223[88],s224[88],s10[15],s11[15],s12[15],s13[15],s14[15],s15[15],s16[15],s17[15],s18[15],s19[15],s20[15],s21[15],s22[15],s23[15],s24[15],s25[15],s26[15],s27[15],s28[15],s29[15],s30[15],s31[15],s32[15],s33[15],s34[15],s35[15],s36[15],s37[15],s38[15],s39[15],s40[15],s41[15],s42[15],s43[15],s44[15],s45[15],s46[15],s47[15],s48[15],s49[15],s50[15],s51[15],s52[15],s53[15],s54[15],s55[15],s56[15],s57[15],s58[15],s59[15],s60[15],s61[15],s62[15],s63[15],s64[15],s65[15],s66[15],s67[15],s68[15],s69[15],s70[15],s71[15],s72[15],s73[15],s74[15],s75[15],s76[15],s77[15],s78[15],s79[15],s80[15],s81[15],s82[15],s83[15],s84[15],s85[15],s85[16],s85[17],s85[18],s85[19],s85[20],s85[21],s85[22],s85[23],s85[24],s85[25],s85[26],s85[27],s85[28],s85[29],s85[30],s85[31],s85[32],s85[33],s85[34],s85[35],s85[36],s85[37],s85[38],s85[39],s85[40],s85[41],s85[42],s85[43],s85[44],s83[47],s81[50],s79[53],s77[56],s76[58],s76[59],s76[60],s76[61],s76[62],s76[63],s76[64],s76[65],s76[66],s76[67],s76[68],s76[69],s76[70],s76[71],s76[72],s76[73],s76[74],s76[75],s76[76],s76[77],s76[78],s76[79],s76[80],s76[81],s76[82],s75[84],s74[86],s73[88],s72[90],s71[92],s70[94],s69[96],s68[98],s9[158],s7[161],s5[164],s3[167],s1[170],s71[101],s70[103],s69[105],s68[107],s67[109],s66[111],s65[113],s64[115],s63[117],s62[119],s61[121],s60[123],s59[125],s58[127],s57[129],s56[131],s55[133],s54[135],s53[137],s52[139],s51[141],s50[143],s49[145],s48[147],s47[149],s46[151],s45[153],s44[155],s43[157],s42[159],s41[161],s40[163],s39[165],s38[167],s37[169],s36[171],s35[173],s34[175],s33[177],s32[179],s31[181],s30[183],s29[185],s28[187],s27[189],s26[191],s25[193],s24[195],s23[197],s22[199],s21[201],s20[203],s19[205],s18[207],s17[209],s16[211],s15[213],s14[215],s13[217],s12[219],s11[221],s10[223],s230[340],s229[342],s228[344],s227[346],s226[348],s225[350],s224[304],s223[306],s222[308],s221[310],s220[312],s219[314],s218[316],s217[318],s216[320],s215[322],s214[324],s213[326],s212[328],s211[330],s210[332],s209[334],s208[336],s207[338],s207[339],s207[340],s207[341],s207[342],s207[343],s207[344],s207[345],s207[346],s207[347],s207[348],s207[349],s207[350],s207[351],s207[352],s207[353],s207[354],s207[355],s207[356],s207[357],s207[358],s207[359],s207[360],s207[361],s207[362],s207[363],s207[364],s207[365],s207[366],s207[367],s207[368],s207[369],s207[370],s207[371],s207[372],s207[373],s207[374],s207[375],s207[376],s207[377],s207[378],s207[379],s207[380],s207[381],s207[382],s207[383],s207[384],s207[385],s207[386],s207[387],s207[388],s207[389],s207[390],s207[391],s207[392],s207[393],s207[394],s207[395],s207[396],s207[397],s207[398],s207[399],s207[400],s207[401],s207[402],s206[404],s205[406],s204[408],s203[410],s202[412],s201[414],s200[416],s199[418],s198[420],s197[422],s196[424],s195[426],s194[428],s193[430],pp255[208],pp254[210],pp253[212],pp252[214],pp251[216],pp250[218],pp249[220],pp248[222],pp247[224],pp246[226],pp245[228],pp244[230],pp243[232],pp242[234],pp241[236],pp240[238],pp239[240],pp238[242],pp239[242],pp240[242],pp241[242],pp242[242],pp243[242],pp244[242],pp245[242],pp246[242],pp247[242]};
    CLA_468 KS_231(s231, c231, in231_1, in231_2);
    wire[465:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {pp14[9],pp9[15],pp8[17],pp6[20],pp4[23],pp2[26],pp0[29],s228[11],s227[13],s228[13],s229[13],s230[13],s231[13],s231[14],s231[15],s231[16],s231[17],s231[18],s231[19],s231[20],s231[21],s231[22],s231[23],s231[24],s231[25],s231[26],s231[27],s231[28],s231[29],s231[30],s231[31],s231[32],s231[33],s231[34],s231[35],s231[36],s231[37],s231[38],s231[39],s231[40],s231[41],s231[42],s231[43],s231[44],s231[45],s231[46],s231[47],s231[48],s231[49],s231[50],s231[51],s231[52],s231[53],s231[54],s231[55],s231[56],s231[57],s231[58],s231[59],s231[60],s231[61],s231[62],s231[63],s231[64],s231[65],s231[66],s231[67],s231[68],s231[69],s231[70],s231[71],s231[72],s231[73],s231[74],s231[75],s231[76],s231[77],s231[78],s231[79],s231[80],s229[83],s227[86],s225[89],s223[44],s221[47],s219[50],s217[53],s217[54],s217[55],s217[56],s217[57],s217[58],s217[59],s216[61],s215[63],s214[65],s213[67],s212[69],s211[71],s231[100],s231[101],s231[102],s231[103],s231[104],s231[105],s231[106],s231[107],s231[108],s231[109],s231[110],s231[111],s231[112],s231[113],s231[114],s231[115],s231[116],s231[117],s231[118],s231[119],s231[120],s231[121],s231[122],s231[123],s231[124],s231[125],s231[126],s231[127],s231[128],s231[129],s231[130],s231[131],s231[132],s231[133],s231[134],s231[135],s231[136],s231[137],s231[138],s231[139],s231[140],s231[141],s231[142],s231[143],s231[144],s231[145],s231[146],s231[147],s231[148],s231[149],s231[150],s231[151],s231[152],s231[153],s231[154],s231[155],s231[156],s231[157],s231[158],s231[159],s231[160],s231[161],s231[162],s231[163],s231[164],s231[165],s231[166],s231[167],s231[168],s231[169],s231[170],s231[171],s231[172],s231[173],s231[174],s231[175],s231[176],s231[177],s231[178],s231[179],s231[180],s231[181],s231[182],s231[183],s231[184],s231[185],s231[186],s231[187],s231[188],s231[189],s231[190],s231[191],s231[192],s231[193],s231[194],s231[195],s231[196],s231[197],s231[198],s231[199],s231[200],s231[201],s231[202],s231[203],s231[204],s231[205],s231[206],s231[207],s231[208],s231[209],s231[210],s231[211],s231[212],s231[213],s231[214],s231[215],s231[216],s231[217],s231[218],s231[219],s231[220],s231[221],s231[222],s231[223],s231[224],s231[225],s231[226],s231[227],s231[228],s231[229],s231[230],s231[231],s231[232],s231[233],s231[234],s231[235],s231[236],s231[237],s231[238],s231[239],s231[240],s231[241],s231[242],s231[243],s231[244],s231[245],s231[246],s231[247],s231[248],s231[249],s231[250],s231[251],s231[252],s231[253],s231[254],s231[255],s231[256],s231[257],s231[258],s231[259],s231[260],s231[261],s231[262],s231[263],s231[264],s231[265],s231[266],s231[267],s231[268],s231[269],s231[270],s231[271],s231[272],s231[273],s231[274],s231[275],s231[276],s231[277],s231[278],s231[279],s231[280],s231[281],s231[282],s231[283],s231[284],s231[285],s231[286],s231[287],s231[288],s231[289],s231[290],s231[291],s231[292],s231[293],s231[294],s231[295],s231[296],s231[297],s231[298],s231[299],s231[300],s231[301],s231[302],s231[303],s231[304],s231[305],s231[306],s231[307],s231[308],s231[309],s231[310],s231[311],s231[312],s231[313],s231[314],s231[315],s231[316],s231[317],s231[318],s231[319],s231[320],s231[321],s231[322],s231[323],s231[324],s231[325],s231[326],s231[327],s231[328],s231[329],s231[330],s231[331],s231[332],s231[333],s231[334],s231[335],s231[336],s231[337],s231[338],s231[339],s230[341],s229[343],s228[345],s227[347],s226[349],s225[351],s224[305],s223[307],s222[309],s221[311],s220[313],s219[315],s218[317],s217[319],s216[321],s215[323],s214[325],s213[327],s212[329],s211[331],s210[333],s209[335],s208[337],s208[338],s208[339],s208[340],s208[341],s208[342],s208[343],s208[344],s208[345],s208[346],s208[347],s208[348],s208[349],s208[350],s208[351],s208[352],s208[353],s208[354],s208[355],s208[356],s208[357],s208[358],s208[359],s208[360],s208[361],s208[362],s208[363],s208[364],s208[365],s208[366],s208[367],s208[368],s208[369],s208[370],s208[371],s208[372],s208[373],s208[374],s208[375],s208[376],s208[377],s208[378],s208[379],s208[380],s208[381],s208[382],s208[383],s208[384],s208[385],s208[386],s208[387],s208[388],s208[389],s208[390],s208[391],s208[392],s208[393],s208[394],s208[395],s208[396],s208[397],s208[398],s208[399],s208[400],s208[401],s207[403],s206[405],s205[407],s204[409],s203[411],s202[413],s201[415],s200[417],s199[419],s198[421],s197[423],s196[425],s195[427],s194[429],s193[431],pp255[209],pp254[211],pp253[213],pp252[215],pp251[217],pp250[219],pp249[221],pp248[223],pp247[225],pp246[227],pp245[229],pp244[231],pp243[233],pp242[235],pp241[237],pp240[239],pp239[241],pp240[241],pp241[241],pp242[241],pp243[241],pp244[241],pp245[241],pp246[241],pp247[241]};
    assign in232_2 = {pp15[8],pp15[9],pp9[16],pp7[19],pp5[22],pp3[25],pp1[28],s229[10],s228[12],s229[12],s230[12],s231[12],pp0[35],pp1[35],pp2[35],pp3[35],pp4[35],pp5[35],pp6[35],pp6[36],pp6[37],pp6[38],pp6[39],pp6[40],pp6[41],pp6[42],pp6[43],pp6[44],pp6[45],pp6[46],pp6[47],pp6[48],pp6[49],pp6[50],pp6[51],pp6[52],pp6[53],pp6[54],pp6[55],pp6[56],pp6[57],pp6[58],pp6[59],pp6[60],pp6[61],pp6[62],pp6[63],pp6[64],pp6[65],pp6[66],pp6[67],pp6[68],pp6[69],pp6[70],pp6[71],pp6[72],pp6[73],pp6[74],pp6[75],pp6[76],pp6[77],pp6[78],pp6[79],pp6[80],pp6[81],pp6[82],pp6[83],pp6[84],pp6[85],pp6[86],pp6[87],pp6[88],pp6[89],pp6[90],pp6[91],pp6[92],pp6[93],pp5[95],pp4[97],pp3[99],s230[82],s228[85],s226[88],s224[43],s222[46],s220[49],s218[52],s218[53],s218[54],s218[55],s218[56],s218[57],s218[58],s217[60],s216[62],s215[64],s214[66],s213[68],s212[70],s211[72],s211[73],s211[74],s211[75],s211[76],s211[77],s211[78],s211[79],s211[80],s211[81],s211[82],s211[83],s211[84],s211[85],s211[86],s211[87],s212[87],s213[87],s214[87],s215[87],s216[87],s217[87],s218[87],s219[87],s220[87],s221[87],s222[87],s223[87],s224[87],s10[14],s11[14],s12[14],s13[14],s14[14],s15[14],s16[14],s17[14],s18[14],s19[14],s20[14],s21[14],s22[14],s23[14],s24[14],s25[14],s26[14],s27[14],s28[14],s29[14],s30[14],s31[14],s32[14],s33[14],s34[14],s35[14],s36[14],s37[14],s38[14],s39[14],s40[14],s41[14],s42[14],s43[14],s44[14],s45[14],s46[14],s47[14],s48[14],s49[14],s50[14],s51[14],s52[14],s53[14],s54[14],s55[14],s56[14],s57[14],s58[14],s59[14],s60[14],s61[14],s62[14],s63[14],s64[14],s65[14],s66[14],s67[14],s68[14],s69[14],s70[14],s71[14],s72[14],s73[14],s74[14],s75[14],s76[14],s77[14],s78[14],s79[14],s80[14],s81[14],s82[14],s83[14],s84[14],s85[14],s86[14],s86[15],s86[16],s86[17],s86[18],s86[19],s86[20],s86[21],s86[22],s86[23],s86[24],s86[25],s86[26],s86[27],s86[28],s86[29],s86[30],s86[31],s86[32],s86[33],s86[34],s86[35],s86[36],s86[37],s86[38],s86[39],s86[40],s86[41],s86[42],s86[43],s84[46],s82[49],s80[52],s78[55],s77[57],s77[58],s77[59],s77[60],s77[61],s77[62],s77[63],s77[64],s77[65],s77[66],s77[67],s77[68],s77[69],s77[70],s77[71],s77[72],s77[73],s77[74],s77[75],s77[76],s77[77],s77[78],s77[79],s77[80],s77[81],s76[83],s75[85],s74[87],s73[89],s72[91],s71[93],s70[95],s69[97],s68[99],s8[160],s6[163],s4[166],s2[169],s72[100],s71[102],s70[104],s69[106],s68[108],s67[110],s66[112],s65[114],s64[116],s63[118],s62[120],s61[122],s60[124],s59[126],s58[128],s57[130],s56[132],s55[134],s54[136],s53[138],s52[140],s51[142],s50[144],s49[146],s48[148],s47[150],s46[152],s45[154],s44[156],s43[158],s42[160],s41[162],s40[164],s39[166],s38[168],s37[170],s36[172],s35[174],s34[176],s33[178],s32[180],s31[182],s30[184],s29[186],s28[188],s27[190],s26[192],s25[194],s24[196],s23[198],s22[200],s21[202],s20[204],s19[206],s18[208],s17[210],s16[212],s15[214],s14[216],s13[218],s12[220],s11[222],s10[224],s231[340],s230[342],s229[344],s228[346],s227[348],s226[350],s225[352],s224[306],s223[308],s222[310],s221[312],s220[314],s219[316],s218[318],s217[320],s216[322],s215[324],s214[326],s213[328],s212[330],s211[332],s210[334],s209[336],s209[337],s209[338],s209[339],s209[340],s209[341],s209[342],s209[343],s209[344],s209[345],s209[346],s209[347],s209[348],s209[349],s209[350],s209[351],s209[352],s209[353],s209[354],s209[355],s209[356],s209[357],s209[358],s209[359],s209[360],s209[361],s209[362],s209[363],s209[364],s209[365],s209[366],s209[367],s209[368],s209[369],s209[370],s209[371],s209[372],s209[373],s209[374],s209[375],s209[376],s209[377],s209[378],s209[379],s209[380],s209[381],s209[382],s209[383],s209[384],s209[385],s209[386],s209[387],s209[388],s209[389],s209[390],s209[391],s209[392],s209[393],s209[394],s209[395],s209[396],s209[397],s209[398],s209[399],s209[400],s208[402],s207[404],s206[406],s205[408],s204[410],s203[412],s202[414],s201[416],s200[418],s199[420],s198[422],s197[424],s196[426],s195[428],s194[430],s193[432],pp255[210],pp254[212],pp253[214],pp252[216],pp251[218],pp250[220],pp249[222],pp248[224],pp247[226],pp246[228],pp245[230],pp244[232],pp243[234],pp242[236],pp241[238],pp240[240],pp241[240],pp242[240],pp243[240],pp244[240],pp245[240],pp246[240],pp247[240],pp248[240]};
    CLA_466 KS_232(s232, c232, in232_1, in232_2);
    wire[463:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {pp16[8],pp16[9],pp8[18],pp6[21],pp4[24],pp2[27],pp0[30],s229[11],s230[11],s231[11],s232[11],s232[12],s232[13],s232[14],s232[15],s232[16],s232[17],s232[18],s232[19],s232[20],s232[21],s232[22],s232[23],s232[24],s232[25],s232[26],s232[27],s232[28],s232[29],s232[30],s232[31],s232[32],s232[33],s232[34],s232[35],s232[36],s232[37],s232[38],s232[39],s232[40],s232[41],s232[42],s232[43],s232[44],s232[45],s232[46],s232[47],s232[48],s232[49],s232[50],s232[51],s232[52],s232[53],s232[54],s232[55],s232[56],s232[57],s232[58],s232[59],s232[60],s232[61],s232[62],s232[63],s232[64],s232[65],s232[66],s232[67],s232[68],s232[69],s232[70],s232[71],s232[72],s232[73],s232[74],s232[75],s232[76],s232[77],s232[78],s232[79],s231[81],s229[84],s227[87],s225[90],s223[45],s221[48],s219[51],s219[52],s219[53],s219[54],s219[55],s219[56],s219[57],s218[59],s217[61],s216[63],s215[65],s214[67],s213[69],s212[71],s232[100],s232[101],s232[102],s232[103],s232[104],s232[105],s232[106],s232[107],s232[108],s232[109],s232[110],s232[111],s232[112],s232[113],s232[114],s232[115],s232[116],s232[117],s232[118],s232[119],s232[120],s232[121],s232[122],s232[123],s232[124],s232[125],s232[126],s232[127],s232[128],s232[129],s232[130],s232[131],s232[132],s232[133],s232[134],s232[135],s232[136],s232[137],s232[138],s232[139],s232[140],s232[141],s232[142],s232[143],s232[144],s232[145],s232[146],s232[147],s232[148],s232[149],s232[150],s232[151],s232[152],s232[153],s232[154],s232[155],s232[156],s232[157],s232[158],s232[159],s232[160],s232[161],s232[162],s232[163],s232[164],s232[165],s232[166],s232[167],s232[168],s232[169],s232[170],s232[171],s232[172],s232[173],s232[174],s232[175],s232[176],s232[177],s232[178],s232[179],s232[180],s232[181],s232[182],s232[183],s232[184],s232[185],s232[186],s232[187],s232[188],s232[189],s232[190],s232[191],s232[192],s232[193],s232[194],s232[195],s232[196],s232[197],s232[198],s232[199],s232[200],s232[201],s232[202],s232[203],s232[204],s232[205],s232[206],s232[207],s232[208],s232[209],s232[210],s232[211],s232[212],s232[213],s232[214],s232[215],s232[216],s232[217],s232[218],s232[219],s232[220],s232[221],s232[222],s232[223],s232[224],s232[225],s232[226],s232[227],s232[228],s232[229],s232[230],s232[231],s232[232],s232[233],s232[234],s232[235],s232[236],s232[237],s232[238],s232[239],s232[240],s232[241],s232[242],s232[243],s232[244],s232[245],s232[246],s232[247],s232[248],s232[249],s232[250],s232[251],s232[252],s232[253],s232[254],s232[255],s232[256],s232[257],s232[258],s232[259],s232[260],s232[261],s232[262],s232[263],s232[264],s232[265],s232[266],s232[267],s232[268],s232[269],s232[270],s232[271],s232[272],s232[273],s232[274],s232[275],s232[276],s232[277],s232[278],s232[279],s232[280],s232[281],s232[282],s232[283],s232[284],s232[285],s232[286],s232[287],s232[288],s232[289],s232[290],s232[291],s232[292],s232[293],s232[294],s232[295],s232[296],s232[297],s232[298],s232[299],s232[300],s232[301],s232[302],s232[303],s232[304],s232[305],s232[306],s232[307],s232[308],s232[309],s232[310],s232[311],s232[312],s232[313],s232[314],s232[315],s232[316],s232[317],s232[318],s232[319],s232[320],s232[321],s232[322],s232[323],s232[324],s232[325],s232[326],s232[327],s232[328],s232[329],s232[330],s232[331],s232[332],s232[333],s232[334],s232[335],s232[336],s232[337],s232[338],s232[339],s231[341],s230[343],s229[345],s228[347],s227[349],s226[351],s225[353],s224[307],s223[309],s222[311],s221[313],s220[315],s219[317],s218[319],s217[321],s216[323],s215[325],s214[327],s213[329],s212[331],s211[333],s210[335],s210[336],s210[337],s210[338],s210[339],s210[340],s210[341],s210[342],s210[343],s210[344],s210[345],s210[346],s210[347],s210[348],s210[349],s210[350],s210[351],s210[352],s210[353],s210[354],s210[355],s210[356],s210[357],s210[358],s210[359],s210[360],s210[361],s210[362],s210[363],s210[364],s210[365],s210[366],s210[367],s210[368],s210[369],s210[370],s210[371],s210[372],s210[373],s210[374],s210[375],s210[376],s210[377],s210[378],s210[379],s210[380],s210[381],s210[382],s210[383],s210[384],s210[385],s210[386],s210[387],s210[388],s210[389],s210[390],s210[391],s210[392],s210[393],s210[394],s210[395],s210[396],s210[397],s210[398],s210[399],s209[401],s208[403],s207[405],s206[407],s205[409],s204[411],s203[413],s202[415],s201[417],s200[419],s199[421],s198[423],s197[425],s196[427],s195[429],s194[431],s193[433],pp255[211],pp254[213],pp253[215],pp252[217],pp251[219],pp250[221],pp249[223],pp248[225],pp247[227],pp246[229],pp245[231],pp244[233],pp243[235],pp242[237],pp241[239],pp242[239],pp243[239],pp244[239],pp245[239],pp246[239],pp247[239],pp248[239]};
    assign in233_2 = {pp17[7],pp17[8],pp9[17],pp7[20],pp5[23],pp3[26],pp1[29],s230[10],s231[10],s232[10],pp0[34],pp1[34],pp2[34],pp3[34],pp4[34],pp5[34],pp6[34],pp7[34],pp7[35],pp7[36],pp7[37],pp7[38],pp7[39],pp7[40],pp7[41],pp7[42],pp7[43],pp7[44],pp7[45],pp7[46],pp7[47],pp7[48],pp7[49],pp7[50],pp7[51],pp7[52],pp7[53],pp7[54],pp7[55],pp7[56],pp7[57],pp7[58],pp7[59],pp7[60],pp7[61],pp7[62],pp7[63],pp7[64],pp7[65],pp7[66],pp7[67],pp7[68],pp7[69],pp7[70],pp7[71],pp7[72],pp7[73],pp7[74],pp7[75],pp7[76],pp7[77],pp7[78],pp7[79],pp7[80],pp7[81],pp7[82],pp7[83],pp7[84],pp7[85],pp7[86],pp7[87],pp7[88],pp7[89],pp7[90],pp7[91],pp7[92],pp6[94],pp5[96],pp4[98],s232[80],s230[83],s228[86],s226[89],s224[44],s222[47],s220[50],s220[51],s220[52],s220[53],s220[54],s220[55],s220[56],s219[58],s218[60],s217[62],s216[64],s215[66],s214[68],s213[70],s212[72],s212[73],s212[74],s212[75],s212[76],s212[77],s212[78],s212[79],s212[80],s212[81],s212[82],s212[83],s212[84],s212[85],s212[86],s213[86],s214[86],s215[86],s216[86],s217[86],s218[86],s219[86],s220[86],s221[86],s222[86],s223[86],s224[86],s10[13],s11[13],s12[13],s13[13],s14[13],s15[13],s16[13],s17[13],s18[13],s19[13],s20[13],s21[13],s22[13],s23[13],s24[13],s25[13],s26[13],s27[13],s28[13],s29[13],s30[13],s31[13],s32[13],s33[13],s34[13],s35[13],s36[13],s37[13],s38[13],s39[13],s40[13],s41[13],s42[13],s43[13],s44[13],s45[13],s46[13],s47[13],s48[13],s49[13],s50[13],s51[13],s52[13],s53[13],s54[13],s55[13],s56[13],s57[13],s58[13],s59[13],s60[13],s61[13],s62[13],s63[13],s64[13],s65[13],s66[13],s67[13],s68[13],s69[13],s70[13],s71[13],s72[13],s73[13],s74[13],s75[13],s76[13],s77[13],s78[13],s79[13],s80[13],s81[13],s82[13],s83[13],s84[13],s85[13],s86[13],s87[13],s87[14],s87[15],s87[16],s87[17],s87[18],s87[19],s87[20],s87[21],s87[22],s87[23],s87[24],s87[25],s87[26],s87[27],s87[28],s87[29],s87[30],s87[31],s87[32],s87[33],s87[34],s87[35],s87[36],s87[37],s87[38],s87[39],s87[40],s87[41],s87[42],s85[45],s83[48],s81[51],s79[54],s78[56],s78[57],s78[58],s78[59],s78[60],s78[61],s78[62],s78[63],s78[64],s78[65],s78[66],s78[67],s78[68],s78[69],s78[70],s78[71],s78[72],s78[73],s78[74],s78[75],s78[76],s78[77],s78[78],s78[79],s78[80],s77[82],s76[84],s75[86],s74[88],s73[90],s72[92],s71[94],s70[96],s69[98],s9[159],s7[162],s5[165],s3[168],s1[171],s72[101],s71[103],s70[105],s69[107],s68[109],s67[111],s66[113],s65[115],s64[117],s63[119],s62[121],s61[123],s60[125],s59[127],s58[129],s57[131],s56[133],s55[135],s54[137],s53[139],s52[141],s51[143],s50[145],s49[147],s48[149],s47[151],s46[153],s45[155],s44[157],s43[159],s42[161],s41[163],s40[165],s39[167],s38[169],s37[171],s36[173],s35[175],s34[177],s33[179],s32[181],s31[183],s30[185],s29[187],s28[189],s27[191],s26[193],s25[195],s24[197],s23[199],s22[201],s21[203],s20[205],s19[207],s18[209],s17[211],s16[213],s15[215],s14[217],s13[219],s12[221],s11[223],s10[225],s232[340],s231[342],s230[344],s229[346],s228[348],s227[350],s226[352],s225[354],s224[308],s223[310],s222[312],s221[314],s220[316],s219[318],s218[320],s217[322],s216[324],s215[326],s214[328],s213[330],s212[332],s211[334],s211[335],s211[336],s211[337],s211[338],s211[339],s211[340],s211[341],s211[342],s211[343],s211[344],s211[345],s211[346],s211[347],s211[348],s211[349],s211[350],s211[351],s211[352],s211[353],s211[354],s211[355],s211[356],s211[357],s211[358],s211[359],s211[360],s211[361],s211[362],s211[363],s211[364],s211[365],s211[366],s211[367],s211[368],s211[369],s211[370],s211[371],s211[372],s211[373],s211[374],s211[375],s211[376],s211[377],s211[378],s211[379],s211[380],s211[381],s211[382],s211[383],s211[384],s211[385],s211[386],s211[387],s211[388],s211[389],s211[390],s211[391],s211[392],s211[393],s211[394],s211[395],s211[396],s211[397],s211[398],s210[400],s209[402],s208[404],s207[406],s206[408],s205[410],s204[412],s203[414],s202[416],s201[418],s200[420],s199[422],s198[424],s197[426],s196[428],s195[430],s194[432],s193[434],pp255[212],pp254[214],pp253[216],pp252[218],pp251[220],pp250[222],pp249[224],pp248[226],pp247[228],pp246[230],pp245[232],pp244[234],pp243[236],pp242[238],pp243[238],pp244[238],pp245[238],pp246[238],pp247[238],pp248[238],pp249[238]};
    CLA_464 KS_233(s233, c233, in233_1, in233_2);
    wire[461:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {pp18[7],pp17[9],pp8[19],pp6[22],pp4[25],pp2[28],pp0[31],pp0[32],pp0[33],s233[10],s233[11],s233[12],s233[13],s233[14],s233[15],s233[16],s233[17],s233[18],s233[19],s233[20],s233[21],s233[22],s233[23],s233[24],s233[25],s233[26],s233[27],s233[28],s233[29],s233[30],s233[31],s233[32],s233[33],s233[34],s233[35],s233[36],s233[37],s233[38],s233[39],s233[40],s233[41],s233[42],s233[43],s233[44],s233[45],s233[46],s233[47],s233[48],s233[49],s233[50],s233[51],s233[52],s233[53],s233[54],s233[55],s233[56],s233[57],s233[58],s233[59],s233[60],s233[61],s233[62],s233[63],s233[64],s233[65],s233[66],s233[67],s233[68],s233[69],s233[70],s233[71],s233[72],s233[73],s233[74],s233[75],s233[76],s233[77],s233[78],s233[79],s231[82],s229[85],s227[88],s225[91],s223[46],s221[49],s221[50],s221[51],s221[52],s221[53],s221[54],s221[55],s220[57],s219[59],s218[61],s217[63],s216[65],s215[67],s214[69],s213[71],s233[100],s233[101],s233[102],s233[103],s233[104],s233[105],s233[106],s233[107],s233[108],s233[109],s233[110],s233[111],s233[112],s233[113],s233[114],s233[115],s233[116],s233[117],s233[118],s233[119],s233[120],s233[121],s233[122],s233[123],s233[124],s233[125],s233[126],s233[127],s233[128],s233[129],s233[130],s233[131],s233[132],s233[133],s233[134],s233[135],s233[136],s233[137],s233[138],s233[139],s233[140],s233[141],s233[142],s233[143],s233[144],s233[145],s233[146],s233[147],s233[148],s233[149],s233[150],s233[151],s233[152],s233[153],s233[154],s233[155],s233[156],s233[157],s233[158],s233[159],s233[160],s233[161],s233[162],s233[163],s233[164],s233[165],s233[166],s233[167],s233[168],s233[169],s233[170],s233[171],s233[172],s233[173],s233[174],s233[175],s233[176],s233[177],s233[178],s233[179],s233[180],s233[181],s233[182],s233[183],s233[184],s233[185],s233[186],s233[187],s233[188],s233[189],s233[190],s233[191],s233[192],s233[193],s233[194],s233[195],s233[196],s233[197],s233[198],s233[199],s233[200],s233[201],s233[202],s233[203],s233[204],s233[205],s233[206],s233[207],s233[208],s233[209],s233[210],s233[211],s233[212],s233[213],s233[214],s233[215],s233[216],s233[217],s233[218],s233[219],s233[220],s233[221],s233[222],s233[223],s233[224],s233[225],s233[226],s233[227],s233[228],s233[229],s233[230],s233[231],s233[232],s233[233],s233[234],s233[235],s233[236],s233[237],s233[238],s233[239],s233[240],s233[241],s233[242],s233[243],s233[244],s233[245],s233[246],s233[247],s233[248],s233[249],s233[250],s233[251],s233[252],s233[253],s233[254],s233[255],s233[256],s233[257],s233[258],s233[259],s233[260],s233[261],s233[262],s233[263],s233[264],s233[265],s233[266],s233[267],s233[268],s233[269],s233[270],s233[271],s233[272],s233[273],s233[274],s233[275],s233[276],s233[277],s233[278],s233[279],s233[280],s233[281],s233[282],s233[283],s233[284],s233[285],s233[286],s233[287],s233[288],s233[289],s233[290],s233[291],s233[292],s233[293],s233[294],s233[295],s233[296],s233[297],s233[298],s233[299],s233[300],s233[301],s233[302],s233[303],s233[304],s233[305],s233[306],s233[307],s233[308],s233[309],s233[310],s233[311],s233[312],s233[313],s233[314],s233[315],s233[316],s233[317],s233[318],s233[319],s233[320],s233[321],s233[322],s233[323],s233[324],s233[325],s233[326],s233[327],s233[328],s233[329],s233[330],s233[331],s233[332],s233[333],s233[334],s233[335],s233[336],s233[337],s233[338],s233[339],s232[341],s231[343],s230[345],s229[347],s228[349],s227[351],s226[353],s225[355],s224[309],s223[311],s222[313],s221[315],s220[317],s219[319],s218[321],s217[323],s216[325],s215[327],s214[329],s213[331],s212[333],s212[334],s212[335],s212[336],s212[337],s212[338],s212[339],s212[340],s212[341],s212[342],s212[343],s212[344],s212[345],s212[346],s212[347],s212[348],s212[349],s212[350],s212[351],s212[352],s212[353],s212[354],s212[355],s212[356],s212[357],s212[358],s212[359],s212[360],s212[361],s212[362],s212[363],s212[364],s212[365],s212[366],s212[367],s212[368],s212[369],s212[370],s212[371],s212[372],s212[373],s212[374],s212[375],s212[376],s212[377],s212[378],s212[379],s212[380],s212[381],s212[382],s212[383],s212[384],s212[385],s212[386],s212[387],s212[388],s212[389],s212[390],s212[391],s212[392],s212[393],s212[394],s212[395],s212[396],s212[397],s211[399],s210[401],s209[403],s208[405],s207[407],s206[409],s205[411],s204[413],s203[415],s202[417],s201[419],s200[421],s199[423],s198[425],s197[427],s196[429],s195[431],s194[433],s193[435],pp255[213],pp254[215],pp253[217],pp252[219],pp251[221],pp250[223],pp249[225],pp248[227],pp247[229],pp246[231],pp245[233],pp244[235],pp243[237],pp244[237],pp245[237],pp246[237],pp247[237],pp248[237],pp249[237]};
    assign in234_2 = {pp19[6],pp18[8],pp9[18],pp7[21],pp5[24],pp3[27],pp1[30],pp1[31],pp1[32],pp1[33],pp2[33],pp3[33],pp4[33],pp5[33],pp6[33],pp7[33],pp8[33],pp8[34],pp8[35],pp8[36],pp8[37],pp8[38],pp8[39],pp8[40],pp8[41],pp8[42],pp8[43],pp8[44],pp8[45],pp8[46],pp8[47],pp8[48],pp8[49],pp8[50],pp8[51],pp8[52],pp8[53],pp8[54],pp8[55],pp8[56],pp8[57],pp8[58],pp8[59],pp8[60],pp8[61],pp8[62],pp8[63],pp8[64],pp8[65],pp8[66],pp8[67],pp8[68],pp8[69],pp8[70],pp8[71],pp8[72],pp8[73],pp8[74],pp8[75],pp8[76],pp8[77],pp8[78],pp8[79],pp8[80],pp8[81],pp8[82],pp8[83],pp8[84],pp8[85],pp8[86],pp8[87],pp8[88],pp8[89],pp8[90],pp8[91],pp7[93],pp6[95],pp5[97],pp4[99],s232[81],s230[84],s228[87],s226[90],s224[45],s222[48],s222[49],s222[50],s222[51],s222[52],s222[53],s222[54],s221[56],s220[58],s219[60],s218[62],s217[64],s216[66],s215[68],s214[70],s213[72],s213[73],s213[74],s213[75],s213[76],s213[77],s213[78],s213[79],s213[80],s213[81],s213[82],s213[83],s213[84],s213[85],s214[85],s215[85],s216[85],s217[85],s218[85],s219[85],s220[85],s221[85],s222[85],s223[85],s224[85],s10[12],s11[12],s12[12],s13[12],s14[12],s15[12],s16[12],s17[12],s18[12],s19[12],s20[12],s21[12],s22[12],s23[12],s24[12],s25[12],s26[12],s27[12],s28[12],s29[12],s30[12],s31[12],s32[12],s33[12],s34[12],s35[12],s36[12],s37[12],s38[12],s39[12],s40[12],s41[12],s42[12],s43[12],s44[12],s45[12],s46[12],s47[12],s48[12],s49[12],s50[12],s51[12],s52[12],s53[12],s54[12],s55[12],s56[12],s57[12],s58[12],s59[12],s60[12],s61[12],s62[12],s63[12],s64[12],s65[12],s66[12],s67[12],s68[12],s69[12],s70[12],s71[12],s72[12],s73[12],s74[12],s75[12],s76[12],s77[12],s78[12],s79[12],s80[12],s81[12],s82[12],s83[12],s84[12],s85[12],s86[12],s87[12],s88[12],s88[13],s88[14],s88[15],s88[16],s88[17],s88[18],s88[19],s88[20],s88[21],s88[22],s88[23],s88[24],s88[25],s88[26],s88[27],s88[28],s88[29],s88[30],s88[31],s88[32],s88[33],s88[34],s88[35],s88[36],s88[37],s88[38],s88[39],s88[40],s88[41],s86[44],s84[47],s82[50],s80[53],s79[55],s79[56],s79[57],s79[58],s79[59],s79[60],s79[61],s79[62],s79[63],s79[64],s79[65],s79[66],s79[67],s79[68],s79[69],s79[70],s79[71],s79[72],s79[73],s79[74],s79[75],s79[76],s79[77],s79[78],s79[79],s78[81],s77[83],s76[85],s75[87],s74[89],s73[91],s72[93],s71[95],s70[97],s69[99],s8[161],s6[164],s4[167],s2[170],s73[100],s72[102],s71[104],s70[106],s69[108],s68[110],s67[112],s66[114],s65[116],s64[118],s63[120],s62[122],s61[124],s60[126],s59[128],s58[130],s57[132],s56[134],s55[136],s54[138],s53[140],s52[142],s51[144],s50[146],s49[148],s48[150],s47[152],s46[154],s45[156],s44[158],s43[160],s42[162],s41[164],s40[166],s39[168],s38[170],s37[172],s36[174],s35[176],s34[178],s33[180],s32[182],s31[184],s30[186],s29[188],s28[190],s27[192],s26[194],s25[196],s24[198],s23[200],s22[202],s21[204],s20[206],s19[208],s18[210],s17[212],s16[214],s15[216],s14[218],s13[220],s12[222],s11[224],s10[226],s233[340],s232[342],s231[344],s230[346],s229[348],s228[350],s227[352],s226[354],s225[356],s224[310],s223[312],s222[314],s221[316],s220[318],s219[320],s218[322],s217[324],s216[326],s215[328],s214[330],s213[332],s213[333],s213[334],s213[335],s213[336],s213[337],s213[338],s213[339],s213[340],s213[341],s213[342],s213[343],s213[344],s213[345],s213[346],s213[347],s213[348],s213[349],s213[350],s213[351],s213[352],s213[353],s213[354],s213[355],s213[356],s213[357],s213[358],s213[359],s213[360],s213[361],s213[362],s213[363],s213[364],s213[365],s213[366],s213[367],s213[368],s213[369],s213[370],s213[371],s213[372],s213[373],s213[374],s213[375],s213[376],s213[377],s213[378],s213[379],s213[380],s213[381],s213[382],s213[383],s213[384],s213[385],s213[386],s213[387],s213[388],s213[389],s213[390],s213[391],s213[392],s213[393],s213[394],s213[395],s213[396],s212[398],s211[400],s210[402],s209[404],s208[406],s207[408],s206[410],s205[412],s204[414],s203[416],s202[418],s201[420],s200[422],s199[424],s198[426],s197[428],s196[430],s195[432],s194[434],s193[436],pp255[214],pp254[216],pp253[218],pp252[220],pp251[222],pp250[224],pp249[226],pp248[228],pp247[230],pp246[232],pp245[234],pp244[236],pp245[236],pp246[236],pp247[236],pp248[236],pp249[236],pp250[236]};
    CLA_462 KS_234(s234, c234, in234_1, in234_2);
    wire[459:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {pp19[7],pp18[9],pp8[20],pp6[23],pp4[26],pp2[29],pp2[30],pp2[31],pp2[32],s234[10],s234[11],s234[12],s234[13],s234[14],s234[15],s234[16],s234[17],s234[18],s234[19],s234[20],s234[21],s234[22],s234[23],s234[24],s234[25],s234[26],s234[27],s234[28],s234[29],s234[30],s234[31],s234[32],s234[33],s234[34],s234[35],s234[36],s234[37],s234[38],s234[39],s234[40],s234[41],s234[42],s234[43],s234[44],s234[45],s234[46],s234[47],s234[48],s234[49],s234[50],s234[51],s234[52],s234[53],s234[54],s234[55],s234[56],s234[57],s234[58],s234[59],s234[60],s234[61],s234[62],s234[63],s234[64],s234[65],s234[66],s234[67],s234[68],s234[69],s234[70],s234[71],s234[72],s234[73],s234[74],s234[75],s234[76],s234[77],s234[78],s233[80],s231[83],s229[86],s227[89],s225[92],s223[47],s223[48],s223[49],s223[50],s223[51],s223[52],s223[53],s222[55],s221[57],s220[59],s219[61],s218[63],s217[65],s216[67],s215[69],s214[71],s234[100],s234[101],s234[102],s234[103],s234[104],s234[105],s234[106],s234[107],s234[108],s234[109],s234[110],s234[111],s234[112],s234[113],s234[114],s234[115],s234[116],s234[117],s234[118],s234[119],s234[120],s234[121],s234[122],s234[123],s234[124],s234[125],s234[126],s234[127],s234[128],s234[129],s234[130],s234[131],s234[132],s234[133],s234[134],s234[135],s234[136],s234[137],s234[138],s234[139],s234[140],s234[141],s234[142],s234[143],s234[144],s234[145],s234[146],s234[147],s234[148],s234[149],s234[150],s234[151],s234[152],s234[153],s234[154],s234[155],s234[156],s234[157],s234[158],s234[159],s234[160],s234[161],s234[162],s234[163],s234[164],s234[165],s234[166],s234[167],s234[168],s234[169],s234[170],s234[171],s234[172],s234[173],s234[174],s234[175],s234[176],s234[177],s234[178],s234[179],s234[180],s234[181],s234[182],s234[183],s234[184],s234[185],s234[186],s234[187],s234[188],s234[189],s234[190],s234[191],s234[192],s234[193],s234[194],s234[195],s234[196],s234[197],s234[198],s234[199],s234[200],s234[201],s234[202],s234[203],s234[204],s234[205],s234[206],s234[207],s234[208],s234[209],s234[210],s234[211],s234[212],s234[213],s234[214],s234[215],s234[216],s234[217],s234[218],s234[219],s234[220],s234[221],s234[222],s234[223],s234[224],s234[225],s234[226],s234[227],s234[228],s234[229],s234[230],s234[231],s234[232],s234[233],s234[234],s234[235],s234[236],s234[237],s234[238],s234[239],s234[240],s234[241],s234[242],s234[243],s234[244],s234[245],s234[246],s234[247],s234[248],s234[249],s234[250],s234[251],s234[252],s234[253],s234[254],s234[255],s234[256],s234[257],s234[258],s234[259],s234[260],s234[261],s234[262],s234[263],s234[264],s234[265],s234[266],s234[267],s234[268],s234[269],s234[270],s234[271],s234[272],s234[273],s234[274],s234[275],s234[276],s234[277],s234[278],s234[279],s234[280],s234[281],s234[282],s234[283],s234[284],s234[285],s234[286],s234[287],s234[288],s234[289],s234[290],s234[291],s234[292],s234[293],s234[294],s234[295],s234[296],s234[297],s234[298],s234[299],s234[300],s234[301],s234[302],s234[303],s234[304],s234[305],s234[306],s234[307],s234[308],s234[309],s234[310],s234[311],s234[312],s234[313],s234[314],s234[315],s234[316],s234[317],s234[318],s234[319],s234[320],s234[321],s234[322],s234[323],s234[324],s234[325],s234[326],s234[327],s234[328],s234[329],s234[330],s234[331],s234[332],s234[333],s234[334],s234[335],s234[336],s234[337],s234[338],s234[339],s233[341],s232[343],s231[345],s230[347],s229[349],s228[351],s227[353],s226[355],s225[357],s224[311],s223[313],s222[315],s221[317],s220[319],s219[321],s218[323],s217[325],s216[327],s215[329],s214[331],s214[332],s214[333],s214[334],s214[335],s214[336],s214[337],s214[338],s214[339],s214[340],s214[341],s214[342],s214[343],s214[344],s214[345],s214[346],s214[347],s214[348],s214[349],s214[350],s214[351],s214[352],s214[353],s214[354],s214[355],s214[356],s214[357],s214[358],s214[359],s214[360],s214[361],s214[362],s214[363],s214[364],s214[365],s214[366],s214[367],s214[368],s214[369],s214[370],s214[371],s214[372],s214[373],s214[374],s214[375],s214[376],s214[377],s214[378],s214[379],s214[380],s214[381],s214[382],s214[383],s214[384],s214[385],s214[386],s214[387],s214[388],s214[389],s214[390],s214[391],s214[392],s214[393],s214[394],s214[395],s213[397],s212[399],s211[401],s210[403],s209[405],s208[407],s207[409],s206[411],s205[413],s204[415],s203[417],s202[419],s201[421],s200[423],s199[425],s198[427],s197[429],s196[431],s195[433],s194[435],s193[437],pp255[215],pp254[217],pp253[219],pp252[221],pp251[223],pp250[225],pp249[227],pp248[229],pp247[231],pp246[233],pp245[235],pp246[235],pp247[235],pp248[235],pp249[235],pp250[235]};
    assign in235_2 = {pp20[6],pp19[8],pp9[19],pp7[22],pp5[25],pp3[28],pp3[29],pp3[30],pp3[31],pp3[32],pp4[32],pp5[32],pp6[32],pp7[32],pp8[32],pp9[32],pp9[33],pp9[34],pp9[35],pp9[36],pp9[37],pp9[38],pp9[39],pp9[40],pp9[41],pp9[42],pp9[43],pp9[44],pp9[45],pp9[46],pp9[47],pp9[48],pp9[49],pp9[50],pp9[51],pp9[52],pp9[53],pp9[54],pp9[55],pp9[56],pp9[57],pp9[58],pp9[59],pp9[60],pp9[61],pp9[62],pp9[63],pp9[64],pp9[65],pp9[66],pp9[67],pp9[68],pp9[69],pp9[70],pp9[71],pp9[72],pp9[73],pp9[74],pp9[75],pp9[76],pp9[77],pp9[78],pp9[79],pp9[80],pp9[81],pp9[82],pp9[83],pp9[84],pp9[85],pp9[86],pp9[87],pp9[88],pp9[89],pp9[90],pp8[92],pp7[94],pp6[96],pp5[98],s234[79],s232[82],s230[85],s228[88],s226[91],s224[46],s224[47],s224[48],s224[49],s224[50],s224[51],s224[52],s223[54],s222[56],s221[58],s220[60],s219[62],s218[64],s217[66],s216[68],s215[70],s214[72],s214[73],s214[74],s214[75],s214[76],s214[77],s214[78],s214[79],s214[80],s214[81],s214[82],s214[83],s214[84],s215[84],s216[84],s217[84],s218[84],s219[84],s220[84],s221[84],s222[84],s223[84],s224[84],s10[11],s11[11],s12[11],s13[11],s14[11],s15[11],s16[11],s17[11],s18[11],s19[11],s20[11],s21[11],s22[11],s23[11],s24[11],s25[11],s26[11],s27[11],s28[11],s29[11],s30[11],s31[11],s32[11],s33[11],s34[11],s35[11],s36[11],s37[11],s38[11],s39[11],s40[11],s41[11],s42[11],s43[11],s44[11],s45[11],s46[11],s47[11],s48[11],s49[11],s50[11],s51[11],s52[11],s53[11],s54[11],s55[11],s56[11],s57[11],s58[11],s59[11],s60[11],s61[11],s62[11],s63[11],s64[11],s65[11],s66[11],s67[11],s68[11],s69[11],s70[11],s71[11],s72[11],s73[11],s74[11],s75[11],s76[11],s77[11],s78[11],s79[11],s80[11],s81[11],s82[11],s83[11],s84[11],s85[11],s86[11],s87[11],s88[11],s89[11],s89[12],s89[13],s89[14],s89[15],s89[16],s89[17],s89[18],s89[19],s89[20],s89[21],s89[22],s89[23],s89[24],s89[25],s89[26],s89[27],s89[28],s89[29],s89[30],s89[31],s89[32],s89[33],s89[34],s89[35],s89[36],s89[37],s89[38],s89[39],s89[40],s87[43],s85[46],s83[49],s81[52],s80[54],s80[55],s80[56],s80[57],s80[58],s80[59],s80[60],s80[61],s80[62],s80[63],s80[64],s80[65],s80[66],s80[67],s80[68],s80[69],s80[70],s80[71],s80[72],s80[73],s80[74],s80[75],s80[76],s80[77],s80[78],s79[80],s78[82],s77[84],s76[86],s75[88],s74[90],s73[92],s72[94],s71[96],s70[98],s9[160],s7[163],s5[166],s3[169],s1[172],s73[101],s72[103],s71[105],s70[107],s69[109],s68[111],s67[113],s66[115],s65[117],s64[119],s63[121],s62[123],s61[125],s60[127],s59[129],s58[131],s57[133],s56[135],s55[137],s54[139],s53[141],s52[143],s51[145],s50[147],s49[149],s48[151],s47[153],s46[155],s45[157],s44[159],s43[161],s42[163],s41[165],s40[167],s39[169],s38[171],s37[173],s36[175],s35[177],s34[179],s33[181],s32[183],s31[185],s30[187],s29[189],s28[191],s27[193],s26[195],s25[197],s24[199],s23[201],s22[203],s21[205],s20[207],s19[209],s18[211],s17[213],s16[215],s15[217],s14[219],s13[221],s12[223],s11[225],s10[227],s234[340],s233[342],s232[344],s231[346],s230[348],s229[350],s228[352],s227[354],s226[356],s225[358],s224[312],s223[314],s222[316],s221[318],s220[320],s219[322],s218[324],s217[326],s216[328],s215[330],s215[331],s215[332],s215[333],s215[334],s215[335],s215[336],s215[337],s215[338],s215[339],s215[340],s215[341],s215[342],s215[343],s215[344],s215[345],s215[346],s215[347],s215[348],s215[349],s215[350],s215[351],s215[352],s215[353],s215[354],s215[355],s215[356],s215[357],s215[358],s215[359],s215[360],s215[361],s215[362],s215[363],s215[364],s215[365],s215[366],s215[367],s215[368],s215[369],s215[370],s215[371],s215[372],s215[373],s215[374],s215[375],s215[376],s215[377],s215[378],s215[379],s215[380],s215[381],s215[382],s215[383],s215[384],s215[385],s215[386],s215[387],s215[388],s215[389],s215[390],s215[391],s215[392],s215[393],s215[394],s214[396],s213[398],s212[400],s211[402],s210[404],s209[406],s208[408],s207[410],s206[412],s205[414],s204[416],s203[418],s202[420],s201[422],s200[424],s199[426],s198[428],s197[430],s196[432],s195[434],s194[436],s193[438],pp255[216],pp254[218],pp253[220],pp252[222],pp251[224],pp250[226],pp249[228],pp248[230],pp247[232],pp246[234],pp247[234],pp248[234],pp249[234],pp250[234],pp251[234]};
    CLA_460 KS_235(s235, c235, in235_1, in235_2);
    wire[457:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {pp20[7],pp19[9],pp8[21],pp6[24],pp4[27],pp4[28],pp4[29],pp4[30],pp4[31],s235[10],s235[11],s235[12],s235[13],s235[14],s235[15],s235[16],s235[17],s235[18],s235[19],s235[20],s235[21],s235[22],s235[23],s235[24],s235[25],s235[26],s235[27],s235[28],s235[29],s235[30],s235[31],s235[32],s235[33],s235[34],s235[35],s235[36],s235[37],s235[38],s235[39],s235[40],s235[41],s235[42],s235[43],s235[44],s235[45],s235[46],s235[47],s235[48],s235[49],s235[50],s235[51],s235[52],s235[53],s235[54],s235[55],s235[56],s235[57],s235[58],s235[59],s235[60],s235[61],s235[62],s235[63],s235[64],s235[65],s235[66],s235[67],s235[68],s235[69],s235[70],s235[71],s235[72],s235[73],s235[74],s235[75],s235[76],s235[77],s235[78],s233[81],s231[84],s229[87],s227[90],s225[93],s225[94],s225[95],s225[96],s225[97],s225[98],s225[99],s224[53],s223[55],s222[57],s221[59],s220[61],s219[63],s218[65],s217[67],s216[69],s215[71],s235[100],s235[101],s235[102],s235[103],s235[104],s235[105],s235[106],s235[107],s235[108],s235[109],s235[110],s235[111],s235[112],s235[113],s235[114],s235[115],s235[116],s235[117],s235[118],s235[119],s235[120],s235[121],s235[122],s235[123],s235[124],s235[125],s235[126],s235[127],s235[128],s235[129],s235[130],s235[131],s235[132],s235[133],s235[134],s235[135],s235[136],s235[137],s235[138],s235[139],s235[140],s235[141],s235[142],s235[143],s235[144],s235[145],s235[146],s235[147],s235[148],s235[149],s235[150],s235[151],s235[152],s235[153],s235[154],s235[155],s235[156],s235[157],s235[158],s235[159],s235[160],s235[161],s235[162],s235[163],s235[164],s235[165],s235[166],s235[167],s235[168],s235[169],s235[170],s235[171],s235[172],s235[173],s235[174],s235[175],s235[176],s235[177],s235[178],s235[179],s235[180],s235[181],s235[182],s235[183],s235[184],s235[185],s235[186],s235[187],s235[188],s235[189],s235[190],s235[191],s235[192],s235[193],s235[194],s235[195],s235[196],s235[197],s235[198],s235[199],s235[200],s235[201],s235[202],s235[203],s235[204],s235[205],s235[206],s235[207],s235[208],s235[209],s235[210],s235[211],s235[212],s235[213],s235[214],s235[215],s235[216],s235[217],s235[218],s235[219],s235[220],s235[221],s235[222],s235[223],s235[224],s235[225],s235[226],s235[227],s235[228],s235[229],s235[230],s235[231],s235[232],s235[233],s235[234],s235[235],s235[236],s235[237],s235[238],s235[239],s235[240],s235[241],s235[242],s235[243],s235[244],s235[245],s235[246],s235[247],s235[248],s235[249],s235[250],s235[251],s235[252],s235[253],s235[254],s235[255],s235[256],s235[257],s235[258],s235[259],s235[260],s235[261],s235[262],s235[263],s235[264],s235[265],s235[266],s235[267],s235[268],s235[269],s235[270],s235[271],s235[272],s235[273],s235[274],s235[275],s235[276],s235[277],s235[278],s235[279],s235[280],s235[281],s235[282],s235[283],s235[284],s235[285],s235[286],s235[287],s235[288],s235[289],s235[290],s235[291],s235[292],s235[293],s235[294],s235[295],s235[296],s235[297],s235[298],s235[299],s235[300],s235[301],s235[302],s235[303],s235[304],s235[305],s235[306],s235[307],s235[308],s235[309],s235[310],s235[311],s235[312],s235[313],s235[314],s235[315],s235[316],s235[317],s235[318],s235[319],s235[320],s235[321],s235[322],s235[323],s235[324],s235[325],s235[326],s235[327],s235[328],s235[329],s235[330],s235[331],s235[332],s235[333],s235[334],s235[335],s235[336],s235[337],s235[338],s235[339],s234[341],s233[343],s232[345],s231[347],s230[349],s229[351],s228[353],s227[355],s226[357],s225[359],s224[313],s223[315],s222[317],s221[319],s220[321],s219[323],s218[325],s217[327],s216[329],s216[330],s216[331],s216[332],s216[333],s216[334],s216[335],s216[336],s216[337],s216[338],s216[339],s216[340],s216[341],s216[342],s216[343],s216[344],s216[345],s216[346],s216[347],s216[348],s216[349],s216[350],s216[351],s216[352],s216[353],s216[354],s216[355],s216[356],s216[357],s216[358],s216[359],s216[360],s216[361],s216[362],s216[363],s216[364],s216[365],s216[366],s216[367],s216[368],s216[369],s216[370],s216[371],s216[372],s216[373],s216[374],s216[375],s216[376],s216[377],s216[378],s216[379],s216[380],s216[381],s216[382],s216[383],s216[384],s216[385],s216[386],s216[387],s216[388],s216[389],s216[390],s216[391],s216[392],s216[393],s215[395],s214[397],s213[399],s212[401],s211[403],s210[405],s209[407],s208[409],s207[411],s206[413],s205[415],s204[417],s203[419],s202[421],s201[423],s200[425],s199[427],s198[429],s197[431],s196[433],s195[435],s194[437],s193[439],pp255[217],pp254[219],pp253[221],pp252[223],pp251[225],pp250[227],pp249[229],pp248[231],pp247[233],pp248[233],pp249[233],pp250[233],pp251[233]};
    assign in236_2 = {pp21[6],pp20[8],pp9[20],pp7[23],pp5[26],pp5[27],pp5[28],pp5[29],pp5[30],pp5[31],pp6[31],pp7[31],pp8[31],pp9[31],pp32[9],pp33[9],pp34[9],pp35[9],pp36[9],pp37[9],pp38[9],pp39[9],pp40[9],pp41[9],pp42[9],pp43[9],pp44[9],pp45[9],pp46[9],pp47[9],pp48[9],pp49[9],pp50[9],pp51[9],pp52[9],pp53[9],pp54[9],pp55[9],pp56[9],pp57[9],pp58[9],pp59[9],pp60[9],pp61[9],pp62[9],pp63[9],pp64[9],pp65[9],pp66[9],pp67[9],pp68[9],pp69[9],pp70[9],pp71[9],pp72[9],pp73[9],pp74[9],pp75[9],pp76[9],pp77[9],pp78[9],pp79[9],pp80[9],pp81[9],pp82[9],pp83[9],pp84[9],pp85[9],pp86[9],pp87[9],pp88[9],pp89[9],pp90[9],pp9[91],pp8[93],pp7[95],pp6[97],pp5[99],s234[80],s232[83],s230[86],s228[89],s226[92],s226[93],s226[94],s226[95],s226[96],s226[97],s226[98],s226[99],s224[54],s223[56],s222[58],s221[60],s220[62],s219[64],s218[66],s217[68],s216[70],s215[72],s215[73],s215[74],s215[75],s215[76],s215[77],s215[78],s215[79],s215[80],s215[81],s215[82],s215[83],s216[83],s217[83],s218[83],s219[83],s220[83],s221[83],s222[83],s223[83],s224[83],s10[10],s11[10],s12[10],s13[10],s14[10],s15[10],s16[10],s17[10],s18[10],s19[10],s20[10],s21[10],s22[10],s23[10],s24[10],s25[10],s26[10],s27[10],s28[10],s29[10],s30[10],s31[10],s32[10],s33[10],s34[10],s35[10],s36[10],s37[10],s38[10],s39[10],s40[10],s41[10],s42[10],s43[10],s44[10],s45[10],s46[10],s47[10],s48[10],s49[10],s50[10],s51[10],s52[10],s53[10],s54[10],s55[10],s56[10],s57[10],s58[10],s59[10],s60[10],s61[10],s62[10],s63[10],s64[10],s65[10],s66[10],s67[10],s68[10],s69[10],s70[10],s71[10],s72[10],s73[10],s74[10],s75[10],s76[10],s77[10],s78[10],s79[10],s80[10],s81[10],s82[10],s83[10],s84[10],s85[10],s86[10],s87[10],s88[10],s89[10],s90[10],s90[11],s90[12],s90[13],s90[14],s90[15],s90[16],s90[17],s90[18],s90[19],s90[20],s90[21],s90[22],s90[23],s90[24],s90[25],s90[26],s90[27],s90[28],s90[29],s90[30],s90[31],s90[32],s90[33],s90[34],s90[35],s90[36],s90[37],s90[38],s90[39],s88[42],s86[45],s84[48],s82[51],s81[53],s81[54],s81[55],s81[56],s81[57],s81[58],s81[59],s81[60],s81[61],s81[62],s81[63],s81[64],s81[65],s81[66],s81[67],s81[68],s81[69],s81[70],s81[71],s81[72],s81[73],s81[74],s81[75],s81[76],s81[77],s80[79],s79[81],s78[83],s77[85],s76[87],s75[89],s74[91],s73[93],s72[95],s71[97],s70[99],s8[162],s6[165],s4[168],s2[171],s74[100],s73[102],s72[104],s71[106],s70[108],s69[110],s68[112],s67[114],s66[116],s65[118],s64[120],s63[122],s62[124],s61[126],s60[128],s59[130],s58[132],s57[134],s56[136],s55[138],s54[140],s53[142],s52[144],s51[146],s50[148],s49[150],s48[152],s47[154],s46[156],s45[158],s44[160],s43[162],s42[164],s41[166],s40[168],s39[170],s38[172],s37[174],s36[176],s35[178],s34[180],s33[182],s32[184],s31[186],s30[188],s29[190],s28[192],s27[194],s26[196],s25[198],s24[200],s23[202],s22[204],s21[206],s20[208],s19[210],s18[212],s17[214],s16[216],s15[218],s14[220],s13[222],s12[224],s11[226],s10[228],s235[340],s234[342],s233[344],s232[346],s231[348],s230[350],s229[352],s228[354],s227[356],s226[358],s225[360],s224[314],s223[316],s222[318],s221[320],s220[322],s219[324],s218[326],s217[328],s217[329],s217[330],s217[331],s217[332],s217[333],s217[334],s217[335],s217[336],s217[337],s217[338],s217[339],s217[340],s217[341],s217[342],s217[343],s217[344],s217[345],s217[346],s217[347],s217[348],s217[349],s217[350],s217[351],s217[352],s217[353],s217[354],s217[355],s217[356],s217[357],s217[358],s217[359],s217[360],s217[361],s217[362],s217[363],s217[364],s217[365],s217[366],s217[367],s217[368],s217[369],s217[370],s217[371],s217[372],s217[373],s217[374],s217[375],s217[376],s217[377],s217[378],s217[379],s217[380],s217[381],s217[382],s217[383],s217[384],s217[385],s217[386],s217[387],s217[388],s217[389],s217[390],s217[391],s217[392],s216[394],s215[396],s214[398],s213[400],s212[402],s211[404],s210[406],s209[408],s208[410],s207[412],s206[414],s205[416],s204[418],s203[420],s202[422],s201[424],s200[426],s199[428],s198[430],s197[432],s196[434],s195[436],s194[438],s193[440],pp255[218],pp254[220],pp253[222],pp252[224],pp251[226],pp250[228],pp249[230],pp248[232],pp249[232],pp250[232],pp251[232],pp252[232]};
    CLA_458 KS_236(s236, c236, in236_1, in236_2);
    wire[455:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {pp21[7],pp20[9],pp8[22],pp6[25],pp6[26],pp6[27],pp6[28],pp6[29],pp6[30],s236[10],s236[11],s236[12],s236[13],s236[14],s236[15],s236[16],s236[17],s236[18],s236[19],s236[20],s236[21],s236[22],s236[23],s236[24],s236[25],s236[26],s236[27],s236[28],s236[29],s236[30],s236[31],s236[32],s236[33],s236[34],s236[35],s236[36],s236[37],s236[38],s236[39],s236[40],s236[41],s236[42],s236[43],s236[44],s236[45],s236[46],s236[47],s236[48],s236[49],s236[50],s236[51],s236[52],s236[53],s236[54],s236[55],s236[56],s236[57],s236[58],s236[59],s236[60],s236[61],s236[62],s236[63],s236[64],s236[65],s236[66],s236[67],s236[68],s236[69],s236[70],s236[71],s236[72],s236[73],s236[74],s236[75],s236[76],s236[77],s235[79],s233[82],s231[85],s229[88],s227[91],s227[92],s227[93],s227[94],s227[95],s227[96],s227[97],s227[98],s227[99],s224[55],s223[57],s222[59],s221[61],s220[63],s219[65],s218[67],s217[69],s216[71],s236[100],s236[101],s236[102],s236[103],s236[104],s236[105],s236[106],s236[107],s236[108],s236[109],s236[110],s236[111],s236[112],s236[113],s236[114],s236[115],s236[116],s236[117],s236[118],s236[119],s236[120],s236[121],s236[122],s236[123],s236[124],s236[125],s236[126],s236[127],s236[128],s236[129],s236[130],s236[131],s236[132],s236[133],s236[134],s236[135],s236[136],s236[137],s236[138],s236[139],s236[140],s236[141],s236[142],s236[143],s236[144],s236[145],s236[146],s236[147],s236[148],s236[149],s236[150],s236[151],s236[152],s236[153],s236[154],s236[155],s236[156],s236[157],s236[158],s236[159],s236[160],s236[161],s236[162],s236[163],s236[164],s236[165],s236[166],s236[167],s236[168],s236[169],s236[170],s236[171],s236[172],s236[173],s236[174],s236[175],s236[176],s236[177],s236[178],s236[179],s236[180],s236[181],s236[182],s236[183],s236[184],s236[185],s236[186],s236[187],s236[188],s236[189],s236[190],s236[191],s236[192],s236[193],s236[194],s236[195],s236[196],s236[197],s236[198],s236[199],s236[200],s236[201],s236[202],s236[203],s236[204],s236[205],s236[206],s236[207],s236[208],s236[209],s236[210],s236[211],s236[212],s236[213],s236[214],s236[215],s236[216],s236[217],s236[218],s236[219],s236[220],s236[221],s236[222],s236[223],s236[224],s236[225],s236[226],s236[227],s236[228],s236[229],s236[230],s236[231],s236[232],s236[233],s236[234],s236[235],s236[236],s236[237],s236[238],s236[239],s236[240],s236[241],s236[242],s236[243],s236[244],s236[245],s236[246],s236[247],s236[248],s236[249],s236[250],s236[251],s236[252],s236[253],s236[254],s236[255],s236[256],s236[257],s236[258],s236[259],s236[260],s236[261],s236[262],s236[263],s236[264],s236[265],s236[266],s236[267],s236[268],s236[269],s236[270],s236[271],s236[272],s236[273],s236[274],s236[275],s236[276],s236[277],s236[278],s236[279],s236[280],s236[281],s236[282],s236[283],s236[284],s236[285],s236[286],s236[287],s236[288],s236[289],s236[290],s236[291],s236[292],s236[293],s236[294],s236[295],s236[296],s236[297],s236[298],s236[299],s236[300],s236[301],s236[302],s236[303],s236[304],s236[305],s236[306],s236[307],s236[308],s236[309],s236[310],s236[311],s236[312],s236[313],s236[314],s236[315],s236[316],s236[317],s236[318],s236[319],s236[320],s236[321],s236[322],s236[323],s236[324],s236[325],s236[326],s236[327],s236[328],s236[329],s236[330],s236[331],s236[332],s236[333],s236[334],s236[335],s236[336],s236[337],s236[338],s236[339],s235[341],s234[343],s233[345],s232[347],s231[349],s230[351],s229[353],s228[355],s227[357],s226[359],s225[361],s224[315],s223[317],s222[319],s221[321],s220[323],s219[325],s218[327],s218[328],s218[329],s218[330],s218[331],s218[332],s218[333],s218[334],s218[335],s218[336],s218[337],s218[338],s218[339],s218[340],s218[341],s218[342],s218[343],s218[344],s218[345],s218[346],s218[347],s218[348],s218[349],s218[350],s218[351],s218[352],s218[353],s218[354],s218[355],s218[356],s218[357],s218[358],s218[359],s218[360],s218[361],s218[362],s218[363],s218[364],s218[365],s218[366],s218[367],s218[368],s218[369],s218[370],s218[371],s218[372],s218[373],s218[374],s218[375],s218[376],s218[377],s218[378],s218[379],s218[380],s218[381],s218[382],s218[383],s218[384],s218[385],s218[386],s218[387],s218[388],s218[389],s218[390],s218[391],s217[393],s216[395],s215[397],s214[399],s213[401],s212[403],s211[405],s210[407],s209[409],s208[411],s207[413],s206[415],s205[417],s204[419],s203[421],s202[423],s201[425],s200[427],s199[429],s198[431],s197[433],s196[435],s195[437],s194[439],s193[441],pp255[219],pp254[221],pp253[223],pp252[225],pp251[227],pp250[229],pp249[231],pp250[231],pp251[231],pp252[231]};
    assign in237_2 = {pp22[6],pp21[8],pp9[21],pp7[24],pp7[25],pp7[26],pp7[27],pp7[28],pp7[29],pp7[30],pp8[30],pp9[30],pp31[9],pp33[8],pp34[8],pp35[8],pp36[8],pp37[8],pp38[8],pp39[8],pp40[8],pp41[8],pp42[8],pp43[8],pp44[8],pp45[8],pp46[8],pp47[8],pp48[8],pp49[8],pp50[8],pp51[8],pp52[8],pp53[8],pp54[8],pp55[8],pp56[8],pp57[8],pp58[8],pp59[8],pp60[8],pp61[8],pp62[8],pp63[8],pp64[8],pp65[8],pp66[8],pp67[8],pp68[8],pp69[8],pp70[8],pp71[8],pp72[8],pp73[8],pp74[8],pp75[8],pp76[8],pp77[8],pp78[8],pp79[8],pp80[8],pp81[8],pp82[8],pp83[8],pp84[8],pp85[8],pp86[8],pp87[8],pp88[8],pp89[8],pp90[8],pp91[8],pp91[9],pp9[92],pp8[94],pp7[96],pp6[98],s236[78],s234[81],s232[84],s230[87],s228[90],s228[91],s228[92],s228[93],s228[94],s228[95],s228[96],s228[97],s228[98],s228[99],s224[56],s223[58],s222[60],s221[62],s220[64],s219[66],s218[68],s217[70],s216[72],s216[73],s216[74],s216[75],s216[76],s216[77],s216[78],s216[79],s216[80],s216[81],s216[82],s217[82],s218[82],s219[82],s220[82],s221[82],s222[82],s223[82],s224[82],s1[18],s1[19],s1[20],s1[21],s1[22],s1[23],s1[24],s1[25],s1[26],s1[27],s1[28],s1[29],s1[30],s1[31],s1[32],s1[33],s1[34],s1[35],s1[36],s1[37],s1[38],s1[39],s1[40],s1[41],s1[42],s1[43],s1[44],s1[45],s1[46],s1[47],s1[48],s1[49],s1[50],s1[51],s1[52],s1[53],s1[54],s1[55],s1[56],s1[57],s1[58],s1[59],s1[60],s1[61],s1[62],s1[63],s1[64],s1[65],s1[66],s1[67],s1[68],s1[69],s1[70],s1[71],s1[72],s1[73],s1[74],s1[75],s1[76],s1[77],s1[78],s1[79],s1[80],s1[81],s1[82],s1[83],s1[84],s1[85],s1[86],s1[87],s1[88],s1[89],s1[90],s1[91],s1[92],s1[93],s1[94],s1[95],s1[96],s1[97],s1[98],s100[0],s91[10],s91[11],s91[12],s91[13],s91[14],s91[15],s91[16],s91[17],s91[18],s91[19],s91[20],s91[21],s91[22],s91[23],s91[24],s91[25],s91[26],s91[27],s91[28],s91[29],s91[30],s91[31],s91[32],s91[33],s91[34],s91[35],s91[36],s91[37],s91[38],s89[41],s87[44],s85[47],s83[50],s82[52],s82[53],s82[54],s82[55],s82[56],s82[57],s82[58],s82[59],s82[60],s82[61],s82[62],s82[63],s82[64],s82[65],s82[66],s82[67],s82[68],s82[69],s82[70],s82[71],s82[72],s82[73],s82[74],s82[75],s82[76],s81[78],s80[80],s79[82],s78[84],s77[86],s76[88],s75[90],s74[92],s73[94],s72[96],s71[98],s9[161],s7[164],s5[167],s3[170],s1[173],s74[101],s73[103],s72[105],s71[107],s70[109],s69[111],s68[113],s67[115],s66[117],s65[119],s64[121],s63[123],s62[125],s61[127],s60[129],s59[131],s58[133],s57[135],s56[137],s55[139],s54[141],s53[143],s52[145],s51[147],s50[149],s49[151],s48[153],s47[155],s46[157],s45[159],s44[161],s43[163],s42[165],s41[167],s40[169],s39[171],s38[173],s37[175],s36[177],s35[179],s34[181],s33[183],s32[185],s31[187],s30[189],s29[191],s28[193],s27[195],s26[197],s25[199],s24[201],s23[203],s22[205],s21[207],s20[209],s19[211],s18[213],s17[215],s16[217],s15[219],s14[221],s13[223],s12[225],s11[227],s10[229],s236[340],s235[342],s234[344],s233[346],s232[348],s231[350],s230[352],s229[354],s228[356],s227[358],s226[360],s225[362],s224[316],s223[318],s222[320],s221[322],s220[324],s219[326],s219[327],s219[328],s219[329],s219[330],s219[331],s219[332],s219[333],s219[334],s219[335],s219[336],s219[337],s219[338],s219[339],s219[340],s219[341],s219[342],s219[343],s219[344],s219[345],s219[346],s219[347],s219[348],s219[349],s219[350],s219[351],s219[352],s219[353],s219[354],s219[355],s219[356],s219[357],s219[358],s219[359],s219[360],s219[361],s219[362],s219[363],s219[364],s219[365],s219[366],s219[367],s219[368],s219[369],s219[370],s219[371],s219[372],s219[373],s219[374],s219[375],s219[376],s219[377],s219[378],s219[379],s219[380],s219[381],s219[382],s219[383],s219[384],s219[385],s219[386],s219[387],s219[388],s219[389],s219[390],s218[392],s217[394],s216[396],s215[398],s214[400],s213[402],s212[404],s211[406],s210[408],s209[410],s208[412],s207[414],s206[416],s205[418],s204[420],s203[422],s202[424],s201[426],s200[428],s199[430],s198[432],s197[434],s196[436],s195[438],s194[440],s193[442],pp255[220],pp254[222],pp253[224],pp252[226],pp251[228],pp250[230],pp251[230],pp252[230],pp253[230]};
    CLA_456 KS_237(s237, c237, in237_1, in237_2);
    wire[453:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {pp22[7],pp21[9],pp8[23],pp8[24],pp8[25],pp8[26],pp8[27],pp8[28],pp8[29],s237[10],s237[11],s237[12],s237[13],s237[14],s237[15],s237[16],s237[17],s237[18],s237[19],s237[20],s237[21],s237[22],s237[23],s237[24],s237[25],s237[26],s237[27],s237[28],s237[29],s237[30],s237[31],s237[32],s237[33],s237[34],s237[35],s237[36],s237[37],s237[38],s237[39],s237[40],s237[41],s237[42],s237[43],s237[44],s237[45],s237[46],s237[47],s237[48],s237[49],s237[50],s237[51],s237[52],s237[53],s237[54],s237[55],s237[56],s237[57],s237[58],s237[59],s237[60],s237[61],s237[62],s237[63],s237[64],s237[65],s237[66],s237[67],s237[68],s237[69],s237[70],s237[71],s237[72],s237[73],s237[74],s237[75],s237[76],s237[77],s235[80],s233[83],s231[86],s229[89],s229[90],s229[91],s229[92],s229[93],s229[94],s229[95],s229[96],s229[97],s229[98],s229[99],s224[57],s223[59],s222[61],s221[63],s220[65],s219[67],s218[69],s217[71],s237[100],s237[101],s237[102],s237[103],s237[104],s237[105],s237[106],s237[107],s237[108],s237[109],s237[110],s237[111],s237[112],s237[113],s237[114],s237[115],s237[116],s237[117],s237[118],s237[119],s237[120],s237[121],s237[122],s237[123],s237[124],s237[125],s237[126],s237[127],s237[128],s237[129],s237[130],s237[131],s237[132],s237[133],s237[134],s237[135],s237[136],s237[137],s237[138],s237[139],s237[140],s237[141],s237[142],s237[143],s237[144],s237[145],s237[146],s237[147],s237[148],s237[149],s237[150],s237[151],s237[152],s237[153],s237[154],s237[155],s237[156],s237[157],s237[158],s237[159],s237[160],s237[161],s237[162],s237[163],s237[164],s237[165],s237[166],s237[167],s237[168],s237[169],s237[170],s237[171],s237[172],s237[173],s237[174],s237[175],s237[176],s237[177],s237[178],s237[179],s237[180],s237[181],s237[182],s237[183],s237[184],s237[185],s237[186],s237[187],s237[188],s237[189],s237[190],s237[191],s237[192],s237[193],s237[194],s237[195],s237[196],s237[197],s237[198],s237[199],s237[200],s237[201],s237[202],s237[203],s237[204],s237[205],s237[206],s237[207],s237[208],s237[209],s237[210],s237[211],s237[212],s237[213],s237[214],s237[215],s237[216],s237[217],s237[218],s237[219],s237[220],s237[221],s237[222],s237[223],s237[224],s237[225],s237[226],s237[227],s237[228],s237[229],s237[230],s237[231],s237[232],s237[233],s237[234],s237[235],s237[236],s237[237],s237[238],s237[239],s237[240],s237[241],s237[242],s237[243],s237[244],s237[245],s237[246],s237[247],s237[248],s237[249],s237[250],s237[251],s237[252],s237[253],s237[254],s237[255],s237[256],s237[257],s237[258],s237[259],s237[260],s237[261],s237[262],s237[263],s237[264],s237[265],s237[266],s237[267],s237[268],s237[269],s237[270],s237[271],s237[272],s237[273],s237[274],s237[275],s237[276],s237[277],s237[278],s237[279],s237[280],s237[281],s237[282],s237[283],s237[284],s237[285],s237[286],s237[287],s237[288],s237[289],s237[290],s237[291],s237[292],s237[293],s237[294],s237[295],s237[296],s237[297],s237[298],s237[299],s237[300],s237[301],s237[302],s237[303],s237[304],s237[305],s237[306],s237[307],s237[308],s237[309],s237[310],s237[311],s237[312],s237[313],s237[314],s237[315],s237[316],s237[317],s237[318],s237[319],s237[320],s237[321],s237[322],s237[323],s237[324],s237[325],s237[326],s237[327],s237[328],s237[329],s237[330],s237[331],s237[332],s237[333],s237[334],s237[335],s237[336],s237[337],s237[338],s237[339],s236[341],s235[343],s234[345],s233[347],s232[349],s231[351],s230[353],s229[355],s228[357],s227[359],s226[361],s225[363],s224[317],s223[319],s222[321],s221[323],s220[325],s220[326],s220[327],s220[328],s220[329],s220[330],s220[331],s220[332],s220[333],s220[334],s220[335],s220[336],s220[337],s220[338],s220[339],s220[340],s220[341],s220[342],s220[343],s220[344],s220[345],s220[346],s220[347],s220[348],s220[349],s220[350],s220[351],s220[352],s220[353],s220[354],s220[355],s220[356],s220[357],s220[358],s220[359],s220[360],s220[361],s220[362],s220[363],s220[364],s220[365],s220[366],s220[367],s220[368],s220[369],s220[370],s220[371],s220[372],s220[373],s220[374],s220[375],s220[376],s220[377],s220[378],s220[379],s220[380],s220[381],s220[382],s220[383],s220[384],s220[385],s220[386],s220[387],s220[388],s220[389],s219[391],s218[393],s217[395],s216[397],s215[399],s214[401],s213[403],s212[405],s211[407],s210[409],s209[411],s208[413],s207[415],s206[417],s205[419],s204[421],s203[423],s202[425],s201[427],s200[429],s199[431],s198[433],s197[435],s196[437],s195[439],s194[441],s193[443],pp255[221],pp254[223],pp253[225],pp252[227],pp251[229],pp252[229],pp253[229]};
    assign in238_2 = {pp23[6],pp22[8],pp9[22],pp9[23],pp9[24],pp9[25],pp9[26],pp9[27],pp9[28],pp9[29],pp30[9],pp32[8],pp34[7],pp35[7],pp36[7],pp37[7],pp38[7],pp39[7],pp40[7],pp41[7],pp42[7],pp43[7],pp44[7],pp45[7],pp46[7],pp47[7],pp48[7],pp49[7],pp50[7],pp51[7],pp52[7],pp53[7],pp54[7],pp55[7],pp56[7],pp57[7],pp58[7],pp59[7],pp60[7],pp61[7],pp62[7],pp63[7],pp64[7],pp65[7],pp66[7],pp67[7],pp68[7],pp69[7],pp70[7],pp71[7],pp72[7],pp73[7],pp74[7],pp75[7],pp76[7],pp77[7],pp78[7],pp79[7],pp80[7],pp81[7],pp82[7],pp83[7],pp84[7],pp85[7],pp86[7],pp87[7],pp88[7],pp89[7],pp90[7],pp91[7],pp92[7],pp92[8],pp92[9],pp9[93],pp8[95],pp7[97],pp6[99],s236[79],s234[82],s232[85],s230[88],s230[89],s230[90],s230[91],s230[92],s230[93],s230[94],s230[95],s230[96],s230[97],s230[98],s230[99],s224[58],s223[60],s222[62],s221[64],s220[66],s219[68],s218[70],s217[72],s217[73],s217[74],s217[75],s217[76],s217[77],s217[78],s217[79],s217[80],s217[81],s218[81],s219[81],s220[81],s221[81],s222[81],s223[81],s224[81],s1[17],s2[17],s2[18],s2[19],s2[20],s2[21],s2[22],s2[23],s2[24],s2[25],s2[26],s2[27],s2[28],s2[29],s2[30],s2[31],s2[32],s2[33],s2[34],s2[35],s2[36],s2[37],s2[38],s2[39],s2[40],s2[41],s2[42],s2[43],s2[44],s2[45],s2[46],s2[47],s2[48],s2[49],s2[50],s2[51],s2[52],s2[53],s2[54],s2[55],s2[56],s2[57],s2[58],s2[59],s2[60],s2[61],s2[62],s2[63],s2[64],s2[65],s2[66],s2[67],s2[68],s2[69],s2[70],s2[71],s2[72],s2[73],s2[74],s2[75],s2[76],s2[77],s2[78],s2[79],s2[80],s2[81],s2[82],s2[83],s2[84],s2[85],s2[86],s2[87],s2[88],s2[89],s2[90],s2[91],s2[92],s2[93],s2[94],s2[95],s2[96],s2[97],s1[99],s100[1],s92[10],s92[11],s92[12],s92[13],s92[14],s92[15],s92[16],s92[17],s92[18],s92[19],s92[20],s92[21],s92[22],s92[23],s92[24],s92[25],s92[26],s92[27],s92[28],s92[29],s92[30],s92[31],s92[32],s92[33],s92[34],s92[35],s92[36],s92[37],s90[40],s88[43],s86[46],s84[49],s83[51],s83[52],s83[53],s83[54],s83[55],s83[56],s83[57],s83[58],s83[59],s83[60],s83[61],s83[62],s83[63],s83[64],s83[65],s83[66],s83[67],s83[68],s83[69],s83[70],s83[71],s83[72],s83[73],s83[74],s83[75],s82[77],s81[79],s80[81],s79[83],s78[85],s77[87],s76[89],s75[91],s74[93],s73[95],s72[97],s71[99],s8[163],s6[166],s4[169],s2[172],s75[100],s74[102],s73[104],s72[106],s71[108],s70[110],s69[112],s68[114],s67[116],s66[118],s65[120],s64[122],s63[124],s62[126],s61[128],s60[130],s59[132],s58[134],s57[136],s56[138],s55[140],s54[142],s53[144],s52[146],s51[148],s50[150],s49[152],s48[154],s47[156],s46[158],s45[160],s44[162],s43[164],s42[166],s41[168],s40[170],s39[172],s38[174],s37[176],s36[178],s35[180],s34[182],s33[184],s32[186],s31[188],s30[190],s29[192],s28[194],s27[196],s26[198],s25[200],s24[202],s23[204],s22[206],s21[208],s20[210],s19[212],s18[214],s17[216],s16[218],s15[220],s14[222],s13[224],s12[226],s11[228],s10[230],s237[340],s236[342],s235[344],s234[346],s233[348],s232[350],s231[352],s230[354],s229[356],s228[358],s227[360],s226[362],s225[364],s224[318],s223[320],s222[322],s221[324],s221[325],s221[326],s221[327],s221[328],s221[329],s221[330],s221[331],s221[332],s221[333],s221[334],s221[335],s221[336],s221[337],s221[338],s221[339],s221[340],s221[341],s221[342],s221[343],s221[344],s221[345],s221[346],s221[347],s221[348],s221[349],s221[350],s221[351],s221[352],s221[353],s221[354],s221[355],s221[356],s221[357],s221[358],s221[359],s221[360],s221[361],s221[362],s221[363],s221[364],s221[365],s221[366],s221[367],s221[368],s221[369],s221[370],s221[371],s221[372],s221[373],s221[374],s221[375],s221[376],s221[377],s221[378],s221[379],s221[380],s221[381],s221[382],s221[383],s221[384],s221[385],s221[386],s221[387],s221[388],s220[390],s219[392],s218[394],s217[396],s216[398],s215[400],s214[402],s213[404],s212[406],s211[408],s210[410],s209[412],s208[414],s207[416],s206[418],s205[420],s204[422],s203[424],s202[426],s201[428],s200[430],s199[432],s198[434],s197[436],s196[438],s195[440],s194[442],s193[444],pp255[222],pp254[224],pp253[226],pp252[228],pp253[228],pp254[228]};
    CLA_454 KS_238(s238, c238, in238_1, in238_2);
    wire[451:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {pp23[7],pp22[9],pp23[9],pp24[9],pp25[9],pp26[9],pp27[9],pp28[9],pp29[9],s238[10],s238[11],s238[12],s238[13],s238[14],s238[15],s238[16],s238[17],s238[18],s238[19],s238[20],s238[21],s238[22],s238[23],s238[24],s238[25],s238[26],s238[27],s238[28],s238[29],s238[30],s238[31],s238[32],s238[33],s238[34],s238[35],s238[36],s238[37],s238[38],s238[39],s238[40],s238[41],s238[42],s238[43],s238[44],s238[45],s238[46],s238[47],s238[48],s238[49],s238[50],s238[51],s238[52],s238[53],s238[54],s238[55],s238[56],s238[57],s238[58],s238[59],s238[60],s238[61],s238[62],s238[63],s238[64],s238[65],s238[66],s238[67],s238[68],s238[69],s238[70],s238[71],s238[72],s238[73],s238[74],s238[75],s238[76],s237[78],s235[81],s233[84],s231[87],s231[88],s231[89],s231[90],s231[91],s231[92],s231[93],s231[94],s231[95],s231[96],s231[97],s231[98],s231[99],s224[59],s223[61],s222[63],s221[65],s220[67],s219[69],s218[71],s238[100],s238[101],s238[102],s238[103],s238[104],s238[105],s238[106],s238[107],s238[108],s238[109],s238[110],s238[111],s238[112],s238[113],s238[114],s238[115],s238[116],s238[117],s238[118],s238[119],s238[120],s238[121],s238[122],s238[123],s238[124],s238[125],s238[126],s238[127],s238[128],s238[129],s238[130],s238[131],s238[132],s238[133],s238[134],s238[135],s238[136],s238[137],s238[138],s238[139],s238[140],s238[141],s238[142],s238[143],s238[144],s238[145],s238[146],s238[147],s238[148],s238[149],s238[150],s238[151],s238[152],s238[153],s238[154],s238[155],s238[156],s238[157],s238[158],s238[159],s238[160],s238[161],s238[162],s238[163],s238[164],s238[165],s238[166],s238[167],s238[168],s238[169],s238[170],s238[171],s238[172],s238[173],s238[174],s238[175],s238[176],s238[177],s238[178],s238[179],s238[180],s238[181],s238[182],s238[183],s238[184],s238[185],s238[186],s238[187],s238[188],s238[189],s238[190],s238[191],s238[192],s238[193],s238[194],s238[195],s238[196],s238[197],s238[198],s238[199],s238[200],s238[201],s238[202],s238[203],s238[204],s238[205],s238[206],s238[207],s238[208],s238[209],s238[210],s238[211],s238[212],s238[213],s238[214],s238[215],s238[216],s238[217],s238[218],s238[219],s238[220],s238[221],s238[222],s238[223],s238[224],s238[225],s238[226],s238[227],s238[228],s238[229],s238[230],s238[231],s238[232],s238[233],s238[234],s238[235],s238[236],s238[237],s238[238],s238[239],s238[240],s238[241],s238[242],s238[243],s238[244],s238[245],s238[246],s238[247],s238[248],s238[249],s238[250],s238[251],s238[252],s238[253],s238[254],s238[255],s238[256],s238[257],s238[258],s238[259],s238[260],s238[261],s238[262],s238[263],s238[264],s238[265],s238[266],s238[267],s238[268],s238[269],s238[270],s238[271],s238[272],s238[273],s238[274],s238[275],s238[276],s238[277],s238[278],s238[279],s238[280],s238[281],s238[282],s238[283],s238[284],s238[285],s238[286],s238[287],s238[288],s238[289],s238[290],s238[291],s238[292],s238[293],s238[294],s238[295],s238[296],s238[297],s238[298],s238[299],s238[300],s238[301],s238[302],s238[303],s238[304],s238[305],s238[306],s238[307],s238[308],s238[309],s238[310],s238[311],s238[312],s238[313],s238[314],s238[315],s238[316],s238[317],s238[318],s238[319],s238[320],s238[321],s238[322],s238[323],s238[324],s238[325],s238[326],s238[327],s238[328],s238[329],s238[330],s238[331],s238[332],s238[333],s238[334],s238[335],s238[336],s238[337],s238[338],s238[339],s237[341],s236[343],s235[345],s234[347],s233[349],s232[351],s231[353],s230[355],s229[357],s228[359],s227[361],s226[363],s225[365],s224[319],s223[321],s222[323],s222[324],s222[325],s222[326],s222[327],s222[328],s222[329],s222[330],s222[331],s222[332],s222[333],s222[334],s222[335],s222[336],s222[337],s222[338],s222[339],s222[340],s222[341],s222[342],s222[343],s222[344],s222[345],s222[346],s222[347],s222[348],s222[349],s222[350],s222[351],s222[352],s222[353],s222[354],s222[355],s222[356],s222[357],s222[358],s222[359],s222[360],s222[361],s222[362],s222[363],s222[364],s222[365],s222[366],s222[367],s222[368],s222[369],s222[370],s222[371],s222[372],s222[373],s222[374],s222[375],s222[376],s222[377],s222[378],s222[379],s222[380],s222[381],s222[382],s222[383],s222[384],s222[385],s222[386],s222[387],s221[389],s220[391],s219[393],s218[395],s217[397],s216[399],s215[401],s214[403],s213[405],s212[407],s211[409],s210[411],s209[413],s208[415],s207[417],s206[419],s205[421],s204[423],s203[425],s202[427],s201[429],s200[431],s199[433],s198[435],s197[437],s196[439],s195[441],s194[443],s193[445],pp255[223],pp254[225],pp253[227],pp254[227]};
    assign in239_2 = {pp24[6],pp23[8],pp24[8],pp25[8],pp26[8],pp27[8],pp28[8],pp29[8],pp30[8],pp31[8],pp33[7],pp35[6],pp36[6],pp37[6],pp38[6],pp39[6],pp40[6],pp41[6],pp42[6],pp43[6],pp44[6],pp45[6],pp46[6],pp47[6],pp48[6],pp49[6],pp50[6],pp51[6],pp52[6],pp53[6],pp54[6],pp55[6],pp56[6],pp57[6],pp58[6],pp59[6],pp60[6],pp61[6],pp62[6],pp63[6],pp64[6],pp65[6],pp66[6],pp67[6],pp68[6],pp69[6],pp70[6],pp71[6],pp72[6],pp73[6],pp74[6],pp75[6],pp76[6],pp77[6],pp78[6],pp79[6],pp80[6],pp81[6],pp82[6],pp83[6],pp84[6],pp85[6],pp86[6],pp87[6],pp88[6],pp89[6],pp90[6],pp91[6],pp92[6],pp93[6],pp93[7],pp93[8],pp93[9],pp9[94],pp8[96],pp7[98],s238[77],s236[80],s234[83],s232[86],s232[87],s232[88],s232[89],s232[90],s232[91],s232[92],s232[93],s232[94],s232[95],s232[96],s232[97],s232[98],s232[99],s224[60],s223[62],s222[64],s221[66],s220[68],s219[70],s218[72],s218[73],s218[74],s218[75],s218[76],s218[77],s218[78],s218[79],s218[80],s219[80],s220[80],s221[80],s222[80],s223[80],s224[80],s1[16],s2[16],s3[16],s3[17],s3[18],s3[19],s3[20],s3[21],s3[22],s3[23],s3[24],s3[25],s3[26],s3[27],s3[28],s3[29],s3[30],s3[31],s3[32],s3[33],s3[34],s3[35],s3[36],s3[37],s3[38],s3[39],s3[40],s3[41],s3[42],s3[43],s3[44],s3[45],s3[46],s3[47],s3[48],s3[49],s3[50],s3[51],s3[52],s3[53],s3[54],s3[55],s3[56],s3[57],s3[58],s3[59],s3[60],s3[61],s3[62],s3[63],s3[64],s3[65],s3[66],s3[67],s3[68],s3[69],s3[70],s3[71],s3[72],s3[73],s3[74],s3[75],s3[76],s3[77],s3[78],s3[79],s3[80],s3[81],s3[82],s3[83],s3[84],s3[85],s3[86],s3[87],s3[88],s3[89],s3[90],s3[91],s3[92],s3[93],s3[94],s3[95],s3[96],s2[98],s101[0],s100[2],s93[10],s93[11],s93[12],s93[13],s93[14],s93[15],s93[16],s93[17],s93[18],s93[19],s93[20],s93[21],s93[22],s93[23],s93[24],s93[25],s93[26],s93[27],s93[28],s93[29],s93[30],s93[31],s93[32],s93[33],s93[34],s93[35],s93[36],s91[39],s89[42],s87[45],s85[48],s84[50],s84[51],s84[52],s84[53],s84[54],s84[55],s84[56],s84[57],s84[58],s84[59],s84[60],s84[61],s84[62],s84[63],s84[64],s84[65],s84[66],s84[67],s84[68],s84[69],s84[70],s84[71],s84[72],s84[73],s84[74],s83[76],s82[78],s81[80],s80[82],s79[84],s78[86],s77[88],s76[90],s75[92],s74[94],s73[96],s72[98],s9[162],s7[165],s5[168],s3[171],s1[174],s75[101],s74[103],s73[105],s72[107],s71[109],s70[111],s69[113],s68[115],s67[117],s66[119],s65[121],s64[123],s63[125],s62[127],s61[129],s60[131],s59[133],s58[135],s57[137],s56[139],s55[141],s54[143],s53[145],s52[147],s51[149],s50[151],s49[153],s48[155],s47[157],s46[159],s45[161],s44[163],s43[165],s42[167],s41[169],s40[171],s39[173],s38[175],s37[177],s36[179],s35[181],s34[183],s33[185],s32[187],s31[189],s30[191],s29[193],s28[195],s27[197],s26[199],s25[201],s24[203],s23[205],s22[207],s21[209],s20[211],s19[213],s18[215],s17[217],s16[219],s15[221],s14[223],s13[225],s12[227],s11[229],s10[231],s238[340],s237[342],s236[344],s235[346],s234[348],s233[350],s232[352],s231[354],s230[356],s229[358],s228[360],s227[362],s226[364],s225[366],s224[320],s223[322],s223[323],s223[324],s223[325],s223[326],s223[327],s223[328],s223[329],s223[330],s223[331],s223[332],s223[333],s223[334],s223[335],s223[336],s223[337],s223[338],s223[339],s223[340],s223[341],s223[342],s223[343],s223[344],s223[345],s223[346],s223[347],s223[348],s223[349],s223[350],s223[351],s223[352],s223[353],s223[354],s223[355],s223[356],s223[357],s223[358],s223[359],s223[360],s223[361],s223[362],s223[363],s223[364],s223[365],s223[366],s223[367],s223[368],s223[369],s223[370],s223[371],s223[372],s223[373],s223[374],s223[375],s223[376],s223[377],s223[378],s223[379],s223[380],s223[381],s223[382],s223[383],s223[384],s223[385],s223[386],s222[388],s221[390],s220[392],s219[394],s218[396],s217[398],s216[400],s215[402],s214[404],s213[406],s212[408],s211[410],s210[412],s209[414],s208[416],s207[418],s206[420],s205[422],s204[424],s203[426],s202[428],s201[430],s200[432],s199[434],s198[436],s197[438],s196[440],s195[442],s194[444],s193[446],pp255[224],pp254[226],pp255[226]};
    CLA_452 KS_239(s239, c239, in239_1, in239_2);
    wire[449:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {pp24[7],pp25[7],pp26[7],pp27[7],pp28[7],pp29[7],pp30[7],pp31[7],pp32[7],s239[10],s239[11],s239[12],s239[13],s239[14],s239[15],s239[16],s239[17],s239[18],s239[19],s239[20],s239[21],s239[22],s239[23],s239[24],s239[25],s239[26],s239[27],s239[28],s239[29],s239[30],s239[31],s239[32],s239[33],s239[34],s239[35],s239[36],s239[37],s239[38],s239[39],s239[40],s239[41],s239[42],s239[43],s239[44],s239[45],s239[46],s239[47],s239[48],s239[49],s239[50],s239[51],s239[52],s239[53],s239[54],s239[55],s239[56],s239[57],s239[58],s239[59],s239[60],s239[61],s239[62],s239[63],s239[64],s239[65],s239[66],s239[67],s239[68],s239[69],s239[70],s239[71],s239[72],s239[73],s239[74],s239[75],s239[76],s237[79],s235[82],s233[85],s233[86],s233[87],s233[88],s233[89],s233[90],s233[91],s233[92],s233[93],s233[94],s233[95],s233[96],s233[97],s233[98],s233[99],s224[61],s223[63],s222[65],s221[67],s220[69],s219[71],s239[100],s239[101],s239[102],s239[103],s239[104],s239[105],s239[106],s239[107],s239[108],s239[109],s239[110],s239[111],s239[112],s239[113],s239[114],s239[115],s239[116],s239[117],s239[118],s239[119],s239[120],s239[121],s239[122],s239[123],s239[124],s239[125],s239[126],s239[127],s239[128],s239[129],s239[130],s239[131],s239[132],s239[133],s239[134],s239[135],s239[136],s239[137],s239[138],s239[139],s239[140],s239[141],s239[142],s239[143],s239[144],s239[145],s239[146],s239[147],s239[148],s239[149],s239[150],s239[151],s239[152],s239[153],s239[154],s239[155],s239[156],s239[157],s239[158],s239[159],s239[160],s239[161],s239[162],s239[163],s239[164],s239[165],s239[166],s239[167],s239[168],s239[169],s239[170],s239[171],s239[172],s239[173],s239[174],s239[175],s239[176],s239[177],s239[178],s239[179],s239[180],s239[181],s239[182],s239[183],s239[184],s239[185],s239[186],s239[187],s239[188],s239[189],s239[190],s239[191],s239[192],s239[193],s239[194],s239[195],s239[196],s239[197],s239[198],s239[199],s239[200],s239[201],s239[202],s239[203],s239[204],s239[205],s239[206],s239[207],s239[208],s239[209],s239[210],s239[211],s239[212],s239[213],s239[214],s239[215],s239[216],s239[217],s239[218],s239[219],s239[220],s239[221],s239[222],s239[223],s239[224],s239[225],s239[226],s239[227],s239[228],s239[229],s239[230],s239[231],s239[232],s239[233],s239[234],s239[235],s239[236],s239[237],s239[238],s239[239],s239[240],s239[241],s239[242],s239[243],s239[244],s239[245],s239[246],s239[247],s239[248],s239[249],s239[250],s239[251],s239[252],s239[253],s239[254],s239[255],s239[256],s239[257],s239[258],s239[259],s239[260],s239[261],s239[262],s239[263],s239[264],s239[265],s239[266],s239[267],s239[268],s239[269],s239[270],s239[271],s239[272],s239[273],s239[274],s239[275],s239[276],s239[277],s239[278],s239[279],s239[280],s239[281],s239[282],s239[283],s239[284],s239[285],s239[286],s239[287],s239[288],s239[289],s239[290],s239[291],s239[292],s239[293],s239[294],s239[295],s239[296],s239[297],s239[298],s239[299],s239[300],s239[301],s239[302],s239[303],s239[304],s239[305],s239[306],s239[307],s239[308],s239[309],s239[310],s239[311],s239[312],s239[313],s239[314],s239[315],s239[316],s239[317],s239[318],s239[319],s239[320],s239[321],s239[322],s239[323],s239[324],s239[325],s239[326],s239[327],s239[328],s239[329],s239[330],s239[331],s239[332],s239[333],s239[334],s239[335],s239[336],s239[337],s239[338],s239[339],s238[341],s237[343],s236[345],s235[347],s234[349],s233[351],s232[353],s231[355],s230[357],s229[359],s228[361],s227[363],s226[365],s225[367],s224[321],s224[322],s224[323],s224[324],s224[325],s224[326],s224[327],s224[328],s224[329],s224[330],s224[331],s224[332],s224[333],s224[334],s224[335],s224[336],s224[337],s224[338],s224[339],s224[340],s224[341],s224[342],s224[343],s224[344],s224[345],s224[346],s224[347],s224[348],s224[349],s224[350],s224[351],s224[352],s224[353],s224[354],s224[355],s224[356],s224[357],s224[358],s224[359],s224[360],s224[361],s224[362],s224[363],s224[364],s224[365],s224[366],s224[367],s224[368],s224[369],s224[370],s224[371],s224[372],s224[373],s224[374],s224[375],s224[376],s224[377],s224[378],s224[379],s224[380],s224[381],s224[382],s224[383],s224[384],s224[385],s223[387],s222[389],s221[391],s220[393],s219[395],s218[397],s217[399],s216[401],s215[403],s214[405],s213[407],s212[409],s211[411],s210[413],s209[415],s208[417],s207[419],s206[421],s205[423],s204[425],s203[427],s202[429],s201[431],s200[433],s199[435],s198[437],s197[439],s196[441],s195[443],s194[445],s193[447],pp255[225]};
    assign in240_2 = {pp25[6],pp26[6],pp27[6],pp28[6],pp29[6],pp30[6],pp31[6],pp32[6],pp33[6],pp34[6],pp36[5],pp37[5],pp38[5],pp39[5],pp40[5],pp41[5],pp42[5],pp43[5],pp44[5],pp45[5],pp46[5],pp47[5],pp48[5],pp49[5],pp50[5],pp51[5],pp52[5],pp53[5],pp54[5],pp55[5],pp56[5],pp57[5],pp58[5],pp59[5],pp60[5],pp61[5],pp62[5],pp63[5],pp64[5],pp65[5],pp66[5],pp67[5],pp68[5],pp69[5],pp70[5],pp71[5],pp72[5],pp73[5],pp74[5],pp75[5],pp76[5],pp77[5],pp78[5],pp79[5],pp80[5],pp81[5],pp82[5],pp83[5],pp84[5],pp85[5],pp86[5],pp87[5],pp88[5],pp89[5],pp90[5],pp91[5],pp92[5],pp93[5],pp94[5],pp94[6],pp94[7],pp94[8],pp94[9],pp9[95],pp8[97],pp7[99],s238[78],s236[81],s234[84],s234[85],s234[86],s234[87],s234[88],s234[89],s234[90],s234[91],s234[92],s234[93],s234[94],s234[95],s234[96],s234[97],s234[98],s234[99],s224[62],s223[64],s222[66],s221[68],s220[70],s219[72],s219[73],s219[74],s219[75],s219[76],s219[77],s219[78],s219[79],s220[79],s221[79],s222[79],s223[79],s224[79],s1[15],s2[15],s3[15],s4[15],s4[16],s4[17],s4[18],s4[19],s4[20],s4[21],s4[22],s4[23],s4[24],s4[25],s4[26],s4[27],s4[28],s4[29],s4[30],s4[31],s4[32],s4[33],s4[34],s4[35],s4[36],s4[37],s4[38],s4[39],s4[40],s4[41],s4[42],s4[43],s4[44],s4[45],s4[46],s4[47],s4[48],s4[49],s4[50],s4[51],s4[52],s4[53],s4[54],s4[55],s4[56],s4[57],s4[58],s4[59],s4[60],s4[61],s4[62],s4[63],s4[64],s4[65],s4[66],s4[67],s4[68],s4[69],s4[70],s4[71],s4[72],s4[73],s4[74],s4[75],s4[76],s4[77],s4[78],s4[79],s4[80],s4[81],s4[82],s4[83],s4[84],s4[85],s4[86],s4[87],s4[88],s4[89],s4[90],s4[91],s4[92],s4[93],s4[94],s4[95],s3[97],s2[99],s101[1],s100[3],s94[10],s94[11],s94[12],s94[13],s94[14],s94[15],s94[16],s94[17],s94[18],s94[19],s94[20],s94[21],s94[22],s94[23],s94[24],s94[25],s94[26],s94[27],s94[28],s94[29],s94[30],s94[31],s94[32],s94[33],s94[34],s94[35],s92[38],s90[41],s88[44],s86[47],s85[49],s85[50],s85[51],s85[52],s85[53],s85[54],s85[55],s85[56],s85[57],s85[58],s85[59],s85[60],s85[61],s85[62],s85[63],s85[64],s85[65],s85[66],s85[67],s85[68],s85[69],s85[70],s85[71],s85[72],s85[73],s84[75],s83[77],s82[79],s81[81],s80[83],s79[85],s78[87],s77[89],s76[91],s75[93],s74[95],s73[97],s72[99],s8[164],s6[167],s4[170],s2[173],s76[100],s75[102],s74[104],s73[106],s72[108],s71[110],s70[112],s69[114],s68[116],s67[118],s66[120],s65[122],s64[124],s63[126],s62[128],s61[130],s60[132],s59[134],s58[136],s57[138],s56[140],s55[142],s54[144],s53[146],s52[148],s51[150],s50[152],s49[154],s48[156],s47[158],s46[160],s45[162],s44[164],s43[166],s42[168],s41[170],s40[172],s39[174],s38[176],s37[178],s36[180],s35[182],s34[184],s33[186],s32[188],s31[190],s30[192],s29[194],s28[196],s27[198],s26[200],s25[202],s24[204],s23[206],s22[208],s21[210],s20[212],s19[214],s18[216],s17[218],s16[220],s15[222],s14[224],s13[226],s12[228],s11[230],s10[232],s239[340],s238[342],s237[344],s236[346],s235[348],s234[350],s233[352],s232[354],s231[356],s230[358],s229[360],s228[362],s227[364],s226[366],s225[368],s225[369],s225[370],s225[371],s225[372],s225[373],s225[374],s225[375],s225[376],s225[377],s225[378],s225[379],s225[380],s225[381],s225[382],s225[383],s225[384],s225[385],s225[386],s225[387],s225[388],s225[389],s225[390],s225[391],s225[392],s225[393],s225[394],s225[395],s225[396],s225[397],s225[398],s225[399],s225[400],s225[401],s225[402],s225[403],s225[404],s225[405],s225[406],s225[407],s225[408],s225[409],s225[410],s225[411],s225[412],s225[413],s225[414],s225[415],s225[416],s225[417],s225[418],s225[419],s225[420],s225[421],s225[422],s225[423],s225[424],s225[425],s225[426],s225[427],s225[428],s225[429],s225[430],s225[431],s225[432],s225[433],s225[434],s225[435],s225[436],s225[437],s225[438],s225[439],s225[440],s225[441],s225[442],s225[443],s225[444],s225[445],s225[446],s225[447],s225[448],s225[449],s225[450],s225[451],s225[452],s225[453],s225[454],s225[455],s225[456],s225[457],s225[458],s225[459],s225[460],s225[461],s225[462],s225[463],s225[464]};
    CLA_450 KS_240(s240, c240, in240_1, in240_2);

    /*Stage 5*/
    wire[495:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {pp0[8],pp0[9],pp0[10],pp0[11],pp0[12],pp0[13],pp0[14],pp0[15],pp2[14],pp4[13],pp6[12],pp8[11],pp9[11],pp12[9],pp14[8],pp16[7],pp18[6],pp20[5],pp21[5],pp22[5],pp23[5],pp24[5],pp25[5],pp26[5],pp27[5],pp28[5],pp29[5],pp30[5],pp31[5],pp32[5],pp33[5],pp34[5],pp35[5],s240[10],s240[11],s240[12],s240[13],s240[14],s240[15],s240[16],s240[17],s240[18],s240[19],s240[20],s240[21],s240[22],s240[23],s240[24],s240[25],s240[26],s240[27],s240[28],s240[29],s240[30],s240[31],s240[32],s240[33],s240[34],s240[35],s240[36],s240[37],s240[38],s240[39],s240[40],s240[41],s240[42],s240[43],s240[44],s240[45],s240[46],s240[47],s240[48],s240[49],s240[50],s240[51],s240[52],s240[53],s240[54],s240[55],s240[56],s240[57],s240[58],s240[59],s240[60],s240[61],s240[62],s240[63],s240[64],s240[65],s240[66],s240[67],s240[68],s240[69],s240[70],s240[71],s240[72],s240[73],s240[74],s240[75],s239[77],s237[80],s235[83],s235[84],s235[85],s235[86],s235[87],s235[88],s235[89],s235[90],s235[91],s235[92],s235[93],s235[94],s235[95],s235[96],s235[97],s235[98],s235[99],s224[63],s223[65],s222[67],s221[69],s220[71],s240[100],s240[101],s240[102],s240[103],s240[104],s240[105],s240[106],s240[107],s240[108],s240[109],s240[110],s240[111],s240[112],s240[113],s240[114],s240[115],s240[116],s240[117],s240[118],s240[119],s240[120],s240[121],s240[122],s240[123],s240[124],s240[125],s240[126],s240[127],s240[128],s240[129],s240[130],s240[131],s240[132],s240[133],s240[134],s240[135],s240[136],s240[137],s240[138],s240[139],s240[140],s240[141],s240[142],s240[143],s240[144],s240[145],s240[146],s240[147],s240[148],s240[149],s240[150],s240[151],s240[152],s240[153],s240[154],s240[155],s240[156],s240[157],s240[158],s240[159],s240[160],s240[161],s240[162],s240[163],s240[164],s240[165],s240[166],s240[167],s240[168],s240[169],s240[170],s240[171],s240[172],s240[173],s240[174],s240[175],s240[176],s240[177],s240[178],s240[179],s240[180],s240[181],s240[182],s240[183],s240[184],s240[185],s240[186],s240[187],s240[188],s240[189],s240[190],s240[191],s240[192],s240[193],s240[194],s240[195],s240[196],s240[197],s240[198],s240[199],s240[200],s240[201],s240[202],s240[203],s240[204],s240[205],s240[206],s240[207],s240[208],s240[209],s240[210],s240[211],s240[212],s240[213],s240[214],s240[215],s240[216],s240[217],s240[218],s240[219],s240[220],s240[221],s240[222],s240[223],s240[224],s240[225],s240[226],s240[227],s240[228],s240[229],s240[230],s240[231],s240[232],s240[233],s240[234],s240[235],s240[236],s240[237],s240[238],s240[239],s240[240],s240[241],s240[242],s240[243],s240[244],s240[245],s240[246],s240[247],s240[248],s240[249],s240[250],s240[251],s240[252],s240[253],s240[254],s240[255],s240[256],s240[257],s240[258],s240[259],s240[260],s240[261],s240[262],s240[263],s240[264],s240[265],s240[266],s240[267],s240[268],s240[269],s240[270],s240[271],s240[272],s240[273],s240[274],s240[275],s240[276],s240[277],s240[278],s240[279],s240[280],s240[281],s240[282],s240[283],s240[284],s240[285],s240[286],s240[287],s240[288],s240[289],s240[290],s240[291],s240[292],s240[293],s240[294],s240[295],s240[296],s240[297],s240[298],s240[299],s240[300],s240[301],s240[302],s240[303],s240[304],s240[305],s240[306],s240[307],s240[308],s240[309],s240[310],s240[311],s240[312],s240[313],s240[314],s240[315],s240[316],s240[317],s240[318],s240[319],s240[320],s240[321],s240[322],s240[323],s240[324],s240[325],s240[326],s240[327],s240[328],s240[329],s240[330],s240[331],s240[332],s240[333],s240[334],s240[335],s240[336],s240[337],s240[338],s240[339],s239[341],s238[343],s237[345],s236[347],s235[349],s234[351],s233[353],s232[355],s231[357],s230[359],s229[361],s228[363],s227[365],s226[367],s226[368],s226[369],s226[370],s226[371],s226[372],s226[373],s226[374],s226[375],s226[376],s226[377],s226[378],s226[379],s226[380],s226[381],s226[382],s226[383],s226[384],s226[385],s226[386],s226[387],s226[388],s226[389],s226[390],s226[391],s226[392],s226[393],s226[394],s226[395],s226[396],s226[397],s226[398],s226[399],s226[400],s226[401],s226[402],s226[403],s226[404],s226[405],s226[406],s226[407],s226[408],s226[409],s226[410],s226[411],s226[412],s226[413],s226[414],s226[415],s226[416],s226[417],s226[418],s226[419],s226[420],s226[421],s226[422],s226[423],s226[424],s226[425],s226[426],s226[427],s226[428],s226[429],s226[430],s226[431],s226[432],s226[433],s226[434],s226[435],s226[436],s226[437],s226[438],s226[439],s226[440],s226[441],s226[442],s226[443],s226[444],s226[445],s226[446],s226[447],s226[448],s226[449],s226[450],s226[451],s226[452],s226[453],s226[454],s226[455],s226[456],s226[457],s226[458],s226[459],s226[460],s226[461],s226[462],s226[463],s225[465],pp255[227],pp254[229],pp253[231],pp252[233],pp251[235],pp250[237],pp249[239],pp248[241],pp247[243],pp246[245],pp245[247],pp244[249],pp243[251],pp242[253],pp241[255],pp242[255],pp243[255],pp244[255],pp245[255],pp246[255],pp247[255],pp248[255]};
    assign in241_2 = {pp1[7],pp1[8],pp10[0],pp1[10],pp1[11],pp1[12],pp1[13],pp1[14],pp3[13],pp5[12],pp7[11],pp9[10],pp11[9],pp13[8],pp15[7],pp17[6],pp19[5],pp21[4],pp22[4],pp23[4],pp24[4],pp25[4],pp26[4],pp27[4],pp28[4],pp29[4],pp30[4],pp31[4],pp32[4],pp33[4],pp34[4],pp35[4],pp36[4],pp37[4],pp38[4],pp39[4],pp40[4],pp41[4],pp42[4],pp43[4],pp44[4],pp45[4],pp46[4],pp47[4],pp48[4],pp49[4],pp50[4],pp51[4],pp52[4],pp53[4],pp54[4],pp55[4],pp56[4],pp57[4],pp58[4],pp59[4],pp60[4],pp61[4],pp62[4],pp63[4],pp64[4],pp65[4],pp66[4],pp67[4],pp68[4],pp69[4],pp70[4],pp71[4],pp72[4],pp73[4],pp74[4],pp75[4],pp76[4],pp77[4],pp78[4],pp79[4],pp80[4],pp81[4],pp82[4],pp83[4],pp84[4],pp85[4],pp86[4],pp87[4],pp88[4],pp89[4],pp90[4],pp91[4],pp92[4],pp93[4],pp94[4],pp95[4],pp95[5],pp95[6],pp95[7],pp95[8],pp95[9],pp9[96],pp8[98],s240[76],s238[79],s236[82],s236[83],s236[84],s236[85],s236[86],s236[87],s236[88],s236[89],s236[90],s236[91],s236[92],s236[93],s236[94],s236[95],s236[96],s236[97],s236[98],s236[99],s224[64],s223[66],s222[68],s221[70],s220[72],s220[73],s220[74],s220[75],s220[76],s220[77],s220[78],s221[78],s222[78],s223[78],s224[78],s1[14],s2[14],s3[14],s4[14],s5[14],s5[15],s5[16],s5[17],s5[18],s5[19],s5[20],s5[21],s5[22],s5[23],s5[24],s5[25],s5[26],s5[27],s5[28],s5[29],s5[30],s5[31],s5[32],s5[33],s5[34],s5[35],s5[36],s5[37],s5[38],s5[39],s5[40],s5[41],s5[42],s5[43],s5[44],s5[45],s5[46],s5[47],s5[48],s5[49],s5[50],s5[51],s5[52],s5[53],s5[54],s5[55],s5[56],s5[57],s5[58],s5[59],s5[60],s5[61],s5[62],s5[63],s5[64],s5[65],s5[66],s5[67],s5[68],s5[69],s5[70],s5[71],s5[72],s5[73],s5[74],s5[75],s5[76],s5[77],s5[78],s5[79],s5[80],s5[81],s5[82],s5[83],s5[84],s5[85],s5[86],s5[87],s5[88],s5[89],s5[90],s5[91],s5[92],s5[93],s5[94],s4[96],s3[98],s102[0],s101[2],s100[4],s95[10],s95[11],s95[12],s95[13],s95[14],s95[15],s95[16],s95[17],s95[18],s95[19],s95[20],s95[21],s95[22],s95[23],s95[24],s95[25],s95[26],s95[27],s95[28],s95[29],s95[30],s95[31],s95[32],s95[33],s95[34],s93[37],s91[40],s89[43],s87[46],s86[48],s86[49],s86[50],s86[51],s86[52],s86[53],s86[54],s86[55],s86[56],s86[57],s86[58],s86[59],s86[60],s86[61],s86[62],s86[63],s86[64],s86[65],s86[66],s86[67],s86[68],s86[69],s86[70],s86[71],s86[72],s85[74],s84[76],s83[78],s82[80],s81[82],s80[84],s79[86],s78[88],s77[90],s76[92],s75[94],s74[96],s73[98],s9[163],s7[166],s5[169],s3[172],s1[175],s76[101],s75[103],s74[105],s73[107],s72[109],s71[111],s70[113],s69[115],s68[117],s67[119],s66[121],s65[123],s64[125],s63[127],s62[129],s61[131],s60[133],s59[135],s58[137],s57[139],s56[141],s55[143],s54[145],s53[147],s52[149],s51[151],s50[153],s49[155],s48[157],s47[159],s46[161],s45[163],s44[165],s43[167],s42[169],s41[171],s40[173],s39[175],s38[177],s37[179],s36[181],s35[183],s34[185],s33[187],s32[189],s31[191],s30[193],s29[195],s28[197],s27[199],s26[201],s25[203],s24[205],s23[207],s22[209],s21[211],s20[213],s19[215],s18[217],s17[219],s16[221],s15[223],s14[225],s13[227],s12[229],s11[231],s10[233],s240[340],s239[342],s238[344],s237[346],s236[348],s235[350],s234[352],s233[354],s232[356],s231[358],s230[360],s229[362],s228[364],s227[366],s227[367],s227[368],s227[369],s227[370],s227[371],s227[372],s227[373],s227[374],s227[375],s227[376],s227[377],s227[378],s227[379],s227[380],s227[381],s227[382],s227[383],s227[384],s227[385],s227[386],s227[387],s227[388],s227[389],s227[390],s227[391],s227[392],s227[393],s227[394],s227[395],s227[396],s227[397],s227[398],s227[399],s227[400],s227[401],s227[402],s227[403],s227[404],s227[405],s227[406],s227[407],s227[408],s227[409],s227[410],s227[411],s227[412],s227[413],s227[414],s227[415],s227[416],s227[417],s227[418],s227[419],s227[420],s227[421],s227[422],s227[423],s227[424],s227[425],s227[426],s227[427],s227[428],s227[429],s227[430],s227[431],s227[432],s227[433],s227[434],s227[435],s227[436],s227[437],s227[438],s227[439],s227[440],s227[441],s227[442],s227[443],s227[444],s227[445],s227[446],s227[447],s227[448],s227[449],s227[450],s227[451],s227[452],s227[453],s227[454],s227[455],s227[456],s227[457],s227[458],s227[459],s227[460],s227[461],s227[462],s226[464],s225[466],pp255[228],pp254[230],pp253[232],pp252[234],pp251[236],pp250[238],pp249[240],pp248[242],pp247[244],pp246[246],pp245[248],pp244[250],pp243[252],pp242[254],pp243[254],pp244[254],pp245[254],pp246[254],pp247[254],pp248[254],pp249[254]};
    CLA_496 KS_241(s241, c241, in241_1, in241_2);
    wire[493:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {pp2[7],s241[2],pp10[1],pp2[10],pp2[11],pp2[12],pp2[13],pp4[12],pp6[11],s241[10],s241[11],s241[12],s241[13],s241[14],s241[15],s241[16],s241[17],s241[18],s241[19],s241[20],s241[21],s241[22],s241[23],s241[24],s241[25],s241[26],s241[27],s241[28],s241[29],s241[30],s241[31],s241[32],s241[33],s241[34],s241[35],s241[36],s241[37],s241[38],s241[39],s241[40],s241[41],s241[42],s241[43],s241[44],s241[45],s241[46],s241[47],s241[48],s241[49],s241[50],s241[51],s241[52],s241[53],s241[54],s241[55],s241[56],s241[57],s241[58],s241[59],s241[60],s241[61],s241[62],s241[63],s241[64],s241[65],s241[66],s241[67],s241[68],s241[69],s241[70],s241[71],s241[72],s241[73],s241[74],s241[75],s241[76],s241[77],s241[78],s241[79],s241[80],s241[81],s241[82],s241[83],s241[84],s241[85],s241[86],s241[87],s241[88],s241[89],s241[90],s241[91],s241[92],s241[93],s241[94],s241[95],s241[96],s241[97],s241[98],s241[99],s241[100],s241[101],s241[102],s241[103],s241[104],s241[105],s241[106],s241[107],s241[108],s241[109],s241[110],s241[111],s241[112],s241[113],s241[114],s241[115],s241[116],s241[117],s241[118],s241[119],s241[120],s241[121],s241[122],s241[123],s241[124],s241[125],s241[126],s241[127],s241[128],s241[129],s241[130],s241[131],s241[132],s241[133],s241[134],s241[135],s241[136],s241[137],s241[138],s241[139],s241[140],s241[141],s241[142],s241[143],s241[144],s241[145],s241[146],s241[147],s241[148],s241[149],s241[150],s241[151],s241[152],s241[153],s241[154],s241[155],s241[156],s241[157],s241[158],s241[159],s241[160],s241[161],s241[162],s241[163],s241[164],s241[165],s241[166],s241[167],s241[168],s241[169],s241[170],s241[171],s241[172],s241[173],s241[174],s241[175],s241[176],s241[177],s241[178],s241[179],s241[180],s241[181],s241[182],s241[183],s241[184],s241[185],s241[186],s241[187],s241[188],s241[189],s241[190],s241[191],s241[192],s241[193],s241[194],s241[195],s241[196],s241[197],s241[198],s241[199],s241[200],s241[201],s241[202],s241[203],s241[204],s241[205],s241[206],s241[207],s241[208],s241[209],s241[210],s241[211],s241[212],s241[213],s241[214],s241[215],s241[216],s241[217],s241[218],s241[219],s241[220],s241[221],s241[222],s241[223],s241[224],s241[225],s241[226],s241[227],s241[228],s241[229],s241[230],s241[231],s241[232],s241[233],s241[234],s241[235],s241[236],s241[237],s241[238],s241[239],s241[240],s241[241],s241[242],s241[243],s241[244],s241[245],s241[246],s241[247],s241[248],s241[249],s241[250],s241[251],s241[252],s241[253],s241[254],s241[255],s241[256],s241[257],s241[258],s241[259],s241[260],s241[261],s241[262],s241[263],s241[264],s241[265],s241[266],s241[267],s241[268],s241[269],s241[270],s241[271],s241[272],s241[273],s241[274],s241[275],s241[276],s241[277],s241[278],s241[279],s241[280],s241[281],s241[282],s241[283],s241[284],s241[285],s241[286],s241[287],s241[288],s241[289],s241[290],s241[291],s241[292],s241[293],s241[294],s241[295],s241[296],s241[297],s241[298],s241[299],s241[300],s241[301],s241[302],s241[303],s241[304],s241[305],s241[306],s241[307],s241[308],s241[309],s241[310],s241[311],s241[312],s241[313],s241[314],s241[315],s241[316],s241[317],s241[318],s241[319],s241[320],s241[321],s241[322],s241[323],s241[324],s241[325],s241[326],s241[327],s241[328],s241[329],s241[330],s241[331],s241[332],s241[333],s241[334],s241[335],s241[336],s241[337],s241[338],s241[339],s241[340],s241[341],s241[342],s241[343],s241[344],s241[345],s241[346],s241[347],s241[348],s241[349],s241[350],s241[351],s241[352],s241[353],s241[354],s241[355],s241[356],s241[357],s241[358],s241[359],s241[360],s241[361],s241[362],s241[363],s240[341],s239[343],s238[345],s237[347],s236[349],s235[351],s234[353],s233[355],s232[357],s231[359],s230[361],s229[363],s228[365],s228[366],s228[367],s228[368],s228[369],s228[370],s228[371],s228[372],s228[373],s228[374],s228[375],s228[376],s228[377],s228[378],s228[379],s228[380],s228[381],s228[382],s228[383],s228[384],s228[385],s228[386],s228[387],s228[388],s228[389],s228[390],s228[391],s228[392],s228[393],s228[394],s228[395],s228[396],s228[397],s228[398],s228[399],s228[400],s228[401],s228[402],s228[403],s228[404],s228[405],s228[406],s228[407],s228[408],s228[409],s228[410],s228[411],s228[412],s228[413],s228[414],s228[415],s228[416],s228[417],s228[418],s228[419],s228[420],s228[421],s228[422],s228[423],s228[424],s228[425],s228[426],s228[427],s228[428],s228[429],s228[430],s228[431],s228[432],s228[433],s228[434],s228[435],s228[436],s228[437],s228[438],s228[439],s228[440],s228[441],s228[442],s228[443],s228[444],s228[445],s228[446],s228[447],s228[448],s228[449],s228[450],s228[451],s228[452],s228[453],s228[454],s228[455],s228[456],s228[457],s228[458],s228[459],s228[460],s228[461],s227[463],s226[465],s225[467],pp255[229],pp254[231],pp253[233],pp252[235],pp251[237],pp250[239],pp249[241],pp248[243],pp247[245],pp246[247],pp245[249],pp244[251],pp243[253],pp244[253],pp245[253],pp246[253],pp247[253],pp248[253],pp249[253]};
    assign in242_2 = {pp3[6],pp1[9],pp11[0],pp10[2],pp3[10],pp3[11],pp3[12],pp5[11],pp7[10],pp8[10],pp10[9],pp12[8],pp14[7],pp16[6],pp18[5],pp20[4],pp22[3],pp23[3],pp24[3],pp25[3],pp26[3],pp27[3],pp28[3],pp29[3],pp30[3],pp31[3],pp32[3],pp33[3],pp34[3],pp35[3],pp36[3],pp37[3],pp38[3],pp39[3],pp40[3],pp41[3],pp42[3],pp43[3],pp44[3],pp45[3],pp46[3],pp47[3],pp48[3],pp49[3],pp50[3],pp51[3],pp52[3],pp53[3],pp54[3],pp55[3],pp56[3],pp57[3],pp58[3],pp59[3],pp60[3],pp61[3],pp62[3],pp63[3],pp64[3],pp65[3],pp66[3],pp67[3],pp68[3],pp69[3],pp70[3],pp71[3],pp72[3],pp73[3],pp74[3],pp75[3],pp76[3],pp77[3],pp78[3],pp79[3],pp80[3],pp81[3],pp82[3],pp83[3],pp84[3],pp85[3],pp86[3],pp87[3],pp88[3],pp89[3],pp90[3],pp91[3],pp92[3],pp93[3],pp94[3],pp95[3],pp96[3],pp96[4],pp96[5],pp96[6],pp96[7],pp96[8],pp96[9],pp9[97],pp8[99],s239[78],s237[81],s237[82],s237[83],s237[84],s237[85],s237[86],s237[87],s237[88],s237[89],s237[90],s237[91],s237[92],s237[93],s237[94],s237[95],s237[96],s237[97],s237[98],s237[99],s224[65],s223[67],s222[69],s221[71],s221[72],s221[73],s221[74],s221[75],s221[76],s221[77],s222[77],s223[77],s224[77],s1[13],s2[13],s3[13],s4[13],s5[13],s6[13],s6[14],s6[15],s6[16],s6[17],s6[18],s6[19],s6[20],s6[21],s6[22],s6[23],s6[24],s6[25],s6[26],s6[27],s6[28],s6[29],s6[30],s6[31],s6[32],s6[33],s6[34],s6[35],s6[36],s6[37],s6[38],s6[39],s6[40],s6[41],s6[42],s6[43],s6[44],s6[45],s6[46],s6[47],s6[48],s6[49],s6[50],s6[51],s6[52],s6[53],s6[54],s6[55],s6[56],s6[57],s6[58],s6[59],s6[60],s6[61],s6[62],s6[63],s6[64],s6[65],s6[66],s6[67],s6[68],s6[69],s6[70],s6[71],s6[72],s6[73],s6[74],s6[75],s6[76],s6[77],s6[78],s6[79],s6[80],s6[81],s6[82],s6[83],s6[84],s6[85],s6[86],s6[87],s6[88],s6[89],s6[90],s6[91],s6[92],s6[93],s5[95],s4[97],s3[99],s102[1],s101[3],s100[5],s96[10],s96[11],s96[12],s96[13],s96[14],s96[15],s96[16],s96[17],s96[18],s96[19],s96[20],s96[21],s96[22],s96[23],s96[24],s96[25],s96[26],s96[27],s96[28],s96[29],s96[30],s96[31],s96[32],s96[33],s94[36],s92[39],s90[42],s88[45],s87[47],s87[48],s87[49],s87[50],s87[51],s87[52],s87[53],s87[54],s87[55],s87[56],s87[57],s87[58],s87[59],s87[60],s87[61],s87[62],s87[63],s87[64],s87[65],s87[66],s87[67],s87[68],s87[69],s87[70],s87[71],s86[73],s85[75],s84[77],s83[79],s82[81],s81[83],s80[85],s79[87],s78[89],s77[91],s76[93],s75[95],s74[97],s73[99],s8[165],s6[168],s4[171],s2[174],s77[100],s76[102],s75[104],s74[106],s73[108],s72[110],s71[112],s70[114],s69[116],s68[118],s67[120],s66[122],s65[124],s64[126],s63[128],s62[130],s61[132],s60[134],s59[136],s58[138],s57[140],s56[142],s55[144],s54[146],s53[148],s52[150],s51[152],s50[154],s49[156],s48[158],s47[160],s46[162],s45[164],s44[166],s43[168],s42[170],s41[172],s40[174],s39[176],s38[178],s37[180],s36[182],s35[184],s34[186],s33[188],s32[190],s31[192],s30[194],s29[196],s28[198],s27[200],s26[202],s25[204],s24[206],s23[208],s22[210],s21[212],s20[214],s19[216],s18[218],s17[220],s16[222],s15[224],s14[226],s13[228],s12[230],s11[232],s10[234],s241[364],s240[342],s239[344],s238[346],s237[348],s236[350],s235[352],s234[354],s233[356],s232[358],s231[360],s230[362],s229[364],s229[365],s229[366],s229[367],s229[368],s229[369],s229[370],s229[371],s229[372],s229[373],s229[374],s229[375],s229[376],s229[377],s229[378],s229[379],s229[380],s229[381],s229[382],s229[383],s229[384],s229[385],s229[386],s229[387],s229[388],s229[389],s229[390],s229[391],s229[392],s229[393],s229[394],s229[395],s229[396],s229[397],s229[398],s229[399],s229[400],s229[401],s229[402],s229[403],s229[404],s229[405],s229[406],s229[407],s229[408],s229[409],s229[410],s229[411],s229[412],s229[413],s229[414],s229[415],s229[416],s229[417],s229[418],s229[419],s229[420],s229[421],s229[422],s229[423],s229[424],s229[425],s229[426],s229[427],s229[428],s229[429],s229[430],s229[431],s229[432],s229[433],s229[434],s229[435],s229[436],s229[437],s229[438],s229[439],s229[440],s229[441],s229[442],s229[443],s229[444],s229[445],s229[446],s229[447],s229[448],s229[449],s229[450],s229[451],s229[452],s229[453],s229[454],s229[455],s229[456],s229[457],s229[458],s229[459],s229[460],s228[462],s227[464],s226[466],s225[468],pp255[230],pp254[232],pp253[234],pp252[236],pp251[238],pp250[240],pp249[242],pp248[244],pp247[246],pp246[248],pp245[250],pp244[252],pp245[252],pp246[252],pp247[252],pp248[252],pp249[252],pp250[252]};
    CLA_494 KS_242(s242, c242, in242_1, in242_2);
    wire[491:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {pp2[8],s241[3],pp11[1],pp10[3],pp4[10],pp4[11],pp6[10],pp10[7],pp10[8],s242[10],s242[11],s242[12],s242[13],s242[14],s242[15],s242[16],s242[17],s242[18],s242[19],s242[20],s242[21],s242[22],s242[23],s242[24],s242[25],s242[26],s242[27],s242[28],s242[29],s242[30],s242[31],s242[32],s242[33],s242[34],s242[35],s242[36],s242[37],s242[38],s242[39],s242[40],s242[41],s242[42],s242[43],s242[44],s242[45],s242[46],s242[47],s242[48],s242[49],s242[50],s242[51],s242[52],s242[53],s242[54],s242[55],s242[56],s242[57],s242[58],s242[59],s242[60],s242[61],s242[62],s242[63],s242[64],s242[65],s242[66],s242[67],s242[68],s242[69],s242[70],s242[71],s242[72],s242[73],s242[74],s242[75],s242[76],s242[77],s242[78],s242[79],s242[80],s242[81],s242[82],s242[83],s242[84],s242[85],s242[86],s242[87],s242[88],s242[89],s242[90],s242[91],s242[92],s242[93],s242[94],s242[95],s242[96],s242[97],s242[98],s240[77],s242[100],s242[101],s242[102],s242[103],s242[104],s242[105],s242[106],s242[107],s242[108],s242[109],s242[110],s242[111],s242[112],s242[113],s242[114],s242[115],s242[116],s242[117],s242[118],s242[119],s242[120],s242[121],s242[122],s242[123],s242[124],s242[125],s242[126],s242[127],s242[128],s242[129],s242[130],s242[131],s242[132],s242[133],s242[134],s242[135],s242[136],s242[137],s242[138],s242[139],s242[140],s242[141],s242[142],s242[143],s242[144],s242[145],s242[146],s242[147],s242[148],s242[149],s242[150],s242[151],s242[152],s242[153],s242[154],s242[155],s242[156],s242[157],s242[158],s242[159],s242[160],s242[161],s242[162],s242[163],s242[164],s242[165],s242[166],s242[167],s242[168],s242[169],s242[170],s242[171],s242[172],s242[173],s242[174],s242[175],s242[176],s242[177],s242[178],s242[179],s242[180],s242[181],s242[182],s242[183],s242[184],s242[185],s242[186],s242[187],s242[188],s242[189],s242[190],s242[191],s242[192],s242[193],s242[194],s242[195],s242[196],s242[197],s242[198],s242[199],s242[200],s242[201],s242[202],s242[203],s242[204],s242[205],s242[206],s242[207],s242[208],s242[209],s242[210],s242[211],s242[212],s242[213],s242[214],s242[215],s242[216],s242[217],s242[218],s242[219],s242[220],s242[221],s242[222],s242[223],s242[224],s242[225],s242[226],s242[227],s242[228],s242[229],s242[230],s242[231],s242[232],s242[233],s242[234],s242[235],s242[236],s242[237],s242[238],s242[239],s242[240],s242[241],s242[242],s242[243],s242[244],s242[245],s242[246],s242[247],s242[248],s242[249],s242[250],s242[251],s242[252],s242[253],s242[254],s242[255],s242[256],s242[257],s242[258],s242[259],s242[260],s242[261],s242[262],s242[263],s242[264],s242[265],s242[266],s242[267],s242[268],s242[269],s242[270],s242[271],s242[272],s242[273],s242[274],s242[275],s242[276],s242[277],s242[278],s242[279],s242[280],s242[281],s242[282],s242[283],s242[284],s242[285],s242[286],s242[287],s242[288],s242[289],s242[290],s242[291],s242[292],s242[293],s242[294],s242[295],s242[296],s242[297],s242[298],s242[299],s242[300],s242[301],s242[302],s242[303],s242[304],s242[305],s242[306],s242[307],s242[308],s242[309],s242[310],s242[311],s242[312],s242[313],s242[314],s242[315],s242[316],s242[317],s242[318],s242[319],s242[320],s242[321],s242[322],s242[323],s242[324],s242[325],s242[326],s242[327],s242[328],s242[329],s242[330],s242[331],s242[332],s242[333],s242[334],s242[335],s242[336],s242[337],s242[338],s242[339],s242[340],s242[341],s242[342],s242[343],s242[344],s242[345],s242[346],s242[347],s242[348],s242[349],s242[350],s242[351],s242[352],s242[353],s242[354],s242[355],s242[356],s242[357],s242[358],s242[359],s242[360],s242[361],s242[362],s242[363],s241[365],s240[343],s239[345],s238[347],s237[349],s236[351],s235[353],s234[355],s233[357],s232[359],s231[361],s230[363],s230[364],s230[365],s230[366],s230[367],s230[368],s230[369],s230[370],s230[371],s230[372],s230[373],s230[374],s230[375],s230[376],s230[377],s230[378],s230[379],s230[380],s230[381],s230[382],s230[383],s230[384],s230[385],s230[386],s230[387],s230[388],s230[389],s230[390],s230[391],s230[392],s230[393],s230[394],s230[395],s230[396],s230[397],s230[398],s230[399],s230[400],s230[401],s230[402],s230[403],s230[404],s230[405],s230[406],s230[407],s230[408],s230[409],s230[410],s230[411],s230[412],s230[413],s230[414],s230[415],s230[416],s230[417],s230[418],s230[419],s230[420],s230[421],s230[422],s230[423],s230[424],s230[425],s230[426],s230[427],s230[428],s230[429],s230[430],s230[431],s230[432],s230[433],s230[434],s230[435],s230[436],s230[437],s230[438],s230[439],s230[440],s230[441],s230[442],s230[443],s230[444],s230[445],s230[446],s230[447],s230[448],s230[449],s230[450],s230[451],s230[452],s230[453],s230[454],s230[455],s230[456],s230[457],s230[458],s230[459],s229[461],s228[463],s227[465],s226[467],s225[469],pp255[231],pp254[233],pp253[235],pp252[237],pp251[239],pp250[241],pp249[243],pp248[245],pp247[247],pp246[249],pp245[251],pp246[251],pp247[251],pp248[251],pp249[251],pp250[251]};
    assign in243_2 = {pp3[7],s242[2],pp12[0],pp11[2],pp10[4],pp5[10],pp10[6],pp11[6],pp11[7],pp11[8],pp13[7],pp15[6],pp17[5],pp19[4],pp21[3],pp23[2],pp24[2],pp25[2],pp26[2],pp27[2],pp28[2],pp29[2],pp30[2],pp31[2],pp32[2],pp33[2],pp34[2],pp35[2],pp36[2],pp37[2],pp38[2],pp39[2],pp40[2],pp41[2],pp42[2],pp43[2],pp44[2],pp45[2],pp46[2],pp47[2],pp48[2],pp49[2],pp50[2],pp51[2],pp52[2],pp53[2],pp54[2],pp55[2],pp56[2],pp57[2],pp58[2],pp59[2],pp60[2],pp61[2],pp62[2],pp63[2],pp64[2],pp65[2],pp66[2],pp67[2],pp68[2],pp69[2],pp70[2],pp71[2],pp72[2],pp73[2],pp74[2],pp75[2],pp76[2],pp77[2],pp78[2],pp79[2],pp80[2],pp81[2],pp82[2],pp83[2],pp84[2],pp85[2],pp86[2],pp87[2],pp88[2],pp89[2],pp90[2],pp91[2],pp92[2],pp93[2],pp94[2],pp95[2],pp96[2],pp97[2],pp97[3],pp97[4],pp97[5],pp97[6],pp97[7],pp97[8],pp97[9],pp9[98],s242[99],s238[80],s238[81],s238[82],s238[83],s238[84],s238[85],s238[86],s238[87],s238[88],s238[89],s238[90],s238[91],s238[92],s238[93],s238[94],s238[95],s238[96],s238[97],s238[98],s238[99],s224[66],s223[68],s222[70],s222[71],s222[72],s222[73],s222[74],s222[75],s222[76],s223[76],s224[76],s1[12],s2[12],s3[12],s4[12],s5[12],s6[12],s7[12],s7[13],s7[14],s7[15],s7[16],s7[17],s7[18],s7[19],s7[20],s7[21],s7[22],s7[23],s7[24],s7[25],s7[26],s7[27],s7[28],s7[29],s7[30],s7[31],s7[32],s7[33],s7[34],s7[35],s7[36],s7[37],s7[38],s7[39],s7[40],s7[41],s7[42],s7[43],s7[44],s7[45],s7[46],s7[47],s7[48],s7[49],s7[50],s7[51],s7[52],s7[53],s7[54],s7[55],s7[56],s7[57],s7[58],s7[59],s7[60],s7[61],s7[62],s7[63],s7[64],s7[65],s7[66],s7[67],s7[68],s7[69],s7[70],s7[71],s7[72],s7[73],s7[74],s7[75],s7[76],s7[77],s7[78],s7[79],s7[80],s7[81],s7[82],s7[83],s7[84],s7[85],s7[86],s7[87],s7[88],s7[89],s7[90],s7[91],s7[92],s6[94],s5[96],s4[98],s103[0],s102[2],s101[4],s100[6],s97[10],s97[11],s97[12],s97[13],s97[14],s97[15],s97[16],s97[17],s97[18],s97[19],s97[20],s97[21],s97[22],s97[23],s97[24],s97[25],s97[26],s97[27],s97[28],s97[29],s97[30],s97[31],s97[32],s95[35],s93[38],s91[41],s89[44],s88[46],s88[47],s88[48],s88[49],s88[50],s88[51],s88[52],s88[53],s88[54],s88[55],s88[56],s88[57],s88[58],s88[59],s88[60],s88[61],s88[62],s88[63],s88[64],s88[65],s88[66],s88[67],s88[68],s88[69],s88[70],s87[72],s86[74],s85[76],s84[78],s83[80],s82[82],s81[84],s80[86],s79[88],s78[90],s77[92],s76[94],s75[96],s74[98],s9[164],s7[167],s5[170],s3[173],s1[176],s77[101],s76[103],s75[105],s74[107],s73[109],s72[111],s71[113],s70[115],s69[117],s68[119],s67[121],s66[123],s65[125],s64[127],s63[129],s62[131],s61[133],s60[135],s59[137],s58[139],s57[141],s56[143],s55[145],s54[147],s53[149],s52[151],s51[153],s50[155],s49[157],s48[159],s47[161],s46[163],s45[165],s44[167],s43[169],s42[171],s41[173],s40[175],s39[177],s38[179],s37[181],s36[183],s35[185],s34[187],s33[189],s32[191],s31[193],s30[195],s29[197],s28[199],s27[201],s26[203],s25[205],s24[207],s23[209],s22[211],s21[213],s20[215],s19[217],s18[219],s17[221],s16[223],s15[225],s14[227],s13[229],s12[231],s11[233],s10[235],s242[364],s241[366],s240[344],s239[346],s238[348],s237[350],s236[352],s235[354],s234[356],s233[358],s232[360],s231[362],s231[363],s231[364],s231[365],s231[366],s231[367],s231[368],s231[369],s231[370],s231[371],s231[372],s231[373],s231[374],s231[375],s231[376],s231[377],s231[378],s231[379],s231[380],s231[381],s231[382],s231[383],s231[384],s231[385],s231[386],s231[387],s231[388],s231[389],s231[390],s231[391],s231[392],s231[393],s231[394],s231[395],s231[396],s231[397],s231[398],s231[399],s231[400],s231[401],s231[402],s231[403],s231[404],s231[405],s231[406],s231[407],s231[408],s231[409],s231[410],s231[411],s231[412],s231[413],s231[414],s231[415],s231[416],s231[417],s231[418],s231[419],s231[420],s231[421],s231[422],s231[423],s231[424],s231[425],s231[426],s231[427],s231[428],s231[429],s231[430],s231[431],s231[432],s231[433],s231[434],s231[435],s231[436],s231[437],s231[438],s231[439],s231[440],s231[441],s231[442],s231[443],s231[444],s231[445],s231[446],s231[447],s231[448],s231[449],s231[450],s231[451],s231[452],s231[453],s231[454],s231[455],s231[456],s231[457],s231[458],s230[460],s229[462],s228[464],s227[466],s226[468],s225[470],pp255[232],pp254[234],pp253[236],pp252[238],pp251[240],pp250[242],pp249[244],pp248[246],pp247[248],pp246[250],pp247[250],pp248[250],pp249[250],pp250[250],pp251[250]};
    CLA_492 KS_243(s243, c243, in243_1, in243_2);
    wire[489:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp2[9],s241[4],pp12[1],pp11[3],pp10[5],pp11[5],pp12[5],pp12[6],pp12[7],s243[10],s243[11],s243[12],s243[13],s243[14],s243[15],s243[16],s243[17],s243[18],s243[19],s243[20],s243[21],s243[22],s243[23],s243[24],s243[25],s243[26],s243[27],s243[28],s243[29],s243[30],s243[31],s243[32],s243[33],s243[34],s243[35],s243[36],s243[37],s243[38],s243[39],s243[40],s243[41],s243[42],s243[43],s243[44],s243[45],s243[46],s243[47],s243[48],s243[49],s243[50],s243[51],s243[52],s243[53],s243[54],s243[55],s243[56],s243[57],s243[58],s243[59],s243[60],s243[61],s243[62],s243[63],s243[64],s243[65],s243[66],s243[67],s243[68],s243[69],s243[70],s243[71],s243[72],s243[73],s243[74],s243[75],s243[76],s243[77],s243[78],s243[79],s243[80],s243[81],s243[82],s243[83],s243[84],s243[85],s243[86],s243[87],s243[88],s243[89],s243[90],s243[91],s243[92],s243[93],s243[94],s243[95],s243[96],s243[97],s243[98],s239[79],s243[100],s243[101],s243[102],s243[103],s243[104],s243[105],s243[106],s243[107],s243[108],s243[109],s243[110],s243[111],s243[112],s243[113],s243[114],s243[115],s243[116],s243[117],s243[118],s243[119],s243[120],s243[121],s243[122],s243[123],s243[124],s243[125],s243[126],s243[127],s243[128],s243[129],s243[130],s243[131],s243[132],s243[133],s243[134],s243[135],s243[136],s243[137],s243[138],s243[139],s243[140],s243[141],s243[142],s243[143],s243[144],s243[145],s243[146],s243[147],s243[148],s243[149],s243[150],s243[151],s243[152],s243[153],s243[154],s243[155],s243[156],s243[157],s243[158],s243[159],s243[160],s243[161],s243[162],s243[163],s243[164],s243[165],s243[166],s243[167],s243[168],s243[169],s243[170],s243[171],s243[172],s243[173],s243[174],s243[175],s243[176],s243[177],s243[178],s243[179],s243[180],s243[181],s243[182],s243[183],s243[184],s243[185],s243[186],s243[187],s243[188],s243[189],s243[190],s243[191],s243[192],s243[193],s243[194],s243[195],s243[196],s243[197],s243[198],s243[199],s243[200],s243[201],s243[202],s243[203],s243[204],s243[205],s243[206],s243[207],s243[208],s243[209],s243[210],s243[211],s243[212],s243[213],s243[214],s243[215],s243[216],s243[217],s243[218],s243[219],s243[220],s243[221],s243[222],s243[223],s243[224],s243[225],s243[226],s243[227],s243[228],s243[229],s243[230],s243[231],s243[232],s243[233],s243[234],s243[235],s243[236],s243[237],s243[238],s243[239],s243[240],s243[241],s243[242],s243[243],s243[244],s243[245],s243[246],s243[247],s243[248],s243[249],s243[250],s243[251],s243[252],s243[253],s243[254],s243[255],s243[256],s243[257],s243[258],s243[259],s243[260],s243[261],s243[262],s243[263],s243[264],s243[265],s243[266],s243[267],s243[268],s243[269],s243[270],s243[271],s243[272],s243[273],s243[274],s243[275],s243[276],s243[277],s243[278],s243[279],s243[280],s243[281],s243[282],s243[283],s243[284],s243[285],s243[286],s243[287],s243[288],s243[289],s243[290],s243[291],s243[292],s243[293],s243[294],s243[295],s243[296],s243[297],s243[298],s243[299],s243[300],s243[301],s243[302],s243[303],s243[304],s243[305],s243[306],s243[307],s243[308],s243[309],s243[310],s243[311],s243[312],s243[313],s243[314],s243[315],s243[316],s243[317],s243[318],s243[319],s243[320],s243[321],s243[322],s243[323],s243[324],s243[325],s243[326],s243[327],s243[328],s243[329],s243[330],s243[331],s243[332],s243[333],s243[334],s243[335],s243[336],s243[337],s243[338],s243[339],s243[340],s243[341],s243[342],s243[343],s243[344],s243[345],s243[346],s243[347],s243[348],s243[349],s243[350],s243[351],s243[352],s243[353],s243[354],s243[355],s243[356],s243[357],s243[358],s243[359],s243[360],s243[361],s243[362],s243[363],s242[365],s241[367],s240[345],s239[347],s238[349],s237[351],s236[353],s235[355],s234[357],s233[359],s232[361],s232[362],s232[363],s232[364],s232[365],s232[366],s232[367],s232[368],s232[369],s232[370],s232[371],s232[372],s232[373],s232[374],s232[375],s232[376],s232[377],s232[378],s232[379],s232[380],s232[381],s232[382],s232[383],s232[384],s232[385],s232[386],s232[387],s232[388],s232[389],s232[390],s232[391],s232[392],s232[393],s232[394],s232[395],s232[396],s232[397],s232[398],s232[399],s232[400],s232[401],s232[402],s232[403],s232[404],s232[405],s232[406],s232[407],s232[408],s232[409],s232[410],s232[411],s232[412],s232[413],s232[414],s232[415],s232[416],s232[417],s232[418],s232[419],s232[420],s232[421],s232[422],s232[423],s232[424],s232[425],s232[426],s232[427],s232[428],s232[429],s232[430],s232[431],s232[432],s232[433],s232[434],s232[435],s232[436],s232[437],s232[438],s232[439],s232[440],s232[441],s232[442],s232[443],s232[444],s232[445],s232[446],s232[447],s232[448],s232[449],s232[450],s232[451],s232[452],s232[453],s232[454],s232[455],s232[456],s232[457],s231[459],s230[461],s229[463],s228[465],s227[467],s226[469],s225[471],pp255[233],pp254[235],pp253[237],pp252[239],pp251[241],pp250[243],pp249[245],pp248[247],pp247[249],pp248[249],pp249[249],pp250[249],pp251[249]};
    assign in244_2 = {pp3[8],s242[3],pp13[0],pp12[2],pp11[4],pp12[4],pp13[4],pp13[5],pp13[6],pp14[6],pp16[5],pp18[4],pp20[3],pp22[2],pp24[1],pp25[1],pp26[1],pp27[1],pp28[1],pp29[1],pp30[1],pp31[1],pp32[1],pp33[1],pp34[1],pp35[1],pp36[1],pp37[1],pp38[1],pp39[1],pp40[1],pp41[1],pp42[1],pp43[1],pp44[1],pp45[1],pp46[1],pp47[1],pp48[1],pp49[1],pp50[1],pp51[1],pp52[1],pp53[1],pp54[1],pp55[1],pp56[1],pp57[1],pp58[1],pp59[1],pp60[1],pp61[1],pp62[1],pp63[1],pp64[1],pp65[1],pp66[1],pp67[1],pp68[1],pp69[1],pp70[1],pp71[1],pp72[1],pp73[1],pp74[1],pp75[1],pp76[1],pp77[1],pp78[1],pp79[1],pp80[1],pp81[1],pp82[1],pp83[1],pp84[1],pp85[1],pp86[1],pp87[1],pp88[1],pp89[1],pp90[1],pp91[1],pp92[1],pp93[1],pp94[1],pp95[1],pp96[1],pp97[1],pp98[1],pp98[2],pp98[3],pp98[4],pp98[5],pp98[6],pp98[7],pp98[8],pp98[9],pp9[99],s240[78],s239[80],s239[81],s239[82],s239[83],s239[84],s239[85],s239[86],s239[87],s239[88],s239[89],s239[90],s239[91],s239[92],s239[93],s239[94],s239[95],s239[96],s239[97],s239[98],s239[99],s224[67],s223[69],s223[70],s223[71],s223[72],s223[73],s223[74],s223[75],s224[75],s1[11],s2[11],s3[11],s4[11],s5[11],s6[11],s7[11],s8[11],s8[12],s8[13],s8[14],s8[15],s8[16],s8[17],s8[18],s8[19],s8[20],s8[21],s8[22],s8[23],s8[24],s8[25],s8[26],s8[27],s8[28],s8[29],s8[30],s8[31],s8[32],s8[33],s8[34],s8[35],s8[36],s8[37],s8[38],s8[39],s8[40],s8[41],s8[42],s8[43],s8[44],s8[45],s8[46],s8[47],s8[48],s8[49],s8[50],s8[51],s8[52],s8[53],s8[54],s8[55],s8[56],s8[57],s8[58],s8[59],s8[60],s8[61],s8[62],s8[63],s8[64],s8[65],s8[66],s8[67],s8[68],s8[69],s8[70],s8[71],s8[72],s8[73],s8[74],s8[75],s8[76],s8[77],s8[78],s8[79],s8[80],s8[81],s8[82],s8[83],s8[84],s8[85],s8[86],s8[87],s8[88],s8[89],s8[90],s8[91],s7[93],s6[95],s5[97],s4[99],s103[1],s102[3],s101[5],s100[7],s98[10],s98[11],s98[12],s98[13],s98[14],s98[15],s98[16],s98[17],s98[18],s98[19],s98[20],s98[21],s98[22],s98[23],s98[24],s98[25],s98[26],s98[27],s98[28],s98[29],s98[30],s98[31],s96[34],s94[37],s92[40],s90[43],s89[45],s89[46],s89[47],s89[48],s89[49],s89[50],s89[51],s89[52],s89[53],s89[54],s89[55],s89[56],s89[57],s89[58],s89[59],s89[60],s89[61],s89[62],s89[63],s89[64],s89[65],s89[66],s89[67],s89[68],s89[69],s88[71],s87[73],s86[75],s85[77],s84[79],s83[81],s82[83],s81[85],s80[87],s79[89],s78[91],s77[93],s76[95],s75[97],s74[99],s8[166],s6[169],s4[172],s2[175],s78[100],s77[102],s76[104],s75[106],s74[108],s73[110],s72[112],s71[114],s70[116],s69[118],s68[120],s67[122],s66[124],s65[126],s64[128],s63[130],s62[132],s61[134],s60[136],s59[138],s58[140],s57[142],s56[144],s55[146],s54[148],s53[150],s52[152],s51[154],s50[156],s49[158],s48[160],s47[162],s46[164],s45[166],s44[168],s43[170],s42[172],s41[174],s40[176],s39[178],s38[180],s37[182],s36[184],s35[186],s34[188],s33[190],s32[192],s31[194],s30[196],s29[198],s28[200],s27[202],s26[204],s25[206],s24[208],s23[210],s22[212],s21[214],s20[216],s19[218],s18[220],s17[222],s16[224],s15[226],s14[228],s13[230],s12[232],s11[234],s10[236],s243[364],s242[366],s241[368],s240[346],s239[348],s238[350],s237[352],s236[354],s235[356],s234[358],s233[360],s233[361],s233[362],s233[363],s233[364],s233[365],s233[366],s233[367],s233[368],s233[369],s233[370],s233[371],s233[372],s233[373],s233[374],s233[375],s233[376],s233[377],s233[378],s233[379],s233[380],s233[381],s233[382],s233[383],s233[384],s233[385],s233[386],s233[387],s233[388],s233[389],s233[390],s233[391],s233[392],s233[393],s233[394],s233[395],s233[396],s233[397],s233[398],s233[399],s233[400],s233[401],s233[402],s233[403],s233[404],s233[405],s233[406],s233[407],s233[408],s233[409],s233[410],s233[411],s233[412],s233[413],s233[414],s233[415],s233[416],s233[417],s233[418],s233[419],s233[420],s233[421],s233[422],s233[423],s233[424],s233[425],s233[426],s233[427],s233[428],s233[429],s233[430],s233[431],s233[432],s233[433],s233[434],s233[435],s233[436],s233[437],s233[438],s233[439],s233[440],s233[441],s233[442],s233[443],s233[444],s233[445],s233[446],s233[447],s233[448],s233[449],s233[450],s233[451],s233[452],s233[453],s233[454],s233[455],s233[456],s232[458],s231[460],s230[462],s229[464],s228[466],s227[468],s226[470],s225[472],pp255[234],pp254[236],pp253[238],pp252[240],pp251[242],pp250[244],pp249[246],pp248[248],pp249[248],pp250[248],pp251[248],pp252[248]};
    CLA_490 KS_244(s244, c244, in244_1, in244_2);
    wire[487:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {s243[2],s241[5],pp13[1],pp12[3],pp13[3],pp14[3],pp14[4],pp14[5],pp15[5],s244[10],s244[11],s244[12],s244[13],s244[14],s244[15],s244[16],s244[17],s244[18],s244[19],s244[20],s244[21],s244[22],s244[23],s244[24],s244[25],s244[26],s244[27],s244[28],s244[29],s244[30],s244[31],s244[32],s244[33],s244[34],s244[35],s244[36],s244[37],s244[38],s244[39],s244[40],s244[41],s244[42],s244[43],s244[44],s244[45],s244[46],s244[47],s244[48],s244[49],s244[50],s244[51],s244[52],s244[53],s244[54],s244[55],s244[56],s244[57],s244[58],s244[59],s244[60],s244[61],s244[62],s244[63],s244[64],s244[65],s244[66],s244[67],s244[68],s244[69],s244[70],s244[71],s244[72],s244[73],s244[74],s244[75],s244[76],s244[77],s244[78],s244[79],s244[80],s244[81],s244[82],s244[83],s244[84],s244[85],s244[86],s244[87],s244[88],s244[89],s244[90],s244[91],s244[92],s244[93],s244[94],s244[95],s244[96],s244[97],s243[99],s240[79],s244[100],s244[101],s244[102],s244[103],s244[104],s244[105],s244[106],s244[107],s244[108],s244[109],s244[110],s244[111],s244[112],s244[113],s244[114],s244[115],s244[116],s244[117],s244[118],s244[119],s244[120],s244[121],s244[122],s244[123],s244[124],s244[125],s244[126],s244[127],s244[128],s244[129],s244[130],s244[131],s244[132],s244[133],s244[134],s244[135],s244[136],s244[137],s244[138],s244[139],s244[140],s244[141],s244[142],s244[143],s244[144],s244[145],s244[146],s244[147],s244[148],s244[149],s244[150],s244[151],s244[152],s244[153],s244[154],s244[155],s244[156],s244[157],s244[158],s244[159],s244[160],s244[161],s244[162],s244[163],s244[164],s244[165],s244[166],s244[167],s244[168],s244[169],s244[170],s244[171],s244[172],s244[173],s244[174],s244[175],s244[176],s244[177],s244[178],s244[179],s244[180],s244[181],s244[182],s244[183],s244[184],s244[185],s244[186],s244[187],s244[188],s244[189],s244[190],s244[191],s244[192],s244[193],s244[194],s244[195],s244[196],s244[197],s244[198],s244[199],s244[200],s244[201],s244[202],s244[203],s244[204],s244[205],s244[206],s244[207],s244[208],s244[209],s244[210],s244[211],s244[212],s244[213],s244[214],s244[215],s244[216],s244[217],s244[218],s244[219],s244[220],s244[221],s244[222],s244[223],s244[224],s244[225],s244[226],s244[227],s244[228],s244[229],s244[230],s244[231],s244[232],s244[233],s244[234],s244[235],s244[236],s244[237],s244[238],s244[239],s244[240],s244[241],s244[242],s244[243],s244[244],s244[245],s244[246],s244[247],s244[248],s244[249],s244[250],s244[251],s244[252],s244[253],s244[254],s244[255],s244[256],s244[257],s244[258],s244[259],s244[260],s244[261],s244[262],s244[263],s244[264],s244[265],s244[266],s244[267],s244[268],s244[269],s244[270],s244[271],s244[272],s244[273],s244[274],s244[275],s244[276],s244[277],s244[278],s244[279],s244[280],s244[281],s244[282],s244[283],s244[284],s244[285],s244[286],s244[287],s244[288],s244[289],s244[290],s244[291],s244[292],s244[293],s244[294],s244[295],s244[296],s244[297],s244[298],s244[299],s244[300],s244[301],s244[302],s244[303],s244[304],s244[305],s244[306],s244[307],s244[308],s244[309],s244[310],s244[311],s244[312],s244[313],s244[314],s244[315],s244[316],s244[317],s244[318],s244[319],s244[320],s244[321],s244[322],s244[323],s244[324],s244[325],s244[326],s244[327],s244[328],s244[329],s244[330],s244[331],s244[332],s244[333],s244[334],s244[335],s244[336],s244[337],s244[338],s244[339],s244[340],s244[341],s244[342],s244[343],s244[344],s244[345],s244[346],s244[347],s244[348],s244[349],s244[350],s244[351],s244[352],s244[353],s244[354],s244[355],s244[356],s244[357],s244[358],s244[359],s244[360],s244[361],s244[362],s244[363],s243[365],s242[367],s241[369],s240[347],s239[349],s238[351],s237[353],s236[355],s235[357],s234[359],s234[360],s234[361],s234[362],s234[363],s234[364],s234[365],s234[366],s234[367],s234[368],s234[369],s234[370],s234[371],s234[372],s234[373],s234[374],s234[375],s234[376],s234[377],s234[378],s234[379],s234[380],s234[381],s234[382],s234[383],s234[384],s234[385],s234[386],s234[387],s234[388],s234[389],s234[390],s234[391],s234[392],s234[393],s234[394],s234[395],s234[396],s234[397],s234[398],s234[399],s234[400],s234[401],s234[402],s234[403],s234[404],s234[405],s234[406],s234[407],s234[408],s234[409],s234[410],s234[411],s234[412],s234[413],s234[414],s234[415],s234[416],s234[417],s234[418],s234[419],s234[420],s234[421],s234[422],s234[423],s234[424],s234[425],s234[426],s234[427],s234[428],s234[429],s234[430],s234[431],s234[432],s234[433],s234[434],s234[435],s234[436],s234[437],s234[438],s234[439],s234[440],s234[441],s234[442],s234[443],s234[444],s234[445],s234[446],s234[447],s234[448],s234[449],s234[450],s234[451],s234[452],s234[453],s234[454],s234[455],s233[457],s232[459],s231[461],s230[463],s229[465],s228[467],s227[469],s226[471],s225[473],pp255[235],pp254[237],pp253[239],pp252[241],pp251[243],pp250[245],pp249[247],pp250[247],pp251[247],pp252[247]};
    assign in245_2 = {pp3[9],s242[4],pp14[0],pp13[2],pp14[2],pp15[2],pp15[3],pp15[4],pp16[4],pp17[4],pp19[3],pp21[2],pp23[1],pp25[0],pp26[0],pp27[0],pp28[0],pp29[0],pp30[0],pp31[0],pp32[0],pp33[0],pp34[0],pp35[0],pp36[0],pp37[0],pp38[0],pp39[0],pp40[0],pp41[0],pp42[0],pp43[0],pp44[0],pp45[0],pp46[0],pp47[0],pp48[0],pp49[0],pp50[0],pp51[0],pp52[0],pp53[0],pp54[0],pp55[0],pp56[0],pp57[0],pp58[0],pp59[0],pp60[0],pp61[0],pp62[0],pp63[0],pp64[0],pp65[0],pp66[0],pp67[0],pp68[0],pp69[0],pp70[0],pp71[0],pp72[0],pp73[0],pp74[0],pp75[0],pp76[0],pp77[0],pp78[0],pp79[0],pp80[0],pp81[0],pp82[0],pp83[0],pp84[0],pp85[0],pp86[0],pp87[0],pp88[0],pp89[0],pp90[0],pp91[0],pp92[0],pp93[0],pp94[0],pp95[0],pp96[0],pp97[0],pp98[0],pp99[0],pp99[1],pp99[2],pp99[3],pp99[4],pp99[5],pp99[6],pp99[7],pp99[8],pp99[9],s244[98],s244[99],s240[80],s240[81],s240[82],s240[83],s240[84],s240[85],s240[86],s240[87],s240[88],s240[89],s240[90],s240[91],s240[92],s240[93],s240[94],s240[95],s240[96],s240[97],s240[98],s240[99],s224[68],s224[69],s224[70],s224[71],s224[72],s224[73],s224[74],s1[10],s2[10],s3[10],s4[10],s5[10],s6[10],s7[10],s8[10],s9[10],s9[11],s9[12],s9[13],s9[14],s9[15],s9[16],s9[17],s9[18],s9[19],s9[20],s9[21],s9[22],s9[23],s9[24],s9[25],s9[26],s9[27],s9[28],s9[29],s9[30],s9[31],s9[32],s9[33],s9[34],s9[35],s9[36],s9[37],s9[38],s9[39],s9[40],s9[41],s9[42],s9[43],s9[44],s9[45],s9[46],s9[47],s9[48],s9[49],s9[50],s9[51],s9[52],s9[53],s9[54],s9[55],s9[56],s9[57],s9[58],s9[59],s9[60],s9[61],s9[62],s9[63],s9[64],s9[65],s9[66],s9[67],s9[68],s9[69],s9[70],s9[71],s9[72],s9[73],s9[74],s9[75],s9[76],s9[77],s9[78],s9[79],s9[80],s9[81],s9[82],s9[83],s9[84],s9[85],s9[86],s9[87],s9[88],s9[89],s9[90],s8[92],s7[94],s6[96],s5[98],s104[0],s103[2],s102[4],s101[6],s100[8],s99[10],s99[11],s99[12],s99[13],s99[14],s99[15],s99[16],s99[17],s99[18],s99[19],s99[20],s99[21],s99[22],s99[23],s99[24],s99[25],s99[26],s99[27],s99[28],s99[29],s99[30],s97[33],s95[36],s93[39],s91[42],s90[44],s90[45],s90[46],s90[47],s90[48],s90[49],s90[50],s90[51],s90[52],s90[53],s90[54],s90[55],s90[56],s90[57],s90[58],s90[59],s90[60],s90[61],s90[62],s90[63],s90[64],s90[65],s90[66],s90[67],s90[68],s89[70],s88[72],s87[74],s86[76],s85[78],s84[80],s83[82],s82[84],s81[86],s80[88],s79[90],s78[92],s77[94],s76[96],s75[98],s9[165],s7[168],s5[171],s3[174],s1[177],s78[101],s77[103],s76[105],s75[107],s74[109],s73[111],s72[113],s71[115],s70[117],s69[119],s68[121],s67[123],s66[125],s65[127],s64[129],s63[131],s62[133],s61[135],s60[137],s59[139],s58[141],s57[143],s56[145],s55[147],s54[149],s53[151],s52[153],s51[155],s50[157],s49[159],s48[161],s47[163],s46[165],s45[167],s44[169],s43[171],s42[173],s41[175],s40[177],s39[179],s38[181],s37[183],s36[185],s35[187],s34[189],s33[191],s32[193],s31[195],s30[197],s29[199],s28[201],s27[203],s26[205],s25[207],s24[209],s23[211],s22[213],s21[215],s20[217],s19[219],s18[221],s17[223],s16[225],s15[227],s14[229],s13[231],s12[233],s11[235],s10[237],s244[364],s243[366],s242[368],s241[370],s240[348],s239[350],s238[352],s237[354],s236[356],s235[358],s235[359],s235[360],s235[361],s235[362],s235[363],s235[364],s235[365],s235[366],s235[367],s235[368],s235[369],s235[370],s235[371],s235[372],s235[373],s235[374],s235[375],s235[376],s235[377],s235[378],s235[379],s235[380],s235[381],s235[382],s235[383],s235[384],s235[385],s235[386],s235[387],s235[388],s235[389],s235[390],s235[391],s235[392],s235[393],s235[394],s235[395],s235[396],s235[397],s235[398],s235[399],s235[400],s235[401],s235[402],s235[403],s235[404],s235[405],s235[406],s235[407],s235[408],s235[409],s235[410],s235[411],s235[412],s235[413],s235[414],s235[415],s235[416],s235[417],s235[418],s235[419],s235[420],s235[421],s235[422],s235[423],s235[424],s235[425],s235[426],s235[427],s235[428],s235[429],s235[430],s235[431],s235[432],s235[433],s235[434],s235[435],s235[436],s235[437],s235[438],s235[439],s235[440],s235[441],s235[442],s235[443],s235[444],s235[445],s235[446],s235[447],s235[448],s235[449],s235[450],s235[451],s235[452],s235[453],s235[454],s234[456],s233[458],s232[460],s231[462],s230[464],s229[466],s228[468],s227[470],s226[472],s225[474],pp255[236],pp254[238],pp253[240],pp252[242],pp251[244],pp250[246],pp251[246],pp252[246],pp253[246]};
    CLA_488 KS_245(s245, c245, in245_1, in245_2);
    wire[485:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {s243[3],s241[6],pp14[1],pp15[1],pp16[1],pp16[2],pp16[3],pp17[3],pp18[3],s245[10],s245[11],s245[12],s245[13],s245[14],s245[15],s245[16],s245[17],s245[18],s245[19],s245[20],s245[21],s245[22],s245[23],s245[24],s245[25],s245[26],s245[27],s245[28],s245[29],s245[30],s245[31],s245[32],s245[33],s245[34],s245[35],s245[36],s245[37],s245[38],s245[39],s245[40],s245[41],s245[42],s245[43],s245[44],s245[45],s245[46],s245[47],s245[48],s245[49],s245[50],s245[51],s245[52],s245[53],s245[54],s245[55],s245[56],s245[57],s245[58],s245[59],s245[60],s245[61],s245[62],s245[63],s245[64],s245[65],s245[66],s245[67],s245[68],s245[69],s245[70],s245[71],s245[72],s245[73],s245[74],s245[75],s245[76],s245[77],s245[78],s245[79],s245[80],s245[81],s245[82],s245[83],s245[84],s245[85],s245[86],s245[87],s245[88],s245[89],s245[90],s245[91],s245[92],s245[93],s245[94],s245[95],s245[96],s245[97],s245[98],s245[99],s245[100],s245[101],s245[102],s245[103],s245[104],s245[105],s245[106],s245[107],s245[108],s245[109],s245[110],s245[111],s245[112],s245[113],s245[114],s245[115],s245[116],s245[117],s245[118],s245[119],s245[120],s245[121],s245[122],s245[123],s245[124],s245[125],s245[126],s245[127],s245[128],s245[129],s245[130],s245[131],s245[132],s245[133],s245[134],s245[135],s245[136],s245[137],s245[138],s245[139],s245[140],s245[141],s245[142],s245[143],s245[144],s245[145],s245[146],s245[147],s245[148],s245[149],s245[150],s245[151],s245[152],s245[153],s245[154],s245[155],s245[156],s245[157],s245[158],s245[159],s245[160],s245[161],s245[162],s245[163],s245[164],s245[165],s245[166],s245[167],s245[168],s245[169],s245[170],s245[171],s245[172],s245[173],s245[174],s245[175],s245[176],s245[177],s245[178],s245[179],s245[180],s245[181],s245[182],s245[183],s245[184],s245[185],s245[186],s245[187],s245[188],s245[189],s245[190],s245[191],s245[192],s245[193],s245[194],s245[195],s245[196],s245[197],s245[198],s245[199],s245[200],s245[201],s245[202],s245[203],s245[204],s245[205],s245[206],s245[207],s245[208],s245[209],s245[210],s245[211],s245[212],s245[213],s245[214],s245[215],s245[216],s245[217],s245[218],s245[219],s245[220],s245[221],s245[222],s245[223],s245[224],s245[225],s245[226],s245[227],s245[228],s245[229],s245[230],s245[231],s245[232],s245[233],s245[234],s245[235],s245[236],s245[237],s245[238],s245[239],s245[240],s245[241],s245[242],s245[243],s245[244],s245[245],s245[246],s245[247],s245[248],s245[249],s245[250],s245[251],s245[252],s245[253],s245[254],s245[255],s245[256],s245[257],s245[258],s245[259],s245[260],s245[261],s245[262],s245[263],s245[264],s245[265],s245[266],s245[267],s245[268],s245[269],s245[270],s245[271],s245[272],s245[273],s245[274],s245[275],s245[276],s245[277],s245[278],s245[279],s245[280],s245[281],s245[282],s245[283],s245[284],s245[285],s245[286],s245[287],s245[288],s245[289],s245[290],s245[291],s245[292],s245[293],s245[294],s245[295],s245[296],s245[297],s245[298],s245[299],s245[300],s245[301],s245[302],s245[303],s245[304],s245[305],s245[306],s245[307],s245[308],s245[309],s245[310],s245[311],s245[312],s245[313],s245[314],s245[315],s245[316],s245[317],s245[318],s245[319],s245[320],s245[321],s245[322],s245[323],s245[324],s245[325],s245[326],s245[327],s245[328],s245[329],s245[330],s245[331],s245[332],s245[333],s245[334],s245[335],s245[336],s245[337],s245[338],s245[339],s245[340],s245[341],s245[342],s245[343],s245[344],s245[345],s245[346],s245[347],s245[348],s245[349],s245[350],s245[351],s245[352],s245[353],s245[354],s245[355],s245[356],s245[357],s245[358],s245[359],s245[360],s245[361],s245[362],s245[363],s244[365],s243[367],s242[369],s241[371],s240[349],s239[351],s238[353],s237[355],s236[357],s236[358],s236[359],s236[360],s236[361],s236[362],s236[363],s236[364],s236[365],s236[366],s236[367],s236[368],s236[369],s236[370],s236[371],s236[372],s236[373],s236[374],s236[375],s236[376],s236[377],s236[378],s236[379],s236[380],s236[381],s236[382],s236[383],s236[384],s236[385],s236[386],s236[387],s236[388],s236[389],s236[390],s236[391],s236[392],s236[393],s236[394],s236[395],s236[396],s236[397],s236[398],s236[399],s236[400],s236[401],s236[402],s236[403],s236[404],s236[405],s236[406],s236[407],s236[408],s236[409],s236[410],s236[411],s236[412],s236[413],s236[414],s236[415],s236[416],s236[417],s236[418],s236[419],s236[420],s236[421],s236[422],s236[423],s236[424],s236[425],s236[426],s236[427],s236[428],s236[429],s236[430],s236[431],s236[432],s236[433],s236[434],s236[435],s236[436],s236[437],s236[438],s236[439],s236[440],s236[441],s236[442],s236[443],s236[444],s236[445],s236[446],s236[447],s236[448],s236[449],s236[450],s236[451],s236[452],s236[453],s235[455],s234[457],s233[459],s232[461],s231[463],s230[465],s229[467],s228[469],s227[471],s226[473],s225[475],pp255[237],pp254[239],pp253[241],pp252[243],pp251[245],pp252[245],pp253[245]};
    assign in246_2 = {s244[2],s242[5],pp15[0],pp16[0],pp17[0],pp17[1],pp17[2],pp18[2],pp19[2],pp20[2],pp22[1],pp24[0],s225[9],s226[9],s227[9],s228[9],s229[9],s230[9],s231[9],s193[0],s193[1],s193[2],s193[3],s193[4],s193[5],s193[6],s193[7],s193[8],s193[9],s194[9],s195[9],s196[9],s197[9],s198[9],s199[9],s200[9],s201[9],s202[9],s203[9],s204[9],s205[9],s206[9],s207[9],s208[9],s209[9],s210[9],s211[9],s212[9],s213[9],s214[9],s215[9],s129[0],s129[1],s129[2],s129[3],s129[4],s129[5],s129[6],s129[7],s129[8],s129[9],s130[9],s131[9],s132[9],s133[9],s134[9],s135[9],s136[9],s137[9],s138[9],s139[9],s140[9],s141[9],s142[9],s143[9],s144[9],s145[9],s146[9],s147[9],s148[9],s149[9],s150[9],s151[9],s152[9],s153[9],s154[9],s155[9],s156[9],s157[9],s158[9],s159[9],s160[9],s161[9],s162[9],s163[9],s164[9],s165[9],s166[9],s167[9],s168[9],s169[9],s170[9],s171[9],s172[9],s173[9],s174[9],s175[9],s176[9],s177[9],s178[9],s179[9],s180[9],s181[9],s182[9],s183[9],s184[9],s185[9],s186[9],s187[9],s188[9],s189[9],s190[9],s191[9],s192[9],s10[0],s10[1],s10[2],s10[3],s10[4],s10[5],s10[6],s10[7],s10[8],s10[9],s11[9],s12[9],s13[9],s14[9],s15[9],s16[9],s17[9],s18[9],s19[9],s20[9],s21[9],s22[9],s23[9],s24[9],s25[9],s26[9],s27[9],s28[9],s29[9],s30[9],s31[9],s32[9],s33[9],s34[9],s35[9],s36[9],s37[9],s38[9],s39[9],s40[9],s41[9],s42[9],s43[9],s44[9],s45[9],s46[9],s47[9],s48[9],s49[9],s50[9],s51[9],s52[9],s53[9],s54[9],s55[9],s56[9],s57[9],s58[9],s59[9],s60[9],s61[9],s62[9],s63[9],s64[9],s65[9],s66[9],s67[9],s68[9],s69[9],s70[9],s71[9],s72[9],s73[9],s74[9],s75[9],s76[9],s77[9],s78[9],s79[9],s80[9],s81[9],s82[9],s83[9],s84[9],s85[9],s86[9],s87[9],s88[9],s89[9],s90[9],s9[91],s8[93],s7[95],s6[97],s5[99],s104[1],s103[3],s102[5],s101[7],s100[9],s101[9],s102[9],s103[9],s104[9],s105[9],s106[9],s107[9],s108[9],s109[9],s110[9],s111[9],s112[9],s113[9],s114[9],s115[9],s116[9],s117[9],s118[9],s119[9],s120[9],s98[32],s96[35],s94[38],s92[41],s91[43],s91[44],s91[45],s91[46],s91[47],s91[48],s91[49],s91[50],s91[51],s91[52],s91[53],s91[54],s91[55],s91[56],s91[57],s91[58],s91[59],s91[60],s91[61],s91[62],s91[63],s91[64],s91[65],s91[66],s91[67],s90[69],s89[71],s88[73],s87[75],s86[77],s85[79],s84[81],s83[83],s82[85],s81[87],s80[89],s79[91],s78[93],s77[95],s76[97],s75[99],s8[167],s6[170],s4[173],s2[176],s1[178],s1[179],s1[180],s1[181],s1[182],s1[183],s1[184],s1[185],s1[186],s1[187],s1[188],s1[189],s1[190],s1[191],s1[192],s1[193],s1[194],s1[195],s1[196],s1[197],s1[198],s1[199],s1[200],s1[201],s1[202],s1[203],s1[204],s1[205],s1[206],s1[207],s1[208],s1[209],s1[210],s1[211],s1[212],s1[213],s1[214],s1[215],s1[216],s1[217],s1[218],s1[219],s1[220],s1[221],s1[222],s1[223],s1[224],s1[225],s1[226],s1[227],s1[228],s1[229],s1[230],s1[231],s1[232],s1[233],s1[234],s1[235],s1[236],s1[237],s1[238],s1[239],s1[240],s1[241],s1[242],s1[243],s1[244],s1[245],s1[246],s1[247],s245[364],s244[366],s243[368],s242[370],s241[372],s240[350],s239[352],s238[354],s237[356],s237[357],s237[358],s237[359],s237[360],s237[361],s237[362],s237[363],s237[364],s237[365],s237[366],s237[367],s237[368],s237[369],s237[370],s237[371],s237[372],s237[373],s237[374],s237[375],s237[376],s237[377],s237[378],s237[379],s237[380],s237[381],s237[382],s237[383],s237[384],s237[385],s237[386],s237[387],s237[388],s237[389],s237[390],s237[391],s237[392],s237[393],s237[394],s237[395],s237[396],s237[397],s237[398],s237[399],s237[400],s237[401],s237[402],s237[403],s237[404],s237[405],s237[406],s237[407],s237[408],s237[409],s237[410],s237[411],s237[412],s237[413],s237[414],s237[415],s237[416],s237[417],s237[418],s237[419],s237[420],s237[421],s237[422],s237[423],s237[424],s237[425],s237[426],s237[427],s237[428],s237[429],s237[430],s237[431],s237[432],s237[433],s237[434],s237[435],s237[436],s237[437],s237[438],s237[439],s237[440],s237[441],s237[442],s237[443],s237[444],s237[445],s237[446],s237[447],s237[448],s237[449],s237[450],s237[451],s237[452],s236[454],s235[456],s234[458],s233[460],s232[462],s231[464],s230[466],s229[468],s228[470],s227[472],s226[474],s225[476],pp255[238],pp254[240],pp253[242],pp252[244],pp253[244],pp254[244]};
    CLA_486 KS_246(s246, c246, in246_1, in246_2);
    wire[483:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {s243[4],s241[7],s225[0],s225[1],pp18[0],pp18[1],pp19[1],pp20[1],pp21[1],s246[10],s246[11],s246[12],s246[13],s246[14],s246[15],s246[16],s246[17],s246[18],s246[19],s246[20],s246[21],s246[22],s246[23],s246[24],s246[25],s246[26],s246[27],s246[28],s246[29],s246[30],s246[31],s246[32],s246[33],s246[34],s246[35],s246[36],s246[37],s246[38],s246[39],s246[40],s246[41],s246[42],s246[43],s246[44],s246[45],s246[46],s246[47],s246[48],s246[49],s246[50],s246[51],s246[52],s246[53],s246[54],s246[55],s246[56],s246[57],s246[58],s246[59],s246[60],s246[61],s246[62],s246[63],s246[64],s246[65],s246[66],s246[67],s246[68],s246[69],s246[70],s246[71],s246[72],s246[73],s246[74],s246[75],s246[76],s246[77],s246[78],s246[79],s246[80],s246[81],s246[82],s246[83],s246[84],s246[85],s246[86],s246[87],s246[88],s246[89],s246[90],s246[91],s246[92],s246[93],s246[94],s246[95],s246[96],s246[97],s246[98],s246[99],s246[100],s246[101],s246[102],s246[103],s246[104],s246[105],s246[106],s246[107],s246[108],s246[109],s246[110],s246[111],s246[112],s246[113],s246[114],s246[115],s246[116],s246[117],s246[118],s246[119],s246[120],s246[121],s246[122],s246[123],s246[124],s246[125],s246[126],s246[127],s246[128],s246[129],s246[130],s246[131],s246[132],s246[133],s246[134],s246[135],s246[136],s246[137],s246[138],s246[139],s246[140],s246[141],s246[142],s246[143],s246[144],s246[145],s246[146],s246[147],s246[148],s246[149],s246[150],s246[151],s246[152],s246[153],s246[154],s246[155],s246[156],s246[157],s246[158],s246[159],s246[160],s246[161],s246[162],s246[163],s246[164],s246[165],s246[166],s246[167],s246[168],s246[169],s246[170],s246[171],s246[172],s246[173],s246[174],s246[175],s246[176],s246[177],s246[178],s246[179],s246[180],s246[181],s246[182],s246[183],s246[184],s246[185],s246[186],s246[187],s246[188],s246[189],s246[190],s246[191],s246[192],s246[193],s246[194],s246[195],s246[196],s246[197],s246[198],s246[199],s246[200],s246[201],s246[202],s246[203],s246[204],s246[205],s246[206],s246[207],s246[208],s246[209],s246[210],s246[211],s246[212],s246[213],s246[214],s246[215],s246[216],s246[217],s246[218],s246[219],s246[220],s246[221],s246[222],s246[223],s246[224],s246[225],s246[226],s246[227],s246[228],s246[229],s246[230],s246[231],s246[232],s246[233],s246[234],s246[235],s246[236],s246[237],s246[238],s246[239],s246[240],s246[241],s246[242],s246[243],s246[244],s246[245],s246[246],s246[247],s246[248],s246[249],s246[250],s246[251],s246[252],s246[253],s246[254],s246[255],s246[256],s246[257],s246[258],s246[259],s246[260],s246[261],s246[262],s246[263],s246[264],s246[265],s246[266],s246[267],s246[268],s246[269],s246[270],s246[271],s246[272],s246[273],s246[274],s246[275],s246[276],s246[277],s246[278],s246[279],s246[280],s246[281],s246[282],s246[283],s246[284],s246[285],s246[286],s246[287],s246[288],s246[289],s246[290],s246[291],s246[292],s246[293],s246[294],s246[295],s246[296],s246[297],s246[298],s246[299],s246[300],s246[301],s246[302],s246[303],s246[304],s246[305],s246[306],s246[307],s246[308],s246[309],s246[310],s246[311],s246[312],s246[313],s246[314],s246[315],s246[316],s246[317],s246[318],s246[319],s246[320],s246[321],s246[322],s246[323],s246[324],s246[325],s246[326],s246[327],s246[328],s246[329],s246[330],s246[331],s246[332],s246[333],s246[334],s246[335],s246[336],s246[337],s246[338],s246[339],s246[340],s246[341],s246[342],s246[343],s246[344],s246[345],s246[346],s246[347],s246[348],s246[349],s246[350],s246[351],s246[352],s246[353],s246[354],s246[355],s246[356],s246[357],s246[358],s246[359],s246[360],s246[361],s246[362],s246[363],s245[365],s244[367],s243[369],s242[371],s241[373],s240[351],s239[353],s238[355],s238[356],s238[357],s238[358],s238[359],s238[360],s238[361],s238[362],s238[363],s238[364],s238[365],s238[366],s238[367],s238[368],s238[369],s238[370],s238[371],s238[372],s238[373],s238[374],s238[375],s238[376],s238[377],s238[378],s238[379],s238[380],s238[381],s238[382],s238[383],s238[384],s238[385],s238[386],s238[387],s238[388],s238[389],s238[390],s238[391],s238[392],s238[393],s238[394],s238[395],s238[396],s238[397],s238[398],s238[399],s238[400],s238[401],s238[402],s238[403],s238[404],s238[405],s238[406],s238[407],s238[408],s238[409],s238[410],s238[411],s238[412],s238[413],s238[414],s238[415],s238[416],s238[417],s238[418],s238[419],s238[420],s238[421],s238[422],s238[423],s238[424],s238[425],s238[426],s238[427],s238[428],s238[429],s238[430],s238[431],s238[432],s238[433],s238[434],s238[435],s238[436],s238[437],s238[438],s238[439],s238[440],s238[441],s238[442],s238[443],s238[444],s238[445],s238[446],s238[447],s238[448],s238[449],s238[450],s238[451],s237[453],s236[455],s235[457],s234[459],s233[461],s232[463],s231[465],s230[467],s229[469],s228[471],s227[473],s226[475],s225[477],pp255[239],pp254[241],pp253[243],pp254[243]};
    assign in247_2 = {s244[3],s242[6],s241[8],s226[0],s225[2],pp19[0],pp20[0],pp21[0],pp22[0],pp23[0],s225[8],s226[8],s227[8],s228[8],s229[8],s230[8],s231[8],s232[8],s232[9],s194[0],s194[1],s194[2],s194[3],s194[4],s194[5],s194[6],s194[7],s194[8],s195[8],s196[8],s197[8],s198[8],s199[8],s200[8],s201[8],s202[8],s203[8],s204[8],s205[8],s206[8],s207[8],s208[8],s209[8],s210[8],s211[8],s212[8],s213[8],s214[8],s215[8],s216[8],s216[9],s130[0],s130[1],s130[2],s130[3],s130[4],s130[5],s130[6],s130[7],s130[8],s131[8],s132[8],s133[8],s134[8],s135[8],s136[8],s137[8],s138[8],s139[8],s140[8],s141[8],s142[8],s143[8],s144[8],s145[8],s146[8],s147[8],s148[8],s149[8],s150[8],s151[8],s152[8],s153[8],s154[8],s155[8],s156[8],s157[8],s158[8],s159[8],s160[8],s161[8],s162[8],s163[8],s164[8],s165[8],s166[8],s167[8],s168[8],s169[8],s170[8],s171[8],s172[8],s173[8],s174[8],s175[8],s176[8],s177[8],s178[8],s179[8],s180[8],s181[8],s182[8],s183[8],s184[8],s185[8],s186[8],s187[8],s188[8],s189[8],s190[8],s191[8],s192[8],s1[8],s1[9],s11[0],s11[1],s11[2],s11[3],s11[4],s11[5],s11[6],s11[7],s11[8],s12[8],s13[8],s14[8],s15[8],s16[8],s17[8],s18[8],s19[8],s20[8],s21[8],s22[8],s23[8],s24[8],s25[8],s26[8],s27[8],s28[8],s29[8],s30[8],s31[8],s32[8],s33[8],s34[8],s35[8],s36[8],s37[8],s38[8],s39[8],s40[8],s41[8],s42[8],s43[8],s44[8],s45[8],s46[8],s47[8],s48[8],s49[8],s50[8],s51[8],s52[8],s53[8],s54[8],s55[8],s56[8],s57[8],s58[8],s59[8],s60[8],s61[8],s62[8],s63[8],s64[8],s65[8],s66[8],s67[8],s68[8],s69[8],s70[8],s71[8],s72[8],s73[8],s74[8],s75[8],s76[8],s77[8],s78[8],s79[8],s80[8],s81[8],s82[8],s83[8],s84[8],s85[8],s86[8],s87[8],s88[8],s89[8],s90[8],s91[8],s91[9],s9[92],s8[94],s7[96],s6[98],s105[0],s104[2],s103[4],s102[6],s101[8],s102[8],s103[8],s104[8],s105[8],s106[8],s107[8],s108[8],s109[8],s110[8],s111[8],s112[8],s113[8],s114[8],s115[8],s116[8],s117[8],s118[8],s119[8],s120[8],s121[8],s99[31],s97[34],s95[37],s93[40],s92[42],s92[43],s92[44],s92[45],s92[46],s92[47],s92[48],s92[49],s92[50],s92[51],s92[52],s92[53],s92[54],s92[55],s92[56],s92[57],s92[58],s92[59],s92[60],s92[61],s92[62],s92[63],s92[64],s92[65],s92[66],s91[68],s90[70],s89[72],s88[74],s87[76],s86[78],s85[80],s84[82],s83[84],s82[86],s81[88],s80[90],s79[92],s78[94],s77[96],s76[98],s9[166],s7[169],s5[172],s3[175],s2[177],s2[178],s2[179],s2[180],s2[181],s2[182],s2[183],s2[184],s2[185],s2[186],s2[187],s2[188],s2[189],s2[190],s2[191],s2[192],s2[193],s2[194],s2[195],s2[196],s2[197],s2[198],s2[199],s2[200],s2[201],s2[202],s2[203],s2[204],s2[205],s2[206],s2[207],s2[208],s2[209],s2[210],s2[211],s2[212],s2[213],s2[214],s2[215],s2[216],s2[217],s2[218],s2[219],s2[220],s2[221],s2[222],s2[223],s2[224],s2[225],s2[226],s2[227],s2[228],s2[229],s2[230],s2[231],s2[232],s2[233],s2[234],s2[235],s2[236],s2[237],s2[238],s2[239],s2[240],s2[241],s2[242],s2[243],s2[244],s2[245],s2[246],s1[248],s246[364],s245[366],s244[368],s243[370],s242[372],s241[374],s240[352],s239[354],s239[355],s239[356],s239[357],s239[358],s239[359],s239[360],s239[361],s239[362],s239[363],s239[364],s239[365],s239[366],s239[367],s239[368],s239[369],s239[370],s239[371],s239[372],s239[373],s239[374],s239[375],s239[376],s239[377],s239[378],s239[379],s239[380],s239[381],s239[382],s239[383],s239[384],s239[385],s239[386],s239[387],s239[388],s239[389],s239[390],s239[391],s239[392],s239[393],s239[394],s239[395],s239[396],s239[397],s239[398],s239[399],s239[400],s239[401],s239[402],s239[403],s239[404],s239[405],s239[406],s239[407],s239[408],s239[409],s239[410],s239[411],s239[412],s239[413],s239[414],s239[415],s239[416],s239[417],s239[418],s239[419],s239[420],s239[421],s239[422],s239[423],s239[424],s239[425],s239[426],s239[427],s239[428],s239[429],s239[430],s239[431],s239[432],s239[433],s239[434],s239[435],s239[436],s239[437],s239[438],s239[439],s239[440],s239[441],s239[442],s239[443],s239[444],s239[445],s239[446],s239[447],s239[448],s239[449],s239[450],s238[452],s237[454],s236[456],s235[458],s234[460],s233[462],s232[464],s231[466],s230[468],s229[470],s228[472],s227[474],s226[476],s225[478],pp255[240],pp254[242],pp255[242]};
    CLA_484 KS_247(s247, c247, in247_1, in247_2);
    wire[481:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {s243[5],s242[7],s241[9],s226[1],s225[3],s225[4],s225[5],s225[6],s225[7],s247[10],s247[11],s247[12],s247[13],s247[14],s247[15],s247[16],s247[17],s247[18],s247[19],s247[20],s247[21],s247[22],s247[23],s247[24],s247[25],s247[26],s247[27],s247[28],s247[29],s247[30],s247[31],s247[32],s247[33],s247[34],s247[35],s247[36],s247[37],s247[38],s247[39],s247[40],s247[41],s247[42],s247[43],s247[44],s247[45],s247[46],s247[47],s247[48],s247[49],s247[50],s247[51],s247[52],s247[53],s247[54],s247[55],s247[56],s247[57],s247[58],s247[59],s247[60],s247[61],s247[62],s247[63],s247[64],s247[65],s247[66],s247[67],s247[68],s247[69],s247[70],s247[71],s247[72],s247[73],s247[74],s247[75],s247[76],s247[77],s247[78],s247[79],s247[80],s247[81],s247[82],s247[83],s247[84],s247[85],s247[86],s247[87],s247[88],s247[89],s247[90],s247[91],s247[92],s247[93],s247[94],s247[95],s247[96],s247[97],s247[98],s247[99],s247[100],s247[101],s247[102],s247[103],s247[104],s247[105],s247[106],s247[107],s247[108],s247[109],s247[110],s247[111],s247[112],s247[113],s247[114],s247[115],s247[116],s247[117],s247[118],s247[119],s247[120],s247[121],s247[122],s247[123],s247[124],s247[125],s247[126],s247[127],s247[128],s247[129],s247[130],s247[131],s247[132],s247[133],s247[134],s247[135],s247[136],s247[137],s247[138],s247[139],s247[140],s247[141],s247[142],s247[143],s247[144],s247[145],s247[146],s247[147],s247[148],s247[149],s247[150],s247[151],s247[152],s247[153],s247[154],s247[155],s247[156],s247[157],s247[158],s247[159],s247[160],s247[161],s247[162],s247[163],s247[164],s247[165],s247[166],s247[167],s247[168],s247[169],s247[170],s247[171],s247[172],s247[173],s247[174],s247[175],s247[176],s247[177],s247[178],s247[179],s247[180],s247[181],s247[182],s247[183],s247[184],s247[185],s247[186],s247[187],s247[188],s247[189],s247[190],s247[191],s247[192],s247[193],s247[194],s247[195],s247[196],s247[197],s247[198],s247[199],s247[200],s247[201],s247[202],s247[203],s247[204],s247[205],s247[206],s247[207],s247[208],s247[209],s247[210],s247[211],s247[212],s247[213],s247[214],s247[215],s247[216],s247[217],s247[218],s247[219],s247[220],s247[221],s247[222],s247[223],s247[224],s247[225],s247[226],s247[227],s247[228],s247[229],s247[230],s247[231],s247[232],s247[233],s247[234],s247[235],s247[236],s247[237],s247[238],s247[239],s247[240],s247[241],s247[242],s247[243],s247[244],s247[245],s247[246],s247[247],s247[248],s247[249],s247[250],s247[251],s247[252],s247[253],s247[254],s247[255],s247[256],s247[257],s247[258],s247[259],s247[260],s247[261],s247[262],s247[263],s247[264],s247[265],s247[266],s247[267],s247[268],s247[269],s247[270],s247[271],s247[272],s247[273],s247[274],s247[275],s247[276],s247[277],s247[278],s247[279],s247[280],s247[281],s247[282],s247[283],s247[284],s247[285],s247[286],s247[287],s247[288],s247[289],s247[290],s247[291],s247[292],s247[293],s247[294],s247[295],s247[296],s247[297],s247[298],s247[299],s247[300],s247[301],s247[302],s247[303],s247[304],s247[305],s247[306],s247[307],s247[308],s247[309],s247[310],s247[311],s247[312],s247[313],s247[314],s247[315],s247[316],s247[317],s247[318],s247[319],s247[320],s247[321],s247[322],s247[323],s247[324],s247[325],s247[326],s247[327],s247[328],s247[329],s247[330],s247[331],s247[332],s247[333],s247[334],s247[335],s247[336],s247[337],s247[338],s247[339],s247[340],s247[341],s247[342],s247[343],s247[344],s247[345],s247[346],s247[347],s247[348],s247[349],s247[350],s247[351],s247[352],s247[353],s247[354],s247[355],s247[356],s247[357],s247[358],s247[359],s247[360],s247[361],s247[362],s247[363],s246[365],s245[367],s244[369],s243[371],s242[373],s241[375],s240[353],s240[354],s240[355],s240[356],s240[357],s240[358],s240[359],s240[360],s240[361],s240[362],s240[363],s240[364],s240[365],s240[366],s240[367],s240[368],s240[369],s240[370],s240[371],s240[372],s240[373],s240[374],s240[375],s240[376],s240[377],s240[378],s240[379],s240[380],s240[381],s240[382],s240[383],s240[384],s240[385],s240[386],s240[387],s240[388],s240[389],s240[390],s240[391],s240[392],s240[393],s240[394],s240[395],s240[396],s240[397],s240[398],s240[399],s240[400],s240[401],s240[402],s240[403],s240[404],s240[405],s240[406],s240[407],s240[408],s240[409],s240[410],s240[411],s240[412],s240[413],s240[414],s240[415],s240[416],s240[417],s240[418],s240[419],s240[420],s240[421],s240[422],s240[423],s240[424],s240[425],s240[426],s240[427],s240[428],s240[429],s240[430],s240[431],s240[432],s240[433],s240[434],s240[435],s240[436],s240[437],s240[438],s240[439],s240[440],s240[441],s240[442],s240[443],s240[444],s240[445],s240[446],s240[447],s240[448],s240[449],s239[451],s238[453],s237[455],s236[457],s235[459],s234[461],s233[463],s232[465],s231[467],s230[469],s229[471],s228[473],s227[475],s226[477],s225[479],pp255[241]};
    assign in248_2 = {s244[4],s243[6],s242[8],s227[0],s226[2],s226[3],s226[4],s226[5],s226[6],s226[7],s227[7],s228[7],s229[7],s230[7],s231[7],s232[7],s233[7],s233[8],s233[9],s195[0],s195[1],s195[2],s195[3],s195[4],s195[5],s195[6],s195[7],s196[7],s197[7],s198[7],s199[7],s200[7],s201[7],s202[7],s203[7],s204[7],s205[7],s206[7],s207[7],s208[7],s209[7],s210[7],s211[7],s212[7],s213[7],s214[7],s215[7],s216[7],s217[7],s217[8],s217[9],s131[0],s131[1],s131[2],s131[3],s131[4],s131[5],s131[6],s131[7],s132[7],s133[7],s134[7],s135[7],s136[7],s137[7],s138[7],s139[7],s140[7],s141[7],s142[7],s143[7],s144[7],s145[7],s146[7],s147[7],s148[7],s149[7],s150[7],s151[7],s152[7],s153[7],s154[7],s155[7],s156[7],s157[7],s158[7],s159[7],s160[7],s161[7],s162[7],s163[7],s164[7],s165[7],s166[7],s167[7],s168[7],s169[7],s170[7],s171[7],s172[7],s173[7],s174[7],s175[7],s176[7],s177[7],s178[7],s179[7],s180[7],s181[7],s182[7],s183[7],s184[7],s185[7],s186[7],s187[7],s188[7],s189[7],s190[7],s191[7],s192[7],s1[7],s2[7],s2[8],s2[9],s12[0],s12[1],s12[2],s12[3],s12[4],s12[5],s12[6],s12[7],s13[7],s14[7],s15[7],s16[7],s17[7],s18[7],s19[7],s20[7],s21[7],s22[7],s23[7],s24[7],s25[7],s26[7],s27[7],s28[7],s29[7],s30[7],s31[7],s32[7],s33[7],s34[7],s35[7],s36[7],s37[7],s38[7],s39[7],s40[7],s41[7],s42[7],s43[7],s44[7],s45[7],s46[7],s47[7],s48[7],s49[7],s50[7],s51[7],s52[7],s53[7],s54[7],s55[7],s56[7],s57[7],s58[7],s59[7],s60[7],s61[7],s62[7],s63[7],s64[7],s65[7],s66[7],s67[7],s68[7],s69[7],s70[7],s71[7],s72[7],s73[7],s74[7],s75[7],s76[7],s77[7],s78[7],s79[7],s80[7],s81[7],s82[7],s83[7],s84[7],s85[7],s86[7],s87[7],s88[7],s89[7],s90[7],s91[7],s92[7],s92[8],s92[9],s9[93],s8[95],s7[97],s6[99],s105[1],s104[3],s103[5],s102[7],s103[7],s104[7],s105[7],s106[7],s107[7],s108[7],s109[7],s110[7],s111[7],s112[7],s113[7],s114[7],s115[7],s116[7],s117[7],s118[7],s119[7],s120[7],s121[7],s122[7],s121[9],s98[33],s96[36],s94[39],s93[41],s93[42],s93[43],s93[44],s93[45],s93[46],s93[47],s93[48],s93[49],s93[50],s93[51],s93[52],s93[53],s93[54],s93[55],s93[56],s93[57],s93[58],s93[59],s93[60],s93[61],s93[62],s93[63],s93[64],s93[65],s92[67],s91[69],s90[71],s89[73],s88[75],s87[77],s86[79],s85[81],s84[83],s83[85],s82[87],s81[89],s80[91],s79[93],s78[95],s77[97],s76[99],s8[168],s6[171],s4[174],s3[176],s3[177],s3[178],s3[179],s3[180],s3[181],s3[182],s3[183],s3[184],s3[185],s3[186],s3[187],s3[188],s3[189],s3[190],s3[191],s3[192],s3[193],s3[194],s3[195],s3[196],s3[197],s3[198],s3[199],s3[200],s3[201],s3[202],s3[203],s3[204],s3[205],s3[206],s3[207],s3[208],s3[209],s3[210],s3[211],s3[212],s3[213],s3[214],s3[215],s3[216],s3[217],s3[218],s3[219],s3[220],s3[221],s3[222],s3[223],s3[224],s3[225],s3[226],s3[227],s3[228],s3[229],s3[230],s3[231],s3[232],s3[233],s3[234],s3[235],s3[236],s3[237],s3[238],s3[239],s3[240],s3[241],s3[242],s3[243],s3[244],s3[245],s2[247],s1[249],s247[364],s246[366],s245[368],s244[370],s243[372],s242[374],s241[376],s241[377],s241[378],s241[379],s241[380],s241[381],s241[382],s241[383],s241[384],s241[385],s241[386],s241[387],s241[388],s241[389],s241[390],s241[391],s241[392],s241[393],s241[394],s241[395],s241[396],s241[397],s241[398],s241[399],s241[400],s241[401],s241[402],s241[403],s241[404],s241[405],s241[406],s241[407],s241[408],s241[409],s241[410],s241[411],s241[412],s241[413],s241[414],s241[415],s241[416],s241[417],s241[418],s241[419],s241[420],s241[421],s241[422],s241[423],s241[424],s241[425],s241[426],s241[427],s241[428],s241[429],s241[430],s241[431],s241[432],s241[433],s241[434],s241[435],s241[436],s241[437],s241[438],s241[439],s241[440],s241[441],s241[442],s241[443],s241[444],s241[445],s241[446],s241[447],s241[448],s241[449],s241[450],s241[451],s241[452],s241[453],s241[454],s241[455],s241[456],s241[457],s241[458],s241[459],s241[460],s241[461],s241[462],s241[463],s241[464],s241[465],s241[466],s241[467],s241[468],s241[469],s241[470],s241[471],s241[472],s241[473],s241[474],s241[475],s241[476],s241[477],s241[478],s241[479],s241[480],s241[481],s241[482],s241[483],s241[484],s241[485],s241[486],s241[487],s241[488]};
    CLA_482 KS_248(s248, c248, in248_1, in248_2);

    /*Stage 6*/
    wire[503:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {pp0[4],pp0[5],pp0[6],pp0[7],s241[0],s241[1],s242[1],s243[1],s244[1],s245[1],s245[2],s245[3],s244[5],s243[7],s242[9],s227[1],s227[2],s227[3],s227[4],s227[5],s227[6],s248[10],s248[11],s248[12],s248[13],s248[14],s248[15],s248[16],s248[17],s248[18],s248[19],s248[20],s248[21],s248[22],s248[23],s248[24],s248[25],s248[26],s248[27],s248[28],s248[29],s248[30],s248[31],s248[32],s248[33],s248[34],s248[35],s248[36],s248[37],s248[38],s248[39],s248[40],s248[41],s248[42],s248[43],s248[44],s248[45],s248[46],s248[47],s248[48],s248[49],s248[50],s248[51],s248[52],s248[53],s248[54],s248[55],s248[56],s248[57],s248[58],s248[59],s248[60],s248[61],s248[62],s248[63],s248[64],s248[65],s248[66],s248[67],s248[68],s248[69],s248[70],s248[71],s248[72],s248[73],s248[74],s248[75],s248[76],s248[77],s248[78],s248[79],s248[80],s248[81],s248[82],s248[83],s248[84],s248[85],s248[86],s248[87],s248[88],s248[89],s248[90],s248[91],s248[92],s248[93],s248[94],s248[95],s248[96],s248[97],s248[98],s248[99],s248[100],s248[101],s248[102],s248[103],s248[104],s248[105],s248[106],s248[107],s248[108],s248[109],s248[110],s248[111],s248[112],s248[113],s248[114],s248[115],s248[116],s248[117],s248[118],s248[119],s248[120],s248[121],s248[122],s248[123],s248[124],s248[125],s248[126],s248[127],s248[128],s248[129],s248[130],s248[131],s248[132],s248[133],s248[134],s248[135],s248[136],s248[137],s248[138],s248[139],s248[140],s248[141],s248[142],s248[143],s248[144],s248[145],s248[146],s248[147],s248[148],s248[149],s248[150],s248[151],s248[152],s248[153],s248[154],s248[155],s248[156],s248[157],s248[158],s248[159],s248[160],s248[161],s248[162],s248[163],s248[164],s248[165],s248[166],s248[167],s248[168],s248[169],s248[170],s248[171],s248[172],s248[173],s248[174],s248[175],s248[176],s248[177],s248[178],s248[179],s248[180],s248[181],s248[182],s248[183],s248[184],s248[185],s248[186],s248[187],s248[188],s248[189],s248[190],s248[191],s248[192],s248[193],s248[194],s248[195],s248[196],s248[197],s248[198],s248[199],s248[200],s248[201],s248[202],s248[203],s248[204],s248[205],s248[206],s248[207],s248[208],s248[209],s248[210],s248[211],s248[212],s248[213],s248[214],s248[215],s248[216],s248[217],s248[218],s248[219],s248[220],s248[221],s248[222],s248[223],s248[224],s248[225],s248[226],s248[227],s248[228],s248[229],s248[230],s248[231],s248[232],s248[233],s248[234],s248[235],s248[236],s248[237],s248[238],s248[239],s248[240],s248[241],s248[242],s248[243],s248[244],s248[245],s248[246],s248[247],s248[248],s248[249],s248[250],s248[251],s248[252],s248[253],s248[254],s248[255],s248[256],s248[257],s248[258],s248[259],s248[260],s248[261],s248[262],s248[263],s248[264],s248[265],s248[266],s248[267],s248[268],s248[269],s248[270],s248[271],s248[272],s248[273],s248[274],s248[275],s248[276],s248[277],s248[278],s248[279],s248[280],s248[281],s248[282],s248[283],s248[284],s248[285],s248[286],s248[287],s248[288],s248[289],s248[290],s248[291],s248[292],s248[293],s248[294],s248[295],s248[296],s248[297],s248[298],s248[299],s248[300],s248[301],s248[302],s248[303],s248[304],s248[305],s248[306],s248[307],s248[308],s248[309],s248[310],s248[311],s248[312],s248[313],s248[314],s248[315],s248[316],s248[317],s248[318],s248[319],s248[320],s248[321],s248[322],s248[323],s248[324],s248[325],s248[326],s248[327],s248[328],s248[329],s248[330],s248[331],s248[332],s248[333],s248[334],s248[335],s248[336],s248[337],s248[338],s248[339],s248[340],s248[341],s248[342],s248[343],s248[344],s248[345],s248[346],s248[347],s248[348],s248[349],s248[350],s248[351],s248[352],s248[353],s248[354],s248[355],s248[356],s248[357],s248[358],s248[359],s248[360],s248[361],s248[362],s248[363],s247[365],s246[367],s245[369],s244[371],s243[373],s242[375],s242[376],s242[377],s242[378],s242[379],s242[380],s242[381],s242[382],s242[383],s242[384],s242[385],s242[386],s242[387],s242[388],s242[389],s242[390],s242[391],s242[392],s242[393],s242[394],s242[395],s242[396],s242[397],s242[398],s242[399],s242[400],s242[401],s242[402],s242[403],s242[404],s242[405],s242[406],s242[407],s242[408],s242[409],s242[410],s242[411],s242[412],s242[413],s242[414],s242[415],s242[416],s242[417],s242[418],s242[419],s242[420],s242[421],s242[422],s242[423],s242[424],s242[425],s242[426],s242[427],s242[428],s242[429],s242[430],s242[431],s242[432],s242[433],s242[434],s242[435],s242[436],s242[437],s242[438],s242[439],s242[440],s242[441],s242[442],s242[443],s242[444],s242[445],s242[446],s242[447],s242[448],s242[449],s242[450],s242[451],s242[452],s242[453],s242[454],s242[455],s242[456],s242[457],s242[458],s242[459],s242[460],s242[461],s242[462],s242[463],s242[464],s242[465],s242[466],s242[467],s242[468],s242[469],s242[470],s242[471],s242[472],s242[473],s242[474],s242[475],s242[476],s242[477],s242[478],s242[479],s242[480],s242[481],s242[482],s242[483],s242[484],s242[485],s242[486],s242[487],s241[489],pp255[243],pp254[245],pp253[247],pp252[249],pp251[251],pp250[253],pp249[255],pp250[255],pp251[255],pp252[255]};
    assign in249_2 = {pp1[3],pp1[4],pp1[5],pp1[6],pp2[6],s242[0],s243[0],s244[0],s245[0],s246[0],s246[1],s246[2],s245[4],s244[6],s243[8],s228[0],s228[1],s228[2],s228[3],s228[4],s228[5],s228[6],s229[6],s230[6],s231[6],s232[6],s233[6],s234[6],s234[7],s234[8],s234[9],s196[0],s196[1],s196[2],s196[3],s196[4],s196[5],s196[6],s197[6],s198[6],s199[6],s200[6],s201[6],s202[6],s203[6],s204[6],s205[6],s206[6],s207[6],s208[6],s209[6],s210[6],s211[6],s212[6],s213[6],s214[6],s215[6],s216[6],s217[6],s218[6],s218[7],s218[8],s218[9],s132[0],s132[1],s132[2],s132[3],s132[4],s132[5],s132[6],s133[6],s134[6],s135[6],s136[6],s137[6],s138[6],s139[6],s140[6],s141[6],s142[6],s143[6],s144[6],s145[6],s146[6],s147[6],s148[6],s149[6],s150[6],s151[6],s152[6],s153[6],s154[6],s155[6],s156[6],s157[6],s158[6],s159[6],s160[6],s161[6],s162[6],s163[6],s164[6],s165[6],s166[6],s167[6],s168[6],s169[6],s170[6],s171[6],s172[6],s173[6],s174[6],s175[6],s176[6],s177[6],s178[6],s179[6],s180[6],s181[6],s182[6],s183[6],s184[6],s185[6],s186[6],s187[6],s188[6],s189[6],s190[6],s191[6],s192[6],s1[6],s2[6],s3[6],s3[7],s3[8],s3[9],s13[0],s13[1],s13[2],s13[3],s13[4],s13[5],s13[6],s14[6],s15[6],s16[6],s17[6],s18[6],s19[6],s20[6],s21[6],s22[6],s23[6],s24[6],s25[6],s26[6],s27[6],s28[6],s29[6],s30[6],s31[6],s32[6],s33[6],s34[6],s35[6],s36[6],s37[6],s38[6],s39[6],s40[6],s41[6],s42[6],s43[6],s44[6],s45[6],s46[6],s47[6],s48[6],s49[6],s50[6],s51[6],s52[6],s53[6],s54[6],s55[6],s56[6],s57[6],s58[6],s59[6],s60[6],s61[6],s62[6],s63[6],s64[6],s65[6],s66[6],s67[6],s68[6],s69[6],s70[6],s71[6],s72[6],s73[6],s74[6],s75[6],s76[6],s77[6],s78[6],s79[6],s80[6],s81[6],s82[6],s83[6],s84[6],s85[6],s86[6],s87[6],s88[6],s89[6],s90[6],s91[6],s92[6],s93[6],s93[7],s93[8],s93[9],s9[94],s8[96],s7[98],s106[0],s105[2],s104[4],s103[6],s104[6],s105[6],s106[6],s107[6],s108[6],s109[6],s110[6],s111[6],s112[6],s113[6],s114[6],s115[6],s116[6],s117[6],s118[6],s119[6],s120[6],s121[6],s122[6],s123[6],s122[8],s99[32],s97[35],s95[38],s94[40],s94[41],s94[42],s94[43],s94[44],s94[45],s94[46],s94[47],s94[48],s94[49],s94[50],s94[51],s94[52],s94[53],s94[54],s94[55],s94[56],s94[57],s94[58],s94[59],s94[60],s94[61],s94[62],s94[63],s94[64],s93[66],s92[68],s91[70],s90[72],s89[74],s88[76],s87[78],s86[80],s85[82],s84[84],s83[86],s82[88],s81[90],s80[92],s79[94],s78[96],s77[98],s9[167],s7[170],s5[173],s4[175],s4[176],s4[177],s4[178],s4[179],s4[180],s4[181],s4[182],s4[183],s4[184],s4[185],s4[186],s4[187],s4[188],s4[189],s4[190],s4[191],s4[192],s4[193],s4[194],s4[195],s4[196],s4[197],s4[198],s4[199],s4[200],s4[201],s4[202],s4[203],s4[204],s4[205],s4[206],s4[207],s4[208],s4[209],s4[210],s4[211],s4[212],s4[213],s4[214],s4[215],s4[216],s4[217],s4[218],s4[219],s4[220],s4[221],s4[222],s4[223],s4[224],s4[225],s4[226],s4[227],s4[228],s4[229],s4[230],s4[231],s4[232],s4[233],s4[234],s4[235],s4[236],s4[237],s4[238],s4[239],s4[240],s4[241],s4[242],s4[243],s4[244],s3[246],s2[248],s1[250],s248[364],s247[366],s246[368],s245[370],s244[372],s243[374],s243[375],s243[376],s243[377],s243[378],s243[379],s243[380],s243[381],s243[382],s243[383],s243[384],s243[385],s243[386],s243[387],s243[388],s243[389],s243[390],s243[391],s243[392],s243[393],s243[394],s243[395],s243[396],s243[397],s243[398],s243[399],s243[400],s243[401],s243[402],s243[403],s243[404],s243[405],s243[406],s243[407],s243[408],s243[409],s243[410],s243[411],s243[412],s243[413],s243[414],s243[415],s243[416],s243[417],s243[418],s243[419],s243[420],s243[421],s243[422],s243[423],s243[424],s243[425],s243[426],s243[427],s243[428],s243[429],s243[430],s243[431],s243[432],s243[433],s243[434],s243[435],s243[436],s243[437],s243[438],s243[439],s243[440],s243[441],s243[442],s243[443],s243[444],s243[445],s243[446],s243[447],s243[448],s243[449],s243[450],s243[451],s243[452],s243[453],s243[454],s243[455],s243[456],s243[457],s243[458],s243[459],s243[460],s243[461],s243[462],s243[463],s243[464],s243[465],s243[466],s243[467],s243[468],s243[469],s243[470],s243[471],s243[472],s243[473],s243[474],s243[475],s243[476],s243[477],s243[478],s243[479],s243[480],s243[481],s243[482],s243[483],s243[484],s243[485],s243[486],s242[488],s241[490],pp255[244],pp254[246],pp253[248],pp252[250],pp251[252],pp250[254],pp251[254],pp252[254],pp253[254]};
    CLA_504 KS_249(s249, c249, in249_1, in249_2);
    wire[501:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {pp2[3],s249[2],s249[3],s249[4],s249[5],s249[6],s249[7],s249[8],s249[9],s249[10],s249[11],s249[12],s249[13],s249[14],s249[15],s249[16],s249[17],s249[18],s249[19],s249[20],s249[21],s249[22],s249[23],s249[24],s249[25],s249[26],s249[27],s249[28],s249[29],s249[30],s249[31],s249[32],s249[33],s249[34],s249[35],s249[36],s249[37],s249[38],s249[39],s249[40],s249[41],s249[42],s249[43],s249[44],s249[45],s249[46],s249[47],s249[48],s249[49],s249[50],s249[51],s249[52],s249[53],s249[54],s249[55],s249[56],s249[57],s249[58],s249[59],s249[60],s249[61],s249[62],s249[63],s249[64],s249[65],s249[66],s249[67],s249[68],s249[69],s249[70],s249[71],s249[72],s249[73],s249[74],s249[75],s249[76],s249[77],s249[78],s249[79],s249[80],s249[81],s249[82],s249[83],s249[84],s249[85],s249[86],s249[87],s249[88],s249[89],s249[90],s249[91],s249[92],s249[93],s249[94],s249[95],s249[96],s249[97],s249[98],s249[99],s249[100],s249[101],s249[102],s249[103],s249[104],s249[105],s249[106],s249[107],s249[108],s249[109],s249[110],s249[111],s249[112],s249[113],s249[114],s249[115],s249[116],s249[117],s249[118],s249[119],s249[120],s249[121],s249[122],s249[123],s249[124],s249[125],s249[126],s249[127],s249[128],s249[129],s249[130],s249[131],s249[132],s249[133],s249[134],s249[135],s249[136],s249[137],s249[138],s249[139],s249[140],s249[141],s249[142],s249[143],s249[144],s249[145],s249[146],s249[147],s249[148],s249[149],s249[150],s249[151],s249[152],s249[153],s249[154],s249[155],s249[156],s249[157],s249[158],s249[159],s249[160],s249[161],s249[162],s249[163],s249[164],s249[165],s249[166],s249[167],s249[168],s249[169],s249[170],s249[171],s249[172],s249[173],s249[174],s249[175],s249[176],s249[177],s249[178],s249[179],s249[180],s249[181],s249[182],s249[183],s249[184],s249[185],s249[186],s249[187],s249[188],s249[189],s249[190],s249[191],s249[192],s249[193],s249[194],s249[195],s249[196],s249[197],s249[198],s249[199],s249[200],s249[201],s249[202],s249[203],s249[204],s249[205],s249[206],s249[207],s249[208],s249[209],s249[210],s249[211],s249[212],s249[213],s249[214],s249[215],s249[216],s249[217],s249[218],s249[219],s249[220],s249[221],s249[222],s249[223],s249[224],s249[225],s249[226],s249[227],s249[228],s249[229],s249[230],s249[231],s249[232],s249[233],s249[234],s249[235],s249[236],s249[237],s249[238],s249[239],s249[240],s249[241],s249[242],s249[243],s249[244],s249[245],s249[246],s249[247],s249[248],s249[249],s249[250],s249[251],s249[252],s249[253],s249[254],s249[255],s249[256],s249[257],s249[258],s249[259],s249[260],s249[261],s249[262],s249[263],s249[264],s249[265],s249[266],s249[267],s249[268],s249[269],s249[270],s249[271],s249[272],s249[273],s249[274],s249[275],s249[276],s249[277],s249[278],s249[279],s249[280],s249[281],s249[282],s249[283],s249[284],s249[285],s249[286],s249[287],s249[288],s249[289],s249[290],s249[291],s249[292],s249[293],s249[294],s249[295],s249[296],s249[297],s249[298],s249[299],s249[300],s249[301],s249[302],s249[303],s249[304],s249[305],s249[306],s249[307],s249[308],s249[309],s249[310],s249[311],s249[312],s249[313],s249[314],s249[315],s249[316],s249[317],s249[318],s249[319],s249[320],s249[321],s249[322],s249[323],s249[324],s249[325],s249[326],s249[327],s249[328],s249[329],s249[330],s249[331],s249[332],s249[333],s249[334],s249[335],s249[336],s249[337],s249[338],s249[339],s249[340],s249[341],s249[342],s249[343],s249[344],s249[345],s249[346],s249[347],s249[348],s249[349],s249[350],s249[351],s249[352],s249[353],s249[354],s249[355],s249[356],s249[357],s249[358],s249[359],s249[360],s249[361],s249[362],s249[363],s249[364],s249[365],s249[366],s249[367],s249[368],s249[369],s249[370],s249[371],s249[372],s249[373],s249[374],s249[375],s248[365],s247[367],s246[369],s245[371],s244[373],s244[374],s244[375],s244[376],s244[377],s244[378],s244[379],s244[380],s244[381],s244[382],s244[383],s244[384],s244[385],s244[386],s244[387],s244[388],s244[389],s244[390],s244[391],s244[392],s244[393],s244[394],s244[395],s244[396],s244[397],s244[398],s244[399],s244[400],s244[401],s244[402],s244[403],s244[404],s244[405],s244[406],s244[407],s244[408],s244[409],s244[410],s244[411],s244[412],s244[413],s244[414],s244[415],s244[416],s244[417],s244[418],s244[419],s244[420],s244[421],s244[422],s244[423],s244[424],s244[425],s244[426],s244[427],s244[428],s244[429],s244[430],s244[431],s244[432],s244[433],s244[434],s244[435],s244[436],s244[437],s244[438],s244[439],s244[440],s244[441],s244[442],s244[443],s244[444],s244[445],s244[446],s244[447],s244[448],s244[449],s244[450],s244[451],s244[452],s244[453],s244[454],s244[455],s244[456],s244[457],s244[458],s244[459],s244[460],s244[461],s244[462],s244[463],s244[464],s244[465],s244[466],s244[467],s244[468],s244[469],s244[470],s244[471],s244[472],s244[473],s244[474],s244[475],s244[476],s244[477],s244[478],s244[479],s244[480],s244[481],s244[482],s244[483],s244[484],s244[485],s243[487],s242[489],s241[491],pp255[245],pp254[247],pp253[249],pp252[251],pp251[253],pp252[253],pp253[253]};
    assign in250_2 = {pp3[2],pp2[4],pp2[5],pp3[5],pp4[5],pp4[6],pp4[7],pp4[8],pp4[9],s247[0],s247[1],s246[3],s245[5],s244[7],s243[9],s229[0],s229[1],s229[2],s229[3],s229[4],s229[5],s230[5],s231[5],s232[5],s233[5],s234[5],s235[5],s235[6],s235[7],s235[8],s235[9],s197[0],s197[1],s197[2],s197[3],s197[4],s197[5],s198[5],s199[5],s200[5],s201[5],s202[5],s203[5],s204[5],s205[5],s206[5],s207[5],s208[5],s209[5],s210[5],s211[5],s212[5],s213[5],s214[5],s215[5],s216[5],s217[5],s218[5],s219[5],s219[6],s219[7],s219[8],s219[9],s133[0],s133[1],s133[2],s133[3],s133[4],s133[5],s134[5],s135[5],s136[5],s137[5],s138[5],s139[5],s140[5],s141[5],s142[5],s143[5],s144[5],s145[5],s146[5],s147[5],s148[5],s149[5],s150[5],s151[5],s152[5],s153[5],s154[5],s155[5],s156[5],s157[5],s158[5],s159[5],s160[5],s161[5],s162[5],s163[5],s164[5],s165[5],s166[5],s167[5],s168[5],s169[5],s170[5],s171[5],s172[5],s173[5],s174[5],s175[5],s176[5],s177[5],s178[5],s179[5],s180[5],s181[5],s182[5],s183[5],s184[5],s185[5],s186[5],s187[5],s188[5],s189[5],s190[5],s191[5],s192[5],s1[5],s2[5],s3[5],s4[5],s4[6],s4[7],s4[8],s4[9],s14[0],s14[1],s14[2],s14[3],s14[4],s14[5],s15[5],s16[5],s17[5],s18[5],s19[5],s20[5],s21[5],s22[5],s23[5],s24[5],s25[5],s26[5],s27[5],s28[5],s29[5],s30[5],s31[5],s32[5],s33[5],s34[5],s35[5],s36[5],s37[5],s38[5],s39[5],s40[5],s41[5],s42[5],s43[5],s44[5],s45[5],s46[5],s47[5],s48[5],s49[5],s50[5],s51[5],s52[5],s53[5],s54[5],s55[5],s56[5],s57[5],s58[5],s59[5],s60[5],s61[5],s62[5],s63[5],s64[5],s65[5],s66[5],s67[5],s68[5],s69[5],s70[5],s71[5],s72[5],s73[5],s74[5],s75[5],s76[5],s77[5],s78[5],s79[5],s80[5],s81[5],s82[5],s83[5],s84[5],s85[5],s86[5],s87[5],s88[5],s89[5],s90[5],s91[5],s92[5],s93[5],s94[5],s94[6],s94[7],s94[8],s94[9],s9[95],s8[97],s7[99],s106[1],s105[3],s104[5],s105[5],s106[5],s107[5],s108[5],s109[5],s110[5],s111[5],s112[5],s113[5],s114[5],s115[5],s116[5],s117[5],s118[5],s119[5],s120[5],s121[5],s122[5],s123[5],s124[5],s123[7],s122[9],s98[34],s96[37],s95[39],s95[40],s95[41],s95[42],s95[43],s95[44],s95[45],s95[46],s95[47],s95[48],s95[49],s95[50],s95[51],s95[52],s95[53],s95[54],s95[55],s95[56],s95[57],s95[58],s95[59],s95[60],s95[61],s95[62],s95[63],s94[65],s93[67],s92[69],s91[71],s90[73],s89[75],s88[77],s87[79],s86[81],s85[83],s84[85],s83[87],s82[89],s81[91],s80[93],s79[95],s78[97],s77[99],s8[169],s6[172],s5[174],s5[175],s5[176],s5[177],s5[178],s5[179],s5[180],s5[181],s5[182],s5[183],s5[184],s5[185],s5[186],s5[187],s5[188],s5[189],s5[190],s5[191],s5[192],s5[193],s5[194],s5[195],s5[196],s5[197],s5[198],s5[199],s5[200],s5[201],s5[202],s5[203],s5[204],s5[205],s5[206],s5[207],s5[208],s5[209],s5[210],s5[211],s5[212],s5[213],s5[214],s5[215],s5[216],s5[217],s5[218],s5[219],s5[220],s5[221],s5[222],s5[223],s5[224],s5[225],s5[226],s5[227],s5[228],s5[229],s5[230],s5[231],s5[232],s5[233],s5[234],s5[235],s5[236],s5[237],s5[238],s5[239],s5[240],s5[241],s5[242],s5[243],s4[245],s3[247],s2[249],s1[251],s249[376],s248[366],s247[368],s246[370],s245[372],s245[373],s245[374],s245[375],s245[376],s245[377],s245[378],s245[379],s245[380],s245[381],s245[382],s245[383],s245[384],s245[385],s245[386],s245[387],s245[388],s245[389],s245[390],s245[391],s245[392],s245[393],s245[394],s245[395],s245[396],s245[397],s245[398],s245[399],s245[400],s245[401],s245[402],s245[403],s245[404],s245[405],s245[406],s245[407],s245[408],s245[409],s245[410],s245[411],s245[412],s245[413],s245[414],s245[415],s245[416],s245[417],s245[418],s245[419],s245[420],s245[421],s245[422],s245[423],s245[424],s245[425],s245[426],s245[427],s245[428],s245[429],s245[430],s245[431],s245[432],s245[433],s245[434],s245[435],s245[436],s245[437],s245[438],s245[439],s245[440],s245[441],s245[442],s245[443],s245[444],s245[445],s245[446],s245[447],s245[448],s245[449],s245[450],s245[451],s245[452],s245[453],s245[454],s245[455],s245[456],s245[457],s245[458],s245[459],s245[460],s245[461],s245[462],s245[463],s245[464],s245[465],s245[466],s245[467],s245[468],s245[469],s245[470],s245[471],s245[472],s245[473],s245[474],s245[475],s245[476],s245[477],s245[478],s245[479],s245[480],s245[481],s245[482],s245[483],s245[484],s244[486],s243[488],s242[490],s241[492],pp255[246],pp254[248],pp253[250],pp252[252],pp253[252],pp254[252]};
    CLA_502 KS_250(s250, c250, in250_1, in250_2);
    wire[499:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp3[3],s250[2],s250[3],s250[4],s250[5],s250[6],s250[7],s250[8],s250[9],s250[10],s250[11],s250[12],s250[13],s250[14],s250[15],s250[16],s250[17],s250[18],s250[19],s250[20],s250[21],s250[22],s250[23],s250[24],s250[25],s250[26],s250[27],s250[28],s250[29],s250[30],s250[31],s250[32],s250[33],s250[34],s250[35],s250[36],s250[37],s250[38],s250[39],s250[40],s250[41],s250[42],s250[43],s250[44],s250[45],s250[46],s250[47],s250[48],s250[49],s250[50],s250[51],s250[52],s250[53],s250[54],s250[55],s250[56],s250[57],s250[58],s250[59],s250[60],s250[61],s250[62],s250[63],s250[64],s250[65],s250[66],s250[67],s250[68],s250[69],s250[70],s250[71],s250[72],s250[73],s250[74],s250[75],s250[76],s250[77],s250[78],s250[79],s250[80],s250[81],s250[82],s250[83],s250[84],s250[85],s250[86],s250[87],s250[88],s250[89],s250[90],s250[91],s250[92],s250[93],s250[94],s250[95],s250[96],s250[97],s250[98],s250[99],s250[100],s250[101],s250[102],s250[103],s250[104],s250[105],s250[106],s250[107],s250[108],s250[109],s250[110],s250[111],s250[112],s250[113],s250[114],s250[115],s250[116],s250[117],s250[118],s250[119],s250[120],s250[121],s250[122],s250[123],s250[124],s250[125],s250[126],s250[127],s250[128],s250[129],s250[130],s250[131],s250[132],s250[133],s250[134],s250[135],s250[136],s250[137],s250[138],s250[139],s250[140],s250[141],s250[142],s250[143],s250[144],s250[145],s250[146],s250[147],s250[148],s250[149],s250[150],s250[151],s250[152],s250[153],s250[154],s250[155],s250[156],s250[157],s250[158],s250[159],s250[160],s250[161],s250[162],s250[163],s250[164],s250[165],s250[166],s250[167],s250[168],s250[169],s250[170],s250[171],s250[172],s250[173],s250[174],s250[175],s250[176],s250[177],s250[178],s250[179],s250[180],s250[181],s250[182],s250[183],s250[184],s250[185],s250[186],s250[187],s250[188],s250[189],s250[190],s250[191],s250[192],s250[193],s250[194],s250[195],s250[196],s250[197],s250[198],s250[199],s250[200],s250[201],s250[202],s250[203],s250[204],s250[205],s250[206],s250[207],s250[208],s250[209],s250[210],s250[211],s250[212],s250[213],s250[214],s250[215],s250[216],s250[217],s250[218],s250[219],s250[220],s250[221],s250[222],s250[223],s250[224],s250[225],s250[226],s250[227],s250[228],s250[229],s250[230],s250[231],s250[232],s250[233],s250[234],s250[235],s250[236],s250[237],s250[238],s250[239],s250[240],s250[241],s250[242],s250[243],s250[244],s250[245],s250[246],s250[247],s250[248],s250[249],s250[250],s250[251],s250[252],s250[253],s250[254],s250[255],s250[256],s250[257],s250[258],s250[259],s250[260],s250[261],s250[262],s250[263],s250[264],s250[265],s250[266],s250[267],s250[268],s250[269],s250[270],s250[271],s250[272],s250[273],s250[274],s250[275],s250[276],s250[277],s250[278],s250[279],s250[280],s250[281],s250[282],s250[283],s250[284],s250[285],s250[286],s250[287],s250[288],s250[289],s250[290],s250[291],s250[292],s250[293],s250[294],s250[295],s250[296],s250[297],s250[298],s250[299],s250[300],s250[301],s250[302],s250[303],s250[304],s250[305],s250[306],s250[307],s250[308],s250[309],s250[310],s250[311],s250[312],s250[313],s250[314],s250[315],s250[316],s250[317],s250[318],s250[319],s250[320],s250[321],s250[322],s250[323],s250[324],s250[325],s250[326],s250[327],s250[328],s250[329],s250[330],s250[331],s250[332],s250[333],s250[334],s250[335],s250[336],s250[337],s250[338],s250[339],s250[340],s250[341],s250[342],s250[343],s250[344],s250[345],s250[346],s250[347],s250[348],s250[349],s250[350],s250[351],s250[352],s250[353],s250[354],s250[355],s250[356],s250[357],s250[358],s250[359],s250[360],s250[361],s250[362],s250[363],s250[364],s250[365],s250[366],s250[367],s250[368],s250[369],s250[370],s250[371],s250[372],s250[373],s250[374],s250[375],s249[377],s248[367],s247[369],s246[371],s246[372],s246[373],s246[374],s246[375],s246[376],s246[377],s246[378],s246[379],s246[380],s246[381],s246[382],s246[383],s246[384],s246[385],s246[386],s246[387],s246[388],s246[389],s246[390],s246[391],s246[392],s246[393],s246[394],s246[395],s246[396],s246[397],s246[398],s246[399],s246[400],s246[401],s246[402],s246[403],s246[404],s246[405],s246[406],s246[407],s246[408],s246[409],s246[410],s246[411],s246[412],s246[413],s246[414],s246[415],s246[416],s246[417],s246[418],s246[419],s246[420],s246[421],s246[422],s246[423],s246[424],s246[425],s246[426],s246[427],s246[428],s246[429],s246[430],s246[431],s246[432],s246[433],s246[434],s246[435],s246[436],s246[437],s246[438],s246[439],s246[440],s246[441],s246[442],s246[443],s246[444],s246[445],s246[446],s246[447],s246[448],s246[449],s246[450],s246[451],s246[452],s246[453],s246[454],s246[455],s246[456],s246[457],s246[458],s246[459],s246[460],s246[461],s246[462],s246[463],s246[464],s246[465],s246[466],s246[467],s246[468],s246[469],s246[470],s246[471],s246[472],s246[473],s246[474],s246[475],s246[476],s246[477],s246[478],s246[479],s246[480],s246[481],s246[482],s246[483],s245[485],s244[487],s243[489],s242[491],s241[493],pp255[247],pp254[249],pp253[251],pp254[251]};
    assign in251_2 = {pp4[2],pp3[4],pp4[4],pp5[4],pp5[5],pp5[6],pp5[7],pp5[8],pp5[9],s248[0],s247[2],s246[4],s245[6],s244[8],s244[9],s230[0],s230[1],s230[2],s230[3],s230[4],s231[4],s232[4],s233[4],s234[4],s235[4],s236[4],s236[5],s236[6],s236[7],s236[8],s236[9],s198[0],s198[1],s198[2],s198[3],s198[4],s199[4],s200[4],s201[4],s202[4],s203[4],s204[4],s205[4],s206[4],s207[4],s208[4],s209[4],s210[4],s211[4],s212[4],s213[4],s214[4],s215[4],s216[4],s217[4],s218[4],s219[4],s220[4],s220[5],s220[6],s220[7],s220[8],s220[9],s134[0],s134[1],s134[2],s134[3],s134[4],s135[4],s136[4],s137[4],s138[4],s139[4],s140[4],s141[4],s142[4],s143[4],s144[4],s145[4],s146[4],s147[4],s148[4],s149[4],s150[4],s151[4],s152[4],s153[4],s154[4],s155[4],s156[4],s157[4],s158[4],s159[4],s160[4],s161[4],s162[4],s163[4],s164[4],s165[4],s166[4],s167[4],s168[4],s169[4],s170[4],s171[4],s172[4],s173[4],s174[4],s175[4],s176[4],s177[4],s178[4],s179[4],s180[4],s181[4],s182[4],s183[4],s184[4],s185[4],s186[4],s187[4],s188[4],s189[4],s190[4],s191[4],s192[4],s1[4],s2[4],s3[4],s4[4],s5[4],s5[5],s5[6],s5[7],s5[8],s5[9],s15[0],s15[1],s15[2],s15[3],s15[4],s16[4],s17[4],s18[4],s19[4],s20[4],s21[4],s22[4],s23[4],s24[4],s25[4],s26[4],s27[4],s28[4],s29[4],s30[4],s31[4],s32[4],s33[4],s34[4],s35[4],s36[4],s37[4],s38[4],s39[4],s40[4],s41[4],s42[4],s43[4],s44[4],s45[4],s46[4],s47[4],s48[4],s49[4],s50[4],s51[4],s52[4],s53[4],s54[4],s55[4],s56[4],s57[4],s58[4],s59[4],s60[4],s61[4],s62[4],s63[4],s64[4],s65[4],s66[4],s67[4],s68[4],s69[4],s70[4],s71[4],s72[4],s73[4],s74[4],s75[4],s76[4],s77[4],s78[4],s79[4],s80[4],s81[4],s82[4],s83[4],s84[4],s85[4],s86[4],s87[4],s88[4],s89[4],s90[4],s91[4],s92[4],s93[4],s94[4],s95[4],s95[5],s95[6],s95[7],s95[8],s95[9],s9[96],s8[98],s107[0],s106[2],s105[4],s106[4],s107[4],s108[4],s109[4],s110[4],s111[4],s112[4],s113[4],s114[4],s115[4],s116[4],s117[4],s118[4],s119[4],s120[4],s121[4],s122[4],s123[4],s124[4],s125[4],s124[6],s123[8],s99[33],s97[36],s96[38],s96[39],s96[40],s96[41],s96[42],s96[43],s96[44],s96[45],s96[46],s96[47],s96[48],s96[49],s96[50],s96[51],s96[52],s96[53],s96[54],s96[55],s96[56],s96[57],s96[58],s96[59],s96[60],s96[61],s96[62],s95[64],s94[66],s93[68],s92[70],s91[72],s90[74],s89[76],s88[78],s87[80],s86[82],s85[84],s84[86],s83[88],s82[90],s81[92],s80[94],s79[96],s78[98],s9[168],s7[171],s6[173],s6[174],s6[175],s6[176],s6[177],s6[178],s6[179],s6[180],s6[181],s6[182],s6[183],s6[184],s6[185],s6[186],s6[187],s6[188],s6[189],s6[190],s6[191],s6[192],s6[193],s6[194],s6[195],s6[196],s6[197],s6[198],s6[199],s6[200],s6[201],s6[202],s6[203],s6[204],s6[205],s6[206],s6[207],s6[208],s6[209],s6[210],s6[211],s6[212],s6[213],s6[214],s6[215],s6[216],s6[217],s6[218],s6[219],s6[220],s6[221],s6[222],s6[223],s6[224],s6[225],s6[226],s6[227],s6[228],s6[229],s6[230],s6[231],s6[232],s6[233],s6[234],s6[235],s6[236],s6[237],s6[238],s6[239],s6[240],s6[241],s6[242],s5[244],s4[246],s3[248],s2[250],s1[252],s250[376],s249[378],s248[368],s247[370],s247[371],s247[372],s247[373],s247[374],s247[375],s247[376],s247[377],s247[378],s247[379],s247[380],s247[381],s247[382],s247[383],s247[384],s247[385],s247[386],s247[387],s247[388],s247[389],s247[390],s247[391],s247[392],s247[393],s247[394],s247[395],s247[396],s247[397],s247[398],s247[399],s247[400],s247[401],s247[402],s247[403],s247[404],s247[405],s247[406],s247[407],s247[408],s247[409],s247[410],s247[411],s247[412],s247[413],s247[414],s247[415],s247[416],s247[417],s247[418],s247[419],s247[420],s247[421],s247[422],s247[423],s247[424],s247[425],s247[426],s247[427],s247[428],s247[429],s247[430],s247[431],s247[432],s247[433],s247[434],s247[435],s247[436],s247[437],s247[438],s247[439],s247[440],s247[441],s247[442],s247[443],s247[444],s247[445],s247[446],s247[447],s247[448],s247[449],s247[450],s247[451],s247[452],s247[453],s247[454],s247[455],s247[456],s247[457],s247[458],s247[459],s247[460],s247[461],s247[462],s247[463],s247[464],s247[465],s247[466],s247[467],s247[468],s247[469],s247[470],s247[471],s247[472],s247[473],s247[474],s247[475],s247[476],s247[477],s247[478],s247[479],s247[480],s247[481],s247[482],s246[484],s245[486],s244[488],s243[490],s242[492],s241[494],pp255[248],pp254[250],pp255[250]};
    CLA_500 KS_251(s251, c251, in251_1, in251_2);
    wire[497:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp4[3],s251[2],s251[3],s251[4],s251[5],s251[6],s251[7],s251[8],s251[9],s251[10],s251[11],s251[12],s251[13],s251[14],s251[15],s251[16],s251[17],s251[18],s251[19],s251[20],s251[21],s251[22],s251[23],s251[24],s251[25],s251[26],s251[27],s251[28],s251[29],s251[30],s251[31],s251[32],s251[33],s251[34],s251[35],s251[36],s251[37],s251[38],s251[39],s251[40],s251[41],s251[42],s251[43],s251[44],s251[45],s251[46],s251[47],s251[48],s251[49],s251[50],s251[51],s251[52],s251[53],s251[54],s251[55],s251[56],s251[57],s251[58],s251[59],s251[60],s251[61],s251[62],s251[63],s251[64],s251[65],s251[66],s251[67],s251[68],s251[69],s251[70],s251[71],s251[72],s251[73],s251[74],s251[75],s251[76],s251[77],s251[78],s251[79],s251[80],s251[81],s251[82],s251[83],s251[84],s251[85],s251[86],s251[87],s251[88],s251[89],s251[90],s251[91],s251[92],s251[93],s251[94],s251[95],s251[96],s251[97],s251[98],s251[99],s251[100],s251[101],s251[102],s251[103],s251[104],s251[105],s251[106],s251[107],s251[108],s251[109],s251[110],s251[111],s251[112],s251[113],s251[114],s251[115],s251[116],s251[117],s251[118],s251[119],s251[120],s251[121],s251[122],s251[123],s251[124],s251[125],s251[126],s251[127],s251[128],s251[129],s251[130],s251[131],s251[132],s251[133],s251[134],s251[135],s251[136],s251[137],s251[138],s251[139],s251[140],s251[141],s251[142],s251[143],s251[144],s251[145],s251[146],s251[147],s251[148],s251[149],s251[150],s251[151],s251[152],s251[153],s251[154],s251[155],s251[156],s251[157],s251[158],s251[159],s251[160],s251[161],s251[162],s251[163],s251[164],s251[165],s251[166],s251[167],s251[168],s251[169],s251[170],s251[171],s251[172],s251[173],s251[174],s251[175],s251[176],s251[177],s251[178],s251[179],s251[180],s251[181],s251[182],s251[183],s251[184],s251[185],s251[186],s251[187],s251[188],s251[189],s251[190],s251[191],s251[192],s251[193],s251[194],s251[195],s251[196],s251[197],s251[198],s251[199],s251[200],s251[201],s251[202],s251[203],s251[204],s251[205],s251[206],s251[207],s251[208],s251[209],s251[210],s251[211],s251[212],s251[213],s251[214],s251[215],s251[216],s251[217],s251[218],s251[219],s251[220],s251[221],s251[222],s251[223],s251[224],s251[225],s251[226],s251[227],s251[228],s251[229],s251[230],s251[231],s251[232],s251[233],s251[234],s251[235],s251[236],s251[237],s251[238],s251[239],s251[240],s251[241],s251[242],s251[243],s251[244],s251[245],s251[246],s251[247],s251[248],s251[249],s251[250],s251[251],s251[252],s251[253],s251[254],s251[255],s251[256],s251[257],s251[258],s251[259],s251[260],s251[261],s251[262],s251[263],s251[264],s251[265],s251[266],s251[267],s251[268],s251[269],s251[270],s251[271],s251[272],s251[273],s251[274],s251[275],s251[276],s251[277],s251[278],s251[279],s251[280],s251[281],s251[282],s251[283],s251[284],s251[285],s251[286],s251[287],s251[288],s251[289],s251[290],s251[291],s251[292],s251[293],s251[294],s251[295],s251[296],s251[297],s251[298],s251[299],s251[300],s251[301],s251[302],s251[303],s251[304],s251[305],s251[306],s251[307],s251[308],s251[309],s251[310],s251[311],s251[312],s251[313],s251[314],s251[315],s251[316],s251[317],s251[318],s251[319],s251[320],s251[321],s251[322],s251[323],s251[324],s251[325],s251[326],s251[327],s251[328],s251[329],s251[330],s251[331],s251[332],s251[333],s251[334],s251[335],s251[336],s251[337],s251[338],s251[339],s251[340],s251[341],s251[342],s251[343],s251[344],s251[345],s251[346],s251[347],s251[348],s251[349],s251[350],s251[351],s251[352],s251[353],s251[354],s251[355],s251[356],s251[357],s251[358],s251[359],s251[360],s251[361],s251[362],s251[363],s251[364],s251[365],s251[366],s251[367],s251[368],s251[369],s251[370],s251[371],s251[372],s251[373],s251[374],s251[375],s250[377],s249[379],s248[369],s248[370],s248[371],s248[372],s248[373],s248[374],s248[375],s248[376],s248[377],s248[378],s248[379],s248[380],s248[381],s248[382],s248[383],s248[384],s248[385],s248[386],s248[387],s248[388],s248[389],s248[390],s248[391],s248[392],s248[393],s248[394],s248[395],s248[396],s248[397],s248[398],s248[399],s248[400],s248[401],s248[402],s248[403],s248[404],s248[405],s248[406],s248[407],s248[408],s248[409],s248[410],s248[411],s248[412],s248[413],s248[414],s248[415],s248[416],s248[417],s248[418],s248[419],s248[420],s248[421],s248[422],s248[423],s248[424],s248[425],s248[426],s248[427],s248[428],s248[429],s248[430],s248[431],s248[432],s248[433],s248[434],s248[435],s248[436],s248[437],s248[438],s248[439],s248[440],s248[441],s248[442],s248[443],s248[444],s248[445],s248[446],s248[447],s248[448],s248[449],s248[450],s248[451],s248[452],s248[453],s248[454],s248[455],s248[456],s248[457],s248[458],s248[459],s248[460],s248[461],s248[462],s248[463],s248[464],s248[465],s248[466],s248[467],s248[468],s248[469],s248[470],s248[471],s248[472],s248[473],s248[474],s248[475],s248[476],s248[477],s248[478],s248[479],s248[480],s248[481],s247[483],s246[485],s245[487],s244[489],s243[491],s242[493],s241[495],pp255[249]};
    assign in252_2 = {pp5[2],pp5[3],pp6[3],pp6[4],pp6[5],pp6[6],pp6[7],pp6[8],pp6[9],s248[1],s247[3],s246[5],s245[7],s245[8],s245[9],s231[0],s231[1],s231[2],s231[3],s232[3],s233[3],s234[3],s235[3],s236[3],s237[3],s237[4],s237[5],s237[6],s237[7],s237[8],s237[9],s199[0],s199[1],s199[2],s199[3],s200[3],s201[3],s202[3],s203[3],s204[3],s205[3],s206[3],s207[3],s208[3],s209[3],s210[3],s211[3],s212[3],s213[3],s214[3],s215[3],s216[3],s217[3],s218[3],s219[3],s220[3],s221[3],s221[4],s221[5],s221[6],s221[7],s221[8],s221[9],s135[0],s135[1],s135[2],s135[3],s136[3],s137[3],s138[3],s139[3],s140[3],s141[3],s142[3],s143[3],s144[3],s145[3],s146[3],s147[3],s148[3],s149[3],s150[3],s151[3],s152[3],s153[3],s154[3],s155[3],s156[3],s157[3],s158[3],s159[3],s160[3],s161[3],s162[3],s163[3],s164[3],s165[3],s166[3],s167[3],s168[3],s169[3],s170[3],s171[3],s172[3],s173[3],s174[3],s175[3],s176[3],s177[3],s178[3],s179[3],s180[3],s181[3],s182[3],s183[3],s184[3],s185[3],s186[3],s187[3],s188[3],s189[3],s190[3],s191[3],s192[3],s1[3],s2[3],s3[3],s4[3],s5[3],s6[3],s6[4],s6[5],s6[6],s6[7],s6[8],s6[9],s16[0],s16[1],s16[2],s16[3],s17[3],s18[3],s19[3],s20[3],s21[3],s22[3],s23[3],s24[3],s25[3],s26[3],s27[3],s28[3],s29[3],s30[3],s31[3],s32[3],s33[3],s34[3],s35[3],s36[3],s37[3],s38[3],s39[3],s40[3],s41[3],s42[3],s43[3],s44[3],s45[3],s46[3],s47[3],s48[3],s49[3],s50[3],s51[3],s52[3],s53[3],s54[3],s55[3],s56[3],s57[3],s58[3],s59[3],s60[3],s61[3],s62[3],s63[3],s64[3],s65[3],s66[3],s67[3],s68[3],s69[3],s70[3],s71[3],s72[3],s73[3],s74[3],s75[3],s76[3],s77[3],s78[3],s79[3],s80[3],s81[3],s82[3],s83[3],s84[3],s85[3],s86[3],s87[3],s88[3],s89[3],s90[3],s91[3],s92[3],s93[3],s94[3],s95[3],s96[3],s96[4],s96[5],s96[6],s96[7],s96[8],s96[9],s9[97],s8[99],s107[1],s106[3],s107[3],s108[3],s109[3],s110[3],s111[3],s112[3],s113[3],s114[3],s115[3],s116[3],s117[3],s118[3],s119[3],s120[3],s121[3],s122[3],s123[3],s124[3],s125[3],s126[3],s125[5],s124[7],s123[9],s98[35],s97[37],s97[38],s97[39],s97[40],s97[41],s97[42],s97[43],s97[44],s97[45],s97[46],s97[47],s97[48],s97[49],s97[50],s97[51],s97[52],s97[53],s97[54],s97[55],s97[56],s97[57],s97[58],s97[59],s97[60],s97[61],s96[63],s95[65],s94[67],s93[69],s92[71],s91[73],s90[75],s89[77],s88[79],s87[81],s86[83],s85[85],s84[87],s83[89],s82[91],s81[93],s80[95],s79[97],s78[99],s8[170],s7[172],s7[173],s7[174],s7[175],s7[176],s7[177],s7[178],s7[179],s7[180],s7[181],s7[182],s7[183],s7[184],s7[185],s7[186],s7[187],s7[188],s7[189],s7[190],s7[191],s7[192],s7[193],s7[194],s7[195],s7[196],s7[197],s7[198],s7[199],s7[200],s7[201],s7[202],s7[203],s7[204],s7[205],s7[206],s7[207],s7[208],s7[209],s7[210],s7[211],s7[212],s7[213],s7[214],s7[215],s7[216],s7[217],s7[218],s7[219],s7[220],s7[221],s7[222],s7[223],s7[224],s7[225],s7[226],s7[227],s7[228],s7[229],s7[230],s7[231],s7[232],s7[233],s7[234],s7[235],s7[236],s7[237],s7[238],s7[239],s7[240],s7[241],s6[243],s5[245],s4[247],s3[249],s2[251],s1[253],s251[376],s250[378],s249[380],s249[381],s249[382],s249[383],s249[384],s249[385],s249[386],s249[387],s249[388],s249[389],s249[390],s249[391],s249[392],s249[393],s249[394],s249[395],s249[396],s249[397],s249[398],s249[399],s249[400],s249[401],s249[402],s249[403],s249[404],s249[405],s249[406],s249[407],s249[408],s249[409],s249[410],s249[411],s249[412],s249[413],s249[414],s249[415],s249[416],s249[417],s249[418],s249[419],s249[420],s249[421],s249[422],s249[423],s249[424],s249[425],s249[426],s249[427],s249[428],s249[429],s249[430],s249[431],s249[432],s249[433],s249[434],s249[435],s249[436],s249[437],s249[438],s249[439],s249[440],s249[441],s249[442],s249[443],s249[444],s249[445],s249[446],s249[447],s249[448],s249[449],s249[450],s249[451],s249[452],s249[453],s249[454],s249[455],s249[456],s249[457],s249[458],s249[459],s249[460],s249[461],s249[462],s249[463],s249[464],s249[465],s249[466],s249[467],s249[468],s249[469],s249[470],s249[471],s249[472],s249[473],s249[474],s249[475],s249[476],s249[477],s249[478],s249[479],s249[480],s249[481],s249[482],s249[483],s249[484],s249[485],s249[486],s249[487],s249[488],s249[489],s249[490],s249[491],s249[492],s249[493],s249[494],s249[495],s249[496],s249[497],s249[498],s249[499],s249[500]};
    CLA_498 KS_252(s252, c252, in252_1, in252_2);

    /*Stage 7*/
    wire[507:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp0[2],pp0[3],s249[0],s249[1],s250[1],s251[1],s252[1],s252[2],s252[3],s252[4],s252[5],s252[6],s252[7],s252[8],s252[9],s252[10],s252[11],s252[12],s252[13],s252[14],s252[15],s252[16],s252[17],s252[18],s252[19],s252[20],s252[21],s252[22],s252[23],s252[24],s252[25],s252[26],s252[27],s252[28],s252[29],s252[30],s252[31],s252[32],s252[33],s252[34],s252[35],s252[36],s252[37],s252[38],s252[39],s252[40],s252[41],s252[42],s252[43],s252[44],s252[45],s252[46],s252[47],s252[48],s252[49],s252[50],s252[51],s252[52],s252[53],s252[54],s252[55],s252[56],s252[57],s252[58],s252[59],s252[60],s252[61],s252[62],s252[63],s252[64],s252[65],s252[66],s252[67],s252[68],s252[69],s252[70],s252[71],s252[72],s252[73],s252[74],s252[75],s252[76],s252[77],s252[78],s252[79],s252[80],s252[81],s252[82],s252[83],s252[84],s252[85],s252[86],s252[87],s252[88],s252[89],s252[90],s252[91],s252[92],s252[93],s252[94],s252[95],s252[96],s252[97],s252[98],s252[99],s252[100],s252[101],s252[102],s252[103],s252[104],s252[105],s252[106],s252[107],s252[108],s252[109],s252[110],s252[111],s252[112],s252[113],s252[114],s252[115],s252[116],s252[117],s252[118],s252[119],s252[120],s252[121],s252[122],s252[123],s252[124],s252[125],s252[126],s252[127],s252[128],s252[129],s252[130],s252[131],s252[132],s252[133],s252[134],s252[135],s252[136],s252[137],s252[138],s252[139],s252[140],s252[141],s252[142],s252[143],s252[144],s252[145],s252[146],s252[147],s252[148],s252[149],s252[150],s252[151],s252[152],s252[153],s252[154],s252[155],s252[156],s252[157],s252[158],s252[159],s252[160],s252[161],s252[162],s252[163],s252[164],s252[165],s252[166],s252[167],s252[168],s252[169],s252[170],s252[171],s252[172],s252[173],s252[174],s252[175],s252[176],s252[177],s252[178],s252[179],s252[180],s252[181],s252[182],s252[183],s252[184],s252[185],s252[186],s252[187],s252[188],s252[189],s252[190],s252[191],s252[192],s252[193],s252[194],s252[195],s252[196],s252[197],s252[198],s252[199],s252[200],s252[201],s252[202],s252[203],s252[204],s252[205],s252[206],s252[207],s252[208],s252[209],s252[210],s252[211],s252[212],s252[213],s252[214],s252[215],s252[216],s252[217],s252[218],s252[219],s252[220],s252[221],s252[222],s252[223],s252[224],s252[225],s252[226],s252[227],s252[228],s252[229],s252[230],s252[231],s252[232],s252[233],s252[234],s252[235],s252[236],s252[237],s252[238],s252[239],s252[240],s252[241],s252[242],s252[243],s252[244],s252[245],s252[246],s252[247],s252[248],s252[249],s252[250],s252[251],s252[252],s252[253],s252[254],s252[255],s252[256],s252[257],s252[258],s252[259],s252[260],s252[261],s252[262],s252[263],s252[264],s252[265],s252[266],s252[267],s252[268],s252[269],s252[270],s252[271],s252[272],s252[273],s252[274],s252[275],s252[276],s252[277],s252[278],s252[279],s252[280],s252[281],s252[282],s252[283],s252[284],s252[285],s252[286],s252[287],s252[288],s252[289],s252[290],s252[291],s252[292],s252[293],s252[294],s252[295],s252[296],s252[297],s252[298],s252[299],s252[300],s252[301],s252[302],s252[303],s252[304],s252[305],s252[306],s252[307],s252[308],s252[309],s252[310],s252[311],s252[312],s252[313],s252[314],s252[315],s252[316],s252[317],s252[318],s252[319],s252[320],s252[321],s252[322],s252[323],s252[324],s252[325],s252[326],s252[327],s252[328],s252[329],s252[330],s252[331],s252[332],s252[333],s252[334],s252[335],s252[336],s252[337],s252[338],s252[339],s252[340],s252[341],s252[342],s252[343],s252[344],s252[345],s252[346],s252[347],s252[348],s252[349],s252[350],s252[351],s252[352],s252[353],s252[354],s252[355],s252[356],s252[357],s252[358],s252[359],s252[360],s252[361],s252[362],s252[363],s252[364],s252[365],s252[366],s252[367],s252[368],s252[369],s252[370],s252[371],s252[372],s252[373],s252[374],s252[375],s251[377],s250[379],s250[380],s250[381],s250[382],s250[383],s250[384],s250[385],s250[386],s250[387],s250[388],s250[389],s250[390],s250[391],s250[392],s250[393],s250[394],s250[395],s250[396],s250[397],s250[398],s250[399],s250[400],s250[401],s250[402],s250[403],s250[404],s250[405],s250[406],s250[407],s250[408],s250[409],s250[410],s250[411],s250[412],s250[413],s250[414],s250[415],s250[416],s250[417],s250[418],s250[419],s250[420],s250[421],s250[422],s250[423],s250[424],s250[425],s250[426],s250[427],s250[428],s250[429],s250[430],s250[431],s250[432],s250[433],s250[434],s250[435],s250[436],s250[437],s250[438],s250[439],s250[440],s250[441],s250[442],s250[443],s250[444],s250[445],s250[446],s250[447],s250[448],s250[449],s250[450],s250[451],s250[452],s250[453],s250[454],s250[455],s250[456],s250[457],s250[458],s250[459],s250[460],s250[461],s250[462],s250[463],s250[464],s250[465],s250[466],s250[467],s250[468],s250[469],s250[470],s250[471],s250[472],s250[473],s250[474],s250[475],s250[476],s250[477],s250[478],s250[479],s250[480],s250[481],s250[482],s250[483],s250[484],s250[485],s250[486],s250[487],s250[488],s250[489],s250[490],s250[491],s250[492],s250[493],s250[494],s250[495],s250[496],s250[497],s250[498],s250[499],s249[501],pp255[251],pp254[253],pp253[255],pp254[255]};
    assign in253_2 = {pp1[1],pp1[2],pp2[2],s250[0],s251[0],s252[0],pp6[2],pp7[2],pp7[3],pp7[4],pp7[5],pp7[6],pp7[7],pp7[8],pp7[9],s248[2],s247[4],s246[6],s246[7],s246[8],s246[9],s232[0],s232[1],s232[2],s233[2],s234[2],s235[2],s236[2],s237[2],s238[2],s238[3],s238[4],s238[5],s238[6],s238[7],s238[8],s238[9],s200[0],s200[1],s200[2],s201[2],s202[2],s203[2],s204[2],s205[2],s206[2],s207[2],s208[2],s209[2],s210[2],s211[2],s212[2],s213[2],s214[2],s215[2],s216[2],s217[2],s218[2],s219[2],s220[2],s221[2],s222[2],s222[3],s222[4],s222[5],s222[6],s222[7],s222[8],s222[9],s136[0],s136[1],s136[2],s137[2],s138[2],s139[2],s140[2],s141[2],s142[2],s143[2],s144[2],s145[2],s146[2],s147[2],s148[2],s149[2],s150[2],s151[2],s152[2],s153[2],s154[2],s155[2],s156[2],s157[2],s158[2],s159[2],s160[2],s161[2],s162[2],s163[2],s164[2],s165[2],s166[2],s167[2],s168[2],s169[2],s170[2],s171[2],s172[2],s173[2],s174[2],s175[2],s176[2],s177[2],s178[2],s179[2],s180[2],s181[2],s182[2],s183[2],s184[2],s185[2],s186[2],s187[2],s188[2],s189[2],s190[2],s191[2],s192[2],s1[2],s2[2],s3[2],s4[2],s5[2],s6[2],s7[2],s7[3],s7[4],s7[5],s7[6],s7[7],s7[8],s7[9],s17[0],s17[1],s17[2],s18[2],s19[2],s20[2],s21[2],s22[2],s23[2],s24[2],s25[2],s26[2],s27[2],s28[2],s29[2],s30[2],s31[2],s32[2],s33[2],s34[2],s35[2],s36[2],s37[2],s38[2],s39[2],s40[2],s41[2],s42[2],s43[2],s44[2],s45[2],s46[2],s47[2],s48[2],s49[2],s50[2],s51[2],s52[2],s53[2],s54[2],s55[2],s56[2],s57[2],s58[2],s59[2],s60[2],s61[2],s62[2],s63[2],s64[2],s65[2],s66[2],s67[2],s68[2],s69[2],s70[2],s71[2],s72[2],s73[2],s74[2],s75[2],s76[2],s77[2],s78[2],s79[2],s80[2],s81[2],s82[2],s83[2],s84[2],s85[2],s86[2],s87[2],s88[2],s89[2],s90[2],s91[2],s92[2],s93[2],s94[2],s95[2],s96[2],s97[2],s97[3],s97[4],s97[5],s97[6],s97[7],s97[8],s97[9],s9[98],s108[0],s107[2],s108[2],s109[2],s110[2],s111[2],s112[2],s113[2],s114[2],s115[2],s116[2],s117[2],s118[2],s119[2],s120[2],s121[2],s122[2],s123[2],s124[2],s125[2],s126[2],s127[2],s126[4],s125[6],s124[8],s99[34],s98[36],s98[37],s98[38],s98[39],s98[40],s98[41],s98[42],s98[43],s98[44],s98[45],s98[46],s98[47],s98[48],s98[49],s98[50],s98[51],s98[52],s98[53],s98[54],s98[55],s98[56],s98[57],s98[58],s98[59],s98[60],s97[62],s96[64],s95[66],s94[68],s93[70],s92[72],s91[74],s90[76],s89[78],s88[80],s87[82],s86[84],s85[86],s84[88],s83[90],s82[92],s81[94],s80[96],s79[98],s9[169],s8[171],s8[172],s8[173],s8[174],s8[175],s8[176],s8[177],s8[178],s8[179],s8[180],s8[181],s8[182],s8[183],s8[184],s8[185],s8[186],s8[187],s8[188],s8[189],s8[190],s8[191],s8[192],s8[193],s8[194],s8[195],s8[196],s8[197],s8[198],s8[199],s8[200],s8[201],s8[202],s8[203],s8[204],s8[205],s8[206],s8[207],s8[208],s8[209],s8[210],s8[211],s8[212],s8[213],s8[214],s8[215],s8[216],s8[217],s8[218],s8[219],s8[220],s8[221],s8[222],s8[223],s8[224],s8[225],s8[226],s8[227],s8[228],s8[229],s8[230],s8[231],s8[232],s8[233],s8[234],s8[235],s8[236],s8[237],s8[238],s8[239],s8[240],s7[242],s6[244],s5[246],s4[248],s3[250],s2[252],s1[254],s252[376],s251[378],s251[379],s251[380],s251[381],s251[382],s251[383],s251[384],s251[385],s251[386],s251[387],s251[388],s251[389],s251[390],s251[391],s251[392],s251[393],s251[394],s251[395],s251[396],s251[397],s251[398],s251[399],s251[400],s251[401],s251[402],s251[403],s251[404],s251[405],s251[406],s251[407],s251[408],s251[409],s251[410],s251[411],s251[412],s251[413],s251[414],s251[415],s251[416],s251[417],s251[418],s251[419],s251[420],s251[421],s251[422],s251[423],s251[424],s251[425],s251[426],s251[427],s251[428],s251[429],s251[430],s251[431],s251[432],s251[433],s251[434],s251[435],s251[436],s251[437],s251[438],s251[439],s251[440],s251[441],s251[442],s251[443],s251[444],s251[445],s251[446],s251[447],s251[448],s251[449],s251[450],s251[451],s251[452],s251[453],s251[454],s251[455],s251[456],s251[457],s251[458],s251[459],s251[460],s251[461],s251[462],s251[463],s251[464],s251[465],s251[466],s251[467],s251[468],s251[469],s251[470],s251[471],s251[472],s251[473],s251[474],s251[475],s251[476],s251[477],s251[478],s251[479],s251[480],s251[481],s251[482],s251[483],s251[484],s251[485],s251[486],s251[487],s251[488],s251[489],s251[490],s251[491],s251[492],s251[493],s251[494],s251[495],s251[496],s251[497],s251[498],s250[500],s249[502],pp255[252],pp254[254],pp255[254]};
    CLA_508 KS_253(s253, c253, in253_1, in253_2);
    wire[505:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp2[1],s253[2],s253[3],s253[4],s253[5],s253[6],s253[7],s253[8],s253[9],s253[10],s253[11],s253[12],s253[13],s253[14],s253[15],s253[16],s253[17],s253[18],s253[19],s253[20],s253[21],s253[22],s253[23],s253[24],s253[25],s253[26],s253[27],s253[28],s253[29],s253[30],s253[31],s253[32],s253[33],s253[34],s253[35],s253[36],s253[37],s253[38],s253[39],s253[40],s253[41],s253[42],s253[43],s253[44],s253[45],s253[46],s253[47],s253[48],s253[49],s253[50],s253[51],s253[52],s253[53],s253[54],s253[55],s253[56],s253[57],s253[58],s253[59],s253[60],s253[61],s253[62],s253[63],s253[64],s253[65],s253[66],s253[67],s253[68],s253[69],s253[70],s253[71],s253[72],s253[73],s253[74],s253[75],s253[76],s253[77],s253[78],s253[79],s253[80],s253[81],s253[82],s253[83],s253[84],s253[85],s253[86],s253[87],s253[88],s253[89],s253[90],s253[91],s253[92],s253[93],s253[94],s253[95],s253[96],s253[97],s253[98],s253[99],s253[100],s253[101],s253[102],s253[103],s253[104],s253[105],s253[106],s253[107],s253[108],s253[109],s253[110],s253[111],s253[112],s253[113],s253[114],s253[115],s253[116],s253[117],s253[118],s253[119],s253[120],s253[121],s253[122],s253[123],s253[124],s253[125],s253[126],s253[127],s253[128],s253[129],s253[130],s253[131],s253[132],s253[133],s253[134],s253[135],s253[136],s253[137],s253[138],s253[139],s253[140],s253[141],s253[142],s253[143],s253[144],s253[145],s253[146],s253[147],s253[148],s253[149],s253[150],s253[151],s253[152],s253[153],s253[154],s253[155],s253[156],s253[157],s253[158],s253[159],s253[160],s253[161],s253[162],s253[163],s253[164],s253[165],s253[166],s253[167],s253[168],s253[169],s253[170],s253[171],s253[172],s253[173],s253[174],s253[175],s253[176],s253[177],s253[178],s253[179],s253[180],s253[181],s253[182],s253[183],s253[184],s253[185],s253[186],s253[187],s253[188],s253[189],s253[190],s253[191],s253[192],s253[193],s253[194],s253[195],s253[196],s253[197],s253[198],s253[199],s253[200],s253[201],s253[202],s253[203],s253[204],s253[205],s253[206],s253[207],s253[208],s253[209],s253[210],s253[211],s253[212],s253[213],s253[214],s253[215],s253[216],s253[217],s253[218],s253[219],s253[220],s253[221],s253[222],s253[223],s253[224],s253[225],s253[226],s253[227],s253[228],s253[229],s253[230],s253[231],s253[232],s253[233],s253[234],s253[235],s253[236],s253[237],s253[238],s253[239],s253[240],s253[241],s253[242],s253[243],s253[244],s253[245],s253[246],s253[247],s253[248],s253[249],s253[250],s253[251],s253[252],s253[253],s253[254],s253[255],s253[256],s253[257],s253[258],s253[259],s253[260],s253[261],s253[262],s253[263],s253[264],s253[265],s253[266],s253[267],s253[268],s253[269],s253[270],s253[271],s253[272],s253[273],s253[274],s253[275],s253[276],s253[277],s253[278],s253[279],s253[280],s253[281],s253[282],s253[283],s253[284],s253[285],s253[286],s253[287],s253[288],s253[289],s253[290],s253[291],s253[292],s253[293],s253[294],s253[295],s253[296],s253[297],s253[298],s253[299],s253[300],s253[301],s253[302],s253[303],s253[304],s253[305],s253[306],s253[307],s253[308],s253[309],s253[310],s253[311],s253[312],s253[313],s253[314],s253[315],s253[316],s253[317],s253[318],s253[319],s253[320],s253[321],s253[322],s253[323],s253[324],s253[325],s253[326],s253[327],s253[328],s253[329],s253[330],s253[331],s253[332],s253[333],s253[334],s253[335],s253[336],s253[337],s253[338],s253[339],s253[340],s253[341],s253[342],s253[343],s253[344],s253[345],s253[346],s253[347],s253[348],s253[349],s253[350],s253[351],s253[352],s253[353],s253[354],s253[355],s253[356],s253[357],s253[358],s253[359],s253[360],s253[361],s253[362],s253[363],s253[364],s253[365],s253[366],s253[367],s253[368],s253[369],s253[370],s253[371],s253[372],s253[373],s253[374],s253[375],s253[376],s253[377],s253[378],s253[379],s253[380],s253[381],s252[377],s252[378],s252[379],s252[380],s252[381],s252[382],s252[383],s252[384],s252[385],s252[386],s252[387],s252[388],s252[389],s252[390],s252[391],s252[392],s252[393],s252[394],s252[395],s252[396],s252[397],s252[398],s252[399],s252[400],s252[401],s252[402],s252[403],s252[404],s252[405],s252[406],s252[407],s252[408],s252[409],s252[410],s252[411],s252[412],s252[413],s252[414],s252[415],s252[416],s252[417],s252[418],s252[419],s252[420],s252[421],s252[422],s252[423],s252[424],s252[425],s252[426],s252[427],s252[428],s252[429],s252[430],s252[431],s252[432],s252[433],s252[434],s252[435],s252[436],s252[437],s252[438],s252[439],s252[440],s252[441],s252[442],s252[443],s252[444],s252[445],s252[446],s252[447],s252[448],s252[449],s252[450],s252[451],s252[452],s252[453],s252[454],s252[455],s252[456],s252[457],s252[458],s252[459],s252[460],s252[461],s252[462],s252[463],s252[464],s252[465],s252[466],s252[467],s252[468],s252[469],s252[470],s252[471],s252[472],s252[473],s252[474],s252[475],s252[476],s252[477],s252[478],s252[479],s252[480],s252[481],s252[482],s252[483],s252[484],s252[485],s252[486],s252[487],s252[488],s252[489],s252[490],s252[491],s252[492],s252[493],s252[494],s252[495],s252[496],s252[497],s251[499],s250[501],s249[503],pp255[253]};
    assign in254_2 = {pp3[0],pp3[1],pp4[1],pp5[1],pp6[1],pp7[1],pp8[1],pp8[2],pp8[3],pp8[4],pp8[5],pp8[6],pp8[7],pp8[8],pp8[9],s248[3],s247[5],s247[6],s247[7],s247[8],s247[9],s233[0],s233[1],s234[1],s235[1],s236[1],s237[1],s238[1],s239[1],s239[2],s239[3],s239[4],s239[5],s239[6],s239[7],s239[8],s239[9],s201[0],s201[1],s202[1],s203[1],s204[1],s205[1],s206[1],s207[1],s208[1],s209[1],s210[1],s211[1],s212[1],s213[1],s214[1],s215[1],s216[1],s217[1],s218[1],s219[1],s220[1],s221[1],s222[1],s223[1],s223[2],s223[3],s223[4],s223[5],s223[6],s223[7],s223[8],s223[9],s137[0],s137[1],s138[1],s139[1],s140[1],s141[1],s142[1],s143[1],s144[1],s145[1],s146[1],s147[1],s148[1],s149[1],s150[1],s151[1],s152[1],s153[1],s154[1],s155[1],s156[1],s157[1],s158[1],s159[1],s160[1],s161[1],s162[1],s163[1],s164[1],s165[1],s166[1],s167[1],s168[1],s169[1],s170[1],s171[1],s172[1],s173[1],s174[1],s175[1],s176[1],s177[1],s178[1],s179[1],s180[1],s181[1],s182[1],s183[1],s184[1],s185[1],s186[1],s187[1],s188[1],s189[1],s190[1],s191[1],s192[1],s1[1],s2[1],s3[1],s4[1],s5[1],s6[1],s7[1],s8[1],s8[2],s8[3],s8[4],s8[5],s8[6],s8[7],s8[8],s8[9],s18[0],s18[1],s19[1],s20[1],s21[1],s22[1],s23[1],s24[1],s25[1],s26[1],s27[1],s28[1],s29[1],s30[1],s31[1],s32[1],s33[1],s34[1],s35[1],s36[1],s37[1],s38[1],s39[1],s40[1],s41[1],s42[1],s43[1],s44[1],s45[1],s46[1],s47[1],s48[1],s49[1],s50[1],s51[1],s52[1],s53[1],s54[1],s55[1],s56[1],s57[1],s58[1],s59[1],s60[1],s61[1],s62[1],s63[1],s64[1],s65[1],s66[1],s67[1],s68[1],s69[1],s70[1],s71[1],s72[1],s73[1],s74[1],s75[1],s76[1],s77[1],s78[1],s79[1],s80[1],s81[1],s82[1],s83[1],s84[1],s85[1],s86[1],s87[1],s88[1],s89[1],s90[1],s91[1],s92[1],s93[1],s94[1],s95[1],s96[1],s97[1],s98[1],s98[2],s98[3],s98[4],s98[5],s98[6],s98[7],s98[8],s98[9],s9[99],s108[1],s109[1],s110[1],s111[1],s112[1],s113[1],s114[1],s115[1],s116[1],s117[1],s118[1],s119[1],s120[1],s121[1],s122[1],s123[1],s124[1],s125[1],s126[1],s127[1],s128[1],s127[3],s126[5],s125[7],s124[9],s99[35],s99[36],s99[37],s99[38],s99[39],s99[40],s99[41],s99[42],s99[43],s99[44],s99[45],s99[46],s99[47],s99[48],s99[49],s99[50],s99[51],s99[52],s99[53],s99[54],s99[55],s99[56],s99[57],s99[58],s99[59],s98[61],s97[63],s96[65],s95[67],s94[69],s93[71],s92[73],s91[75],s90[77],s89[79],s88[81],s87[83],s86[85],s85[87],s84[89],s83[91],s82[93],s81[95],s80[97],s79[99],s9[170],s9[171],s9[172],s9[173],s9[174],s9[175],s9[176],s9[177],s9[178],s9[179],s9[180],s9[181],s9[182],s9[183],s9[184],s9[185],s9[186],s9[187],s9[188],s9[189],s9[190],s9[191],s9[192],s9[193],s9[194],s9[195],s9[196],s9[197],s9[198],s9[199],s9[200],s9[201],s9[202],s9[203],s9[204],s9[205],s9[206],s9[207],s9[208],s9[209],s9[210],s9[211],s9[212],s9[213],s9[214],s9[215],s9[216],s9[217],s9[218],s9[219],s9[220],s9[221],s9[222],s9[223],s9[224],s9[225],s9[226],s9[227],s9[228],s9[229],s9[230],s9[231],s9[232],s9[233],s9[234],s9[235],s9[236],s9[237],s9[238],s9[239],s8[241],s7[243],s6[245],s5[247],s4[249],s3[251],s2[253],s1[255],s253[382],s253[383],s253[384],s253[385],s253[386],s253[387],s253[388],s253[389],s253[390],s253[391],s253[392],s253[393],s253[394],s253[395],s253[396],s253[397],s253[398],s253[399],s253[400],s253[401],s253[402],s253[403],s253[404],s253[405],s253[406],s253[407],s253[408],s253[409],s253[410],s253[411],s253[412],s253[413],s253[414],s253[415],s253[416],s253[417],s253[418],s253[419],s253[420],s253[421],s253[422],s253[423],s253[424],s253[425],s253[426],s253[427],s253[428],s253[429],s253[430],s253[431],s253[432],s253[433],s253[434],s253[435],s253[436],s253[437],s253[438],s253[439],s253[440],s253[441],s253[442],s253[443],s253[444],s253[445],s253[446],s253[447],s253[448],s253[449],s253[450],s253[451],s253[452],s253[453],s253[454],s253[455],s253[456],s253[457],s253[458],s253[459],s253[460],s253[461],s253[462],s253[463],s253[464],s253[465],s253[466],s253[467],s253[468],s253[469],s253[470],s253[471],s253[472],s253[473],s253[474],s253[475],s253[476],s253[477],s253[478],s253[479],s253[480],s253[481],s253[482],s253[483],s253[484],s253[485],s253[486],s253[487],s253[488],s253[489],s253[490],s253[491],s253[492],s253[493],s253[494],s253[495],s253[496],s253[497],s253[498],s253[499],s253[500],s253[501],s253[502],s253[503],s253[504],s253[505],s253[506]};
    CLA_506 KS_254(s254, c254, in254_1, in254_2);


    /*Final Stage 7*/
    wire[509:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],s253[0],s253[1],pp4[0],pp5[0],pp6[0],pp7[0],pp8[0],pp9[0],pp9[1],pp9[2],pp9[3],pp9[4],pp9[5],pp9[6],pp9[7],pp9[8],pp9[9],s248[4],s248[5],s248[6],s248[7],s248[8],s248[9],s234[0],s235[0],s236[0],s237[0],s238[0],s239[0],s240[0],s240[1],s240[2],s240[3],s240[4],s240[5],s240[6],s240[7],s240[8],s240[9],s202[0],s203[0],s204[0],s205[0],s206[0],s207[0],s208[0],s209[0],s210[0],s211[0],s212[0],s213[0],s214[0],s215[0],s216[0],s217[0],s218[0],s219[0],s220[0],s221[0],s222[0],s223[0],s224[0],s224[1],s224[2],s224[3],s224[4],s224[5],s224[6],s224[7],s224[8],s224[9],s138[0],s139[0],s140[0],s141[0],s142[0],s143[0],s144[0],s145[0],s146[0],s147[0],s148[0],s149[0],s150[0],s151[0],s152[0],s153[0],s154[0],s155[0],s156[0],s157[0],s158[0],s159[0],s160[0],s161[0],s162[0],s163[0],s164[0],s165[0],s166[0],s167[0],s168[0],s169[0],s170[0],s171[0],s172[0],s173[0],s174[0],s175[0],s176[0],s177[0],s178[0],s179[0],s180[0],s181[0],s182[0],s183[0],s184[0],s185[0],s186[0],s187[0],s188[0],s189[0],s190[0],s191[0],s192[0],s1[0],s2[0],s3[0],s4[0],s5[0],s6[0],s7[0],s8[0],s9[0],s9[1],s9[2],s9[3],s9[4],s9[5],s9[6],s9[7],s9[8],s9[9],s19[0],s20[0],s21[0],s22[0],s23[0],s24[0],s25[0],s26[0],s27[0],s28[0],s29[0],s30[0],s31[0],s32[0],s33[0],s34[0],s35[0],s36[0],s37[0],s38[0],s39[0],s40[0],s41[0],s42[0],s43[0],s44[0],s45[0],s46[0],s47[0],s48[0],s49[0],s50[0],s51[0],s52[0],s53[0],s54[0],s55[0],s56[0],s57[0],s58[0],s59[0],s60[0],s61[0],s62[0],s63[0],s64[0],s65[0],s66[0],s67[0],s68[0],s69[0],s70[0],s71[0],s72[0],s73[0],s74[0],s75[0],s76[0],s77[0],s78[0],s79[0],s80[0],s81[0],s82[0],s83[0],s84[0],s85[0],s86[0],s87[0],s88[0],s89[0],s90[0],s91[0],s92[0],s93[0],s94[0],s95[0],s96[0],s97[0],s98[0],s99[0],s99[1],s99[2],s99[3],s99[4],s99[5],s99[6],s99[7],s99[8],s99[9],s109[0],s110[0],s111[0],s112[0],s113[0],s114[0],s115[0],s116[0],s117[0],s118[0],s119[0],s120[0],s121[0],s122[0],s123[0],s124[0],s125[0],s126[0],s127[0],s128[0],1'b0,c128,c127,c126,c125,c124,c123,c122,c121,c120,c119,c118,c117,c116,c115,c114,c113,c112,c111,c110,c109,c108,c107,c106,c105,c104,c103,c102,c101,c100,c99,c98,c97,c96,c95,c94,c93,c92,c91,c90,c89,c88,c87,c86,c85,c84,c83,c82,c81,c80,c79,c78,c77,c76,c75,c74,c73,c72,c71,c70,c69,c68,c67,c66,c65,c64,c63,c62,c61,c60,c59,c58,c57,c56,c55,c54,c53,c52,c51,c50,c49,c48,c47,c46,c45,c44,c43,c42,c41,c40,c39,c38,c37,c36,c35,c34,c33,c32,c31,c30,c29,c28,c27,c26,c25,c24,c23,c22,c21,c20,c19,c18,c17,c16,c15,c14,c13,c12,c11,c10,c9,c8,c7,c6,c5,c4,c3,c2,c1,c192,c191,c190,c189,c188,c187,c186,c185,c184,c183,c182,c181,c180,c179,c178,c177,c176,c175,c174,c173,c172,c171,c170,c169,c168,c167,c166,c165,c164,c163,c162,c161,c160,c159,c158,c157,c156,c155,c154,c153,c152,c151,c150,c149,c148,c147,c146,c145,c144,c143,c142,c141,c140,c139,c138,c137,c136,c135,c134,c133,c132,c131,c130,c129,c224,c223,c222,c221,c220,c219,c218,c217,c216,c215,c214,c213,c212,c211,c210,c209,c208,c207,c206,c205,c204,c203,c202,c201,c200,c199,c198,c197,c196,c195,c194,c193,c240,c239,c238,c237,c236,c235,c234,c233,c232,c231,c230,c229,c228,c227,c226,c225,c248,c247,c246,c245,c244,c243,c242,c241,c252,c251,c250,c249,s253[507],pp255[255]};
    assign in_2 = {pp1[0],pp2[0],s254[0],s254[1],s254[2],s254[3],s254[4],s254[5],s254[6],s254[7],s254[8],s254[9],s254[10],s254[11],s254[12],s254[13],s254[14],s254[15],s254[16],s254[17],s254[18],s254[19],s254[20],s254[21],s254[22],s254[23],s254[24],s254[25],s254[26],s254[27],s254[28],s254[29],s254[30],s254[31],s254[32],s254[33],s254[34],s254[35],s254[36],s254[37],s254[38],s254[39],s254[40],s254[41],s254[42],s254[43],s254[44],s254[45],s254[46],s254[47],s254[48],s254[49],s254[50],s254[51],s254[52],s254[53],s254[54],s254[55],s254[56],s254[57],s254[58],s254[59],s254[60],s254[61],s254[62],s254[63],s254[64],s254[65],s254[66],s254[67],s254[68],s254[69],s254[70],s254[71],s254[72],s254[73],s254[74],s254[75],s254[76],s254[77],s254[78],s254[79],s254[80],s254[81],s254[82],s254[83],s254[84],s254[85],s254[86],s254[87],s254[88],s254[89],s254[90],s254[91],s254[92],s254[93],s254[94],s254[95],s254[96],s254[97],s254[98],s254[99],s254[100],s254[101],s254[102],s254[103],s254[104],s254[105],s254[106],s254[107],s254[108],s254[109],s254[110],s254[111],s254[112],s254[113],s254[114],s254[115],s254[116],s254[117],s254[118],s254[119],s254[120],s254[121],s254[122],s254[123],s254[124],s254[125],s254[126],s254[127],s254[128],s254[129],s254[130],s254[131],s254[132],s254[133],s254[134],s254[135],s254[136],s254[137],s254[138],s254[139],s254[140],s254[141],s254[142],s254[143],s254[144],s254[145],s254[146],s254[147],s254[148],s254[149],s254[150],s254[151],s254[152],s254[153],s254[154],s254[155],s254[156],s254[157],s254[158],s254[159],s254[160],s254[161],s254[162],s254[163],s254[164],s254[165],s254[166],s254[167],s254[168],s254[169],s254[170],s254[171],s254[172],s254[173],s254[174],s254[175],s254[176],s254[177],s254[178],s254[179],s254[180],s254[181],s254[182],s254[183],s254[184],s254[185],s254[186],s254[187],s254[188],s254[189],s254[190],s254[191],s254[192],s254[193],s254[194],s254[195],s254[196],s254[197],s254[198],s254[199],s254[200],s254[201],s254[202],s254[203],s254[204],s254[205],s254[206],s254[207],s254[208],s254[209],s254[210],s254[211],s254[212],s254[213],s254[214],s254[215],s254[216],s254[217],s254[218],s254[219],s254[220],s254[221],s254[222],s254[223],s254[224],s254[225],s254[226],s254[227],s254[228],s254[229],s254[230],s254[231],s254[232],s254[233],s254[234],s254[235],s254[236],s254[237],s254[238],s254[239],s254[240],s254[241],s254[242],s254[243],s254[244],s254[245],s254[246],s254[247],s254[248],s254[249],s254[250],s254[251],s254[252],s254[253],s254[254],s254[255],s254[256],s254[257],s254[258],s254[259],s254[260],s254[261],s254[262],s254[263],s254[264],s254[265],s254[266],s254[267],s254[268],s254[269],s254[270],s254[271],s254[272],s254[273],s254[274],s254[275],s254[276],s254[277],s254[278],s254[279],s254[280],s254[281],s254[282],s254[283],s254[284],s254[285],s254[286],s254[287],s254[288],s254[289],s254[290],s254[291],s254[292],s254[293],s254[294],s254[295],s254[296],s254[297],s254[298],s254[299],s254[300],s254[301],s254[302],s254[303],s254[304],s254[305],s254[306],s254[307],s254[308],s254[309],s254[310],s254[311],s254[312],s254[313],s254[314],s254[315],s254[316],s254[317],s254[318],s254[319],s254[320],s254[321],s254[322],s254[323],s254[324],s254[325],s254[326],s254[327],s254[328],s254[329],s254[330],s254[331],s254[332],s254[333],s254[334],s254[335],s254[336],s254[337],s254[338],s254[339],s254[340],s254[341],s254[342],s254[343],s254[344],s254[345],s254[346],s254[347],s254[348],s254[349],s254[350],s254[351],s254[352],s254[353],s254[354],s254[355],s254[356],s254[357],s254[358],s254[359],s254[360],s254[361],s254[362],s254[363],s254[364],s254[365],s254[366],s254[367],s254[368],s254[369],s254[370],s254[371],s254[372],s254[373],s254[374],s254[375],s254[376],s254[377],s254[378],s254[379],s254[380],s254[381],s254[382],s254[383],s254[384],s254[385],s254[386],s254[387],s254[388],s254[389],s254[390],s254[391],s254[392],s254[393],s254[394],s254[395],s254[396],s254[397],s254[398],s254[399],s254[400],s254[401],s254[402],s254[403],s254[404],s254[405],s254[406],s254[407],s254[408],s254[409],s254[410],s254[411],s254[412],s254[413],s254[414],s254[415],s254[416],s254[417],s254[418],s254[419],s254[420],s254[421],s254[422],s254[423],s254[424],s254[425],s254[426],s254[427],s254[428],s254[429],s254[430],s254[431],s254[432],s254[433],s254[434],s254[435],s254[436],s254[437],s254[438],s254[439],s254[440],s254[441],s254[442],s254[443],s254[444],s254[445],s254[446],s254[447],s254[448],s254[449],s254[450],s254[451],s254[452],s254[453],s254[454],s254[455],s254[456],s254[457],s254[458],s254[459],s254[460],s254[461],s254[462],s254[463],s254[464],s254[465],s254[466],s254[467],s254[468],s254[469],s254[470],s254[471],s254[472],s254[473],s254[474],s254[475],s254[476],s254[477],s254[478],s254[479],s254[480],s254[481],s254[482],s254[483],s254[484],s254[485],s254[486],s254[487],s254[488],s254[489],s254[490],s254[491],s254[492],s254[493],s254[494],s254[495],s254[496],s254[497],s254[498],s254[499],s254[500],s254[501],s254[502],s254[503],s254[504],s254[505],c254,c253};
    CLA_510(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = s[126];
    assign product[128] = s[127];
    assign product[129] = s[128];
    assign product[130] = s[129];
    assign product[131] = s[130];
    assign product[132] = s[131];
    assign product[133] = s[132];
    assign product[134] = s[133];
    assign product[135] = s[134];
    assign product[136] = s[135];
    assign product[137] = s[136];
    assign product[138] = s[137];
    assign product[139] = s[138];
    assign product[140] = s[139];
    assign product[141] = s[140];
    assign product[142] = s[141];
    assign product[143] = s[142];
    assign product[144] = s[143];
    assign product[145] = s[144];
    assign product[146] = s[145];
    assign product[147] = s[146];
    assign product[148] = s[147];
    assign product[149] = s[148];
    assign product[150] = s[149];
    assign product[151] = s[150];
    assign product[152] = s[151];
    assign product[153] = s[152];
    assign product[154] = s[153];
    assign product[155] = s[154];
    assign product[156] = s[155];
    assign product[157] = s[156];
    assign product[158] = s[157];
    assign product[159] = s[158];
    assign product[160] = s[159];
    assign product[161] = s[160];
    assign product[162] = s[161];
    assign product[163] = s[162];
    assign product[164] = s[163];
    assign product[165] = s[164];
    assign product[166] = s[165];
    assign product[167] = s[166];
    assign product[168] = s[167];
    assign product[169] = s[168];
    assign product[170] = s[169];
    assign product[171] = s[170];
    assign product[172] = s[171];
    assign product[173] = s[172];
    assign product[174] = s[173];
    assign product[175] = s[174];
    assign product[176] = s[175];
    assign product[177] = s[176];
    assign product[178] = s[177];
    assign product[179] = s[178];
    assign product[180] = s[179];
    assign product[181] = s[180];
    assign product[182] = s[181];
    assign product[183] = s[182];
    assign product[184] = s[183];
    assign product[185] = s[184];
    assign product[186] = s[185];
    assign product[187] = s[186];
    assign product[188] = s[187];
    assign product[189] = s[188];
    assign product[190] = s[189];
    assign product[191] = s[190];
    assign product[192] = s[191];
    assign product[193] = s[192];
    assign product[194] = s[193];
    assign product[195] = s[194];
    assign product[196] = s[195];
    assign product[197] = s[196];
    assign product[198] = s[197];
    assign product[199] = s[198];
    assign product[200] = s[199];
    assign product[201] = s[200];
    assign product[202] = s[201];
    assign product[203] = s[202];
    assign product[204] = s[203];
    assign product[205] = s[204];
    assign product[206] = s[205];
    assign product[207] = s[206];
    assign product[208] = s[207];
    assign product[209] = s[208];
    assign product[210] = s[209];
    assign product[211] = s[210];
    assign product[212] = s[211];
    assign product[213] = s[212];
    assign product[214] = s[213];
    assign product[215] = s[214];
    assign product[216] = s[215];
    assign product[217] = s[216];
    assign product[218] = s[217];
    assign product[219] = s[218];
    assign product[220] = s[219];
    assign product[221] = s[220];
    assign product[222] = s[221];
    assign product[223] = s[222];
    assign product[224] = s[223];
    assign product[225] = s[224];
    assign product[226] = s[225];
    assign product[227] = s[226];
    assign product[228] = s[227];
    assign product[229] = s[228];
    assign product[230] = s[229];
    assign product[231] = s[230];
    assign product[232] = s[231];
    assign product[233] = s[232];
    assign product[234] = s[233];
    assign product[235] = s[234];
    assign product[236] = s[235];
    assign product[237] = s[236];
    assign product[238] = s[237];
    assign product[239] = s[238];
    assign product[240] = s[239];
    assign product[241] = s[240];
    assign product[242] = s[241];
    assign product[243] = s[242];
    assign product[244] = s[243];
    assign product[245] = s[244];
    assign product[246] = s[245];
    assign product[247] = s[246];
    assign product[248] = s[247];
    assign product[249] = s[248];
    assign product[250] = s[249];
    assign product[251] = s[250];
    assign product[252] = s[251];
    assign product[253] = s[252];
    assign product[254] = s[253];
    assign product[255] = s[254];
    assign product[256] = s[255];
    assign product[257] = s[256];
    assign product[258] = s[257];
    assign product[259] = s[258];
    assign product[260] = s[259];
    assign product[261] = s[260];
    assign product[262] = s[261];
    assign product[263] = s[262];
    assign product[264] = s[263];
    assign product[265] = s[264];
    assign product[266] = s[265];
    assign product[267] = s[266];
    assign product[268] = s[267];
    assign product[269] = s[268];
    assign product[270] = s[269];
    assign product[271] = s[270];
    assign product[272] = s[271];
    assign product[273] = s[272];
    assign product[274] = s[273];
    assign product[275] = s[274];
    assign product[276] = s[275];
    assign product[277] = s[276];
    assign product[278] = s[277];
    assign product[279] = s[278];
    assign product[280] = s[279];
    assign product[281] = s[280];
    assign product[282] = s[281];
    assign product[283] = s[282];
    assign product[284] = s[283];
    assign product[285] = s[284];
    assign product[286] = s[285];
    assign product[287] = s[286];
    assign product[288] = s[287];
    assign product[289] = s[288];
    assign product[290] = s[289];
    assign product[291] = s[290];
    assign product[292] = s[291];
    assign product[293] = s[292];
    assign product[294] = s[293];
    assign product[295] = s[294];
    assign product[296] = s[295];
    assign product[297] = s[296];
    assign product[298] = s[297];
    assign product[299] = s[298];
    assign product[300] = s[299];
    assign product[301] = s[300];
    assign product[302] = s[301];
    assign product[303] = s[302];
    assign product[304] = s[303];
    assign product[305] = s[304];
    assign product[306] = s[305];
    assign product[307] = s[306];
    assign product[308] = s[307];
    assign product[309] = s[308];
    assign product[310] = s[309];
    assign product[311] = s[310];
    assign product[312] = s[311];
    assign product[313] = s[312];
    assign product[314] = s[313];
    assign product[315] = s[314];
    assign product[316] = s[315];
    assign product[317] = s[316];
    assign product[318] = s[317];
    assign product[319] = s[318];
    assign product[320] = s[319];
    assign product[321] = s[320];
    assign product[322] = s[321];
    assign product[323] = s[322];
    assign product[324] = s[323];
    assign product[325] = s[324];
    assign product[326] = s[325];
    assign product[327] = s[326];
    assign product[328] = s[327];
    assign product[329] = s[328];
    assign product[330] = s[329];
    assign product[331] = s[330];
    assign product[332] = s[331];
    assign product[333] = s[332];
    assign product[334] = s[333];
    assign product[335] = s[334];
    assign product[336] = s[335];
    assign product[337] = s[336];
    assign product[338] = s[337];
    assign product[339] = s[338];
    assign product[340] = s[339];
    assign product[341] = s[340];
    assign product[342] = s[341];
    assign product[343] = s[342];
    assign product[344] = s[343];
    assign product[345] = s[344];
    assign product[346] = s[345];
    assign product[347] = s[346];
    assign product[348] = s[347];
    assign product[349] = s[348];
    assign product[350] = s[349];
    assign product[351] = s[350];
    assign product[352] = s[351];
    assign product[353] = s[352];
    assign product[354] = s[353];
    assign product[355] = s[354];
    assign product[356] = s[355];
    assign product[357] = s[356];
    assign product[358] = s[357];
    assign product[359] = s[358];
    assign product[360] = s[359];
    assign product[361] = s[360];
    assign product[362] = s[361];
    assign product[363] = s[362];
    assign product[364] = s[363];
    assign product[365] = s[364];
    assign product[366] = s[365];
    assign product[367] = s[366];
    assign product[368] = s[367];
    assign product[369] = s[368];
    assign product[370] = s[369];
    assign product[371] = s[370];
    assign product[372] = s[371];
    assign product[373] = s[372];
    assign product[374] = s[373];
    assign product[375] = s[374];
    assign product[376] = s[375];
    assign product[377] = s[376];
    assign product[378] = s[377];
    assign product[379] = s[378];
    assign product[380] = s[379];
    assign product[381] = s[380];
    assign product[382] = s[381];
    assign product[383] = s[382];
    assign product[384] = s[383];
    assign product[385] = s[384];
    assign product[386] = s[385];
    assign product[387] = s[386];
    assign product[388] = s[387];
    assign product[389] = s[388];
    assign product[390] = s[389];
    assign product[391] = s[390];
    assign product[392] = s[391];
    assign product[393] = s[392];
    assign product[394] = s[393];
    assign product[395] = s[394];
    assign product[396] = s[395];
    assign product[397] = s[396];
    assign product[398] = s[397];
    assign product[399] = s[398];
    assign product[400] = s[399];
    assign product[401] = s[400];
    assign product[402] = s[401];
    assign product[403] = s[402];
    assign product[404] = s[403];
    assign product[405] = s[404];
    assign product[406] = s[405];
    assign product[407] = s[406];
    assign product[408] = s[407];
    assign product[409] = s[408];
    assign product[410] = s[409];
    assign product[411] = s[410];
    assign product[412] = s[411];
    assign product[413] = s[412];
    assign product[414] = s[413];
    assign product[415] = s[414];
    assign product[416] = s[415];
    assign product[417] = s[416];
    assign product[418] = s[417];
    assign product[419] = s[418];
    assign product[420] = s[419];
    assign product[421] = s[420];
    assign product[422] = s[421];
    assign product[423] = s[422];
    assign product[424] = s[423];
    assign product[425] = s[424];
    assign product[426] = s[425];
    assign product[427] = s[426];
    assign product[428] = s[427];
    assign product[429] = s[428];
    assign product[430] = s[429];
    assign product[431] = s[430];
    assign product[432] = s[431];
    assign product[433] = s[432];
    assign product[434] = s[433];
    assign product[435] = s[434];
    assign product[436] = s[435];
    assign product[437] = s[436];
    assign product[438] = s[437];
    assign product[439] = s[438];
    assign product[440] = s[439];
    assign product[441] = s[440];
    assign product[442] = s[441];
    assign product[443] = s[442];
    assign product[444] = s[443];
    assign product[445] = s[444];
    assign product[446] = s[445];
    assign product[447] = s[446];
    assign product[448] = s[447];
    assign product[449] = s[448];
    assign product[450] = s[449];
    assign product[451] = s[450];
    assign product[452] = s[451];
    assign product[453] = s[452];
    assign product[454] = s[453];
    assign product[455] = s[454];
    assign product[456] = s[455];
    assign product[457] = s[456];
    assign product[458] = s[457];
    assign product[459] = s[458];
    assign product[460] = s[459];
    assign product[461] = s[460];
    assign product[462] = s[461];
    assign product[463] = s[462];
    assign product[464] = s[463];
    assign product[465] = s[464];
    assign product[466] = s[465];
    assign product[467] = s[466];
    assign product[468] = s[467];
    assign product[469] = s[468];
    assign product[470] = s[469];
    assign product[471] = s[470];
    assign product[472] = s[471];
    assign product[473] = s[472];
    assign product[474] = s[473];
    assign product[475] = s[474];
    assign product[476] = s[475];
    assign product[477] = s[476];
    assign product[478] = s[477];
    assign product[479] = s[478];
    assign product[480] = s[479];
    assign product[481] = s[480];
    assign product[482] = s[481];
    assign product[483] = s[482];
    assign product[484] = s[483];
    assign product[485] = s[484];
    assign product[486] = s[485];
    assign product[487] = s[486];
    assign product[488] = s[487];
    assign product[489] = s[488];
    assign product[490] = s[489];
    assign product[491] = s[490];
    assign product[492] = s[491];
    assign product[493] = s[492];
    assign product[494] = s[493];
    assign product[495] = s[494];
    assign product[496] = s[495];
    assign product[497] = s[496];
    assign product[498] = s[497];
    assign product[499] = s[498];
    assign product[500] = s[499];
    assign product[501] = s[500];
    assign product[502] = s[501];
    assign product[503] = s[502];
    assign product[504] = s[503];
    assign product[505] = s[504];
    assign product[506] = s[505];
    assign product[507] = s[506];
    assign product[508] = s[507];
    assign product[509] = s[508];
    assign product[510] = s[509];
    assign product[511] = c;
endmodule


