module russian_peasant_modified_unsigned_multiplier_16(product, A, B);
    /* This implementation uses carry look-ahead adders of
     * variable lengths and can extend upto 15 bits long */

    input  [15:0] A, B;
    output [31:0] product;

    wire [31:0] product;
    wire [15:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;

    assign pp0 = A[0] ? B : 16'b00000000;
    assign pp1 = A[1] ? B : 16'b00000000;
    assign pp2 = A[2] ? B : 16'b00000000;
    assign pp3 = A[3] ? B : 16'b00000000;
    assign pp4 = A[4] ? B : 16'b00000000;
    assign pp5 = A[5] ? B : 16'b00000000;
    assign pp6 = A[6] ? B : 16'b00000000;
    assign pp7 = A[7] ? B : 16'b00000000;
    assign pp8 = A[8] ? B : 16'b00000000;
    assign pp9 = A[9] ? B : 16'b00000000;
    assign pp10 = A[10] ? B : 16'b00000000;
    assign pp11 = A[11] ? B : 16'b00000000;
    assign pp12 = A[12] ? B : 16'b00000000;
    assign pp13 = A[13] ? B : 16'b00000000;
    assign pp14 = A[14] ? B : 16'b00000000;
    assign pp15 = A[15] ? B : 16'b00000000;

    assign product[0] = pp0[0];

    /* 1st CLA */
    wire [15:0] G1, P1, C1;
    assign G1[0]  = pp0[1]  & pp1[0];
    assign G1[1]  = pp0[2]  & pp1[1];
    assign G1[2]  = pp0[3]  & pp1[2];
    assign G1[3]  = pp0[4]  & pp1[3];
    assign G1[4]  = pp0[5]  & pp1[4];
    assign G1[5]  = pp0[6]  & pp1[5];
    assign G1[6]  = pp0[7]  & pp1[6];
    assign G1[7]  = pp0[8]  & pp1[7];
    assign G1[8]  = pp0[9]  & pp1[8];
    assign G1[9]  = pp0[10] & pp1[9];
    assign G1[10] = pp0[11] & pp1[10];
    assign G1[11] = pp0[12] & pp1[11];
    assign G1[12] = pp0[13] & pp1[12];
    assign G1[13] = pp0[14] & pp1[13];
    assign G1[14] = pp0[15] & pp1[14];
    assign G1[15] = 0       & pp1[15];
    assign P1[0]  = pp0[1]  ^ pp1[0];
    assign P1[1]  = pp0[2]  ^ pp1[1];
    assign P1[2]  = pp0[3]  ^ pp1[2];
    assign P1[3]  = pp0[4]  ^ pp1[3];
    assign P1[4]  = pp0[5]  ^ pp1[4];
    assign P1[5]  = pp0[6]  ^ pp1[5];
    assign P1[6]  = pp0[7]  ^ pp1[6];
    assign P1[7]  = pp0[8]  ^ pp1[7];
    assign P1[8]  = pp0[9]  ^ pp1[8];
    assign P1[9]  = pp0[10] ^ pp1[9];
    assign P1[10] = pp0[11] ^ pp1[10];
    assign P1[11] = pp0[12] ^ pp1[11];
    assign P1[12] = pp0[13] ^ pp1[12];
    assign P1[13] = pp0[14] ^ pp1[13];
    assign P1[14] = pp0[15] ^ pp1[14];
    assign P1[15] = 0       ^ pp1[15];
    assign C1[0]  = 0;
    assign C1[1]  = G1[0]  | (P1[0] & C1[0]);
    assign C1[2]  = G1[1]  | (P1[1] & C1[1]);
    assign C1[3]  = G1[2]  | (P1[2] & C1[2]);
    assign C1[4]  = G1[3]  | (P1[3] & C1[3]);
    assign C1[5]  = G1[4]  | (P1[4] & C1[4]);
    assign C1[6]  = G1[5]  | (P1[5] & C1[5]);
    assign C1[7]  = G1[6]  | (P1[6] & C1[6]);
    assign C1[8]  = G1[7]  | (P1[7] & C1[7]);
    assign C1[9]  = G1[8]  | (P1[8] & C1[8]);
    assign C1[10] = G1[9]  | (P1[9] & C1[9]);
    assign C1[11] = G1[10] | (P1[10] & C1[10]);
    assign C1[12] = G1[11] | (P1[11] & C1[11]);
    assign C1[13] = G1[12] | (P1[12] & C1[12]);
    assign C1[14] = G1[13] | (P1[13] & C1[13]);
    assign C1[15] = G1[14] | (P1[14] & C1[14]);
    assign c1     = G1[15] | (P1[15] & C1[15]);
    assign s101   = P1[0];
    assign s102   = P1[1]  ^ C1[1];
    assign s103   = P1[2]  ^ C1[2];
    assign s104   = P1[3]  ^ C1[3];
    assign s105   = P1[4]  ^ C1[4];
    assign s106   = P1[5]  ^ C1[5];
    assign s107   = P1[6]  ^ C1[6];
    assign s108   = P1[7]  ^ C1[7];
    assign s109   = P1[8]  ^ C1[8];
    assign s110   = P1[9]  ^ C1[9];
    assign s111   = P1[10] ^ C1[10];
    assign s112   = P1[11] ^ C1[11];
    assign s113   = P1[12] ^ C1[12];
    assign s114   = P1[13] ^ C1[13];
    assign s115   = P1[14] ^ C1[14];
    assign s116   = P1[15] ^ C1[15];

    assign product[1] = s101;

    /* 2nd CLA */
    wire [14:0] G2, P2, C2;
    assign G2[0]  = pp2[1]  & pp3[0];
    assign G2[1]  = pp2[2]  & pp3[1];
    assign G2[2]  = pp2[3]  & pp3[2];
    assign G2[3]  = pp2[4]  & pp3[3];
    assign G2[4]  = pp2[5]  & pp3[4];
    assign G2[5]  = pp2[6]  & pp3[5];
    assign G2[6]  = pp2[7]  & pp3[6];
    assign G2[7]  = pp2[8]  & pp3[7];
    assign G2[8]  = pp2[9]  & pp3[8];
    assign G2[9]  = pp2[10] & pp3[9];
    assign G2[10] = pp2[11] & pp3[10];
    assign G2[11] = pp2[12] & pp3[11];
    assign G2[12] = pp2[13] & pp3[12];
    assign G2[13] = pp2[14] & pp3[13];
    assign G2[14] = pp2[15] & pp3[14];
    assign P2[0]  = pp2[1]  ^ pp3[0];
    assign P2[1]  = pp2[2]  ^ pp3[1];
    assign P2[2]  = pp2[3]  ^ pp3[2];
    assign P2[3]  = pp2[4]  ^ pp3[3];
    assign P2[4]  = pp2[5]  ^ pp3[4];
    assign P2[5]  = pp2[6]  ^ pp3[5];
    assign P2[6]  = pp2[7]  ^ pp3[6];
    assign P2[7]  = pp2[8]  ^ pp3[7];
    assign P2[8]  = pp2[9]  ^ pp3[8];
    assign P2[9]  = pp2[10] ^ pp3[9];
    assign P2[10] = pp2[11] ^ pp3[10];
    assign P2[11] = pp2[12] ^ pp3[11];
    assign P2[12] = pp2[13] ^ pp3[12];
    assign P2[13] = pp2[14] ^ pp3[13];
    assign P2[14] = pp2[15] ^ pp3[14];
    assign C2[0]  = 0;
    assign C2[1]  = G2[0]  | (P2[0]  & C2[0]);
    assign C2[2]  = G2[1]  | (P2[1]  & C2[1]);
    assign C2[3]  = G2[2]  | (P2[2]  & C2[2]);
    assign C2[4]  = G2[3]  | (P2[3]  & C2[3]);
    assign C2[5]  = G2[4]  | (P2[4]  & C2[4]);
    assign C2[6]  = G2[5]  | (P2[5]  & C2[5]);
    assign C2[7]  = G2[6]  | (P2[6]  & C2[6]);
    assign C2[8]  = G2[7]  | (P2[7]  & C2[7]);
    assign C2[9]  = G2[8]  | (P2[8]  & C2[8]);
    assign C2[10] = G2[9]  | (P2[9]  & C2[9]);
    assign C2[11] = G2[10] | (P2[10] & C2[10]);
    assign C2[12] = G2[11] | (P2[11] & C2[11]);
    assign C2[13] = G2[12] | (P2[12] & C2[12]);
    assign C2[14] = G2[13] | (P2[13] & C2[13]);
    assign c2     = G2[14] | (P2[14] & C2[14]);
    assign s201   = P2[0];
    assign s202   = P2[1]  ^ C2[1];
    assign s203   = P2[2]  ^ C2[2];
    assign s204   = P2[3]  ^ C2[3];
    assign s205   = P2[4]  ^ C2[4];
    assign s206   = P2[5]  ^ C2[5];
    assign s207   = P2[6]  ^ C2[6];
    assign s208   = P2[7]  ^ C2[7];
    assign s209   = P2[8]  ^ C2[8];
    assign s210   = P2[9]  ^ C2[9];
    assign s211   = P2[10] ^ C2[10];
    assign s212   = P2[11] ^ C2[11];
    assign s213   = P2[12] ^ C2[12];
    assign s214   = P2[13] ^ C2[13];
    assign s215   = P2[14] ^ C2[14];



     /* 3rd CLA */
    wire [14:0] G3, P3, C3;
    assign G3[0]  = pp4[1]  & pp5[0];
    assign G3[1]  = pp4[2]  & pp5[1];
    assign G3[2]  = pp4[3]  & pp5[2];
    assign G3[3]  = pp4[4]  & pp5[3];
    assign G3[4]  = pp4[5]  & pp5[4];
    assign G3[5]  = pp4[6]  & pp5[5];
    assign G3[6]  = pp4[7]  & pp5[6];
    assign G3[7]  = pp4[8]  & pp5[7];
    assign G3[8]  = pp4[9]  & pp5[8];
    assign G3[9]  = pp4[10] & pp5[9];
    assign G3[10] = pp4[11] & pp5[10];
    assign G3[11] = pp4[12] & pp5[11];
    assign G3[12] = pp4[13] & pp5[12];
    assign G3[13] = pp4[14] & pp5[13];
    assign G3[14] = pp4[15] & pp5[14];
    assign P3[0]  = pp4[1]  ^ pp5[0];
    assign P3[1]  = pp4[2]  ^ pp5[1];
    assign P3[2]  = pp4[3]  ^ pp5[2];
    assign P3[3]  = pp4[4]  ^ pp5[3];
    assign P3[4]  = pp4[5]  ^ pp5[4];
    assign P3[5]  = pp4[6]  ^ pp5[5];
    assign P3[6]  = pp4[7]  ^ pp5[6];
    assign P3[7]  = pp4[8]  ^ pp5[7];
    assign P3[8]  = pp4[9]  ^ pp5[8];
    assign P3[9]  = pp4[10] ^ pp5[9];
    assign P3[10] = pp4[11] ^ pp5[10];
    assign P3[11] = pp4[12] ^ pp5[11];
    assign P3[12] = pp4[13] ^ pp5[12];
    assign P3[13] = pp4[14] ^ pp5[13];
    assign P3[14] = pp4[15] ^ pp5[14];
    assign C3[0]  = 0;
    assign C3[1]  = G3[0]  | (P3[0] & C3[0]);
    assign C3[2]  = G3[1]  | (P3[1] & C3[1]);
    assign C3[3]  = G3[2]  | (P3[2] & C3[2]);
    assign C3[4]  = G3[3]  | (P3[3] & C3[3]);
    assign C3[5]  = G3[4]  | (P3[4] & C3[4]);
    assign C3[6]  = G3[5]  | (P3[5] & C3[5]);
    assign C3[7]  = G3[6]  | (P3[6] & C3[6]);
    assign C3[8]  = G3[7]  | (P3[7] & C3[7]);
    assign C3[9]  = G3[8]  | (P3[8] & C3[8]);
    assign C3[10] = G3[9]  | (P3[9] & C3[9]);
    assign C3[11] = G3[10] | (P3[10] & C3[10]);
    assign C3[12] = G3[11] | (P3[11] & C3[11]);
    assign C3[13] = G3[12] | (P3[12] & C3[12]);
    assign C3[14] = G3[13] | (P3[13] & C3[13]);
    assign c3     = G3[14] | (P3[14] & C3[14]);
    assign s301   = P3[0];
    assign s302   = P3[1]  ^ C3[1];
    assign s303   = P3[2]  ^ C3[2];
    assign s304   = P3[3]  ^ C3[3];
    assign s305   = P3[4]  ^ C3[4];
    assign s306   = P3[5]  ^ C3[5];
    assign s307   = P3[6]  ^ C3[6];
    assign s308   = P3[7]  ^ C3[7];
    assign s309   = P3[8]  ^ C3[8];
    assign s310   = P3[9]  ^ C3[9];
    assign s311   = P3[10] ^ C3[10];
    assign s312   = P3[11] ^ C3[11];
    assign s313   = P3[12] ^ C3[12];
    assign s314   = P3[13] ^ C3[13];
    assign s315   = P3[14] ^ C3[14];

     /* 4th CLA */
    wire [14:0] G4, P4, C4;
    assign G4[0]  = pp6[1]  & pp7[0];
    assign G4[1]  = pp6[2]  & pp7[1];
    assign G4[2]  = pp6[3]  & pp7[2];
    assign G4[3]  = pp6[4]  & pp7[3];
    assign G4[4]  = pp6[5]  & pp7[4];
    assign G4[5]  = pp6[6]  & pp7[5];
    assign G4[6]  = pp6[7]  & pp7[6];
    assign G4[7]  = pp6[8]  & pp7[7];
    assign G4[8]  = pp6[9]  & pp7[8];
    assign G4[9]  = pp6[10] & pp7[9];
    assign G4[10] = pp6[11] & pp7[10];
    assign G4[11] = pp6[12] & pp7[11];
    assign G4[12] = pp6[13] & pp7[12];
    assign G4[13] = pp6[14] & pp7[13];
    assign G4[14] = pp6[15] & pp7[14];
    assign P4[0]  = pp6[1]  ^ pp7[0];
    assign P4[1]  = pp6[2]  ^ pp7[1];
    assign P4[2]  = pp6[3]  ^ pp7[2];
    assign P4[3]  = pp6[4]  ^ pp7[3];
    assign P4[4]  = pp6[5]  ^ pp7[4];
    assign P4[5]  = pp6[6]  ^ pp7[5];
    assign P4[6]  = pp6[7]  ^ pp7[6];
    assign P4[7]  = pp6[8]  ^ pp7[7];
    assign P4[8]  = pp6[9]  ^ pp7[8];
    assign P4[9]  = pp6[10] ^ pp7[9];
    assign P4[10] = pp6[11] ^ pp7[10];
    assign P4[11] = pp6[12] ^ pp7[11];
    assign P4[12] = pp6[13] ^ pp7[12];
    assign P4[13] = pp6[14] ^ pp7[13];
    assign P4[14] = pp6[15] ^ pp7[14];
    assign C4[0]  = 0;
    assign C4[1]  = G4[0]  | (P4[0] & C4[0]);
    assign C4[2]  = G4[1]  | (P4[1] & C4[1]);
    assign C4[3]  = G4[2]  | (P4[2] & C4[2]);
    assign C4[4]  = G4[3]  | (P4[3] & C4[3]);
    assign C4[5]  = G4[4]  | (P4[4] & C4[4]);
    assign C4[6]  = G4[5]  | (P4[5] & C4[5]);
    assign C4[7]  = G4[6]  | (P4[6] & C4[6]);
    assign C4[8]  = G4[7]  | (P4[7] & C4[7]);
    assign C4[9]  = G4[8]  | (P4[8] & C4[8]);
    assign C4[10] = G4[9]  | (P4[9] & C4[9]);
    assign C4[11] = G4[10] | (P4[10] & C4[10]);
    assign C4[12] = G4[11] | (P4[11] & C4[11]);
    assign C4[13] = G4[12] | (P4[12] & C4[12]);
    assign C4[14] = G4[13] | (P4[13] & C4[13]);
    assign c4     = G4[14] | (P4[14] & C4[14]);
    assign s401   = P4[0];
    assign s402   = P4[1]  ^ C4[1];
    assign s403   = P4[2]  ^ C4[2];
    assign s404   = P4[3]  ^ C4[3];
    assign s405   = P4[4]  ^ C4[4];
    assign s406   = P4[5]  ^ C4[5];
    assign s407   = P4[6]  ^ C4[6];
    assign s408   = P4[7]  ^ C4[7];
    assign s409   = P4[8]  ^ C4[8];
    assign s410   = P4[9]  ^ C4[9];
    assign s411   = P4[10] ^ C4[10];
    assign s412   = P4[11] ^ C4[11];
    assign s413   = P4[12] ^ C4[12];
    assign s414   = P4[13] ^ C4[13];
    assign s415   = P4[14] ^ C4[14];

     /* 5th CLA */
    wire [14:0] G5, P5, C5;
    assign G5[0]  = pp8[1]  & pp9[0];
    assign G5[1]  = pp8[2]  & pp9[1];
    assign G5[2]  = pp8[3]  & pp9[2];
    assign G5[3]  = pp8[4]  & pp9[3];
    assign G5[4]  = pp8[5]  & pp9[4];
    assign G5[5]  = pp8[6]  & pp9[5];
    assign G5[6]  = pp8[7]  & pp9[6];
    assign G5[7]  = pp8[8]  & pp9[7];
    assign G5[8]  = pp8[9]  & pp9[8];
    assign G5[9]  = pp8[10] & pp9[9];
    assign G5[10] = pp8[11] & pp9[10];
    assign G5[11] = pp8[12] & pp9[11];
    assign G5[12] = pp8[13] & pp9[12];
    assign G5[13] = pp8[14] & pp9[13];
    assign G5[14] = pp8[15] & pp9[14];
    assign P5[0]  = pp8[1]  ^ pp9[0];
    assign P5[1]  = pp8[2]  ^ pp9[1];
    assign P5[2]  = pp8[3]  ^ pp9[2];
    assign P5[3]  = pp8[4]  ^ pp9[3];
    assign P5[4]  = pp8[5]  ^ pp9[4];
    assign P5[5]  = pp8[6]  ^ pp9[5];
    assign P5[6]  = pp8[7]  ^ pp9[6];
    assign P5[7]  = pp8[8]  ^ pp9[7];
    assign P5[8]  = pp8[9]  ^ pp9[8];
    assign P5[9]  = pp8[10] ^ pp9[9];
    assign P5[10] = pp8[11] ^ pp9[10];
    assign P5[11] = pp8[12] ^ pp9[11];
    assign P5[12] = pp8[13] ^ pp9[12];
    assign P5[13] = pp8[14] ^ pp9[13];
    assign P5[14] = pp8[15] ^ pp9[14];
    assign C5[0] = 0;
    assign C5[1]  = G5[0]  | (P5[0]  & C5[0]);
    assign C5[2]  = G5[1]  | (P5[1]  & C5[1]);
    assign C5[3]  = G5[2]  | (P5[2]  & C5[2]);
    assign C5[4]  = G5[3]  | (P5[3]  & C5[3]);
    assign C5[5]  = G5[4]  | (P5[4]  & C5[4]);
    assign C5[6]  = G5[5]  | (P5[5]  & C5[5]);
    assign C5[7]  = G5[6]  | (P5[6]  & C5[6]);
    assign C5[8]  = G5[7]  | (P5[7]  & C5[7]);
    assign C5[9]  = G5[8]  | (P5[8]  & C5[8]);
    assign C5[10] = G5[9]  | (P5[9]  & C5[9]);
    assign C5[11] = G5[10] | (P5[10] & C5[10]);
    assign C5[12] = G5[11] | (P5[11] & C5[11]);
    assign C5[13] = G5[12] | (P5[12] & C5[12]);
    assign C5[14] = G5[13] | (P5[13] & C5[13]);
    assign c5     = G5[14] | (P5[14] & C5[14]);
    assign s501   = P5[0];
    assign s502   = P5[1]  ^ C5[1];
    assign s503   = P5[2]  ^ C5[2];
    assign s504   = P5[3]  ^ C5[3];
    assign s505   = P5[4]  ^ C5[4];
    assign s506   = P5[5]  ^ C5[5];
    assign s507   = P5[6]  ^ C5[6];
    assign s508   = P5[7]  ^ C5[7];
    assign s509   = P5[8]  ^ C5[8];
    assign s510   = P5[9]  ^ C5[9];
    assign s511   = P5[10] ^ C5[10];
    assign s512   = P5[11] ^ C5[11];
    assign s513   = P5[12] ^ C5[12];
    assign s514   = P5[13] ^ C5[13];
    assign s515   = P5[14] ^ C5[14];


     /* 6th CLA */
    wire [11:0] G6, P6, C6;
    assign G6[0]  = pp10[1]  & pp11[0];
    assign G6[1]  = pp10[2]  & pp11[1];
    assign G6[2]  = pp10[3]  & pp11[2];
    assign G6[3]  = pp10[4]  & pp11[3];
    assign G6[4]  = pp10[5]  & pp11[4];
    assign G6[5]  = pp10[6]  & pp11[5];
    assign G6[6]  = pp10[7]  & pp11[6];
    assign G6[7]  = pp10[8]  & pp11[7];
    assign G6[8]  = pp10[9]  & pp11[8];
    assign G6[9]  = pp10[10] & pp11[9];
    assign G6[10] = pp10[11] & pp11[10];
    assign G6[11] = pp10[12] & pp11[11];
    assign P6[0]  = pp10[1]  ^ pp11[0];
    assign P6[1]  = pp10[2]  ^ pp11[1];
    assign P6[2]  = pp10[3]  ^ pp11[2];
    assign P6[3]  = pp10[4]  ^ pp11[3];
    assign P6[4]  = pp10[5]  ^ pp11[4];
    assign P6[5]  = pp10[6]  ^ pp11[5];
    assign P6[6]  = pp10[7]  ^ pp11[6];
    assign P6[7]  = pp10[8]  ^ pp11[7];
    assign P6[8]  = pp10[9]  ^ pp11[8];
    assign P6[9]  = pp10[10] ^ pp11[9];
    assign P6[10] = pp10[11] ^ pp11[10];
    assign P6[11] = pp10[12] ^ pp11[11];
    assign C6[0]  = 0;
    assign C6[1]  = G6[0]  | (P6[0] & C6[0]);
    assign C6[2]  = G6[1]  | (P6[1] & C6[1]);
    assign C6[3]  = G6[2]  | (P6[2] & C6[2]);
    assign C6[4]  = G6[3]  | (P6[3] & C6[3]);
    assign C6[5]  = G6[4]  | (P6[4] & C6[4]);
    assign C6[6]  = G6[5]  | (P6[5] & C6[5]);
    assign C6[7]  = G6[6]  | (P6[6] & C6[6]);
    assign C6[8]  = G6[7]  | (P6[7] & C6[7]);
    assign C6[9]  = G6[8]  | (P6[8] & C6[8]);
    assign C6[10] = G6[9]  | (P6[9] & C6[9]);
    assign C6[11] = G6[10] | (P6[10] & C6[10]);
    assign c6     = G6[11] | (P6[11] & C6[11]);
    assign s601   = P6[0];
    assign s602   = P6[1]  ^ C6[1];
    assign s603   = P6[2]  ^ C6[2];
    assign s604   = P6[3]  ^ C6[3];
    assign s605   = P6[4]  ^ C6[4];
    assign s606   = P6[5]  ^ C6[5];
    assign s607   = P6[6]  ^ C6[6];
    assign s608   = P6[7]  ^ C6[7];
    assign s609   = P6[8]  ^ C6[8];
    assign s610   = P6[9]  ^ C6[9];
    assign s611   = P6[10] ^ C6[10];
    assign s612   = P6[11] ^ C6[11];
 
    /* 7th CLA */
    wire [7:0] G7, P7, C7;
    assign G7[0]  = pp12[1]  & pp13[0];
    assign G7[1]  = pp12[2]  & pp13[1];
    assign G7[2]  = pp12[3]  & pp13[2];
    assign G7[3]  = pp12[4]  & pp13[3];
    assign G7[4]  = pp12[5]  & pp13[4];
    assign G7[5]  = pp12[6]  & pp13[5];
    assign G7[6]  = pp12[7]  & pp13[6];
    assign G7[7]  = pp12[8]  & pp13[7];
    assign P7[0]  = pp12[1]  ^ pp13[0];
    assign P7[1]  = pp12[2]  ^ pp13[1];
    assign P7[2]  = pp12[3]  ^ pp13[2];
    assign P7[3]  = pp12[4]  ^ pp13[3];
    assign P7[4]  = pp12[5]  ^ pp13[4];
    assign P7[5]  = pp12[6]  ^ pp13[5];
    assign P7[6]  = pp12[7]  ^ pp13[6];
    assign P7[7]  = pp12[8]  ^ pp13[7];
    assign C7[0]  = 0;
    assign C7[1] = G7[0] | (P7[0] & C7[0]);
    assign C7[2] = G7[1] | (P7[1] & C7[1]);
    assign C7[3] = G7[2] | (P7[2] & C7[2]);
    assign C7[4] = G7[3] | (P7[3] & C7[3]);
    assign C7[5] = G7[4] | (P7[4] & C7[4]);
    assign C7[6] = G7[5] | (P7[5] & C7[5]);
    assign C7[7] = G7[6] | (P7[6] & C7[6]);
    assign c7    = G7[7] | (P7[7] & C7[7]);
    assign s701  = P7[0];
    assign s702  = P7[1]  ^ C7[1];
    assign s703  = P7[2]  ^ C7[2];
    assign s704  = P7[3]  ^ C7[3];
    assign s705  = P7[4]  ^ C7[4];
    assign s706  = P7[5]  ^ C7[5];
    assign s707  = P7[6]  ^ C7[6];
    assign s708  = P7[7]  ^ C7[7];

    /* 8th CLA */
    wire [3:0] G8, P8, C8;
    assign G8[0]  = pp14[1]  & pp15[0];
    assign G8[1]  = pp14[2]  & pp15[1];
    assign G8[2]  = pp14[3]  & pp15[2];
    assign G8[3]  = pp14[4]  & pp15[3];
    assign P8[0]  = pp14[1]  ^ pp15[0];
    assign P8[1]  = pp14[2]  ^ pp15[1];
    assign P8[2]  = pp14[3]  ^ pp15[2];
    assign P8[3]  = pp14[4]  ^ pp15[3];
    assign C8[0]  = 0;
    assign C8[1]  = G8[0] | (P8[0] & C8[0]);
    assign C8[2]  = G8[1] | (P8[1] & C8[1]);
    assign C8[3]  = G8[2] | (P8[2] & C8[2]);
    assign c8     = G8[3] | (P8[3] & C8[3]);
    assign s801   = P8[0];
    assign s802   = P8[1]  ^ C8[1];
    assign s803   = P8[2]  ^ C8[2];
    assign s804   = P8[3]  ^ C8[3];

    /* 9th CLA */
    wire [19:0] G9, P9, C9;
    assign G9[0]  = s108     & s206;
    assign G9[1]  = s109     & s207;
    assign G9[2]  = s110     & s208;
    assign G9[3]  = s111     & s209;
    assign G9[4]  = s112     & s210;
    assign G9[5]  = s113     & s211;
    assign G9[6]  = s114     & s212;
    assign G9[7]  = s115     & s213;
    assign G9[8]  = s116     & s214;
    assign G9[9]  = c1       & s215;
    assign G9[10] = c2       & pp3[15];
    assign G9[11] = pp14[5]  & pp15[4];
    assign G9[12] = pp14[6]  & pp15[5];
    assign G9[13] = pp14[7]  & pp15[6];
    assign G9[14] = pp14[8]  & pp15[7];
    assign G9[15] = pp14[9]  & pp15[8];
    assign G9[16] = pp14[10] & pp15[9];
    assign G9[17] = pp14[11] & pp15[10];
    assign G9[18] = pp14[12] & pp15[11];
    assign G9[19] = pp14[13] & pp15[12];
    assign P9[0]  = s108     ^ s206;
    assign P9[1]  = s109     ^ s207;
    assign P9[2]  = s110     ^ s208;
    assign P9[3]  = s111     ^ s209;
    assign P9[4]  = s112     ^ s210;
    assign P9[5]  = s113     ^ s211;
    assign P9[6]  = s114     ^ s212;
    assign P9[7]  = s115     ^ s213;
    assign P9[8]  = s116     ^ s214;
    assign P9[9]  = c1       ^ s215;
    assign P9[10] = c2       ^ pp3[15];
    assign P9[11] = pp14[5]  ^ pp15[4];
    assign P9[12] = pp14[6]  ^ pp15[5];
    assign P9[13] = pp14[7]  ^ pp15[6];
    assign P9[14] = pp14[8]  ^ pp15[7];
    assign P9[15] = pp14[9]  ^ pp15[8];
    assign P9[16] = pp14[10] ^ pp15[9];
    assign P9[17] = pp14[11] ^ pp15[10];
    assign P9[18] = pp14[12] ^ pp15[11];
    assign P9[19] = pp14[13] ^ pp15[12];
    assign C9[0]  = 0;
    assign C9[1]  = G9[0]  | (P9[0] & C9[0]);
    assign C9[2]  = G9[1]  | (P9[1] & C9[1]);
    assign C9[3]  = G9[2]  | (P9[2] & C9[2]);
    assign C9[4]  = G9[3]  | (P9[3] & C9[3]);
    assign C9[5]  = G9[4]  | (P9[4] & C9[4]);
    assign C9[6]  = G9[5]  | (P9[5] & C9[5]);
    assign C9[7]  = G9[6]  | (P9[6] & C9[6]);
    assign C9[8]  = G9[7]  | (P9[7] & C9[7]);
    assign C9[9]  = G9[8]  | (P9[8] & C9[8]);
    assign C9[10] = G9[9]  | (P9[9] & C9[9]);
    assign C9[11] = G9[10] | (P9[10] & C9[10]);
    assign C9[12] = G9[11] | (P9[11] & C9[11]);
    assign C9[13] = G9[12] | (P9[12] & C9[12]);
    assign C9[14] = G9[13] | (P9[13] & C9[13]);
    assign C9[15] = G9[14] | (P9[14] & C9[14]);
    assign C9[16] = G9[15] | (P9[15] & C9[15]);
    assign C9[17] = G9[16] | (P9[16] & C9[16]);
    assign C9[18] = G9[17] | (P9[17] & C9[17]);
    assign C9[19] = G9[18] | (P9[18] & C9[18]);
    assign c9    = G9[19]  | (P9[19] & C9[19]);
    assign s901  = P9[0];
    assign s902  = P9[1]  ^ C9[1];
    assign s903  = P9[2]  ^ C9[2];
    assign s904  = P9[3]  ^ C9[3];
    assign s905  = P9[4]  ^ C9[4];
    assign s906  = P9[5]  ^ C9[5];
    assign s907  = P9[6]  ^ C9[6];
    assign s908  = P9[7]  ^ C9[7];
    assign s909  = P9[8]  ^ C9[8];
    assign s910  = P9[9]  ^ C9[9];
    assign s911  = P9[10] ^ C9[10];
    assign s912  = P9[11] ^ C9[11];
    assign s913  = P9[12] ^ C9[12];
    assign s914  = P9[13] ^ C9[13];
    assign s915  = P9[14] ^ C9[14];
    assign s916  = P9[15] ^ C9[15];
    assign s917  = P9[16] ^ C9[16];
    assign s918  = P9[17] ^ C9[17];
    assign s919  = P9[18] ^ C9[18];
    assign s920  = P9[19] ^ C9[19];

    /* 10th CLA */ 
    wire [16:0] GA, PA, CA;
    assign GA[0]   = s306     & s404;
    assign GA[1]   = s307     & s405;
    assign GA[2]   = s308     & s406;
    assign GA[3]   = s309     & s407;
    assign GA[4]   = s310     & s408;
    assign GA[5]   = s311     & s409;
    assign GA[6]   = s312     & s410;
    assign GA[7]   = s313     & s411;
    assign GA[8]   = s314     & s412;
    assign GA[9]   = s315     & s413;
    assign GA[10]  = c3       & s414;
    assign GA[11]  = c7       & s415;
    assign GA[12]  = pp7[15]  & c4;
    assign GA[13]  = pp12[11] & pp13[10];
    assign GA[14]  = pp12[12] & pp13[11];
    assign GA[15]  = pp12[13] & pp13[12];
    assign GA[16]  = pp12[14] & pp13[13];
    assign PA[0]   = s306     ^ s404;
    assign PA[1]   = s307     ^ s405;
    assign PA[2]   = s308     ^ s406;
    assign PA[3]   = s309     ^ s407;
    assign PA[4]   = s310     ^ s408;
    assign PA[5]   = s311     ^ s409;
    assign PA[6]   = s312     ^ s410;
    assign PA[7]   = s313     ^ s411;
    assign PA[8]   = s314     ^ s412;
    assign PA[9]   = s315     ^ s413;
    assign PA[10]  = c3       ^ s414;
    assign PA[11]  = c7       ^ s415;
    assign PA[12]  = pp7[15]  ^ c4;
    assign PA[13]  = pp12[11] ^ pp13[10];
    assign PA[14]  = pp12[12] ^ pp13[11];
    assign PA[15]  = pp12[13] ^ pp13[12];
    assign PA[16]  = pp12[14] ^ pp13[13];
    assign CA[0]  = 0;
    assign CA[1]  = GA[0]  | (PA[0] & CA[0]);
    assign CA[2]  = GA[1]  | (PA[1] & CA[1]);
    assign CA[3]  = GA[2]  | (PA[2] & CA[2]);
    assign CA[4]  = GA[3]  | (PA[3] & CA[3]);
    assign CA[5]  = GA[4]  | (PA[4] & CA[4]);
    assign CA[6]  = GA[5]  | (PA[5] & CA[5]);
    assign CA[7]  = GA[6]  | (PA[6] & CA[6]);
    assign CA[8]  = GA[7]  | (PA[7] & CA[7]);
    assign CA[9]  = GA[8]  | (PA[8] & CA[8]);
    assign CA[10] = GA[9]  | (PA[9] & CA[9]);
    assign CA[11] = GA[10] | (PA[10] & CA[10]);
    assign CA[12] = GA[11] | (PA[11] & CA[11]);
    assign CA[13] = GA[12] | (PA[12] & CA[12]);
    assign CA[14] = GA[13] | (PA[13] & CA[13]);
    assign CA[15] = GA[14] | (PA[14] & CA[14]);
    assign CA[16] = GA[15] | (PA[15] & CA[15]);
    assign c10    = GA[16] | (PA[16] & CA[16]);
    assign sA01   = PA[0];
    assign sA02   = PA[1]  ^ CA[1];
    assign sA03   = PA[2]  ^ CA[2];
    assign sA04   = PA[3]  ^ CA[3];
    assign sA05   = PA[4]  ^ CA[4];
    assign sA06   = PA[5]  ^ CA[5];
    assign sA07   = PA[6]  ^ CA[6];
    assign sA08   = PA[7]  ^ CA[7];
    assign sA09   = PA[8]  ^ CA[8];
    assign sA10   = PA[9]  ^ CA[9];
    assign sA11   = PA[10] ^ CA[10];
    assign sA12   = PA[11] ^ CA[11];
    assign sA13   = PA[12] ^ CA[12];
    assign sA14   = PA[13] ^ CA[13];
    assign sA15   = PA[14] ^ CA[14];
    assign sA16   = PA[15] ^ CA[15];
    assign sA17   = PA[16] ^ CA[16];

    /* 11th CLA */
    wire [13:0] GB, PB, CB;
    assign GB[0]  = s504     & s602;
    assign GB[1]  = s505     & s603;
    assign GB[2]  = s506     & s604;
    assign GB[3]  = s507     & s605;
    assign GB[4]  = s508     & s606;
    assign GB[5]  = s509     & s607;
    assign GB[6]  = s510     & s608;
    assign GB[7]  = s511     & s609;
    assign GB[8]  = s512     & s610;
    assign GB[9]  = s513     & s611;
    assign GB[10] = s514     & s612;
    assign GB[11] = s515     & c6;
    assign GB[12] = pp9[15]  & c5;
    assign GB[13] = pp10[15] & pp11[14];
    assign PB[0]  = s504     ^ s602;
    assign PB[1]  = s505     ^ s603;
    assign PB[2]  = s506     ^ s604;
    assign PB[3]  = s507     ^ s605;
    assign PB[4]  = s508     ^ s606;
    assign PB[5]  = s509     ^ s607;
    assign PB[6]  = s510     ^ s608;
    assign PB[7]  = s511     ^ s609;
    assign PB[8]  = s512     ^ s610;
    assign PB[9]  = s513     ^ s611;
    assign PB[10] = s514     ^ s612;
    assign PB[11] = s515     ^ c6;
    assign PB[12] = pp9[15]  ^ c5;
    assign PB[13] = pp10[15] ^ pp11[14];
    assign CB[0]  = 0;
    assign CB[1]  = GB[0]  | (PB[0] & CB[0]);
    assign CB[2]  = GB[1]  | (PB[1] & CB[1]);
    assign CB[3]  = GB[2]  | (PB[2] & CB[2]);
    assign CB[4]  = GB[3]  | (PB[3] & CB[3]);
    assign CB[5]  = GB[4]  | (PB[4] & CB[4]);
    assign CB[6]  = GB[5]  | (PB[5] & CB[5]);
    assign CB[7]  = GB[6]  | (PB[6] & CB[6]);
    assign CB[8]  = GB[7]  | (PB[7] & CB[7]);
    assign CB[9]  = GB[8]  | (PB[8] & CB[8]);
    assign CB[10] = GB[9]  | (PB[9] & CB[9]);
    assign CB[11] = GB[10] | (PB[10] & CB[10]);
    assign CB[12] = GB[11] | (PB[11] & CB[11]);
    assign CB[13] = GB[12] | (PB[12] & CB[12]);
    assign c11    = GB[13] | (PB[13] & CB[13]);
    assign sB01   = PB[0];
    assign sB02   = PB[1]  ^ CB[1];
    assign sB03   = PB[2]  ^ CB[2];
    assign sB04   = PB[3]  ^ CB[3];
    assign sB05   = PB[4]  ^ CB[4];
    assign sB06   = PB[5]  ^ CB[5];
    assign sB07   = PB[6]  ^ CB[6];
    assign sB08   = PB[7]  ^ CB[7];
    assign sB09   = PB[8]  ^ CB[8];
    assign sB10   = PB[9]  ^ CB[9];
    assign sB11   = PB[10] ^ CB[10];
    assign sB12   = PB[11] ^ CB[11];
    assign sB13   = PB[12] ^ CB[12];
    assign sB14   = PB[13] ^ CB[13];

    /* 12th CLA */
    wire [10:0] GC, PC, CC;
    assign GC[0]  = s702     & pp15[0];
    assign GC[1]  = s703     & s801;
    assign GC[2]  = s704     & s802;
    assign GC[3]  = s705     & s803;
    assign GC[4]  = s706     & s804;
    assign GC[5]  = s707     & c8;
    assign GC[6]  = s708     & pp5[15];
    assign GC[7]  = pp12[9]  & pp13[8];
    assign GC[8]  = pp12[10] & pp13[9];
    assign GC[9]  = pp10[13] & pp11[12];
    assign GC[10] = pp10[14] & pp11[13];
    assign PC[0]  = s702     ^ pp15[0];
    assign PC[1]  = s703     ^ s801;
    assign PC[2]  = s704     ^ s802;
    assign PC[3]  = s705     ^ s803;
    assign PC[4]  = s706     ^ s804;
    assign PC[5]  = s707     ^ c8;
    assign PC[6]  = s708     ^ pp5[15];
    assign PC[7]  = pp12[9]  ^ pp13[8];
    assign PC[8]  = pp12[10] ^ pp13[9];
    assign PC[9]  = pp10[13] ^ pp11[12];
    assign PC[10] = pp10[14] ^ pp11[13];
    assign CC[0] = 0;
    assign CC[1]  = GC[0] | (PC[0]  & CC[0]);
    assign CC[2]  = GC[1] | (PC[1]  & CC[1]);
    assign CC[3]  = GC[2] | (PC[2]  & CC[2]);
    assign CC[4]  = GC[3] | (PC[3]  & CC[3]);
    assign CC[5]  = GC[4] | (PC[4]  & CC[4]);
    assign CC[6]  = GC[5] | (PC[5]  & CC[5]);
    assign CC[7]  = GC[6] | (PC[6]  & CC[6]);
    assign CC[8]  = GC[7] | (PC[7]  & CC[7]);
    assign CC[9]  = GC[8] | (PC[8]  & CC[8]);
    assign CC[10] = GC[9] | (PC[9]  & CC[9]);
    assign c12   = GC[10] | (PC[10] & CC[10]);
    assign sC01  = PC[0];
    assign sC02  = PC[1]  ^ CC[1];
    assign sC03  = PC[2]  ^ CC[2];
    assign sC04  = PC[3]  ^ CC[3];
    assign sC05  = PC[4]  ^ CC[4];
    assign sC06  = PC[5]  ^ CC[5];
    assign sC07  = PC[6]  ^ CC[6];
    assign sC08  = PC[7]  ^ CC[7];
    assign sC09  = PC[8]  ^ CC[8];
    assign sC10  = PC[9]  ^ CC[9];
    assign sC11  = PC[10] ^ CC[10];

    /* 13th CLA */
    wire [25:0] GD, PD, CD;
    assign GD[0]  = s104     & s202;
    assign GD[1]  = s105     & s203;
    assign GD[2]  = s106     & s204;
    assign GD[3]  = s107     & s205;
    assign GD[4]  = s901     & s304; 
    assign GD[5]  = s902     & s305;
    assign GD[6]  = s903     & sA01;
    assign GD[7]  = s904     & sA02;
    assign GD[8]  = s905     & sA03;
    assign GD[9]  = s906     & sA04;
    assign GD[10] = s907     & sA05;
    assign GD[11] = s908     & sA06;
    assign GD[12] = s909     & sA07;
    assign GD[13] = s910     & sA08;
    assign GD[14] = s911     & sA09;
    assign GD[15] = s912     & sA10;
    assign GD[16] = s913     & sA11;
    assign GD[17] = s914     & sA12;
    assign GD[18] = s915     & sA13;
    assign GD[19] = s916     & sA14;
    assign GD[20] = s917     & sA15;
    assign GD[21] = s918     & sA16;
    assign GD[22] = s919     & sA17;
    assign GD[23] = s920     & c10;
    assign GD[24] = c9       & pp13[15];
    assign GD[25] = pp14[15] & pp15[14];
    assign PD[0]  = s104     ^ s202;
    assign PD[1]  = s105     ^ s203;
    assign PD[2]  = s106     ^ s204;
    assign PD[3]  = s107     ^ s205;
    assign PD[4]  = s901     ^ s304;
    assign PD[5]  = s902     ^ s305;
    assign PD[6]  = s903     ^ sA01;
    assign PD[7]  = s904     ^ sA02;
    assign PD[8]  = s905     ^ sA03;
    assign PD[9]  = s906     ^ sA04;
    assign PD[10] = s907     ^ sA05;
    assign PD[11] = s908     ^ sA06;
    assign PD[12] = s909     ^ sA07;
    assign PD[13] = s910     ^ sA08;
    assign PD[14] = s911     ^ sA09;
    assign PD[15] = s912     ^ sA10;
    assign PD[16] = s913     ^ sA11;
    assign PD[17] = s914     ^ sA12;
    assign PD[18] = s915     ^ sA13;
    assign PD[19] = s916     ^ sA14;
    assign PD[20] = s917     ^ sA15;
    assign PD[21] = s918     ^ sA16;
    assign PD[22] = s919     ^ sA17;
    assign PD[23] = s920     ^ c10;
    assign PD[24] = c9       ^ pp13[15];
    assign PD[25] = pp14[15] ^ pp15[14];
    assign CD[0]  = 0;
    assign CD[1]  = GD[0]  | (PD[0]  & CD[0]);
    assign CD[2]  = GD[1]  | (PD[1]  & CD[1]);
    assign CD[3]  = GD[2]  | (PD[2]  & CD[2]);
    assign CD[4]  = GD[3]  | (PD[3]  & CD[3]);
    assign CD[5]  = GD[4]  | (PD[4]  & CD[4]);
    assign CD[6]  = GD[5]  | (PD[5]  & CD[5]);
    assign CD[7]  = GD[6]  | (PD[6]  & CD[6]);
    assign CD[8]  = GD[7]  | (PD[7]  & CD[7]);
    assign CD[9]  = GD[8]  | (PD[8]  & CD[8]);
    assign CD[10] = GD[9]  | (PD[9]  & CD[9]);
    assign CD[11] = GD[10] | (PD[10] & CD[10]);
    assign CD[12] = GD[11] | (PD[11] & CD[11]);
    assign CD[13] = GD[12] | (PD[12] & CD[12]);
    assign CD[14] = GD[13] | (PD[13] & CD[13]);
    assign CD[15] = GD[14] | (PD[14] & CD[14]);
    assign CD[16] = GD[15] | (PD[15] & CD[15]);
    assign CD[17] = GD[16] | (PD[16] & CD[16]);
    assign CD[18] = GD[17] | (PD[17] & CD[17]);
    assign CD[19] = GD[18] | (PD[18] & CD[18]);
    assign CD[20] = GD[19] | (PD[19] & CD[19]);
    assign CD[21] = GD[20] | (PD[20] & CD[20]);
    assign CD[22] = GD[21] | (PD[21] & CD[21]);
    assign CD[23] = GD[22] | (PD[22] & CD[22]);
    assign CD[24] = GD[23] | (PD[23] & CD[23]);
    assign CD[25] = GD[24] | (PD[24] & CD[24]);
    assign c13    = GD[25] | (PD[25] & CD[25]);
    assign sD01   = PD[0];
    assign sD02   = PD[1]  ^ CD[1];
    assign sD03   = PD[2]  ^ CD[2];
    assign sD04   = PD[3]  ^ CD[3];
    assign sD05   = PD[4]  ^ CD[4];
    assign sD06   = PD[5]  ^ CD[5];
    assign sD07   = PD[6]  ^ CD[6];
    assign sD08   = PD[7]  ^ CD[7];
    assign sD09   = PD[8]  ^ CD[8];
    assign sD10   = PD[9]  ^ CD[9];
    assign sD11   = PD[10] ^ CD[10];
    assign sD12   = PD[11] ^ CD[11];
    assign sD13   = PD[12] ^ CD[12];
    assign sD14   = PD[13] ^ CD[13];
    assign sD15   = PD[14] ^ CD[14];
    assign sD16   = PD[15] ^ CD[15];
    assign sD17   = PD[16] ^ CD[16];
    assign sD18   = PD[17] ^ CD[17];
    assign sD19   = PD[18] ^ CD[18];
    assign sD20   = PD[19] ^ CD[19];
    assign sD21   = PD[20] ^ CD[20];
    assign sD22   = PD[21] ^ CD[21];
    assign sD23   = PD[22] ^ CD[22];
    assign sD24   = PD[23] ^ CD[23];
    assign sD25   = PD[24] ^ CD[24];
    assign sD26   = PD[25] ^ CD[25];

    /* 14th CLA */
    wire [22:0] GE, PE, CE;
    assign GE[0]  = s302     & pp6[0];
    assign GE[1]  = s303     & s401;
    assign GE[2]  = s402     & pp8[0];
    assign GE[3]  = s403     & s501;
    assign GE[4]  = s502     & pp10[0];
    assign GE[5]  = s503     & s601;
    assign GE[6]  = sB01     & pp12[0];
    assign GE[7]  = sB02     & s701;
    assign GE[8]  = sB03     & sC01;
    assign GE[9]  = sB04     & sC02;
    assign GE[10] = sB05     & sC03;
    assign GE[11] = sB06     & sC04;
    assign GE[12] = sB07     & sC05;
    assign GE[13] = sB08     & sC06;
    assign GE[14] = sB09     & sC07;
    assign GE[15] = sB10     & sC08;
    assign GE[16] = sB11     & sC09;
    assign GE[17] = sB12     & sC10;
    assign GE[18] = sB13     & sC11;
    assign GE[19] = sB14     & c12;
    assign GE[20] = c11      & pp11[15];
    assign GE[21] = pp12[15] & pp13[14];
    assign GE[22] = pp14[14] & pp15[13];
    assign PE[0]  = s302     ^ pp6[0];
    assign PE[1]  = s303     ^ s401;
    assign PE[2]  = s402     ^ pp8[0];
    assign PE[3]  = s403     ^ s501;
    assign PE[4]  = s502     ^ pp10[0];
    assign PE[5]  = s503     ^ s601;
    assign PE[6]  = sB01     ^ pp12[0];
    assign PE[7]  = sB02     ^ s701;
    assign PE[8]  = sB03     ^ sC01;
    assign PE[9]  = sB04     ^ sC02;
    assign PE[10] = sB05     ^ sC03;
    assign PE[11] = sB06     ^ sC04;
    assign PE[12] = sB07     ^ sC05;
    assign PE[13] = sB08     ^ sC06;
    assign PE[14] = sB09     ^ sC07;
    assign PE[15] = sB10     ^ sC08;
    assign PE[16] = sB11     ^ sC09;
    assign PE[17] = sB12     ^ sC10;
    assign PE[18] = sB13     ^ sC11;
    assign PE[19] = sB14     ^ c12;
    assign PE[20] = c11      ^ pp11[15];
    assign PE[21] = pp12[15] ^ pp13[14];
    assign PE[22] = pp14[14] ^ pp15[13];
    assign CE[0]  = 0;
    assign CE[1]  = GE[0]  | (PE[0]  & CE[0]);
    assign CE[2]  = GE[1]  | (PE[1]  & CE[1]);
    assign CE[3]  = GE[2]  | (PE[2]  & CE[2]);
    assign CE[4]  = GE[3]  | (PE[3]  & CE[3]);
    assign CE[5]  = GE[4]  | (PE[4]  & CE[4]);
    assign CE[6]  = GE[5]  | (PE[5]  & CE[5]);
    assign CE[7]  = GE[6]  | (PE[6]  & CE[6]);
    assign CE[8]  = GE[7]  | (PE[7]  & CE[7]);
    assign CE[9]  = GE[8]  | (PE[8]  & CE[8]);
    assign CE[10] = GE[9]  | (PE[9]  & CE[9]);
    assign CE[11] = GE[10] | (PE[10] & CE[10]);
    assign CE[12] = GE[11] | (PE[11] & CE[11]);
    assign CE[13] = GE[12] | (PE[12] & CE[12]);
    assign CE[14] = GE[13] | (PE[13] & CE[13]);
    assign CE[15] = GE[14] | (PE[14] & CE[14]);
    assign CE[16] = GE[15] | (PE[15] & CE[15]);
    assign CE[17] = GE[16] | (PE[16] & CE[16]);
    assign CE[18] = GE[17] | (PE[17] & CE[17]);
    assign CE[19] = GE[18] | (PE[18] & CE[18]);
    assign CE[20] = GE[19] | (PE[19] & CE[19]);
    assign CE[21] = GE[20] | (PE[20] & CE[20]);
    assign CE[22] = GE[21] | (PE[21] & CE[21]);
    assign c14    = GE[22] | (PE[22] & CE[22]);
    assign sE01   = PE[0];
    assign sE02   = PE[1]  ^ CE[1];
    assign sE03   = PE[2]  ^ CE[2];
    assign sE04   = PE[3]  ^ CE[3];
    assign sE05   = PE[4]  ^ CE[4];
    assign sE06   = PE[5]  ^ CE[5];
    assign sE07   = PE[6]  ^ CE[6];
    assign sE08   = PE[7]  ^ CE[7];
    assign sE09   = PE[8]  ^ CE[8];
    assign sE10   = PE[9]  ^ CE[9];
    assign sE11   = PE[10] ^ CE[10];
    assign sE12   = PE[11] ^ CE[11];
    assign sE13   = PE[12] ^ CE[12];
    assign sE14   = PE[13] ^ CE[13];
    assign sE15   = PE[14] ^ CE[14];
    assign sE16   = PE[15] ^ CE[15];
    assign sE17   = PE[16] ^ CE[16];
    assign sE18   = PE[17] ^ CE[17];
    assign sE19   = PE[18] ^ CE[18];
    assign sE20   = PE[19] ^ CE[19];
    assign sE21   = PE[20] ^ CE[20];
    assign sE22   = PE[21] ^ CE[21];
    assign sE23   = PE[22] ^ CE[22];

    /* Final Stage - 15th CLA */
    wire [28:0] G, P, C;
    assign G[0]  = s102     & pp2[0];
    assign G[1]  = s103     & s201;
    assign G[2]  = sD01     & pp4[0];
    assign G[3]  = sD02     & s301;
    assign G[4]  = sD03     & sE01;
    assign G[5]  = sD04     & sE02;
    assign G[6]  = sD05     & sE03;
    assign G[7]  = sD06     & sE04;
    assign G[8]  = sD07     & sE05;
    assign G[9]  = sD08     & sE06;
    assign G[10] = sD09     & sE07;
    assign G[11] = sD10     & sE08;
    assign G[12] = sD11     & sE09;
    assign G[13] = sD12     & sE10;
    assign G[14] = sD13     & sE11;
    assign G[15] = sD14     & sE12;
    assign G[16] = sD15     & sE13;
    assign G[17] = sD16     & sE14;
    assign G[18] = sD17     & sE15;
    assign G[19] = sD18     & sE16;
    assign G[20] = sD19     & sE17;
    assign G[21] = sD20     & sE18;
    assign G[22] = sD21     & sE19;
    assign G[23] = sD22     & sE20;
    assign G[24] = sD23     & sE21;
    assign G[25] = sD24     & sE22;
    assign G[26] = sD25     & sE23;
    assign G[27] = sD26     & c14;
    assign G[28] = pp15[15] & c13;
    assign P[0]  = s102     ^ pp2[0];
    assign P[1]  = s103     ^ s201;
    assign P[2]  = sD01     ^ pp4[0];
    assign P[3]  = sD02     ^ s301;
    assign P[4]  = sD03     ^ sE01;
    assign P[5]  = sD04     ^ sE02;
    assign P[6]  = sD05     ^ sE03;
    assign P[7]  = sD06     ^ sE04;
    assign P[8]  = sD07     ^ sE05;
    assign P[9]  = sD08     ^ sE06;
    assign P[10] = sD09     ^ sE07;
    assign P[11] = sD10     ^ sE08;
    assign P[12] = sD11     ^ sE09;
    assign P[13] = sD12     ^ sE10;
    assign P[14] = sD13     ^ sE11;
    assign P[15] = sD14     ^ sE12;
    assign P[16] = sD15     ^ sE13;
    assign P[17] = sD16     ^ sE14;
    assign P[18] = sD17     ^ sE15;
    assign P[19] = sD18     ^ sE16;
    assign P[20] = sD19     ^ sE17;
    assign P[21] = sD20     ^ sE18;
    assign P[22] = sD21     ^ sE19;
    assign P[23] = sD22     ^ sE20;
    assign P[24] = sD23     ^ sE21;
    assign P[25] = sD24     ^ sE22;
    assign P[26] = sD25     ^ sE23;
    assign P[27] = sD26     ^ c14;
    assign P[28] = pp15[15] ^ c13;
    assign C[0]  = 0;
    assign C[1]  = G[0]  | (P[0]  & C[0]);
    assign C[2]  = G[1]  | (P[1]  & C[1]);
    assign C[3]  = G[2]  | (P[2]  & C[2]);
    assign C[4]  = G[3]  | (P[3]  & C[3]);
    assign C[5]  = G[4]  | (P[4]  & C[4]);
    assign C[6]  = G[5]  | (P[5]  & C[5]);
    assign C[7]  = G[6]  | (P[6]  & C[6]);
    assign C[8]  = G[7]  | (P[7]  & C[7]);
    assign C[9]  = G[8]  | (P[8]  & C[8]);
    assign C[10] = G[9]  | (P[9]  & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign product[31]  = G[28] | (P[28] & C[28]);
    assign product[2]   = P[0];
    assign product[3]   = P[1]  ^ C[1];
    assign product[4]   = P[2]  ^ C[2];
    assign product[5]   = P[3]  ^ C[3];
    assign product[6]   = P[4]  ^ C[4];
    assign product[7]   = P[5]  ^ C[5];
    assign product[8]   = P[6]  ^ C[6];
    assign product[9]   = P[7]  ^ C[7];
    assign product[10]  = P[8]  ^ C[8];
    assign product[11]  = P[9]  ^ C[9];
    assign product[12]  = P[10] ^ C[10];
    assign product[13]  = P[11] ^ C[11];
    assign product[14]  = P[12] ^ C[12];
    assign product[15]  = P[13] ^ C[13];
    assign product[16]  = P[14] ^ C[14];
    assign product[17]  = P[15] ^ C[15];
    assign product[18]  = P[16] ^ C[16];
    assign product[19]  = P[17] ^ C[17];
    assign product[20]  = P[18] ^ C[18];
    assign product[21]  = P[19] ^ C[19];
    assign product[22]  = P[20] ^ C[20];
    assign product[23]  = P[21] ^ C[21];
    assign product[24]  = P[22] ^ C[22];
    assign product[25]  = P[23] ^ C[23];
    assign product[26]  = P[24] ^ C[24];
    assign product[27]  = P[25] ^ C[25];
    assign product[28]  = P[26] ^ C[26]; 
    assign product[29]  = P[27] ^ C[27];
    assign product[30]  = P[28] ^ C[28];

endmodule
