/*
 * Area: 899.648079
 * Power: 0.2020mW
 * Timing: 0.60
 */
module reduced_multiplier_4(output wire [7:0] product,
                            input wire [3:0] A, B);

    assign product[0] = A[0] & B[0];
    assign product[1] = (A[0] | A[1]) & (A[0] | B[0]) & (A[1] | B[1]) & (B[0] | B[1]) & (~A[0] | ~A[1] | ~B[0] | ~B[1]);
    assign product[2] = (A[0] | A[1] | A[2]) & (A[0] | A[1] | B[0]) & (A[0] | A[2] | B[1]) & (A[0] | B[0] | B[1]) & (A[0] | ~A[1] | ~A[2] | ~B[0] | ~B[1]) & (A[1] | B[0] | B[2]) & (A[2] | B[2] | ~A[0] | ~B[0]) & (B[0] | B[1] | B[2]) & (B[0] | ~A[0] | ~A[1] | ~B[1] | ~B[2]) & (~A[0] | ~A[2] | ~B[0] | ~B[2]);
    assign product[3] = (A[0] | A[1] | A[2] | A[3]) & (A[0] | A[1] | A[2] | B[0]) & (A[0] | A[1] | A[3] | B[1]) & (A[0] | A[1] | B[0] | B[1]) & (A[0] | A[1] | ~A[2] | ~A[3] | ~B[0] | ~B[1]) & (A[0] | A[2] | B[0] | B[2]) & (A[0] | A[3] | B[2] | ~A[1] | ~B[0]) & (A[0] | B[0] | B[1] | B[2]) & (A[0] | B[0] | ~A[1] | ~A[2] | ~B[1] | ~B[2]) & (A[0] | ~A[1] | ~A[3] | ~B[0] | ~B[2]) & (A[1] | A[2] | A[3] | B[3]) & (A[1] | A[2] | ~A[0] | ~A[3] | ~B[0] | ~B[3]) & (A[1] | A[3] | B[1] | ~A[2] | ~B[0] | ~B[2] | ~B[3]) & (A[1] | A[3] | B[2] | ~A[0] | ~A[2] | ~B[1] | ~B[3]) & (A[1] | B[0] | B[1] | B[3]) & (A[1] | B[1] | B[3] | ~A[0] | ~A[2] | ~A[3] | ~B[2]) & (A[1] | B[2] | B[3] | ~A[2] | ~A[3] | ~B[0] | ~B[1]) & (A[2] | A[3] | B[1] | ~A[0] | ~A[1] | ~B[2] | ~B[3]) & (A[2] | A[3] | B[2] | ~A[1] | ~B[0] | ~B[1] | ~B[3]) & (A[2] | B[0] | B[3] | ~A[0] | ~B[1]) & (A[2] | B[1] | B[3] | ~A[1] | ~A[3] | ~B[0] | ~B[2]) & (A[2] | B[2] | B[3] | ~A[0] | ~A[1] | ~A[3] | ~B[1]) & (A[3] | B[1] | B[2] | B[3]) & (A[3] | B[3] | ~A[0] | ~A[1] | ~A[2] | ~B[0]) & (A[3] | B[3] | ~A[0] | ~B[0] | ~B[1] | ~B[2]) & (B[0] | B[1] | B[2] | B[3]) & (B[0] | B[1] | ~A[0] | ~A[1] | ~B[2] | ~B[3]) & (B[0] | ~A[0] | ~A[2] | ~B[1] | ~B[3]) & (B[1] | B[2] | ~A[0] | ~A[3] | ~B[0] | ~B[3]) & (~A[0] | ~A[1] | ~A[2] | ~A[3] | ~B[0] | ~B[3]) & (~A[0] | ~A[3] | ~B[0] | ~B[1] | ~B[2] | ~B[3]) & (~A[1] | ~A[3] | ~B[0] | ~B[1] | ~B[2] | ~B[3]);
    assign product[4] = (A[0] | A[1] | A[2] | B[1]) & (A[0] | A[1] | A[3] | B[2]) & (A[0] | A[1] | B[0] | ~A[2] | ~A[3] | ~B[1] | ~B[2]) & (A[0] | A[1] | B[1] | B[2]) & (A[0] | A[1] | B[2] | ~A[2] | ~B[0]) & (A[0] | A[2] | A[3] | B[3]) & (A[0] | A[2] | B[1] | ~A[3] | ~B[0] | ~B[2] | ~B[3]) & (A[0] | A[2] | B[2] | ~A[1] | ~A[3] | ~B[1] | ~B[3]) & (A[0] | A[3] | B[0] | B[3] | ~A[1] | ~B[1]) & (A[0] | A[3] | B[1] | ~A[1] | ~A[2] | ~B[2] | ~B[3]) & (A[0] | A[3] | B[2] | ~A[2] | ~B[0] | ~B[1] | ~B[3]) & (A[0] | B[0] | B[1] | ~A[1] | ~A[2] | ~B[2] | ~B[3]) & (A[0] | B[0] | ~A[1] | ~A[3] | ~B[1] | ~B[3]) & (A[0] | B[3] | ~A[1] | ~B[0] | ~B[1] | ~B[2]) & (A[1] | A[2] | A[3]) & (A[1] | A[2] | B[0] | B[1]) & (A[1] | A[2] | B[1] | B[3]) & (A[1] | A[2] | ~A[0] | ~B[0] | ~B[1] | ~B[3]) & (A[1] | A[3] | B[1] | B[2]) & (A[1] | A[3] | B[1] | ~A[0] | ~B[0] | ~B[3]) & (A[1] | A[3] | B[2] | B[3]) & (A[1] | A[3] | B[3] | ~A[0] | ~B[0] | ~B[1]) & (A[1] | B[0] | B[1] | B[2]) & (A[1] | B[0] | B[2] | ~A[0] | ~A[2] | ~A[3] | ~B[3]) & (A[1] | B[0] | B[3] | ~A[2] | ~A[3] | ~B[1] | ~B[2]) & (A[1] | B[1] | B[3] | ~A[0] | ~A[3] | ~B[0]) & (A[1] | B[2] | B[3] | ~A[2] | ~B[0]) & (A[1] | ~A[0] | ~A[2] | ~B[0] | ~B[2] | ~B[3]) & (A[1] | ~A[0] | ~A[3] | ~B[0] | ~B[1] | ~B[3]) & (A[2] | A[3] | B[1] | B[3]) & (A[2] | A[3] | B[1] | ~A[0] | ~B[2]) & (A[2] | A[3] | B[2] | B[3]) & (A[2] | A[3] | B[2] | ~A[0] | ~B[0] | ~B[1]) & (A[2] | B[0] | B[1] | B[3]) & (A[2] | B[0] | B[1] | ~A[0] | ~B[2]) & (A[2] | B[0] | B[2] | ~A[1] | ~A[3] | ~B[1] | ~B[3]) & (A[2] | B[0] | B[3] | ~A[0] | ~A[1] | ~A[3] | ~B[2]) & (A[2] | B[1] | ~A[0] | ~A[1] | ~B[2] | ~B[3]) & (A[2] | B[2] | B[3] | ~A[0] | ~A[1] | ~B[0]) & (A[3] | B[0] | B[2] | B[3]) & (A[3] | B[0] | ~A[0] | ~A[1] | ~A[2] | ~B[1]) & (A[3] | B[1] | B[3] | ~A[0] | ~A[1] | ~B[0]) & (A[3] | ~A[0] | ~A[1] | ~B[0] | ~B[1] | ~B[3]) & (A[3] | ~A[0] | ~B[1] | ~B[2] | ~B[3]) & (B[1] | B[2] | B[3]) & (B[1] | B[2] | ~A[0] | ~A[1] | ~A[3] | ~B[0]) & (B[3] | ~A[0] | ~A[1] | ~A[3] | ~B[0] | ~B[1]) & (B[3] | ~A[1] | ~A[2] | ~A[3] | ~B[0]) & (~A[0] | ~A[1] | ~A[2] | ~A[3] | ~B[0]) & (~A[0] | ~B[0] | ~B[1] | ~B[2] | ~B[3]);
    assign product[5] = (A[0] | A[1] | A[2] | B[2]) & (A[0] | A[1] | A[3] | B[3]) & (A[0] | A[1] | B[1] | ~A[2] | ~A[3] | ~B[2] | ~B[3]) & (A[0] | A[1] | B[2] | ~A[3] | ~B[0] | ~B[1] | ~B[3]) & (A[0] | A[1] | B[3] | ~A[2] | ~B[1] | ~B[2]) & (A[0] | A[2] | A[3]) & (A[0] | A[2] | B[1] | B[2]) & (A[0] | A[2] | B[1] | ~A[1] | ~B[0] | ~B[3]) & (A[0] | A[2] | B[2] | B[3]) & (A[0] | A[2] | B[3] | ~A[1] | ~B[0] | ~B[1]) & (A[0] | A[3] | B[1] | B[3]) & (A[0] | A[3] | B[1] | ~A[1] | ~B[2]) & (A[0] | A[3] | B[2] | ~A[1] | ~B[0] | ~B[1]) & (A[0] | B[1] | B[3] | ~A[1] | ~A[2] | ~B[0]) & (A[0] | ~A[1] | ~A[2] | ~B[0] | ~B[1] | ~B[3]) & (A[0] | ~A[1] | ~B[1] | ~B[2] | ~B[3]) & (A[1] | A[2] | A[3]) & (A[1] | A[2] | B[0] | B[2]) & (A[1] | A[2] | B[1] | B[2]) & (A[1] | A[2] | B[2] | B[3]) & (A[1] | A[3] | B[0] | B[3]) & (A[1] | A[3] | B[0] | ~A[0] | ~B[1] | ~B[2]) & (A[1] | A[3] | B[1] | B[3]) & (A[1] | A[3] | B[1] | ~A[0] | ~B[0] | ~B[2]) & (A[1] | B[0] | B[1] | ~A[2] | ~A[3] | ~B[2] | ~B[3]) & (A[1] | B[0] | B[2] | ~A[0] | ~A[3] | ~B[1]) & (A[1] | B[0] | B[3] | ~A[2] | ~B[1]) & (A[1] | B[1] | B[3] | ~A[0] | ~A[2] | ~B[0]) & (A[1] | B[2] | ~A[2] | ~A[3] | ~B[0] | ~B[1] | ~B[3]) & (A[1] | B[3] | ~A[2] | ~A[3] | ~B[1] | ~B[2]) & (A[1] | ~A[0] | ~B[0] | ~B[1] | ~B[2] | ~B[3]) & (A[2] | A[3] | B[0] | B[2]) & (A[2] | A[3] | B[1] | B[2]) & (A[2] | A[3] | B[3]) & (A[2] | B[0] | B[1] | B[2]) & (A[2] | B[0] | B[1] | ~A[0] | ~A[1] | ~A[3] | ~B[3]) & (A[2] | B[0] | B[3] | ~A[0] | ~A[1] | ~B[1]) & (A[2] | B[1] | ~A[1] | ~A[3] | ~B[0] | ~B[2] | ~B[3]) & (A[2] | B[3] | ~A[1] | ~B[0] | ~B[1] | ~B[2]) & (A[3] | B[0] | B[1] | B[3]) & (A[3] | B[0] | B[1] | ~A[1] | ~A[2] | ~B[2]) & (A[3] | B[0] | B[2] | ~A[0] | ~A[1] | ~B[1]) & (A[3] | B[1] | ~A[1] | ~A[2] | ~B[2] | ~B[3]) & (A[3] | B[2] | B[3]) & (A[3] | B[2] | ~A[1] | ~A[2] | ~B[0] | ~B[1]) & (B[0] | B[2] | B[3]) & (B[0] | ~A[1] | ~A[2] | ~A[3] | ~B[1]) & (B[0] | ~A[1] | ~A[3] | ~B[1] | ~B[2] | ~B[3]) & (B[1] | B[2] | B[3]) & (B[1] | ~A[0] | ~A[1] | ~A[2] | ~A[3] | ~B[0]);
    assign product[6] = (A[0] | A[1] | A[3]) & (A[0] | A[1] | B[1] | B[3]) & (A[0] | A[1] | ~A[2] | ~B[2] | ~B[3]) & (A[0] | A[2] | B[0] | B[3]) & (A[0] | A[3] | B[0] | B[2]) & (A[0] | B[1] | ~A[2] | ~A[3] | ~B[2] | ~B[3]) & (A[1] | A[2] | B[3]) & (A[1] | A[2] | ~A[0] | ~B[0] | ~B[1] | ~B[2]) & (A[1] | A[3] | B[0] | B[1]) & (A[1] | A[3] | B[2]) & (A[1] | B[0] | ~A[2] | ~A[3] | ~B[2] | ~B[3]) & (A[1] | B[1] | ~A[2] | ~A[3] | ~B[2] | ~B[3]) & (A[1] | B[2] | ~A[0] | ~A[2] | ~B[1]) & (A[1] | B[2] | ~A[2] | ~B[0] | ~B[1]) & (A[2] | A[3]) & (A[2] | B[1] | B[3]) & (A[2] | B[1] | ~A[0] | ~A[1] | ~B[2]) & (A[2] | B[1] | ~A[1] | ~B[0] | ~B[2]) & (A[2] | ~A[1] | ~B[1] | ~B[2] | ~B[3]) & (A[3] | B[1] | B[2]) & (A[3] | B[3]) & (B[0] | B[1] | B[3]) & (B[0] | B[1] | ~A[2] | ~A[3] | ~B[2]) & (B[1] | B[2] | ~A[0] | ~A[1] | ~A[2] | ~B[0]) & (B[2] | B[3]) & (B[2] | ~A[1] | ~A[2] | ~A[3] | ~B[1]);
    assign product[7] = (A[0] | A[1] | A[2]) & (A[0] | A[1] | B[0] | B[2]) & (A[0] | A[2] | B[0] | B[1]) & (A[0] | B[1] | B[2]) & (A[1] | A[2] | B[0]) & (A[1] | A[2] | B[1]) & (A[1] | B[1] | B[2]) & (A[2] | B[2]) & (B[0] | B[1] | B[2]) & A[3] & B[3];


endmodule
