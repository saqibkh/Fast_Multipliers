module dadda_unsigned_multiplier_RCA_32(product, A, B);
    input [31:0] A, B;
    output [63:0] product;

    wire [31:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;
	wire [31:0] pp16, pp17, pp18, pp19, pp20, pp21, pp22, pp23, pp24, pp25, pp26, pp27, pp28, pp29, pp30, pp31;

	assign pp0[0] = A[0] & B[0];
	assign pp0[1] = A[0] & B[1];
	assign pp0[2] = A[0] & B[2];
	assign pp0[3] = A[0] & B[3];
	assign pp0[4] = A[0] & B[4];
	assign pp0[5] = A[0] & B[5];
	assign pp0[6] = A[0] & B[6];
	assign pp0[7] = A[0] & B[7];
	assign pp0[8] = A[0] & B[8];
	assign pp0[9] = A[0] & B[9];
	assign pp0[10] = A[0] & B[10];
	assign pp0[11] = A[0] & B[11];
	assign pp0[12] = A[0] & B[12];
	assign pp0[13] = A[0] & B[13];
	assign pp0[14] = A[0] & B[14];
	assign pp0[15] = A[0] & B[15];
	assign pp0[16] = A[0] & B[16];
	assign pp0[17] = A[0] & B[17];
	assign pp0[18] = A[0] & B[18];
	assign pp0[19] = A[0] & B[19];
	assign pp0[20] = A[0] & B[20];
	assign pp0[21] = A[0] & B[21];
	assign pp0[22] = A[0] & B[22];
	assign pp0[23] = A[0] & B[23];
	assign pp0[24] = A[0] & B[24];
	assign pp0[25] = A[0] & B[25];
	assign pp0[26] = A[0] & B[26];
	assign pp0[27] = A[0] & B[27];
	assign pp0[28] = A[0] & B[28];
	assign pp0[29] = A[0] & B[29];
	assign pp0[30] = A[0] & B[30];
	assign pp0[31] = A[0] & B[31];
	assign pp1[0] = A[1] & B[0];
	assign pp1[1] = A[1] & B[1];
	assign pp1[2] = A[1] & B[2];
	assign pp1[3] = A[1] & B[3];
	assign pp1[4] = A[1] & B[4];
	assign pp1[5] = A[1] & B[5];
	assign pp1[6] = A[1] & B[6];
	assign pp1[7] = A[1] & B[7];
	assign pp1[8] = A[1] & B[8];
	assign pp1[9] = A[1] & B[9];
	assign pp1[10] = A[1] & B[10];
	assign pp1[11] = A[1] & B[11];
	assign pp1[12] = A[1] & B[12];
	assign pp1[13] = A[1] & B[13];
	assign pp1[14] = A[1] & B[14];
	assign pp1[15] = A[1] & B[15];
	assign pp1[16] = A[1] & B[16];
	assign pp1[17] = A[1] & B[17];
	assign pp1[18] = A[1] & B[18];
	assign pp1[19] = A[1] & B[19];
	assign pp1[20] = A[1] & B[20];
	assign pp1[21] = A[1] & B[21];
	assign pp1[22] = A[1] & B[22];
	assign pp1[23] = A[1] & B[23];
	assign pp1[24] = A[1] & B[24];
	assign pp1[25] = A[1] & B[25];
	assign pp1[26] = A[1] & B[26];
	assign pp1[27] = A[1] & B[27];
	assign pp1[28] = A[1] & B[28];
	assign pp1[29] = A[1] & B[29];
	assign pp1[30] = A[1] & B[30];
	assign pp1[31] = A[1] & B[31];
	assign pp2[0] = A[2] & B[0];
	assign pp2[1] = A[2] & B[1];
	assign pp2[2] = A[2] & B[2];
	assign pp2[3] = A[2] & B[3];
	assign pp2[4] = A[2] & B[4];
	assign pp2[5] = A[2] & B[5];
	assign pp2[6] = A[2] & B[6];
	assign pp2[7] = A[2] & B[7];
	assign pp2[8] = A[2] & B[8];
	assign pp2[9] = A[2] & B[9];
	assign pp2[10] = A[2] & B[10];
	assign pp2[11] = A[2] & B[11];
	assign pp2[12] = A[2] & B[12];
	assign pp2[13] = A[2] & B[13];
	assign pp2[14] = A[2] & B[14];
	assign pp2[15] = A[2] & B[15];
	assign pp2[16] = A[2] & B[16];
	assign pp2[17] = A[2] & B[17];
	assign pp2[18] = A[2] & B[18];
	assign pp2[19] = A[2] & B[19];
	assign pp2[20] = A[2] & B[20];
	assign pp2[21] = A[2] & B[21];
	assign pp2[22] = A[2] & B[22];
	assign pp2[23] = A[2] & B[23];
	assign pp2[24] = A[2] & B[24];
	assign pp2[25] = A[2] & B[25];
	assign pp2[26] = A[2] & B[26];
	assign pp2[27] = A[2] & B[27];
	assign pp2[28] = A[2] & B[28];
	assign pp2[29] = A[2] & B[29];
	assign pp2[30] = A[2] & B[30];
	assign pp2[31] = A[2] & B[31];
	assign pp3[0] = A[3] & B[0];
	assign pp3[1] = A[3] & B[1];
	assign pp3[2] = A[3] & B[2];
	assign pp3[3] = A[3] & B[3];
	assign pp3[4] = A[3] & B[4];
	assign pp3[5] = A[3] & B[5];
	assign pp3[6] = A[3] & B[6];
	assign pp3[7] = A[3] & B[7];
	assign pp3[8] = A[3] & B[8];
	assign pp3[9] = A[3] & B[9];
	assign pp3[10] = A[3] & B[10];
	assign pp3[11] = A[3] & B[11];
	assign pp3[12] = A[3] & B[12];
	assign pp3[13] = A[3] & B[13];
	assign pp3[14] = A[3] & B[14];
	assign pp3[15] = A[3] & B[15];
	assign pp3[16] = A[3] & B[16];
	assign pp3[17] = A[3] & B[17];
	assign pp3[18] = A[3] & B[18];
	assign pp3[19] = A[3] & B[19];
	assign pp3[20] = A[3] & B[20];
	assign pp3[21] = A[3] & B[21];
	assign pp3[22] = A[3] & B[22];
	assign pp3[23] = A[3] & B[23];
	assign pp3[24] = A[3] & B[24];
	assign pp3[25] = A[3] & B[25];
	assign pp3[26] = A[3] & B[26];
	assign pp3[27] = A[3] & B[27];
	assign pp3[28] = A[3] & B[28];
	assign pp3[29] = A[3] & B[29];
	assign pp3[30] = A[3] & B[30];
	assign pp3[31] = A[3] & B[31];
	assign pp4[0] = A[4] & B[0];
	assign pp4[1] = A[4] & B[1];
	assign pp4[2] = A[4] & B[2];
	assign pp4[3] = A[4] & B[3];
	assign pp4[4] = A[4] & B[4];
	assign pp4[5] = A[4] & B[5];
	assign pp4[6] = A[4] & B[6];
	assign pp4[7] = A[4] & B[7];
	assign pp4[8] = A[4] & B[8];
	assign pp4[9] = A[4] & B[9];
	assign pp4[10] = A[4] & B[10];
	assign pp4[11] = A[4] & B[11];
	assign pp4[12] = A[4] & B[12];
	assign pp4[13] = A[4] & B[13];
	assign pp4[14] = A[4] & B[14];
	assign pp4[15] = A[4] & B[15];
	assign pp4[16] = A[4] & B[16];
	assign pp4[17] = A[4] & B[17];
	assign pp4[18] = A[4] & B[18];
	assign pp4[19] = A[4] & B[19];
	assign pp4[20] = A[4] & B[20];
	assign pp4[21] = A[4] & B[21];
	assign pp4[22] = A[4] & B[22];
	assign pp4[23] = A[4] & B[23];
	assign pp4[24] = A[4] & B[24];
	assign pp4[25] = A[4] & B[25];
	assign pp4[26] = A[4] & B[26];
	assign pp4[27] = A[4] & B[27];
	assign pp4[28] = A[4] & B[28];
	assign pp4[29] = A[4] & B[29];
	assign pp4[30] = A[4] & B[30];
	assign pp4[31] = A[4] & B[31];
	assign pp5[0] = A[5] & B[0];
	assign pp5[1] = A[5] & B[1];
	assign pp5[2] = A[5] & B[2];
	assign pp5[3] = A[5] & B[3];
	assign pp5[4] = A[5] & B[4];
	assign pp5[5] = A[5] & B[5];
	assign pp5[6] = A[5] & B[6];
	assign pp5[7] = A[5] & B[7];
	assign pp5[8] = A[5] & B[8];
	assign pp5[9] = A[5] & B[9];
	assign pp5[10] = A[5] & B[10];
	assign pp5[11] = A[5] & B[11];
	assign pp5[12] = A[5] & B[12];
	assign pp5[13] = A[5] & B[13];
	assign pp5[14] = A[5] & B[14];
	assign pp5[15] = A[5] & B[15];
	assign pp5[16] = A[5] & B[16];
	assign pp5[17] = A[5] & B[17];
	assign pp5[18] = A[5] & B[18];
	assign pp5[19] = A[5] & B[19];
	assign pp5[20] = A[5] & B[20];
	assign pp5[21] = A[5] & B[21];
	assign pp5[22] = A[5] & B[22];
	assign pp5[23] = A[5] & B[23];
	assign pp5[24] = A[5] & B[24];
	assign pp5[25] = A[5] & B[25];
	assign pp5[26] = A[5] & B[26];
	assign pp5[27] = A[5] & B[27];
	assign pp5[28] = A[5] & B[28];
	assign pp5[29] = A[5] & B[29];
	assign pp5[30] = A[5] & B[30];
	assign pp5[31] = A[5] & B[31];
	assign pp6[0] = A[6] & B[0];
	assign pp6[1] = A[6] & B[1];
	assign pp6[2] = A[6] & B[2];
	assign pp6[3] = A[6] & B[3];
	assign pp6[4] = A[6] & B[4];
	assign pp6[5] = A[6] & B[5];
	assign pp6[6] = A[6] & B[6];
	assign pp6[7] = A[6] & B[7];
	assign pp6[8] = A[6] & B[8];
	assign pp6[9] = A[6] & B[9];
	assign pp6[10] = A[6] & B[10];
	assign pp6[11] = A[6] & B[11];
	assign pp6[12] = A[6] & B[12];
	assign pp6[13] = A[6] & B[13];
	assign pp6[14] = A[6] & B[14];
	assign pp6[15] = A[6] & B[15];
	assign pp6[16] = A[6] & B[16];
	assign pp6[17] = A[6] & B[17];
	assign pp6[18] = A[6] & B[18];
	assign pp6[19] = A[6] & B[19];
	assign pp6[20] = A[6] & B[20];
	assign pp6[21] = A[6] & B[21];
	assign pp6[22] = A[6] & B[22];
	assign pp6[23] = A[6] & B[23];
	assign pp6[24] = A[6] & B[24];
	assign pp6[25] = A[6] & B[25];
	assign pp6[26] = A[6] & B[26];
	assign pp6[27] = A[6] & B[27];
	assign pp6[28] = A[6] & B[28];
	assign pp6[29] = A[6] & B[29];
	assign pp6[30] = A[6] & B[30];
	assign pp6[31] = A[6] & B[31];
	assign pp7[0] = A[7] & B[0];
	assign pp7[1] = A[7] & B[1];
	assign pp7[2] = A[7] & B[2];
	assign pp7[3] = A[7] & B[3];
	assign pp7[4] = A[7] & B[4];
	assign pp7[5] = A[7] & B[5];
	assign pp7[6] = A[7] & B[6];
	assign pp7[7] = A[7] & B[7];
	assign pp7[8] = A[7] & B[8];
	assign pp7[9] = A[7] & B[9];
	assign pp7[10] = A[7] & B[10];
	assign pp7[11] = A[7] & B[11];
	assign pp7[12] = A[7] & B[12];
	assign pp7[13] = A[7] & B[13];
	assign pp7[14] = A[7] & B[14];
	assign pp7[15] = A[7] & B[15];
	assign pp7[16] = A[7] & B[16];
	assign pp7[17] = A[7] & B[17];
	assign pp7[18] = A[7] & B[18];
	assign pp7[19] = A[7] & B[19];
	assign pp7[20] = A[7] & B[20];
	assign pp7[21] = A[7] & B[21];
	assign pp7[22] = A[7] & B[22];
	assign pp7[23] = A[7] & B[23];
	assign pp7[24] = A[7] & B[24];
	assign pp7[25] = A[7] & B[25];
	assign pp7[26] = A[7] & B[26];
	assign pp7[27] = A[7] & B[27];
	assign pp7[28] = A[7] & B[28];
	assign pp7[29] = A[7] & B[29];
	assign pp7[30] = A[7] & B[30];
	assign pp7[31] = A[7] & B[31];
	assign pp8[0] = A[8] & B[0];
	assign pp8[1] = A[8] & B[1];
	assign pp8[2] = A[8] & B[2];
	assign pp8[3] = A[8] & B[3];
	assign pp8[4] = A[8] & B[4];
	assign pp8[5] = A[8] & B[5];
	assign pp8[6] = A[8] & B[6];
	assign pp8[7] = A[8] & B[7];
	assign pp8[8] = A[8] & B[8];
	assign pp8[9] = A[8] & B[9];
	assign pp8[10] = A[8] & B[10];
	assign pp8[11] = A[8] & B[11];
	assign pp8[12] = A[8] & B[12];
	assign pp8[13] = A[8] & B[13];
	assign pp8[14] = A[8] & B[14];
	assign pp8[15] = A[8] & B[15];
	assign pp8[16] = A[8] & B[16];
	assign pp8[17] = A[8] & B[17];
	assign pp8[18] = A[8] & B[18];
	assign pp8[19] = A[8] & B[19];
	assign pp8[20] = A[8] & B[20];
	assign pp8[21] = A[8] & B[21];
	assign pp8[22] = A[8] & B[22];
	assign pp8[23] = A[8] & B[23];
	assign pp8[24] = A[8] & B[24];
	assign pp8[25] = A[8] & B[25];
	assign pp8[26] = A[8] & B[26];
	assign pp8[27] = A[8] & B[27];
	assign pp8[28] = A[8] & B[28];
	assign pp8[29] = A[8] & B[29];
	assign pp8[30] = A[8] & B[30];
	assign pp8[31] = A[8] & B[31];
	assign pp9[0] = A[9] & B[0];
	assign pp9[1] = A[9] & B[1];
	assign pp9[2] = A[9] & B[2];
	assign pp9[3] = A[9] & B[3];
	assign pp9[4] = A[9] & B[4];
	assign pp9[5] = A[9] & B[5];
	assign pp9[6] = A[9] & B[6];
	assign pp9[7] = A[9] & B[7];
	assign pp9[8] = A[9] & B[8];
	assign pp9[9] = A[9] & B[9];
	assign pp9[10] = A[9] & B[10];
	assign pp9[11] = A[9] & B[11];
	assign pp9[12] = A[9] & B[12];
	assign pp9[13] = A[9] & B[13];
	assign pp9[14] = A[9] & B[14];
	assign pp9[15] = A[9] & B[15];
	assign pp9[16] = A[9] & B[16];
	assign pp9[17] = A[9] & B[17];
	assign pp9[18] = A[9] & B[18];
	assign pp9[19] = A[9] & B[19];
	assign pp9[20] = A[9] & B[20];
	assign pp9[21] = A[9] & B[21];
	assign pp9[22] = A[9] & B[22];
	assign pp9[23] = A[9] & B[23];
	assign pp9[24] = A[9] & B[24];
	assign pp9[25] = A[9] & B[25];
	assign pp9[26] = A[9] & B[26];
	assign pp9[27] = A[9] & B[27];
	assign pp9[28] = A[9] & B[28];
	assign pp9[29] = A[9] & B[29];
	assign pp9[30] = A[9] & B[30];
	assign pp9[31] = A[9] & B[31];
	assign pp10[0] = A[10] & B[0];
	assign pp10[1] = A[10] & B[1];
	assign pp10[2] = A[10] & B[2];
	assign pp10[3] = A[10] & B[3];
	assign pp10[4] = A[10] & B[4];
	assign pp10[5] = A[10] & B[5];
	assign pp10[6] = A[10] & B[6];
	assign pp10[7] = A[10] & B[7];
	assign pp10[8] = A[10] & B[8];
	assign pp10[9] = A[10] & B[9];
	assign pp10[10] = A[10] & B[10];
	assign pp10[11] = A[10] & B[11];
	assign pp10[12] = A[10] & B[12];
	assign pp10[13] = A[10] & B[13];
	assign pp10[14] = A[10] & B[14];
	assign pp10[15] = A[10] & B[15];
	assign pp10[16] = A[10] & B[16];
	assign pp10[17] = A[10] & B[17];
	assign pp10[18] = A[10] & B[18];
	assign pp10[19] = A[10] & B[19];
	assign pp10[20] = A[10] & B[20];
	assign pp10[21] = A[10] & B[21];
	assign pp10[22] = A[10] & B[22];
	assign pp10[23] = A[10] & B[23];
	assign pp10[24] = A[10] & B[24];
	assign pp10[25] = A[10] & B[25];
	assign pp10[26] = A[10] & B[26];
	assign pp10[27] = A[10] & B[27];
	assign pp10[28] = A[10] & B[28];
	assign pp10[29] = A[10] & B[29];
	assign pp10[30] = A[10] & B[30];
	assign pp10[31] = A[10] & B[31];
	assign pp11[0] = A[11] & B[0];
	assign pp11[1] = A[11] & B[1];
	assign pp11[2] = A[11] & B[2];
	assign pp11[3] = A[11] & B[3];
	assign pp11[4] = A[11] & B[4];
	assign pp11[5] = A[11] & B[5];
	assign pp11[6] = A[11] & B[6];
	assign pp11[7] = A[11] & B[7];
	assign pp11[8] = A[11] & B[8];
	assign pp11[9] = A[11] & B[9];
	assign pp11[10] = A[11] & B[10];
	assign pp11[11] = A[11] & B[11];
	assign pp11[12] = A[11] & B[12];
	assign pp11[13] = A[11] & B[13];
	assign pp11[14] = A[11] & B[14];
	assign pp11[15] = A[11] & B[15];
	assign pp11[16] = A[11] & B[16];
	assign pp11[17] = A[11] & B[17];
	assign pp11[18] = A[11] & B[18];
	assign pp11[19] = A[11] & B[19];
	assign pp11[20] = A[11] & B[20];
	assign pp11[21] = A[11] & B[21];
	assign pp11[22] = A[11] & B[22];
	assign pp11[23] = A[11] & B[23];
	assign pp11[24] = A[11] & B[24];
	assign pp11[25] = A[11] & B[25];
	assign pp11[26] = A[11] & B[26];
	assign pp11[27] = A[11] & B[27];
	assign pp11[28] = A[11] & B[28];
	assign pp11[29] = A[11] & B[29];
	assign pp11[30] = A[11] & B[30];
	assign pp11[31] = A[11] & B[31];
	assign pp12[0] = A[12] & B[0];
	assign pp12[1] = A[12] & B[1];
	assign pp12[2] = A[12] & B[2];
	assign pp12[3] = A[12] & B[3];
	assign pp12[4] = A[12] & B[4];
	assign pp12[5] = A[12] & B[5];
	assign pp12[6] = A[12] & B[6];
	assign pp12[7] = A[12] & B[7];
	assign pp12[8] = A[12] & B[8];
	assign pp12[9] = A[12] & B[9];
	assign pp12[10] = A[12] & B[10];
	assign pp12[11] = A[12] & B[11];
	assign pp12[12] = A[12] & B[12];
	assign pp12[13] = A[12] & B[13];
	assign pp12[14] = A[12] & B[14];
	assign pp12[15] = A[12] & B[15];
	assign pp12[16] = A[12] & B[16];
	assign pp12[17] = A[12] & B[17];
	assign pp12[18] = A[12] & B[18];
	assign pp12[19] = A[12] & B[19];
	assign pp12[20] = A[12] & B[20];
	assign pp12[21] = A[12] & B[21];
	assign pp12[22] = A[12] & B[22];
	assign pp12[23] = A[12] & B[23];
	assign pp12[24] = A[12] & B[24];
	assign pp12[25] = A[12] & B[25];
	assign pp12[26] = A[12] & B[26];
	assign pp12[27] = A[12] & B[27];
	assign pp12[28] = A[12] & B[28];
	assign pp12[29] = A[12] & B[29];
	assign pp12[30] = A[12] & B[30];
	assign pp12[31] = A[12] & B[31];
	assign pp13[0] = A[13] & B[0];
	assign pp13[1] = A[13] & B[1];
	assign pp13[2] = A[13] & B[2];
	assign pp13[3] = A[13] & B[3];
	assign pp13[4] = A[13] & B[4];
	assign pp13[5] = A[13] & B[5];
	assign pp13[6] = A[13] & B[6];
	assign pp13[7] = A[13] & B[7];
	assign pp13[8] = A[13] & B[8];
	assign pp13[9] = A[13] & B[9];
	assign pp13[10] = A[13] & B[10];
	assign pp13[11] = A[13] & B[11];
	assign pp13[12] = A[13] & B[12];
	assign pp13[13] = A[13] & B[13];
	assign pp13[14] = A[13] & B[14];
	assign pp13[15] = A[13] & B[15];
	assign pp13[16] = A[13] & B[16];
	assign pp13[17] = A[13] & B[17];
	assign pp13[18] = A[13] & B[18];
	assign pp13[19] = A[13] & B[19];
	assign pp13[20] = A[13] & B[20];
	assign pp13[21] = A[13] & B[21];
	assign pp13[22] = A[13] & B[22];
	assign pp13[23] = A[13] & B[23];
	assign pp13[24] = A[13] & B[24];
	assign pp13[25] = A[13] & B[25];
	assign pp13[26] = A[13] & B[26];
	assign pp13[27] = A[13] & B[27];
	assign pp13[28] = A[13] & B[28];
	assign pp13[29] = A[13] & B[29];
	assign pp13[30] = A[13] & B[30];
	assign pp13[31] = A[13] & B[31];
	assign pp14[0] = A[14] & B[0];
	assign pp14[1] = A[14] & B[1];
	assign pp14[2] = A[14] & B[2];
	assign pp14[3] = A[14] & B[3];
	assign pp14[4] = A[14] & B[4];
	assign pp14[5] = A[14] & B[5];
	assign pp14[6] = A[14] & B[6];
	assign pp14[7] = A[14] & B[7];
	assign pp14[8] = A[14] & B[8];
	assign pp14[9] = A[14] & B[9];
	assign pp14[10] = A[14] & B[10];
	assign pp14[11] = A[14] & B[11];
	assign pp14[12] = A[14] & B[12];
	assign pp14[13] = A[14] & B[13];
	assign pp14[14] = A[14] & B[14];
	assign pp14[15] = A[14] & B[15];
	assign pp14[16] = A[14] & B[16];
	assign pp14[17] = A[14] & B[17];
	assign pp14[18] = A[14] & B[18];
	assign pp14[19] = A[14] & B[19];
	assign pp14[20] = A[14] & B[20];
	assign pp14[21] = A[14] & B[21];
	assign pp14[22] = A[14] & B[22];
	assign pp14[23] = A[14] & B[23];
	assign pp14[24] = A[14] & B[24];
	assign pp14[25] = A[14] & B[25];
	assign pp14[26] = A[14] & B[26];
	assign pp14[27] = A[14] & B[27];
	assign pp14[28] = A[14] & B[28];
	assign pp14[29] = A[14] & B[29];
	assign pp14[30] = A[14] & B[30];
	assign pp14[31] = A[14] & B[31];
	assign pp15[0] = A[15] & B[0];
	assign pp15[1] = A[15] & B[1];
	assign pp15[2] = A[15] & B[2];
	assign pp15[3] = A[15] & B[3];
	assign pp15[4] = A[15] & B[4];
	assign pp15[5] = A[15] & B[5];
	assign pp15[6] = A[15] & B[6];
	assign pp15[7] = A[15] & B[7];
	assign pp15[8] = A[15] & B[8];
	assign pp15[9] = A[15] & B[9];
	assign pp15[10] = A[15] & B[10];
	assign pp15[11] = A[15] & B[11];
	assign pp15[12] = A[15] & B[12];
	assign pp15[13] = A[15] & B[13];
	assign pp15[14] = A[15] & B[14];
	assign pp15[15] = A[15] & B[15];
	assign pp15[16] = A[15] & B[16];
	assign pp15[17] = A[15] & B[17];
	assign pp15[18] = A[15] & B[18];
	assign pp15[19] = A[15] & B[19];
	assign pp15[20] = A[15] & B[20];
	assign pp15[21] = A[15] & B[21];
	assign pp15[22] = A[15] & B[22];
	assign pp15[23] = A[15] & B[23];
	assign pp15[24] = A[15] & B[24];
	assign pp15[25] = A[15] & B[25];
	assign pp15[26] = A[15] & B[26];
	assign pp15[27] = A[15] & B[27];
	assign pp15[28] = A[15] & B[28];
	assign pp15[29] = A[15] & B[29];
	assign pp15[30] = A[15] & B[30];
	assign pp15[31] = A[15] & B[31];
	assign pp16[0] = A[16] & B[0];
	assign pp16[1] = A[16] & B[1];
	assign pp16[2] = A[16] & B[2];
	assign pp16[3] = A[16] & B[3];
	assign pp16[4] = A[16] & B[4];
	assign pp16[5] = A[16] & B[5];
	assign pp16[6] = A[16] & B[6];
	assign pp16[7] = A[16] & B[7];
	assign pp16[8] = A[16] & B[8];
	assign pp16[9] = A[16] & B[9];
	assign pp16[10] = A[16] & B[10];
	assign pp16[11] = A[16] & B[11];
	assign pp16[12] = A[16] & B[12];
	assign pp16[13] = A[16] & B[13];
	assign pp16[14] = A[16] & B[14];
	assign pp16[15] = A[16] & B[15];
	assign pp16[16] = A[16] & B[16];
	assign pp16[17] = A[16] & B[17];
	assign pp16[18] = A[16] & B[18];
	assign pp16[19] = A[16] & B[19];
	assign pp16[20] = A[16] & B[20];
	assign pp16[21] = A[16] & B[21];
	assign pp16[22] = A[16] & B[22];
	assign pp16[23] = A[16] & B[23];
	assign pp16[24] = A[16] & B[24];
	assign pp16[25] = A[16] & B[25];
	assign pp16[26] = A[16] & B[26];
	assign pp16[27] = A[16] & B[27];
	assign pp16[28] = A[16] & B[28];
	assign pp16[29] = A[16] & B[29];
	assign pp16[30] = A[16] & B[30];
	assign pp16[31] = A[16] & B[31];
	assign pp17[0] = A[17] & B[0];
	assign pp17[1] = A[17] & B[1];
	assign pp17[2] = A[17] & B[2];
	assign pp17[3] = A[17] & B[3];
	assign pp17[4] = A[17] & B[4];
	assign pp17[5] = A[17] & B[5];
	assign pp17[6] = A[17] & B[6];
	assign pp17[7] = A[17] & B[7];
	assign pp17[8] = A[17] & B[8];
	assign pp17[9] = A[17] & B[9];
	assign pp17[10] = A[17] & B[10];
	assign pp17[11] = A[17] & B[11];
	assign pp17[12] = A[17] & B[12];
	assign pp17[13] = A[17] & B[13];
	assign pp17[14] = A[17] & B[14];
	assign pp17[15] = A[17] & B[15];
	assign pp17[16] = A[17] & B[16];
	assign pp17[17] = A[17] & B[17];
	assign pp17[18] = A[17] & B[18];
	assign pp17[19] = A[17] & B[19];
	assign pp17[20] = A[17] & B[20];
	assign pp17[21] = A[17] & B[21];
	assign pp17[22] = A[17] & B[22];
	assign pp17[23] = A[17] & B[23];
	assign pp17[24] = A[17] & B[24];
	assign pp17[25] = A[17] & B[25];
	assign pp17[26] = A[17] & B[26];
	assign pp17[27] = A[17] & B[27];
	assign pp17[28] = A[17] & B[28];
	assign pp17[29] = A[17] & B[29];
	assign pp17[30] = A[17] & B[30];
	assign pp17[31] = A[17] & B[31];
	assign pp18[0] = A[18] & B[0];
	assign pp18[1] = A[18] & B[1];
	assign pp18[2] = A[18] & B[2];
	assign pp18[3] = A[18] & B[3];
	assign pp18[4] = A[18] & B[4];
	assign pp18[5] = A[18] & B[5];
	assign pp18[6] = A[18] & B[6];
	assign pp18[7] = A[18] & B[7];
	assign pp18[8] = A[18] & B[8];
	assign pp18[9] = A[18] & B[9];
	assign pp18[10] = A[18] & B[10];
	assign pp18[11] = A[18] & B[11];
	assign pp18[12] = A[18] & B[12];
	assign pp18[13] = A[18] & B[13];
	assign pp18[14] = A[18] & B[14];
	assign pp18[15] = A[18] & B[15];
	assign pp18[16] = A[18] & B[16];
	assign pp18[17] = A[18] & B[17];
	assign pp18[18] = A[18] & B[18];
	assign pp18[19] = A[18] & B[19];
	assign pp18[20] = A[18] & B[20];
	assign pp18[21] = A[18] & B[21];
	assign pp18[22] = A[18] & B[22];
	assign pp18[23] = A[18] & B[23];
	assign pp18[24] = A[18] & B[24];
	assign pp18[25] = A[18] & B[25];
	assign pp18[26] = A[18] & B[26];
	assign pp18[27] = A[18] & B[27];
	assign pp18[28] = A[18] & B[28];
	assign pp18[29] = A[18] & B[29];
	assign pp18[30] = A[18] & B[30];
	assign pp18[31] = A[18] & B[31];
	assign pp19[0] = A[19] & B[0];
	assign pp19[1] = A[19] & B[1];
	assign pp19[2] = A[19] & B[2];
	assign pp19[3] = A[19] & B[3];
	assign pp19[4] = A[19] & B[4];
	assign pp19[5] = A[19] & B[5];
	assign pp19[6] = A[19] & B[6];
	assign pp19[7] = A[19] & B[7];
	assign pp19[8] = A[19] & B[8];
	assign pp19[9] = A[19] & B[9];
	assign pp19[10] = A[19] & B[10];
	assign pp19[11] = A[19] & B[11];
	assign pp19[12] = A[19] & B[12];
	assign pp19[13] = A[19] & B[13];
	assign pp19[14] = A[19] & B[14];
	assign pp19[15] = A[19] & B[15];
	assign pp19[16] = A[19] & B[16];
	assign pp19[17] = A[19] & B[17];
	assign pp19[18] = A[19] & B[18];
	assign pp19[19] = A[19] & B[19];
	assign pp19[20] = A[19] & B[20];
	assign pp19[21] = A[19] & B[21];
	assign pp19[22] = A[19] & B[22];
	assign pp19[23] = A[19] & B[23];
	assign pp19[24] = A[19] & B[24];
	assign pp19[25] = A[19] & B[25];
	assign pp19[26] = A[19] & B[26];
	assign pp19[27] = A[19] & B[27];
	assign pp19[28] = A[19] & B[28];
	assign pp19[29] = A[19] & B[29];
	assign pp19[30] = A[19] & B[30];
	assign pp19[31] = A[19] & B[31];
	assign pp20[0] = A[20] & B[0];
	assign pp20[1] = A[20] & B[1];
	assign pp20[2] = A[20] & B[2];
	assign pp20[3] = A[20] & B[3];
	assign pp20[4] = A[20] & B[4];
	assign pp20[5] = A[20] & B[5];
	assign pp20[6] = A[20] & B[6];
	assign pp20[7] = A[20] & B[7];
	assign pp20[8] = A[20] & B[8];
	assign pp20[9] = A[20] & B[9];
	assign pp20[10] = A[20] & B[10];
	assign pp20[11] = A[20] & B[11];
	assign pp20[12] = A[20] & B[12];
	assign pp20[13] = A[20] & B[13];
	assign pp20[14] = A[20] & B[14];
	assign pp20[15] = A[20] & B[15];
	assign pp20[16] = A[20] & B[16];
	assign pp20[17] = A[20] & B[17];
	assign pp20[18] = A[20] & B[18];
	assign pp20[19] = A[20] & B[19];
	assign pp20[20] = A[20] & B[20];
	assign pp20[21] = A[20] & B[21];
	assign pp20[22] = A[20] & B[22];
	assign pp20[23] = A[20] & B[23];
	assign pp20[24] = A[20] & B[24];
	assign pp20[25] = A[20] & B[25];
	assign pp20[26] = A[20] & B[26];
	assign pp20[27] = A[20] & B[27];
	assign pp20[28] = A[20] & B[28];
	assign pp20[29] = A[20] & B[29];
	assign pp20[30] = A[20] & B[30];
	assign pp20[31] = A[20] & B[31];
	assign pp21[0] = A[21] & B[0];
	assign pp21[1] = A[21] & B[1];
	assign pp21[2] = A[21] & B[2];
	assign pp21[3] = A[21] & B[3];
	assign pp21[4] = A[21] & B[4];
	assign pp21[5] = A[21] & B[5];
	assign pp21[6] = A[21] & B[6];
	assign pp21[7] = A[21] & B[7];
	assign pp21[8] = A[21] & B[8];
	assign pp21[9] = A[21] & B[9];
	assign pp21[10] = A[21] & B[10];
	assign pp21[11] = A[21] & B[11];
	assign pp21[12] = A[21] & B[12];
	assign pp21[13] = A[21] & B[13];
	assign pp21[14] = A[21] & B[14];
	assign pp21[15] = A[21] & B[15];
	assign pp21[16] = A[21] & B[16];
	assign pp21[17] = A[21] & B[17];
	assign pp21[18] = A[21] & B[18];
	assign pp21[19] = A[21] & B[19];
	assign pp21[20] = A[21] & B[20];
	assign pp21[21] = A[21] & B[21];
	assign pp21[22] = A[21] & B[22];
	assign pp21[23] = A[21] & B[23];
	assign pp21[24] = A[21] & B[24];
	assign pp21[25] = A[21] & B[25];
	assign pp21[26] = A[21] & B[26];
	assign pp21[27] = A[21] & B[27];
	assign pp21[28] = A[21] & B[28];
	assign pp21[29] = A[21] & B[29];
	assign pp21[30] = A[21] & B[30];
	assign pp21[31] = A[21] & B[31];
	assign pp22[0] = A[22] & B[0];
	assign pp22[1] = A[22] & B[1];
	assign pp22[2] = A[22] & B[2];
	assign pp22[3] = A[22] & B[3];
	assign pp22[4] = A[22] & B[4];
	assign pp22[5] = A[22] & B[5];
	assign pp22[6] = A[22] & B[6];
	assign pp22[7] = A[22] & B[7];
	assign pp22[8] = A[22] & B[8];
	assign pp22[9] = A[22] & B[9];
	assign pp22[10] = A[22] & B[10];
	assign pp22[11] = A[22] & B[11];
	assign pp22[12] = A[22] & B[12];
	assign pp22[13] = A[22] & B[13];
	assign pp22[14] = A[22] & B[14];
	assign pp22[15] = A[22] & B[15];
	assign pp22[16] = A[22] & B[16];
	assign pp22[17] = A[22] & B[17];
	assign pp22[18] = A[22] & B[18];
	assign pp22[19] = A[22] & B[19];
	assign pp22[20] = A[22] & B[20];
	assign pp22[21] = A[22] & B[21];
	assign pp22[22] = A[22] & B[22];
	assign pp22[23] = A[22] & B[23];
	assign pp22[24] = A[22] & B[24];
	assign pp22[25] = A[22] & B[25];
	assign pp22[26] = A[22] & B[26];
	assign pp22[27] = A[22] & B[27];
	assign pp22[28] = A[22] & B[28];
	assign pp22[29] = A[22] & B[29];
	assign pp22[30] = A[22] & B[30];
	assign pp22[31] = A[22] & B[31];
	assign pp23[0] = A[23] & B[0];
	assign pp23[1] = A[23] & B[1];
	assign pp23[2] = A[23] & B[2];
	assign pp23[3] = A[23] & B[3];
	assign pp23[4] = A[23] & B[4];
	assign pp23[5] = A[23] & B[5];
	assign pp23[6] = A[23] & B[6];
	assign pp23[7] = A[23] & B[7];
	assign pp23[8] = A[23] & B[8];
	assign pp23[9] = A[23] & B[9];
	assign pp23[10] = A[23] & B[10];
	assign pp23[11] = A[23] & B[11];
	assign pp23[12] = A[23] & B[12];
	assign pp23[13] = A[23] & B[13];
	assign pp23[14] = A[23] & B[14];
	assign pp23[15] = A[23] & B[15];
	assign pp23[16] = A[23] & B[16];
	assign pp23[17] = A[23] & B[17];
	assign pp23[18] = A[23] & B[18];
	assign pp23[19] = A[23] & B[19];
	assign pp23[20] = A[23] & B[20];
	assign pp23[21] = A[23] & B[21];
	assign pp23[22] = A[23] & B[22];
	assign pp23[23] = A[23] & B[23];
	assign pp23[24] = A[23] & B[24];
	assign pp23[25] = A[23] & B[25];
	assign pp23[26] = A[23] & B[26];
	assign pp23[27] = A[23] & B[27];
	assign pp23[28] = A[23] & B[28];
	assign pp23[29] = A[23] & B[29];
	assign pp23[30] = A[23] & B[30];
	assign pp23[31] = A[23] & B[31];
	assign pp24[0] = A[24] & B[0];
	assign pp24[1] = A[24] & B[1];
	assign pp24[2] = A[24] & B[2];
	assign pp24[3] = A[24] & B[3];
	assign pp24[4] = A[24] & B[4];
	assign pp24[5] = A[24] & B[5];
	assign pp24[6] = A[24] & B[6];
	assign pp24[7] = A[24] & B[7];
	assign pp24[8] = A[24] & B[8];
	assign pp24[9] = A[24] & B[9];
	assign pp24[10] = A[24] & B[10];
	assign pp24[11] = A[24] & B[11];
	assign pp24[12] = A[24] & B[12];
	assign pp24[13] = A[24] & B[13];
	assign pp24[14] = A[24] & B[14];
	assign pp24[15] = A[24] & B[15];
	assign pp24[16] = A[24] & B[16];
	assign pp24[17] = A[24] & B[17];
	assign pp24[18] = A[24] & B[18];
	assign pp24[19] = A[24] & B[19];
	assign pp24[20] = A[24] & B[20];
	assign pp24[21] = A[24] & B[21];
	assign pp24[22] = A[24] & B[22];
	assign pp24[23] = A[24] & B[23];
	assign pp24[24] = A[24] & B[24];
	assign pp24[25] = A[24] & B[25];
	assign pp24[26] = A[24] & B[26];
	assign pp24[27] = A[24] & B[27];
	assign pp24[28] = A[24] & B[28];
	assign pp24[29] = A[24] & B[29];
	assign pp24[30] = A[24] & B[30];
	assign pp24[31] = A[24] & B[31];
	assign pp25[0] = A[25] & B[0];
	assign pp25[1] = A[25] & B[1];
	assign pp25[2] = A[25] & B[2];
	assign pp25[3] = A[25] & B[3];
	assign pp25[4] = A[25] & B[4];
	assign pp25[5] = A[25] & B[5];
	assign pp25[6] = A[25] & B[6];
	assign pp25[7] = A[25] & B[7];
	assign pp25[8] = A[25] & B[8];
	assign pp25[9] = A[25] & B[9];
	assign pp25[10] = A[25] & B[10];
	assign pp25[11] = A[25] & B[11];
	assign pp25[12] = A[25] & B[12];
	assign pp25[13] = A[25] & B[13];
	assign pp25[14] = A[25] & B[14];
	assign pp25[15] = A[25] & B[15];
	assign pp25[16] = A[25] & B[16];
	assign pp25[17] = A[25] & B[17];
	assign pp25[18] = A[25] & B[18];
	assign pp25[19] = A[25] & B[19];
	assign pp25[20] = A[25] & B[20];
	assign pp25[21] = A[25] & B[21];
	assign pp25[22] = A[25] & B[22];
	assign pp25[23] = A[25] & B[23];
	assign pp25[24] = A[25] & B[24];
	assign pp25[25] = A[25] & B[25];
	assign pp25[26] = A[25] & B[26];
	assign pp25[27] = A[25] & B[27];
	assign pp25[28] = A[25] & B[28];
	assign pp25[29] = A[25] & B[29];
	assign pp25[30] = A[25] & B[30];
	assign pp25[31] = A[25] & B[31];
	assign pp26[0] = A[26] & B[0];
	assign pp26[1] = A[26] & B[1];
	assign pp26[2] = A[26] & B[2];
	assign pp26[3] = A[26] & B[3];
	assign pp26[4] = A[26] & B[4];
	assign pp26[5] = A[26] & B[5];
	assign pp26[6] = A[26] & B[6];
	assign pp26[7] = A[26] & B[7];
	assign pp26[8] = A[26] & B[8];
	assign pp26[9] = A[26] & B[9];
	assign pp26[10] = A[26] & B[10];
	assign pp26[11] = A[26] & B[11];
	assign pp26[12] = A[26] & B[12];
	assign pp26[13] = A[26] & B[13];
	assign pp26[14] = A[26] & B[14];
	assign pp26[15] = A[26] & B[15];
	assign pp26[16] = A[26] & B[16];
	assign pp26[17] = A[26] & B[17];
	assign pp26[18] = A[26] & B[18];
	assign pp26[19] = A[26] & B[19];
	assign pp26[20] = A[26] & B[20];
	assign pp26[21] = A[26] & B[21];
	assign pp26[22] = A[26] & B[22];
	assign pp26[23] = A[26] & B[23];
	assign pp26[24] = A[26] & B[24];
	assign pp26[25] = A[26] & B[25];
	assign pp26[26] = A[26] & B[26];
	assign pp26[27] = A[26] & B[27];
	assign pp26[28] = A[26] & B[28];
	assign pp26[29] = A[26] & B[29];
	assign pp26[30] = A[26] & B[30];
	assign pp26[31] = A[26] & B[31];
	assign pp27[0] = A[27] & B[0];
	assign pp27[1] = A[27] & B[1];
	assign pp27[2] = A[27] & B[2];
	assign pp27[3] = A[27] & B[3];
	assign pp27[4] = A[27] & B[4];
	assign pp27[5] = A[27] & B[5];
	assign pp27[6] = A[27] & B[6];
	assign pp27[7] = A[27] & B[7];
	assign pp27[8] = A[27] & B[8];
	assign pp27[9] = A[27] & B[9];
	assign pp27[10] = A[27] & B[10];
	assign pp27[11] = A[27] & B[11];
	assign pp27[12] = A[27] & B[12];
	assign pp27[13] = A[27] & B[13];
	assign pp27[14] = A[27] & B[14];
	assign pp27[15] = A[27] & B[15];
	assign pp27[16] = A[27] & B[16];
	assign pp27[17] = A[27] & B[17];
	assign pp27[18] = A[27] & B[18];
	assign pp27[19] = A[27] & B[19];
	assign pp27[20] = A[27] & B[20];
	assign pp27[21] = A[27] & B[21];
	assign pp27[22] = A[27] & B[22];
	assign pp27[23] = A[27] & B[23];
	assign pp27[24] = A[27] & B[24];
	assign pp27[25] = A[27] & B[25];
	assign pp27[26] = A[27] & B[26];
	assign pp27[27] = A[27] & B[27];
	assign pp27[28] = A[27] & B[28];
	assign pp27[29] = A[27] & B[29];
	assign pp27[30] = A[27] & B[30];
	assign pp27[31] = A[27] & B[31];
	assign pp28[0] = A[28] & B[0];
	assign pp28[1] = A[28] & B[1];
	assign pp28[2] = A[28] & B[2];
	assign pp28[3] = A[28] & B[3];
	assign pp28[4] = A[28] & B[4];
	assign pp28[5] = A[28] & B[5];
	assign pp28[6] = A[28] & B[6];
	assign pp28[7] = A[28] & B[7];
	assign pp28[8] = A[28] & B[8];
	assign pp28[9] = A[28] & B[9];
	assign pp28[10] = A[28] & B[10];
	assign pp28[11] = A[28] & B[11];
	assign pp28[12] = A[28] & B[12];
	assign pp28[13] = A[28] & B[13];
	assign pp28[14] = A[28] & B[14];
	assign pp28[15] = A[28] & B[15];
	assign pp28[16] = A[28] & B[16];
	assign pp28[17] = A[28] & B[17];
	assign pp28[18] = A[28] & B[18];
	assign pp28[19] = A[28] & B[19];
	assign pp28[20] = A[28] & B[20];
	assign pp28[21] = A[28] & B[21];
	assign pp28[22] = A[28] & B[22];
	assign pp28[23] = A[28] & B[23];
	assign pp28[24] = A[28] & B[24];
	assign pp28[25] = A[28] & B[25];
	assign pp28[26] = A[28] & B[26];
	assign pp28[27] = A[28] & B[27];
	assign pp28[28] = A[28] & B[28];
	assign pp28[29] = A[28] & B[29];
	assign pp28[30] = A[28] & B[30];
	assign pp28[31] = A[28] & B[31];
	assign pp29[0] = A[29] & B[0];
	assign pp29[1] = A[29] & B[1];
	assign pp29[2] = A[29] & B[2];
	assign pp29[3] = A[29] & B[3];
	assign pp29[4] = A[29] & B[4];
	assign pp29[5] = A[29] & B[5];
	assign pp29[6] = A[29] & B[6];
	assign pp29[7] = A[29] & B[7];
	assign pp29[8] = A[29] & B[8];
	assign pp29[9] = A[29] & B[9];
	assign pp29[10] = A[29] & B[10];
	assign pp29[11] = A[29] & B[11];
	assign pp29[12] = A[29] & B[12];
	assign pp29[13] = A[29] & B[13];
	assign pp29[14] = A[29] & B[14];
	assign pp29[15] = A[29] & B[15];
	assign pp29[16] = A[29] & B[16];
	assign pp29[17] = A[29] & B[17];
	assign pp29[18] = A[29] & B[18];
	assign pp29[19] = A[29] & B[19];
	assign pp29[20] = A[29] & B[20];
	assign pp29[21] = A[29] & B[21];
	assign pp29[22] = A[29] & B[22];
	assign pp29[23] = A[29] & B[23];
	assign pp29[24] = A[29] & B[24];
	assign pp29[25] = A[29] & B[25];
	assign pp29[26] = A[29] & B[26];
	assign pp29[27] = A[29] & B[27];
	assign pp29[28] = A[29] & B[28];
	assign pp29[29] = A[29] & B[29];
	assign pp29[30] = A[29] & B[30];
	assign pp29[31] = A[29] & B[31];
	assign pp30[0] = A[30] & B[0];
	assign pp30[1] = A[30] & B[1];
	assign pp30[2] = A[30] & B[2];
	assign pp30[3] = A[30] & B[3];
	assign pp30[4] = A[30] & B[4];
	assign pp30[5] = A[30] & B[5];
	assign pp30[6] = A[30] & B[6];
	assign pp30[7] = A[30] & B[7];
	assign pp30[8] = A[30] & B[8];
	assign pp30[9] = A[30] & B[9];
	assign pp30[10] = A[30] & B[10];
	assign pp30[11] = A[30] & B[11];
	assign pp30[12] = A[30] & B[12];
	assign pp30[13] = A[30] & B[13];
	assign pp30[14] = A[30] & B[14];
	assign pp30[15] = A[30] & B[15];
	assign pp30[16] = A[30] & B[16];
	assign pp30[17] = A[30] & B[17];
	assign pp30[18] = A[30] & B[18];
	assign pp30[19] = A[30] & B[19];
	assign pp30[20] = A[30] & B[20];
	assign pp30[21] = A[30] & B[21];
	assign pp30[22] = A[30] & B[22];
	assign pp30[23] = A[30] & B[23];
	assign pp30[24] = A[30] & B[24];
	assign pp30[25] = A[30] & B[25];
	assign pp30[26] = A[30] & B[26];
	assign pp30[27] = A[30] & B[27];
	assign pp30[28] = A[30] & B[28];
	assign pp30[29] = A[30] & B[29];
	assign pp30[30] = A[30] & B[30];
	assign pp30[31] = A[30] & B[31];
	assign pp31[0] = A[31] & B[0];
	assign pp31[1] = A[31] & B[1];
	assign pp31[2] = A[31] & B[2];
	assign pp31[3] = A[31] & B[3];
	assign pp31[4] = A[31] & B[4];
	assign pp31[5] = A[31] & B[5];
	assign pp31[6] = A[31] & B[6];
	assign pp31[7] = A[31] & B[7];
	assign pp31[8] = A[31] & B[8];
	assign pp31[9] = A[31] & B[9];
	assign pp31[10] = A[31] & B[10];
	assign pp31[11] = A[31] & B[11];
	assign pp31[12] = A[31] & B[12];
	assign pp31[13] = A[31] & B[13];
	assign pp31[14] = A[31] & B[14];
	assign pp31[15] = A[31] & B[15];
	assign pp31[16] = A[31] & B[16];
	assign pp31[17] = A[31] & B[17];
	assign pp31[18] = A[31] & B[18];
	assign pp31[19] = A[31] & B[19];
	assign pp31[20] = A[31] & B[20];
	assign pp31[21] = A[31] & B[21];
	assign pp31[22] = A[31] & B[22];
	assign pp31[23] = A[31] & B[23];
	assign pp31[24] = A[31] & B[24];
	assign pp31[25] = A[31] & B[25];
	assign pp31[26] = A[31] & B[26];
	assign pp31[27] = A[31] & B[27];
	assign pp31[28] = A[31] & B[28];
	assign pp31[29] = A[31] & B[29];
	assign pp31[30] = A[31] & B[30];
	assign pp31[31] = A[31] & B[31];

	wire [992:0] S;
	wire [992:0] Cout;
	Half_Adder HA1 (pp0[28], pp1[27], S[1], Cout[1]);
	Full_Adder FA1 (pp0[29], pp1[28], pp2[27], S[2], Cout[2]);
	Half_Adder HA2 (pp3[26], pp4[25], S[3], Cout[3]);
	Full_Adder FA2 (pp0[30], pp1[29], pp2[28], S[4], Cout[4]);
	Full_Adder FA3 (pp3[27], pp4[26], pp5[25], S[5], Cout[5]);
	Half_Adder HA3 (pp6[24], pp7[23], S[6], Cout[6]);
	Full_Adder FA4 (pp0[31], pp1[30], pp2[29], S[7], Cout[7]);
	Full_Adder FA5 (pp3[28], pp4[27], pp5[26], S[8], Cout[8]);
	Full_Adder FA6 (pp6[25], pp7[24], pp8[23], S[9], Cout[9]);
	Half_Adder HA4 (pp9[22], pp10[21], S[10], Cout[10]);
	Full_Adder FA7 (pp1[31], pp2[30], pp3[29], S[11], Cout[11]);
	Full_Adder FA8 (pp4[28], pp5[27], pp6[26], S[12], Cout[12]);
	Full_Adder FA9 (pp7[25], pp8[24], pp9[23], S[13], Cout[13]);
	Half_Adder HA5 (pp10[22], pp11[21], S[14], Cout[14]);
	Full_Adder FA10 (pp2[31], pp3[30], pp4[29], S[15], Cout[15]);
	Full_Adder FA11 (pp5[28], pp6[27], pp7[26], S[16], Cout[16]);
	Full_Adder FA12 (pp8[25], pp9[24], pp10[23], S[17], Cout[17]);
	Full_Adder FA13 (pp3[31], pp4[30], pp5[29], S[18], Cout[18]);
	Full_Adder FA14 (pp6[28], pp7[27], pp8[26], S[19], Cout[19]);
	Full_Adder FA15 (pp4[31], pp5[30], pp6[29], S[20], Cout[20]);
	Half_Adder HA6 (pp0[19], pp1[18], S[21], Cout[21]);
	Full_Adder FA16 (pp0[20], pp1[19], pp2[18], S[22], Cout[22]);
	Half_Adder HA7 (pp3[17], pp4[16], S[23], Cout[23]);
	Full_Adder FA17 (pp0[21], pp1[20], pp2[19], S[24], Cout[24]);
	Full_Adder FA18 (pp3[18], pp4[17], pp5[16], S[25], Cout[25]);
	Half_Adder HA8 (pp6[15], pp7[14], S[26], Cout[26]);
	Full_Adder FA19 (pp0[22], pp1[21], pp2[20], S[27], Cout[27]);
	Full_Adder FA20 (pp3[19], pp4[18], pp5[17], S[28], Cout[28]);
	Full_Adder FA21 (pp6[16], pp7[15], pp8[14], S[29], Cout[29]);
	Half_Adder HA9 (pp9[13], pp10[12], S[30], Cout[30]);
	Full_Adder FA22 (pp0[23], pp1[22], pp2[21], S[31], Cout[31]);
	Full_Adder FA23 (pp3[20], pp4[19], pp5[18], S[32], Cout[32]);
	Full_Adder FA24 (pp6[17], pp7[16], pp8[15], S[33], Cout[33]);
	Full_Adder FA25 (pp9[14], pp10[13], pp11[12], S[34], Cout[34]);
	Half_Adder HA10 (pp12[11], pp13[10], S[35], Cout[35]);
	Full_Adder FA26 (pp0[24], pp1[23], pp2[22], S[36], Cout[36]);
	Full_Adder FA27 (pp3[21], pp4[20], pp5[19], S[37], Cout[37]);
	Full_Adder FA28 (pp6[18], pp7[17], pp8[16], S[38], Cout[38]);
	Full_Adder FA29 (pp9[15], pp10[14], pp11[13], S[39], Cout[39]);
	Full_Adder FA30 (pp12[12], pp13[11], pp14[10], S[40], Cout[40]);
	Half_Adder HA11 (pp15[9], pp16[8], S[41], Cout[41]);
	Full_Adder FA31 (pp0[25], pp1[24], pp2[23], S[42], Cout[42]);
	Full_Adder FA32 (pp3[22], pp4[21], pp5[20], S[43], Cout[43]);
	Full_Adder FA33 (pp6[19], pp7[18], pp8[17], S[44], Cout[44]);
	Full_Adder FA34 (pp9[16], pp10[15], pp11[14], S[45], Cout[45]);
	Full_Adder FA35 (pp12[13], pp13[12], pp14[11], S[46], Cout[46]);
	Full_Adder FA36 (pp15[10], pp16[9], pp17[8], S[47], Cout[47]);
	Half_Adder HA12 (pp18[7], pp19[6], S[48], Cout[48]);
	Full_Adder FA37 (pp0[26], pp1[25], pp2[24], S[49], Cout[49]);
	Full_Adder FA38 (pp3[23], pp4[22], pp5[21], S[50], Cout[50]);
	Full_Adder FA39 (pp6[20], pp7[19], pp8[18], S[51], Cout[51]);
	Full_Adder FA40 (pp9[17], pp10[16], pp11[15], S[52], Cout[52]);
	Full_Adder FA41 (pp12[14], pp13[13], pp14[12], S[53], Cout[53]);
	Full_Adder FA42 (pp15[11], pp16[10], pp17[9], S[54], Cout[54]);
	Full_Adder FA43 (pp18[8], pp19[7], pp20[6], S[55], Cout[55]);
	Half_Adder HA13 (pp21[5], pp22[4], S[56], Cout[56]);
	Full_Adder FA44 (pp0[27], pp1[26], pp2[25], S[57], Cout[57]);
	Full_Adder FA45 (pp3[24], pp4[23], pp5[22], S[58], Cout[58]);
	Full_Adder FA46 (pp6[21], pp7[20], pp8[19], S[59], Cout[59]);
	Full_Adder FA47 (pp9[18], pp10[17], pp11[16], S[60], Cout[60]);
	Full_Adder FA48 (pp12[15], pp13[14], pp14[13], S[61], Cout[61]);
	Full_Adder FA49 (pp15[12], pp16[11], pp17[10], S[62], Cout[62]);
	Full_Adder FA50 (pp18[9], pp19[8], pp20[7], S[63], Cout[63]);
	Full_Adder FA51 (pp21[6], pp22[5], pp23[4], S[64], Cout[64]);
	Half_Adder HA14 (pp24[3], pp25[2], S[65], Cout[65]);
	Full_Adder FA52 (pp2[26], pp3[25], pp4[24], S[66], Cout[66]);
	Full_Adder FA53 (pp5[23], pp6[22], pp7[21], S[67], Cout[67]);
	Full_Adder FA54 (pp8[20], pp9[19], pp10[18], S[68], Cout[68]);
	Full_Adder FA55 (pp11[17], pp12[16], pp13[15], S[69], Cout[69]);
	Full_Adder FA56 (pp14[14], pp15[13], pp16[12], S[70], Cout[70]);
	Full_Adder FA57 (pp17[11], pp18[10], pp19[9], S[71], Cout[71]);
	Full_Adder FA58 (pp20[8], pp21[7], pp22[6], S[72], Cout[72]);
	Full_Adder FA59 (pp23[5], pp24[4], pp25[3], S[73], Cout[73]);
	Full_Adder FA60 (pp26[2], pp27[1], pp28[0], S[74], Cout[74]);
	Full_Adder FA61 (pp5[24], pp6[23], pp7[22], S[75], Cout[75]);
	Full_Adder FA62 (pp8[21], pp9[20], pp10[19], S[76], Cout[76]);
	Full_Adder FA63 (pp11[18], pp12[17], pp13[16], S[77], Cout[77]);
	Full_Adder FA64 (pp14[15], pp15[14], pp16[13], S[78], Cout[78]);
	Full_Adder FA65 (pp17[12], pp18[11], pp19[10], S[79], Cout[79]);
	Full_Adder FA66 (pp20[9], pp21[8], pp22[7], S[80], Cout[80]);
	Full_Adder FA67 (pp23[6], pp24[5], pp25[4], S[81], Cout[81]);
	Full_Adder FA68 (pp26[3], pp27[2], pp28[1], S[82], Cout[82]);
	Full_Adder FA69 (pp29[0], Cout[1], S[2], S[83], Cout[83]);
	Full_Adder FA70 (pp8[22], pp9[21], pp10[20], S[84], Cout[84]);
	Full_Adder FA71 (pp11[19], pp12[18], pp13[17], S[85], Cout[85]);
	Full_Adder FA72 (pp14[16], pp15[15], pp16[14], S[86], Cout[86]);
	Full_Adder FA73 (pp17[13], pp18[12], pp19[11], S[87], Cout[87]);
	Full_Adder FA74 (pp20[10], pp21[9], pp22[8], S[88], Cout[88]);
	Full_Adder FA75 (pp23[7], pp24[6], pp25[5], S[89], Cout[89]);
	Full_Adder FA76 (pp26[4], pp27[3], pp28[2], S[90], Cout[90]);
	Full_Adder FA77 (pp29[1], pp30[0], Cout[2], S[91], Cout[91]);
	Full_Adder FA78 (Cout[3], S[4], S[5], S[92], Cout[92]);
	Full_Adder FA79 (pp11[20], pp12[19], pp13[18], S[93], Cout[93]);
	Full_Adder FA80 (pp14[17], pp15[16], pp16[15], S[94], Cout[94]);
	Full_Adder FA81 (pp17[14], pp18[13], pp19[12], S[95], Cout[95]);
	Full_Adder FA82 (pp20[11], pp21[10], pp22[9], S[96], Cout[96]);
	Full_Adder FA83 (pp23[8], pp24[7], pp25[6], S[97], Cout[97]);
	Full_Adder FA84 (pp26[5], pp27[4], pp28[3], S[98], Cout[98]);
	Full_Adder FA85 (pp29[2], pp30[1], pp31[0], S[99], Cout[99]);
	Full_Adder FA86 (Cout[4], Cout[5], Cout[6], S[100], Cout[100]);
	Full_Adder FA87 (S[7], S[8], S[9], S[101], Cout[101]);
	Full_Adder FA88 (pp12[20], pp13[19], pp14[18], S[102], Cout[102]);
	Full_Adder FA89 (pp15[17], pp16[16], pp17[15], S[103], Cout[103]);
	Full_Adder FA90 (pp18[14], pp19[13], pp20[12], S[104], Cout[104]);
	Full_Adder FA91 (pp21[11], pp22[10], pp23[9], S[105], Cout[105]);
	Full_Adder FA92 (pp24[8], pp25[7], pp26[6], S[106], Cout[106]);
	Full_Adder FA93 (pp27[5], pp28[4], pp29[3], S[107], Cout[107]);
	Full_Adder FA94 (pp30[2], pp31[1], Cout[7], S[108], Cout[108]);
	Full_Adder FA95 (Cout[8], Cout[9], Cout[10], S[109], Cout[109]);
	Full_Adder FA96 (S[11], S[12], S[13], S[110], Cout[110]);
	Full_Adder FA97 (pp11[22], pp12[21], pp13[20], S[111], Cout[111]);
	Full_Adder FA98 (pp14[19], pp15[18], pp16[17], S[112], Cout[112]);
	Full_Adder FA99 (pp17[16], pp18[15], pp19[14], S[113], Cout[113]);
	Full_Adder FA100 (pp20[13], pp21[12], pp22[11], S[114], Cout[114]);
	Full_Adder FA101 (pp23[10], pp24[9], pp25[8], S[115], Cout[115]);
	Full_Adder FA102 (pp26[7], pp27[6], pp28[5], S[116], Cout[116]);
	Full_Adder FA103 (pp29[4], pp30[3], pp31[2], S[117], Cout[117]);
	Full_Adder FA104 (Cout[11], Cout[12], Cout[13], S[118], Cout[118]);
	Full_Adder FA105 (Cout[14], S[15], S[16], S[119], Cout[119]);
	Full_Adder FA106 (pp9[25], pp10[24], pp11[23], S[120], Cout[120]);
	Full_Adder FA107 (pp12[22], pp13[21], pp14[20], S[121], Cout[121]);
	Full_Adder FA108 (pp15[19], pp16[18], pp17[17], S[122], Cout[122]);
	Full_Adder FA109 (pp18[16], pp19[15], pp20[14], S[123], Cout[123]);
	Full_Adder FA110 (pp21[13], pp22[12], pp23[11], S[124], Cout[124]);
	Full_Adder FA111 (pp24[10], pp25[9], pp26[8], S[125], Cout[125]);
	Full_Adder FA112 (pp27[7], pp28[6], pp29[5], S[126], Cout[126]);
	Full_Adder FA113 (pp30[4], pp31[3], Cout[15], S[127], Cout[127]);
	Full_Adder FA114 (Cout[16], Cout[17], S[18], S[128], Cout[128]);
	Full_Adder FA115 (pp7[28], pp8[27], pp9[26], S[129], Cout[129]);
	Full_Adder FA116 (pp10[25], pp11[24], pp12[23], S[130], Cout[130]);
	Full_Adder FA117 (pp13[22], pp14[21], pp15[20], S[131], Cout[131]);
	Full_Adder FA118 (pp16[19], pp17[18], pp18[17], S[132], Cout[132]);
	Full_Adder FA119 (pp19[16], pp20[15], pp21[14], S[133], Cout[133]);
	Full_Adder FA120 (pp22[13], pp23[12], pp24[11], S[134], Cout[134]);
	Full_Adder FA121 (pp25[10], pp26[9], pp27[8], S[135], Cout[135]);
	Full_Adder FA122 (pp28[7], pp29[6], pp30[5], S[136], Cout[136]);
	Full_Adder FA123 (pp31[4], Cout[18], Cout[19], S[137], Cout[137]);
	Full_Adder FA124 (pp5[31], pp6[30], pp7[29], S[138], Cout[138]);
	Full_Adder FA125 (pp8[28], pp9[27], pp10[26], S[139], Cout[139]);
	Full_Adder FA126 (pp11[25], pp12[24], pp13[23], S[140], Cout[140]);
	Full_Adder FA127 (pp14[22], pp15[21], pp16[20], S[141], Cout[141]);
	Full_Adder FA128 (pp17[19], pp18[18], pp19[17], S[142], Cout[142]);
	Full_Adder FA129 (pp20[16], pp21[15], pp22[14], S[143], Cout[143]);
	Full_Adder FA130 (pp23[13], pp24[12], pp25[11], S[144], Cout[144]);
	Full_Adder FA131 (pp26[10], pp27[9], pp28[8], S[145], Cout[145]);
	Full_Adder FA132 (pp29[7], pp30[6], pp31[5], S[146], Cout[146]);
	Full_Adder FA133 (pp6[31], pp7[30], pp8[29], S[147], Cout[147]);
	Full_Adder FA134 (pp9[28], pp10[27], pp11[26], S[148], Cout[148]);
	Full_Adder FA135 (pp12[25], pp13[24], pp14[23], S[149], Cout[149]);
	Full_Adder FA136 (pp15[22], pp16[21], pp17[20], S[150], Cout[150]);
	Full_Adder FA137 (pp18[19], pp19[18], pp20[17], S[151], Cout[151]);
	Full_Adder FA138 (pp21[16], pp22[15], pp23[14], S[152], Cout[152]);
	Full_Adder FA139 (pp24[13], pp25[12], pp26[11], S[153], Cout[153]);
	Full_Adder FA140 (pp27[10], pp28[9], pp29[8], S[154], Cout[154]);
	Full_Adder FA141 (pp7[31], pp8[30], pp9[29], S[155], Cout[155]);
	Full_Adder FA142 (pp10[28], pp11[27], pp12[26], S[156], Cout[156]);
	Full_Adder FA143 (pp13[25], pp14[24], pp15[23], S[157], Cout[157]);
	Full_Adder FA144 (pp16[22], pp17[21], pp18[20], S[158], Cout[158]);
	Full_Adder FA145 (pp19[19], pp20[18], pp21[17], S[159], Cout[159]);
	Full_Adder FA146 (pp22[16], pp23[15], pp24[14], S[160], Cout[160]);
	Full_Adder FA147 (pp25[13], pp26[12], pp27[11], S[161], Cout[161]);
	Full_Adder FA148 (pp8[31], pp9[30], pp10[29], S[162], Cout[162]);
	Full_Adder FA149 (pp11[28], pp12[27], pp13[26], S[163], Cout[163]);
	Full_Adder FA150 (pp14[25], pp15[24], pp16[23], S[164], Cout[164]);
	Full_Adder FA151 (pp17[22], pp18[21], pp19[20], S[165], Cout[165]);
	Full_Adder FA152 (pp20[19], pp21[18], pp22[17], S[166], Cout[166]);
	Full_Adder FA153 (pp23[16], pp24[15], pp25[14], S[167], Cout[167]);
	Full_Adder FA154 (pp9[31], pp10[30], pp11[29], S[168], Cout[168]);
	Full_Adder FA155 (pp12[28], pp13[27], pp14[26], S[169], Cout[169]);
	Full_Adder FA156 (pp15[25], pp16[24], pp17[23], S[170], Cout[170]);
	Full_Adder FA157 (pp18[22], pp19[21], pp20[20], S[171], Cout[171]);
	Full_Adder FA158 (pp21[19], pp22[18], pp23[17], S[172], Cout[172]);
	Full_Adder FA159 (pp10[31], pp11[30], pp12[29], S[173], Cout[173]);
	Full_Adder FA160 (pp13[28], pp14[27], pp15[26], S[174], Cout[174]);
	Full_Adder FA161 (pp16[25], pp17[24], pp18[23], S[175], Cout[175]);
	Full_Adder FA162 (pp19[22], pp20[21], pp21[20], S[176], Cout[176]);
	Full_Adder FA163 (pp11[31], pp12[30], pp13[29], S[177], Cout[177]);
	Full_Adder FA164 (pp14[28], pp15[27], pp16[26], S[178], Cout[178]);
	Full_Adder FA165 (pp17[25], pp18[24], pp19[23], S[179], Cout[179]);
	Full_Adder FA166 (pp12[31], pp13[30], pp14[29], S[180], Cout[180]);
	Full_Adder FA167 (pp15[28], pp16[27], pp17[26], S[181], Cout[181]);
	Full_Adder FA168 (pp13[31], pp14[30], pp15[29], S[182], Cout[182]);
	Half_Adder HA15 (pp0[13], pp1[12], S[183], Cout[183]);
	Full_Adder FA169 (pp0[14], pp1[13], pp2[12], S[184], Cout[184]);
	Half_Adder HA16 (pp3[11], pp4[10], S[185], Cout[185]);
	Full_Adder FA170 (pp0[15], pp1[14], pp2[13], S[186], Cout[186]);
	Full_Adder FA171 (pp3[12], pp4[11], pp5[10], S[187], Cout[187]);
	Half_Adder HA17 (pp6[9], pp7[8], S[188], Cout[188]);
	Full_Adder FA172 (pp0[16], pp1[15], pp2[14], S[189], Cout[189]);
	Full_Adder FA173 (pp3[13], pp4[12], pp5[11], S[190], Cout[190]);
	Full_Adder FA174 (pp6[10], pp7[9], pp8[8], S[191], Cout[191]);
	Half_Adder HA18 (pp9[7], pp10[6], S[192], Cout[192]);
	Full_Adder FA175 (pp0[17], pp1[16], pp2[15], S[193], Cout[193]);
	Full_Adder FA176 (pp3[14], pp4[13], pp5[12], S[194], Cout[194]);
	Full_Adder FA177 (pp6[11], pp7[10], pp8[9], S[195], Cout[195]);
	Full_Adder FA178 (pp9[8], pp10[7], pp11[6], S[196], Cout[196]);
	Half_Adder HA19 (pp12[5], pp13[4], S[197], Cout[197]);
	Full_Adder FA179 (pp0[18], pp1[17], pp2[16], S[198], Cout[198]);
	Full_Adder FA180 (pp3[15], pp4[14], pp5[13], S[199], Cout[199]);
	Full_Adder FA181 (pp6[12], pp7[11], pp8[10], S[200], Cout[200]);
	Full_Adder FA182 (pp9[9], pp10[8], pp11[7], S[201], Cout[201]);
	Full_Adder FA183 (pp12[6], pp13[5], pp14[4], S[202], Cout[202]);
	Half_Adder HA20 (pp15[3], pp16[2], S[203], Cout[203]);
	Full_Adder FA184 (pp2[17], pp3[16], pp4[15], S[204], Cout[204]);
	Full_Adder FA185 (pp5[14], pp6[13], pp7[12], S[205], Cout[205]);
	Full_Adder FA186 (pp8[11], pp9[10], pp10[9], S[206], Cout[206]);
	Full_Adder FA187 (pp11[8], pp12[7], pp13[6], S[207], Cout[207]);
	Full_Adder FA188 (pp14[5], pp15[4], pp16[3], S[208], Cout[208]);
	Full_Adder FA189 (pp17[2], pp18[1], pp19[0], S[209], Cout[209]);
	Full_Adder FA190 (pp5[15], pp6[14], pp7[13], S[210], Cout[210]);
	Full_Adder FA191 (pp8[12], pp9[11], pp10[10], S[211], Cout[211]);
	Full_Adder FA192 (pp11[9], pp12[8], pp13[7], S[212], Cout[212]);
	Full_Adder FA193 (pp14[6], pp15[5], pp16[4], S[213], Cout[213]);
	Full_Adder FA194 (pp17[3], pp18[2], pp19[1], S[214], Cout[214]);
	Full_Adder FA195 (pp20[0], Cout[21], S[22], S[215], Cout[215]);
	Full_Adder FA196 (pp8[13], pp9[12], pp10[11], S[216], Cout[216]);
	Full_Adder FA197 (pp11[10], pp12[9], pp13[8], S[217], Cout[217]);
	Full_Adder FA198 (pp14[7], pp15[6], pp16[5], S[218], Cout[218]);
	Full_Adder FA199 (pp17[4], pp18[3], pp19[2], S[219], Cout[219]);
	Full_Adder FA200 (pp20[1], pp21[0], Cout[22], S[220], Cout[220]);
	Full_Adder FA201 (Cout[23], S[24], S[25], S[221], Cout[221]);
	Full_Adder FA202 (pp11[11], pp12[10], pp13[9], S[222], Cout[222]);
	Full_Adder FA203 (pp14[8], pp15[7], pp16[6], S[223], Cout[223]);
	Full_Adder FA204 (pp17[5], pp18[4], pp19[3], S[224], Cout[224]);
	Full_Adder FA205 (pp20[2], pp21[1], pp22[0], S[225], Cout[225]);
	Full_Adder FA206 (Cout[24], Cout[25], Cout[26], S[226], Cout[226]);
	Full_Adder FA207 (S[27], S[28], S[29], S[227], Cout[227]);
	Full_Adder FA208 (pp14[9], pp15[8], pp16[7], S[228], Cout[228]);
	Full_Adder FA209 (pp17[6], pp18[5], pp19[4], S[229], Cout[229]);
	Full_Adder FA210 (pp20[3], pp21[2], pp22[1], S[230], Cout[230]);
	Full_Adder FA211 (pp23[0], Cout[27], Cout[28], S[231], Cout[231]);
	Full_Adder FA212 (Cout[29], Cout[30], S[31], S[232], Cout[232]);
	Full_Adder FA213 (S[32], S[33], S[34], S[233], Cout[233]);
	Full_Adder FA214 (pp17[7], pp18[6], pp19[5], S[234], Cout[234]);
	Full_Adder FA215 (pp20[4], pp21[3], pp22[2], S[235], Cout[235]);
	Full_Adder FA216 (pp23[1], pp24[0], Cout[31], S[236], Cout[236]);
	Full_Adder FA217 (Cout[32], Cout[33], Cout[34], S[237], Cout[237]);
	Full_Adder FA218 (Cout[35], S[36], S[37], S[238], Cout[238]);
	Full_Adder FA219 (S[38], S[39], S[40], S[239], Cout[239]);
	Full_Adder FA220 (pp20[5], pp21[4], pp22[3], S[240], Cout[240]);
	Full_Adder FA221 (pp23[2], pp24[1], pp25[0], S[241], Cout[241]);
	Full_Adder FA222 (Cout[36], Cout[37], Cout[38], S[242], Cout[242]);
	Full_Adder FA223 (Cout[39], Cout[40], Cout[41], S[243], Cout[243]);
	Full_Adder FA224 (S[42], S[43], S[44], S[244], Cout[244]);
	Full_Adder FA225 (S[45], S[46], S[47], S[245], Cout[245]);
	Full_Adder FA226 (pp23[3], pp24[2], pp25[1], S[246], Cout[246]);
	Full_Adder FA227 (pp26[0], Cout[42], Cout[43], S[247], Cout[247]);
	Full_Adder FA228 (Cout[44], Cout[45], Cout[46], S[248], Cout[248]);
	Full_Adder FA229 (Cout[47], Cout[48], S[49], S[249], Cout[249]);
	Full_Adder FA230 (S[50], S[51], S[52], S[250], Cout[250]);
	Full_Adder FA231 (S[53], S[54], S[55], S[251], Cout[251]);
	Full_Adder FA232 (pp26[1], pp27[0], Cout[49], S[252], Cout[252]);
	Full_Adder FA233 (Cout[50], Cout[51], Cout[52], S[253], Cout[253]);
	Full_Adder FA234 (Cout[53], Cout[54], Cout[55], S[254], Cout[254]);
	Full_Adder FA235 (Cout[56], S[57], S[58], S[255], Cout[255]);
	Full_Adder FA236 (S[59], S[60], S[61], S[256], Cout[256]);
	Full_Adder FA237 (S[62], S[63], S[64], S[257], Cout[257]);
	Full_Adder FA238 (S[1], Cout[57], Cout[58], S[258], Cout[258]);
	Full_Adder FA239 (Cout[59], Cout[60], Cout[61], S[259], Cout[259]);
	Full_Adder FA240 (Cout[62], Cout[63], Cout[64], S[260], Cout[260]);
	Full_Adder FA241 (Cout[65], S[66], S[67], S[261], Cout[261]);
	Full_Adder FA242 (S[68], S[69], S[70], S[262], Cout[262]);
	Full_Adder FA243 (S[71], S[72], S[73], S[263], Cout[263]);
	Full_Adder FA244 (S[3], Cout[66], Cout[67], S[264], Cout[264]);
	Full_Adder FA245 (Cout[68], Cout[69], Cout[70], S[265], Cout[265]);
	Full_Adder FA246 (Cout[71], Cout[72], Cout[73], S[266], Cout[266]);
	Full_Adder FA247 (Cout[74], S[75], S[76], S[267], Cout[267]);
	Full_Adder FA248 (S[77], S[78], S[79], S[268], Cout[268]);
	Full_Adder FA249 (S[80], S[81], S[82], S[269], Cout[269]);
	Full_Adder FA250 (S[6], Cout[75], Cout[76], S[270], Cout[270]);
	Full_Adder FA251 (Cout[77], Cout[78], Cout[79], S[271], Cout[271]);
	Full_Adder FA252 (Cout[80], Cout[81], Cout[82], S[272], Cout[272]);
	Full_Adder FA253 (Cout[83], S[84], S[85], S[273], Cout[273]);
	Full_Adder FA254 (S[86], S[87], S[88], S[274], Cout[274]);
	Full_Adder FA255 (S[89], S[90], S[91], S[275], Cout[275]);
	Full_Adder FA256 (S[10], Cout[84], Cout[85], S[276], Cout[276]);
	Full_Adder FA257 (Cout[86], Cout[87], Cout[88], S[277], Cout[277]);
	Full_Adder FA258 (Cout[89], Cout[90], Cout[91], S[278], Cout[278]);
	Full_Adder FA259 (Cout[92], S[93], S[94], S[279], Cout[279]);
	Full_Adder FA260 (S[95], S[96], S[97], S[280], Cout[280]);
	Full_Adder FA261 (S[98], S[99], S[100], S[281], Cout[281]);
	Full_Adder FA262 (S[14], Cout[93], Cout[94], S[282], Cout[282]);
	Full_Adder FA263 (Cout[95], Cout[96], Cout[97], S[283], Cout[283]);
	Full_Adder FA264 (Cout[98], Cout[99], Cout[100], S[284], Cout[284]);
	Full_Adder FA265 (Cout[101], S[102], S[103], S[285], Cout[285]);
	Full_Adder FA266 (S[104], S[105], S[106], S[286], Cout[286]);
	Full_Adder FA267 (S[107], S[108], S[109], S[287], Cout[287]);
	Full_Adder FA268 (S[17], Cout[102], Cout[103], S[288], Cout[288]);
	Full_Adder FA269 (Cout[104], Cout[105], Cout[106], S[289], Cout[289]);
	Full_Adder FA270 (Cout[107], Cout[108], Cout[109], S[290], Cout[290]);
	Full_Adder FA271 (Cout[110], S[111], S[112], S[291], Cout[291]);
	Full_Adder FA272 (S[113], S[114], S[115], S[292], Cout[292]);
	Full_Adder FA273 (S[116], S[117], S[118], S[293], Cout[293]);
	Full_Adder FA274 (S[19], Cout[111], Cout[112], S[294], Cout[294]);
	Full_Adder FA275 (Cout[113], Cout[114], Cout[115], S[295], Cout[295]);
	Full_Adder FA276 (Cout[116], Cout[117], Cout[118], S[296], Cout[296]);
	Full_Adder FA277 (Cout[119], S[120], S[121], S[297], Cout[297]);
	Full_Adder FA278 (S[122], S[123], S[124], S[298], Cout[298]);
	Full_Adder FA279 (S[125], S[126], S[127], S[299], Cout[299]);
	Full_Adder FA280 (S[20], Cout[120], Cout[121], S[300], Cout[300]);
	Full_Adder FA281 (Cout[122], Cout[123], Cout[124], S[301], Cout[301]);
	Full_Adder FA282 (Cout[125], Cout[126], Cout[127], S[302], Cout[302]);
	Full_Adder FA283 (Cout[128], S[129], S[130], S[303], Cout[303]);
	Full_Adder FA284 (S[131], S[132], S[133], S[304], Cout[304]);
	Full_Adder FA285 (S[134], S[135], S[136], S[305], Cout[305]);
	Full_Adder FA286 (Cout[20], Cout[129], Cout[130], S[306], Cout[306]);
	Full_Adder FA287 (Cout[131], Cout[132], Cout[133], S[307], Cout[307]);
	Full_Adder FA288 (Cout[134], Cout[135], Cout[136], S[308], Cout[308]);
	Full_Adder FA289 (Cout[137], S[138], S[139], S[309], Cout[309]);
	Full_Adder FA290 (S[140], S[141], S[142], S[310], Cout[310]);
	Full_Adder FA291 (S[143], S[144], S[145], S[311], Cout[311]);
	Full_Adder FA292 (pp30[7], pp31[6], Cout[138], S[312], Cout[312]);
	Full_Adder FA293 (Cout[139], Cout[140], Cout[141], S[313], Cout[313]);
	Full_Adder FA294 (Cout[142], Cout[143], Cout[144], S[314], Cout[314]);
	Full_Adder FA295 (Cout[145], Cout[146], S[147], S[315], Cout[315]);
	Full_Adder FA296 (S[148], S[149], S[150], S[316], Cout[316]);
	Full_Adder FA297 (S[151], S[152], S[153], S[317], Cout[317]);
	Full_Adder FA298 (pp28[10], pp29[9], pp30[8], S[318], Cout[318]);
	Full_Adder FA299 (pp31[7], Cout[147], Cout[148], S[319], Cout[319]);
	Full_Adder FA300 (Cout[149], Cout[150], Cout[151], S[320], Cout[320]);
	Full_Adder FA301 (Cout[152], Cout[153], Cout[154], S[321], Cout[321]);
	Full_Adder FA302 (S[155], S[156], S[157], S[322], Cout[322]);
	Full_Adder FA303 (S[158], S[159], S[160], S[323], Cout[323]);
	Full_Adder FA304 (pp26[13], pp27[12], pp28[11], S[324], Cout[324]);
	Full_Adder FA305 (pp29[10], pp30[9], pp31[8], S[325], Cout[325]);
	Full_Adder FA306 (Cout[155], Cout[156], Cout[157], S[326], Cout[326]);
	Full_Adder FA307 (Cout[158], Cout[159], Cout[160], S[327], Cout[327]);
	Full_Adder FA308 (Cout[161], S[162], S[163], S[328], Cout[328]);
	Full_Adder FA309 (S[164], S[165], S[166], S[329], Cout[329]);
	Full_Adder FA310 (pp24[16], pp25[15], pp26[14], S[330], Cout[330]);
	Full_Adder FA311 (pp27[13], pp28[12], pp29[11], S[331], Cout[331]);
	Full_Adder FA312 (pp30[10], pp31[9], Cout[162], S[332], Cout[332]);
	Full_Adder FA313 (Cout[163], Cout[164], Cout[165], S[333], Cout[333]);
	Full_Adder FA314 (Cout[166], Cout[167], S[168], S[334], Cout[334]);
	Full_Adder FA315 (S[169], S[170], S[171], S[335], Cout[335]);
	Full_Adder FA316 (pp22[19], pp23[18], pp24[17], S[336], Cout[336]);
	Full_Adder FA317 (pp25[16], pp26[15], pp27[14], S[337], Cout[337]);
	Full_Adder FA318 (pp28[13], pp29[12], pp30[11], S[338], Cout[338]);
	Full_Adder FA319 (pp31[10], Cout[168], Cout[169], S[339], Cout[339]);
	Full_Adder FA320 (Cout[170], Cout[171], Cout[172], S[340], Cout[340]);
	Full_Adder FA321 (S[173], S[174], S[175], S[341], Cout[341]);
	Full_Adder FA322 (pp20[22], pp21[21], pp22[20], S[342], Cout[342]);
	Full_Adder FA323 (pp23[19], pp24[18], pp25[17], S[343], Cout[343]);
	Full_Adder FA324 (pp26[16], pp27[15], pp28[14], S[344], Cout[344]);
	Full_Adder FA325 (pp29[13], pp30[12], pp31[11], S[345], Cout[345]);
	Full_Adder FA326 (Cout[173], Cout[174], Cout[175], S[346], Cout[346]);
	Full_Adder FA327 (Cout[176], S[177], S[178], S[347], Cout[347]);
	Full_Adder FA328 (pp18[25], pp19[24], pp20[23], S[348], Cout[348]);
	Full_Adder FA329 (pp21[22], pp22[21], pp23[20], S[349], Cout[349]);
	Full_Adder FA330 (pp24[19], pp25[18], pp26[17], S[350], Cout[350]);
	Full_Adder FA331 (pp27[16], pp28[15], pp29[14], S[351], Cout[351]);
	Full_Adder FA332 (pp30[13], pp31[12], Cout[177], S[352], Cout[352]);
	Full_Adder FA333 (Cout[178], Cout[179], S[180], S[353], Cout[353]);
	Full_Adder FA334 (pp16[28], pp17[27], pp18[26], S[354], Cout[354]);
	Full_Adder FA335 (pp19[25], pp20[24], pp21[23], S[355], Cout[355]);
	Full_Adder FA336 (pp22[22], pp23[21], pp24[20], S[356], Cout[356]);
	Full_Adder FA337 (pp25[19], pp26[18], pp27[17], S[357], Cout[357]);
	Full_Adder FA338 (pp28[16], pp29[15], pp30[14], S[358], Cout[358]);
	Full_Adder FA339 (pp31[13], Cout[180], Cout[181], S[359], Cout[359]);
	Full_Adder FA340 (pp14[31], pp15[30], pp16[29], S[360], Cout[360]);
	Full_Adder FA341 (pp17[28], pp18[27], pp19[26], S[361], Cout[361]);
	Full_Adder FA342 (pp20[25], pp21[24], pp22[23], S[362], Cout[362]);
	Full_Adder FA343 (pp23[22], pp24[21], pp25[20], S[363], Cout[363]);
	Full_Adder FA344 (pp26[19], pp27[18], pp28[17], S[364], Cout[364]);
	Full_Adder FA345 (pp29[16], pp30[15], pp31[14], S[365], Cout[365]);
	Full_Adder FA346 (pp15[31], pp16[30], pp17[29], S[366], Cout[366]);
	Full_Adder FA347 (pp18[28], pp19[27], pp20[26], S[367], Cout[367]);
	Full_Adder FA348 (pp21[25], pp22[24], pp23[23], S[368], Cout[368]);
	Full_Adder FA349 (pp24[22], pp25[21], pp26[20], S[369], Cout[369]);
	Full_Adder FA350 (pp27[19], pp28[18], pp29[17], S[370], Cout[370]);
	Full_Adder FA351 (pp16[31], pp17[30], pp18[29], S[371], Cout[371]);
	Full_Adder FA352 (pp19[28], pp20[27], pp21[26], S[372], Cout[372]);
	Full_Adder FA353 (pp22[25], pp23[24], pp24[23], S[373], Cout[373]);
	Full_Adder FA354 (pp25[22], pp26[21], pp27[20], S[374], Cout[374]);
	Full_Adder FA355 (pp17[31], pp18[30], pp19[29], S[375], Cout[375]);
	Full_Adder FA356 (pp20[28], pp21[27], pp22[26], S[376], Cout[376]);
	Full_Adder FA357 (pp23[25], pp24[24], pp25[23], S[377], Cout[377]);
	Full_Adder FA358 (pp18[31], pp19[30], pp20[29], S[378], Cout[378]);
	Full_Adder FA359 (pp21[28], pp22[27], pp23[26], S[379], Cout[379]);
	Full_Adder FA360 (pp19[31], pp20[30], pp21[29], S[380], Cout[380]);
	Half_Adder HA21 (pp0[9], pp1[8], S[381], Cout[381]);
	Full_Adder FA361 (pp0[10], pp1[9], pp2[8], S[382], Cout[382]);
	Half_Adder HA22 (pp3[7], pp4[6], S[383], Cout[383]);
	Full_Adder FA362 (pp0[11], pp1[10], pp2[9], S[384], Cout[384]);
	Full_Adder FA363 (pp3[8], pp4[7], pp5[6], S[385], Cout[385]);
	Half_Adder HA23 (pp6[5], pp7[4], S[386], Cout[386]);
	Full_Adder FA364 (pp0[12], pp1[11], pp2[10], S[387], Cout[387]);
	Full_Adder FA365 (pp3[9], pp4[8], pp5[7], S[388], Cout[388]);
	Full_Adder FA366 (pp6[6], pp7[5], pp8[4], S[389], Cout[389]);
	Half_Adder HA24 (pp9[3], pp10[2], S[390], Cout[390]);
	Full_Adder FA367 (pp2[11], pp3[10], pp4[9], S[391], Cout[391]);
	Full_Adder FA368 (pp5[8], pp6[7], pp7[6], S[392], Cout[392]);
	Full_Adder FA369 (pp8[5], pp9[4], pp10[3], S[393], Cout[393]);
	Full_Adder FA370 (pp11[2], pp12[1], pp13[0], S[394], Cout[394]);
	Full_Adder FA371 (pp5[9], pp6[8], pp7[7], S[395], Cout[395]);
	Full_Adder FA372 (pp8[6], pp9[5], pp10[4], S[396], Cout[396]);
	Full_Adder FA373 (pp11[3], pp12[2], pp13[1], S[397], Cout[397]);
	Full_Adder FA374 (pp14[0], Cout[183], S[184], S[398], Cout[398]);
	Full_Adder FA375 (pp8[7], pp9[6], pp10[5], S[399], Cout[399]);
	Full_Adder FA376 (pp11[4], pp12[3], pp13[2], S[400], Cout[400]);
	Full_Adder FA377 (pp14[1], pp15[0], Cout[184], S[401], Cout[401]);
	Full_Adder FA378 (Cout[185], S[186], S[187], S[402], Cout[402]);
	Full_Adder FA379 (pp11[5], pp12[4], pp13[3], S[403], Cout[403]);
	Full_Adder FA380 (pp14[2], pp15[1], pp16[0], S[404], Cout[404]);
	Full_Adder FA381 (Cout[186], Cout[187], Cout[188], S[405], Cout[405]);
	Full_Adder FA382 (S[189], S[190], S[191], S[406], Cout[406]);
	Full_Adder FA383 (pp14[3], pp15[2], pp16[1], S[407], Cout[407]);
	Full_Adder FA384 (pp17[0], Cout[189], Cout[190], S[408], Cout[408]);
	Full_Adder FA385 (Cout[191], Cout[192], S[193], S[409], Cout[409]);
	Full_Adder FA386 (S[194], S[195], S[196], S[410], Cout[410]);
	Full_Adder FA387 (pp17[1], pp18[0], Cout[193], S[411], Cout[411]);
	Full_Adder FA388 (Cout[194], Cout[195], Cout[196], S[412], Cout[412]);
	Full_Adder FA389 (Cout[197], S[198], S[199], S[413], Cout[413]);
	Full_Adder FA390 (S[200], S[201], S[202], S[414], Cout[414]);
	Full_Adder FA391 (S[21], Cout[198], Cout[199], S[415], Cout[415]);
	Full_Adder FA392 (Cout[200], Cout[201], Cout[202], S[416], Cout[416]);
	Full_Adder FA393 (Cout[203], S[204], S[205], S[417], Cout[417]);
	Full_Adder FA394 (S[206], S[207], S[208], S[418], Cout[418]);
	Full_Adder FA395 (S[23], Cout[204], Cout[205], S[419], Cout[419]);
	Full_Adder FA396 (Cout[206], Cout[207], Cout[208], S[420], Cout[420]);
	Full_Adder FA397 (Cout[209], S[210], S[211], S[421], Cout[421]);
	Full_Adder FA398 (S[212], S[213], S[214], S[422], Cout[422]);
	Full_Adder FA399 (S[26], Cout[210], Cout[211], S[423], Cout[423]);
	Full_Adder FA400 (Cout[212], Cout[213], Cout[214], S[424], Cout[424]);
	Full_Adder FA401 (Cout[215], S[216], S[217], S[425], Cout[425]);
	Full_Adder FA402 (S[218], S[219], S[220], S[426], Cout[426]);
	Full_Adder FA403 (S[30], Cout[216], Cout[217], S[427], Cout[427]);
	Full_Adder FA404 (Cout[218], Cout[219], Cout[220], S[428], Cout[428]);
	Full_Adder FA405 (Cout[221], S[222], S[223], S[429], Cout[429]);
	Full_Adder FA406 (S[224], S[225], S[226], S[430], Cout[430]);
	Full_Adder FA407 (S[35], Cout[222], Cout[223], S[431], Cout[431]);
	Full_Adder FA408 (Cout[224], Cout[225], Cout[226], S[432], Cout[432]);
	Full_Adder FA409 (Cout[227], S[228], S[229], S[433], Cout[433]);
	Full_Adder FA410 (S[230], S[231], S[232], S[434], Cout[434]);
	Full_Adder FA411 (S[41], Cout[228], Cout[229], S[435], Cout[435]);
	Full_Adder FA412 (Cout[230], Cout[231], Cout[232], S[436], Cout[436]);
	Full_Adder FA413 (Cout[233], S[234], S[235], S[437], Cout[437]);
	Full_Adder FA414 (S[236], S[237], S[238], S[438], Cout[438]);
	Full_Adder FA415 (S[48], Cout[234], Cout[235], S[439], Cout[439]);
	Full_Adder FA416 (Cout[236], Cout[237], Cout[238], S[440], Cout[440]);
	Full_Adder FA417 (Cout[239], S[240], S[241], S[441], Cout[441]);
	Full_Adder FA418 (S[242], S[243], S[244], S[442], Cout[442]);
	Full_Adder FA419 (S[56], Cout[240], Cout[241], S[443], Cout[443]);
	Full_Adder FA420 (Cout[242], Cout[243], Cout[244], S[444], Cout[444]);
	Full_Adder FA421 (Cout[245], S[246], S[247], S[445], Cout[445]);
	Full_Adder FA422 (S[248], S[249], S[250], S[446], Cout[446]);
	Full_Adder FA423 (S[65], Cout[246], Cout[247], S[447], Cout[447]);
	Full_Adder FA424 (Cout[248], Cout[249], Cout[250], S[448], Cout[448]);
	Full_Adder FA425 (Cout[251], S[252], S[253], S[449], Cout[449]);
	Full_Adder FA426 (S[254], S[255], S[256], S[450], Cout[450]);
	Full_Adder FA427 (S[74], Cout[252], Cout[253], S[451], Cout[451]);
	Full_Adder FA428 (Cout[254], Cout[255], Cout[256], S[452], Cout[452]);
	Full_Adder FA429 (Cout[257], S[258], S[259], S[453], Cout[453]);
	Full_Adder FA430 (S[260], S[261], S[262], S[454], Cout[454]);
	Full_Adder FA431 (S[83], Cout[258], Cout[259], S[455], Cout[455]);
	Full_Adder FA432 (Cout[260], Cout[261], Cout[262], S[456], Cout[456]);
	Full_Adder FA433 (Cout[263], S[264], S[265], S[457], Cout[457]);
	Full_Adder FA434 (S[266], S[267], S[268], S[458], Cout[458]);
	Full_Adder FA435 (S[92], Cout[264], Cout[265], S[459], Cout[459]);
	Full_Adder FA436 (Cout[266], Cout[267], Cout[268], S[460], Cout[460]);
	Full_Adder FA437 (Cout[269], S[270], S[271], S[461], Cout[461]);
	Full_Adder FA438 (S[272], S[273], S[274], S[462], Cout[462]);
	Full_Adder FA439 (S[101], Cout[270], Cout[271], S[463], Cout[463]);
	Full_Adder FA440 (Cout[272], Cout[273], Cout[274], S[464], Cout[464]);
	Full_Adder FA441 (Cout[275], S[276], S[277], S[465], Cout[465]);
	Full_Adder FA442 (S[278], S[279], S[280], S[466], Cout[466]);
	Full_Adder FA443 (S[110], Cout[276], Cout[277], S[467], Cout[467]);
	Full_Adder FA444 (Cout[278], Cout[279], Cout[280], S[468], Cout[468]);
	Full_Adder FA445 (Cout[281], S[282], S[283], S[469], Cout[469]);
	Full_Adder FA446 (S[284], S[285], S[286], S[470], Cout[470]);
	Full_Adder FA447 (S[119], Cout[282], Cout[283], S[471], Cout[471]);
	Full_Adder FA448 (Cout[284], Cout[285], Cout[286], S[472], Cout[472]);
	Full_Adder FA449 (Cout[287], S[288], S[289], S[473], Cout[473]);
	Full_Adder FA450 (S[290], S[291], S[292], S[474], Cout[474]);
	Full_Adder FA451 (S[128], Cout[288], Cout[289], S[475], Cout[475]);
	Full_Adder FA452 (Cout[290], Cout[291], Cout[292], S[476], Cout[476]);
	Full_Adder FA453 (Cout[293], S[294], S[295], S[477], Cout[477]);
	Full_Adder FA454 (S[296], S[297], S[298], S[478], Cout[478]);
	Full_Adder FA455 (S[137], Cout[294], Cout[295], S[479], Cout[479]);
	Full_Adder FA456 (Cout[296], Cout[297], Cout[298], S[480], Cout[480]);
	Full_Adder FA457 (Cout[299], S[300], S[301], S[481], Cout[481]);
	Full_Adder FA458 (S[302], S[303], S[304], S[482], Cout[482]);
	Full_Adder FA459 (S[146], Cout[300], Cout[301], S[483], Cout[483]);
	Full_Adder FA460 (Cout[302], Cout[303], Cout[304], S[484], Cout[484]);
	Full_Adder FA461 (Cout[305], S[306], S[307], S[485], Cout[485]);
	Full_Adder FA462 (S[308], S[309], S[310], S[486], Cout[486]);
	Full_Adder FA463 (S[154], Cout[306], Cout[307], S[487], Cout[487]);
	Full_Adder FA464 (Cout[308], Cout[309], Cout[310], S[488], Cout[488]);
	Full_Adder FA465 (Cout[311], S[312], S[313], S[489], Cout[489]);
	Full_Adder FA466 (S[314], S[315], S[316], S[490], Cout[490]);
	Full_Adder FA467 (S[161], Cout[312], Cout[313], S[491], Cout[491]);
	Full_Adder FA468 (Cout[314], Cout[315], Cout[316], S[492], Cout[492]);
	Full_Adder FA469 (Cout[317], S[318], S[319], S[493], Cout[493]);
	Full_Adder FA470 (S[320], S[321], S[322], S[494], Cout[494]);
	Full_Adder FA471 (S[167], Cout[318], Cout[319], S[495], Cout[495]);
	Full_Adder FA472 (Cout[320], Cout[321], Cout[322], S[496], Cout[496]);
	Full_Adder FA473 (Cout[323], S[324], S[325], S[497], Cout[497]);
	Full_Adder FA474 (S[326], S[327], S[328], S[498], Cout[498]);
	Full_Adder FA475 (S[172], Cout[324], Cout[325], S[499], Cout[499]);
	Full_Adder FA476 (Cout[326], Cout[327], Cout[328], S[500], Cout[500]);
	Full_Adder FA477 (Cout[329], S[330], S[331], S[501], Cout[501]);
	Full_Adder FA478 (S[332], S[333], S[334], S[502], Cout[502]);
	Full_Adder FA479 (S[176], Cout[330], Cout[331], S[503], Cout[503]);
	Full_Adder FA480 (Cout[332], Cout[333], Cout[334], S[504], Cout[504]);
	Full_Adder FA481 (Cout[335], S[336], S[337], S[505], Cout[505]);
	Full_Adder FA482 (S[338], S[339], S[340], S[506], Cout[506]);
	Full_Adder FA483 (S[179], Cout[336], Cout[337], S[507], Cout[507]);
	Full_Adder FA484 (Cout[338], Cout[339], Cout[340], S[508], Cout[508]);
	Full_Adder FA485 (Cout[341], S[342], S[343], S[509], Cout[509]);
	Full_Adder FA486 (S[344], S[345], S[346], S[510], Cout[510]);
	Full_Adder FA487 (S[181], Cout[342], Cout[343], S[511], Cout[511]);
	Full_Adder FA488 (Cout[344], Cout[345], Cout[346], S[512], Cout[512]);
	Full_Adder FA489 (Cout[347], S[348], S[349], S[513], Cout[513]);
	Full_Adder FA490 (S[350], S[351], S[352], S[514], Cout[514]);
	Full_Adder FA491 (S[182], Cout[348], Cout[349], S[515], Cout[515]);
	Full_Adder FA492 (Cout[350], Cout[351], Cout[352], S[516], Cout[516]);
	Full_Adder FA493 (Cout[353], S[354], S[355], S[517], Cout[517]);
	Full_Adder FA494 (S[356], S[357], S[358], S[518], Cout[518]);
	Full_Adder FA495 (Cout[182], Cout[354], Cout[355], S[519], Cout[519]);
	Full_Adder FA496 (Cout[356], Cout[357], Cout[358], S[520], Cout[520]);
	Full_Adder FA497 (Cout[359], S[360], S[361], S[521], Cout[521]);
	Full_Adder FA498 (S[362], S[363], S[364], S[522], Cout[522]);
	Full_Adder FA499 (pp30[16], pp31[15], Cout[360], S[523], Cout[523]);
	Full_Adder FA500 (Cout[361], Cout[362], Cout[363], S[524], Cout[524]);
	Full_Adder FA501 (Cout[364], Cout[365], S[366], S[525], Cout[525]);
	Full_Adder FA502 (S[367], S[368], S[369], S[526], Cout[526]);
	Full_Adder FA503 (pp28[19], pp29[18], pp30[17], S[527], Cout[527]);
	Full_Adder FA504 (pp31[16], Cout[366], Cout[367], S[528], Cout[528]);
	Full_Adder FA505 (Cout[368], Cout[369], Cout[370], S[529], Cout[529]);
	Full_Adder FA506 (S[371], S[372], S[373], S[530], Cout[530]);
	Full_Adder FA507 (pp26[22], pp27[21], pp28[20], S[531], Cout[531]);
	Full_Adder FA508 (pp29[19], pp30[18], pp31[17], S[532], Cout[532]);
	Full_Adder FA509 (Cout[371], Cout[372], Cout[373], S[533], Cout[533]);
	Full_Adder FA510 (Cout[374], S[375], S[376], S[534], Cout[534]);
	Full_Adder FA511 (pp24[25], pp25[24], pp26[23], S[535], Cout[535]);
	Full_Adder FA512 (pp27[22], pp28[21], pp29[20], S[536], Cout[536]);
	Full_Adder FA513 (pp30[19], pp31[18], Cout[375], S[537], Cout[537]);
	Full_Adder FA514 (Cout[376], Cout[377], S[378], S[538], Cout[538]);
	Full_Adder FA515 (pp22[28], pp23[27], pp24[26], S[539], Cout[539]);
	Full_Adder FA516 (pp25[25], pp26[24], pp27[23], S[540], Cout[540]);
	Full_Adder FA517 (pp28[22], pp29[21], pp30[20], S[541], Cout[541]);
	Full_Adder FA518 (pp31[19], Cout[378], Cout[379], S[542], Cout[542]);
	Full_Adder FA519 (pp20[31], pp21[30], pp22[29], S[543], Cout[543]);
	Full_Adder FA520 (pp23[28], pp24[27], pp25[26], S[544], Cout[544]);
	Full_Adder FA521 (pp26[25], pp27[24], pp28[23], S[545], Cout[545]);
	Full_Adder FA522 (pp29[22], pp30[21], pp31[20], S[546], Cout[546]);
	Full_Adder FA523 (pp21[31], pp22[30], pp23[29], S[547], Cout[547]);
	Full_Adder FA524 (pp24[28], pp25[27], pp26[26], S[548], Cout[548]);
	Full_Adder FA525 (pp27[25], pp28[24], pp29[23], S[549], Cout[549]);
	Full_Adder FA526 (pp22[31], pp23[30], pp24[29], S[550], Cout[550]);
	Full_Adder FA527 (pp25[28], pp26[27], pp27[26], S[551], Cout[551]);
	Full_Adder FA528 (pp23[31], pp24[30], pp25[29], S[552], Cout[552]);
	Half_Adder HA25 (pp0[6], pp1[5], S[553], Cout[553]);
	Full_Adder FA529 (pp0[7], pp1[6], pp2[5], S[554], Cout[554]);
	Half_Adder HA26 (pp3[4], pp4[3], S[555], Cout[555]);
	Full_Adder FA530 (pp0[8], pp1[7], pp2[6], S[556], Cout[556]);
	Full_Adder FA531 (pp3[5], pp4[4], pp5[3], S[557], Cout[557]);
	Half_Adder HA27 (pp6[2], pp7[1], S[558], Cout[558]);
	Full_Adder FA532 (pp2[7], pp3[6], pp4[5], S[559], Cout[559]);
	Full_Adder FA533 (pp5[4], pp6[3], pp7[2], S[560], Cout[560]);
	Full_Adder FA534 (pp8[1], pp9[0], S[381], S[561], Cout[561]);
	Full_Adder FA535 (pp5[5], pp6[4], pp7[3], S[562], Cout[562]);
	Full_Adder FA536 (pp8[2], pp9[1], pp10[0], S[563], Cout[563]);
	Full_Adder FA537 (Cout[381], S[382], S[383], S[564], Cout[564]);
	Full_Adder FA538 (pp8[3], pp9[2], pp10[1], S[565], Cout[565]);
	Full_Adder FA539 (pp11[0], Cout[382], Cout[383], S[566], Cout[566]);
	Full_Adder FA540 (S[384], S[385], S[386], S[567], Cout[567]);
	Full_Adder FA541 (pp11[1], pp12[0], Cout[384], S[568], Cout[568]);
	Full_Adder FA542 (Cout[385], Cout[386], S[387], S[569], Cout[569]);
	Full_Adder FA543 (S[388], S[389], S[390], S[570], Cout[570]);
	Full_Adder FA544 (S[183], Cout[387], Cout[388], S[571], Cout[571]);
	Full_Adder FA545 (Cout[389], Cout[390], S[391], S[572], Cout[572]);
	Full_Adder FA546 (S[392], S[393], S[394], S[573], Cout[573]);
	Full_Adder FA547 (S[185], Cout[391], Cout[392], S[574], Cout[574]);
	Full_Adder FA548 (Cout[393], Cout[394], S[395], S[575], Cout[575]);
	Full_Adder FA549 (S[396], S[397], S[398], S[576], Cout[576]);
	Full_Adder FA550 (S[188], Cout[395], Cout[396], S[577], Cout[577]);
	Full_Adder FA551 (Cout[397], Cout[398], S[399], S[578], Cout[578]);
	Full_Adder FA552 (S[400], S[401], S[402], S[579], Cout[579]);
	Full_Adder FA553 (S[192], Cout[399], Cout[400], S[580], Cout[580]);
	Full_Adder FA554 (Cout[401], Cout[402], S[403], S[581], Cout[581]);
	Full_Adder FA555 (S[404], S[405], S[406], S[582], Cout[582]);
	Full_Adder FA556 (S[197], Cout[403], Cout[404], S[583], Cout[583]);
	Full_Adder FA557 (Cout[405], Cout[406], S[407], S[584], Cout[584]);
	Full_Adder FA558 (S[408], S[409], S[410], S[585], Cout[585]);
	Full_Adder FA559 (S[203], Cout[407], Cout[408], S[586], Cout[586]);
	Full_Adder FA560 (Cout[409], Cout[410], S[411], S[587], Cout[587]);
	Full_Adder FA561 (S[412], S[413], S[414], S[588], Cout[588]);
	Full_Adder FA562 (S[209], Cout[411], Cout[412], S[589], Cout[589]);
	Full_Adder FA563 (Cout[413], Cout[414], S[415], S[590], Cout[590]);
	Full_Adder FA564 (S[416], S[417], S[418], S[591], Cout[591]);
	Full_Adder FA565 (S[215], Cout[415], Cout[416], S[592], Cout[592]);
	Full_Adder FA566 (Cout[417], Cout[418], S[419], S[593], Cout[593]);
	Full_Adder FA567 (S[420], S[421], S[422], S[594], Cout[594]);
	Full_Adder FA568 (S[221], Cout[419], Cout[420], S[595], Cout[595]);
	Full_Adder FA569 (Cout[421], Cout[422], S[423], S[596], Cout[596]);
	Full_Adder FA570 (S[424], S[425], S[426], S[597], Cout[597]);
	Full_Adder FA571 (S[227], Cout[423], Cout[424], S[598], Cout[598]);
	Full_Adder FA572 (Cout[425], Cout[426], S[427], S[599], Cout[599]);
	Full_Adder FA573 (S[428], S[429], S[430], S[600], Cout[600]);
	Full_Adder FA574 (S[233], Cout[427], Cout[428], S[601], Cout[601]);
	Full_Adder FA575 (Cout[429], Cout[430], S[431], S[602], Cout[602]);
	Full_Adder FA576 (S[432], S[433], S[434], S[603], Cout[603]);
	Full_Adder FA577 (S[239], Cout[431], Cout[432], S[604], Cout[604]);
	Full_Adder FA578 (Cout[433], Cout[434], S[435], S[605], Cout[605]);
	Full_Adder FA579 (S[436], S[437], S[438], S[606], Cout[606]);
	Full_Adder FA580 (S[245], Cout[435], Cout[436], S[607], Cout[607]);
	Full_Adder FA581 (Cout[437], Cout[438], S[439], S[608], Cout[608]);
	Full_Adder FA582 (S[440], S[441], S[442], S[609], Cout[609]);
	Full_Adder FA583 (S[251], Cout[439], Cout[440], S[610], Cout[610]);
	Full_Adder FA584 (Cout[441], Cout[442], S[443], S[611], Cout[611]);
	Full_Adder FA585 (S[444], S[445], S[446], S[612], Cout[612]);
	Full_Adder FA586 (S[257], Cout[443], Cout[444], S[613], Cout[613]);
	Full_Adder FA587 (Cout[445], Cout[446], S[447], S[614], Cout[614]);
	Full_Adder FA588 (S[448], S[449], S[450], S[615], Cout[615]);
	Full_Adder FA589 (S[263], Cout[447], Cout[448], S[616], Cout[616]);
	Full_Adder FA590 (Cout[449], Cout[450], S[451], S[617], Cout[617]);
	Full_Adder FA591 (S[452], S[453], S[454], S[618], Cout[618]);
	Full_Adder FA592 (S[269], Cout[451], Cout[452], S[619], Cout[619]);
	Full_Adder FA593 (Cout[453], Cout[454], S[455], S[620], Cout[620]);
	Full_Adder FA594 (S[456], S[457], S[458], S[621], Cout[621]);
	Full_Adder FA595 (S[275], Cout[455], Cout[456], S[622], Cout[622]);
	Full_Adder FA596 (Cout[457], Cout[458], S[459], S[623], Cout[623]);
	Full_Adder FA597 (S[460], S[461], S[462], S[624], Cout[624]);
	Full_Adder FA598 (S[281], Cout[459], Cout[460], S[625], Cout[625]);
	Full_Adder FA599 (Cout[461], Cout[462], S[463], S[626], Cout[626]);
	Full_Adder FA600 (S[464], S[465], S[466], S[627], Cout[627]);
	Full_Adder FA601 (S[287], Cout[463], Cout[464], S[628], Cout[628]);
	Full_Adder FA602 (Cout[465], Cout[466], S[467], S[629], Cout[629]);
	Full_Adder FA603 (S[468], S[469], S[470], S[630], Cout[630]);
	Full_Adder FA604 (S[293], Cout[467], Cout[468], S[631], Cout[631]);
	Full_Adder FA605 (Cout[469], Cout[470], S[471], S[632], Cout[632]);
	Full_Adder FA606 (S[472], S[473], S[474], S[633], Cout[633]);
	Full_Adder FA607 (S[299], Cout[471], Cout[472], S[634], Cout[634]);
	Full_Adder FA608 (Cout[473], Cout[474], S[475], S[635], Cout[635]);
	Full_Adder FA609 (S[476], S[477], S[478], S[636], Cout[636]);
	Full_Adder FA610 (S[305], Cout[475], Cout[476], S[637], Cout[637]);
	Full_Adder FA611 (Cout[477], Cout[478], S[479], S[638], Cout[638]);
	Full_Adder FA612 (S[480], S[481], S[482], S[639], Cout[639]);
	Full_Adder FA613 (S[311], Cout[479], Cout[480], S[640], Cout[640]);
	Full_Adder FA614 (Cout[481], Cout[482], S[483], S[641], Cout[641]);
	Full_Adder FA615 (S[484], S[485], S[486], S[642], Cout[642]);
	Full_Adder FA616 (S[317], Cout[483], Cout[484], S[643], Cout[643]);
	Full_Adder FA617 (Cout[485], Cout[486], S[487], S[644], Cout[644]);
	Full_Adder FA618 (S[488], S[489], S[490], S[645], Cout[645]);
	Full_Adder FA619 (S[323], Cout[487], Cout[488], S[646], Cout[646]);
	Full_Adder FA620 (Cout[489], Cout[490], S[491], S[647], Cout[647]);
	Full_Adder FA621 (S[492], S[493], S[494], S[648], Cout[648]);
	Full_Adder FA622 (S[329], Cout[491], Cout[492], S[649], Cout[649]);
	Full_Adder FA623 (Cout[493], Cout[494], S[495], S[650], Cout[650]);
	Full_Adder FA624 (S[496], S[497], S[498], S[651], Cout[651]);
	Full_Adder FA625 (S[335], Cout[495], Cout[496], S[652], Cout[652]);
	Full_Adder FA626 (Cout[497], Cout[498], S[499], S[653], Cout[653]);
	Full_Adder FA627 (S[500], S[501], S[502], S[654], Cout[654]);
	Full_Adder FA628 (S[341], Cout[499], Cout[500], S[655], Cout[655]);
	Full_Adder FA629 (Cout[501], Cout[502], S[503], S[656], Cout[656]);
	Full_Adder FA630 (S[504], S[505], S[506], S[657], Cout[657]);
	Full_Adder FA631 (S[347], Cout[503], Cout[504], S[658], Cout[658]);
	Full_Adder FA632 (Cout[505], Cout[506], S[507], S[659], Cout[659]);
	Full_Adder FA633 (S[508], S[509], S[510], S[660], Cout[660]);
	Full_Adder FA634 (S[353], Cout[507], Cout[508], S[661], Cout[661]);
	Full_Adder FA635 (Cout[509], Cout[510], S[511], S[662], Cout[662]);
	Full_Adder FA636 (S[512], S[513], S[514], S[663], Cout[663]);
	Full_Adder FA637 (S[359], Cout[511], Cout[512], S[664], Cout[664]);
	Full_Adder FA638 (Cout[513], Cout[514], S[515], S[665], Cout[665]);
	Full_Adder FA639 (S[516], S[517], S[518], S[666], Cout[666]);
	Full_Adder FA640 (S[365], Cout[515], Cout[516], S[667], Cout[667]);
	Full_Adder FA641 (Cout[517], Cout[518], S[519], S[668], Cout[668]);
	Full_Adder FA642 (S[520], S[521], S[522], S[669], Cout[669]);
	Full_Adder FA643 (S[370], Cout[519], Cout[520], S[670], Cout[670]);
	Full_Adder FA644 (Cout[521], Cout[522], S[523], S[671], Cout[671]);
	Full_Adder FA645 (S[524], S[525], S[526], S[672], Cout[672]);
	Full_Adder FA646 (S[374], Cout[523], Cout[524], S[673], Cout[673]);
	Full_Adder FA647 (Cout[525], Cout[526], S[527], S[674], Cout[674]);
	Full_Adder FA648 (S[528], S[529], S[530], S[675], Cout[675]);
	Full_Adder FA649 (S[377], Cout[527], Cout[528], S[676], Cout[676]);
	Full_Adder FA650 (Cout[529], Cout[530], S[531], S[677], Cout[677]);
	Full_Adder FA651 (S[532], S[533], S[534], S[678], Cout[678]);
	Full_Adder FA652 (S[379], Cout[531], Cout[532], S[679], Cout[679]);
	Full_Adder FA653 (Cout[533], Cout[534], S[535], S[680], Cout[680]);
	Full_Adder FA654 (S[536], S[537], S[538], S[681], Cout[681]);
	Full_Adder FA655 (S[380], Cout[535], Cout[536], S[682], Cout[682]);
	Full_Adder FA656 (Cout[537], Cout[538], S[539], S[683], Cout[683]);
	Full_Adder FA657 (S[540], S[541], S[542], S[684], Cout[684]);
	Full_Adder FA658 (Cout[380], Cout[539], Cout[540], S[685], Cout[685]);
	Full_Adder FA659 (Cout[541], Cout[542], S[543], S[686], Cout[686]);
	Full_Adder FA660 (S[544], S[545], S[546], S[687], Cout[687]);
	Full_Adder FA661 (pp30[22], pp31[21], Cout[543], S[688], Cout[688]);
	Full_Adder FA662 (Cout[544], Cout[545], Cout[546], S[689], Cout[689]);
	Full_Adder FA663 (S[547], S[548], S[549], S[690], Cout[690]);
	Full_Adder FA664 (pp28[25], pp29[24], pp30[23], S[691], Cout[691]);
	Full_Adder FA665 (pp31[22], Cout[547], Cout[548], S[692], Cout[692]);
	Full_Adder FA666 (Cout[549], S[550], S[551], S[693], Cout[693]);
	Full_Adder FA667 (pp26[28], pp27[27], pp28[26], S[694], Cout[694]);
	Full_Adder FA668 (pp29[25], pp30[24], pp31[23], S[695], Cout[695]);
	Full_Adder FA669 (Cout[550], Cout[551], S[552], S[696], Cout[696]);
	Full_Adder FA670 (pp24[31], pp25[30], pp26[29], S[697], Cout[697]);
	Full_Adder FA671 (pp27[28], pp28[27], pp29[26], S[698], Cout[698]);
	Full_Adder FA672 (pp30[25], pp31[24], Cout[552], S[699], Cout[699]);
	Full_Adder FA673 (pp25[31], pp26[30], pp27[29], S[700], Cout[700]);
	Full_Adder FA674 (pp28[28], pp29[27], pp30[26], S[701], Cout[701]);
	Full_Adder FA675 (pp26[31], pp27[30], pp28[29], S[702], Cout[702]);
	Half_Adder HA28 (pp0[4], pp1[3], S[703], Cout[703]);
	Full_Adder FA676 (pp0[5], pp1[4], pp2[3], S[704], Cout[704]);
	Half_Adder HA29 (pp3[2], pp4[1], S[705], Cout[705]);
	Full_Adder FA677 (pp2[4], pp3[3], pp4[2], S[706], Cout[706]);
	Full_Adder FA678 (pp5[1], pp6[0], S[553], S[707], Cout[707]);
	Full_Adder FA679 (pp5[2], pp6[1], pp7[0], S[708], Cout[708]);
	Full_Adder FA680 (Cout[553], S[554], S[555], S[709], Cout[709]);
	Full_Adder FA681 (pp8[0], Cout[554], Cout[555], S[710], Cout[710]);
	Full_Adder FA682 (S[556], S[557], S[558], S[711], Cout[711]);
	Full_Adder FA683 (Cout[556], Cout[557], Cout[558], S[712], Cout[712]);
	Full_Adder FA684 (S[559], S[560], S[561], S[713], Cout[713]);
	Full_Adder FA685 (Cout[559], Cout[560], Cout[561], S[714], Cout[714]);
	Full_Adder FA686 (S[562], S[563], S[564], S[715], Cout[715]);
	Full_Adder FA687 (Cout[562], Cout[563], Cout[564], S[716], Cout[716]);
	Full_Adder FA688 (S[565], S[566], S[567], S[717], Cout[717]);
	Full_Adder FA689 (Cout[565], Cout[566], Cout[567], S[718], Cout[718]);
	Full_Adder FA690 (S[568], S[569], S[570], S[719], Cout[719]);
	Full_Adder FA691 (Cout[568], Cout[569], Cout[570], S[720], Cout[720]);
	Full_Adder FA692 (S[571], S[572], S[573], S[721], Cout[721]);
	Full_Adder FA693 (Cout[571], Cout[572], Cout[573], S[722], Cout[722]);
	Full_Adder FA694 (S[574], S[575], S[576], S[723], Cout[723]);
	Full_Adder FA695 (Cout[574], Cout[575], Cout[576], S[724], Cout[724]);
	Full_Adder FA696 (S[577], S[578], S[579], S[725], Cout[725]);
	Full_Adder FA697 (Cout[577], Cout[578], Cout[579], S[726], Cout[726]);
	Full_Adder FA698 (S[580], S[581], S[582], S[727], Cout[727]);
	Full_Adder FA699 (Cout[580], Cout[581], Cout[582], S[728], Cout[728]);
	Full_Adder FA700 (S[583], S[584], S[585], S[729], Cout[729]);
	Full_Adder FA701 (Cout[583], Cout[584], Cout[585], S[730], Cout[730]);
	Full_Adder FA702 (S[586], S[587], S[588], S[731], Cout[731]);
	Full_Adder FA703 (Cout[586], Cout[587], Cout[588], S[732], Cout[732]);
	Full_Adder FA704 (S[589], S[590], S[591], S[733], Cout[733]);
	Full_Adder FA705 (Cout[589], Cout[590], Cout[591], S[734], Cout[734]);
	Full_Adder FA706 (S[592], S[593], S[594], S[735], Cout[735]);
	Full_Adder FA707 (Cout[592], Cout[593], Cout[594], S[736], Cout[736]);
	Full_Adder FA708 (S[595], S[596], S[597], S[737], Cout[737]);
	Full_Adder FA709 (Cout[595], Cout[596], Cout[597], S[738], Cout[738]);
	Full_Adder FA710 (S[598], S[599], S[600], S[739], Cout[739]);
	Full_Adder FA711 (Cout[598], Cout[599], Cout[600], S[740], Cout[740]);
	Full_Adder FA712 (S[601], S[602], S[603], S[741], Cout[741]);
	Full_Adder FA713 (Cout[601], Cout[602], Cout[603], S[742], Cout[742]);
	Full_Adder FA714 (S[604], S[605], S[606], S[743], Cout[743]);
	Full_Adder FA715 (Cout[604], Cout[605], Cout[606], S[744], Cout[744]);
	Full_Adder FA716 (S[607], S[608], S[609], S[745], Cout[745]);
	Full_Adder FA717 (Cout[607], Cout[608], Cout[609], S[746], Cout[746]);
	Full_Adder FA718 (S[610], S[611], S[612], S[747], Cout[747]);
	Full_Adder FA719 (Cout[610], Cout[611], Cout[612], S[748], Cout[748]);
	Full_Adder FA720 (S[613], S[614], S[615], S[749], Cout[749]);
	Full_Adder FA721 (Cout[613], Cout[614], Cout[615], S[750], Cout[750]);
	Full_Adder FA722 (S[616], S[617], S[618], S[751], Cout[751]);
	Full_Adder FA723 (Cout[616], Cout[617], Cout[618], S[752], Cout[752]);
	Full_Adder FA724 (S[619], S[620], S[621], S[753], Cout[753]);
	Full_Adder FA725 (Cout[619], Cout[620], Cout[621], S[754], Cout[754]);
	Full_Adder FA726 (S[622], S[623], S[624], S[755], Cout[755]);
	Full_Adder FA727 (Cout[622], Cout[623], Cout[624], S[756], Cout[756]);
	Full_Adder FA728 (S[625], S[626], S[627], S[757], Cout[757]);
	Full_Adder FA729 (Cout[625], Cout[626], Cout[627], S[758], Cout[758]);
	Full_Adder FA730 (S[628], S[629], S[630], S[759], Cout[759]);
	Full_Adder FA731 (Cout[628], Cout[629], Cout[630], S[760], Cout[760]);
	Full_Adder FA732 (S[631], S[632], S[633], S[761], Cout[761]);
	Full_Adder FA733 (Cout[631], Cout[632], Cout[633], S[762], Cout[762]);
	Full_Adder FA734 (S[634], S[635], S[636], S[763], Cout[763]);
	Full_Adder FA735 (Cout[634], Cout[635], Cout[636], S[764], Cout[764]);
	Full_Adder FA736 (S[637], S[638], S[639], S[765], Cout[765]);
	Full_Adder FA737 (Cout[637], Cout[638], Cout[639], S[766], Cout[766]);
	Full_Adder FA738 (S[640], S[641], S[642], S[767], Cout[767]);
	Full_Adder FA739 (Cout[640], Cout[641], Cout[642], S[768], Cout[768]);
	Full_Adder FA740 (S[643], S[644], S[645], S[769], Cout[769]);
	Full_Adder FA741 (Cout[643], Cout[644], Cout[645], S[770], Cout[770]);
	Full_Adder FA742 (S[646], S[647], S[648], S[771], Cout[771]);
	Full_Adder FA743 (Cout[646], Cout[647], Cout[648], S[772], Cout[772]);
	Full_Adder FA744 (S[649], S[650], S[651], S[773], Cout[773]);
	Full_Adder FA745 (Cout[649], Cout[650], Cout[651], S[774], Cout[774]);
	Full_Adder FA746 (S[652], S[653], S[654], S[775], Cout[775]);
	Full_Adder FA747 (Cout[652], Cout[653], Cout[654], S[776], Cout[776]);
	Full_Adder FA748 (S[655], S[656], S[657], S[777], Cout[777]);
	Full_Adder FA749 (Cout[655], Cout[656], Cout[657], S[778], Cout[778]);
	Full_Adder FA750 (S[658], S[659], S[660], S[779], Cout[779]);
	Full_Adder FA751 (Cout[658], Cout[659], Cout[660], S[780], Cout[780]);
	Full_Adder FA752 (S[661], S[662], S[663], S[781], Cout[781]);
	Full_Adder FA753 (Cout[661], Cout[662], Cout[663], S[782], Cout[782]);
	Full_Adder FA754 (S[664], S[665], S[666], S[783], Cout[783]);
	Full_Adder FA755 (Cout[664], Cout[665], Cout[666], S[784], Cout[784]);
	Full_Adder FA756 (S[667], S[668], S[669], S[785], Cout[785]);
	Full_Adder FA757 (Cout[667], Cout[668], Cout[669], S[786], Cout[786]);
	Full_Adder FA758 (S[670], S[671], S[672], S[787], Cout[787]);
	Full_Adder FA759 (Cout[670], Cout[671], Cout[672], S[788], Cout[788]);
	Full_Adder FA760 (S[673], S[674], S[675], S[789], Cout[789]);
	Full_Adder FA761 (Cout[673], Cout[674], Cout[675], S[790], Cout[790]);
	Full_Adder FA762 (S[676], S[677], S[678], S[791], Cout[791]);
	Full_Adder FA763 (Cout[676], Cout[677], Cout[678], S[792], Cout[792]);
	Full_Adder FA764 (S[679], S[680], S[681], S[793], Cout[793]);
	Full_Adder FA765 (Cout[679], Cout[680], Cout[681], S[794], Cout[794]);
	Full_Adder FA766 (S[682], S[683], S[684], S[795], Cout[795]);
	Full_Adder FA767 (Cout[682], Cout[683], Cout[684], S[796], Cout[796]);
	Full_Adder FA768 (S[685], S[686], S[687], S[797], Cout[797]);
	Full_Adder FA769 (Cout[685], Cout[686], Cout[687], S[798], Cout[798]);
	Full_Adder FA770 (S[688], S[689], S[690], S[799], Cout[799]);
	Full_Adder FA771 (Cout[688], Cout[689], Cout[690], S[800], Cout[800]);
	Full_Adder FA772 (S[691], S[692], S[693], S[801], Cout[801]);
	Full_Adder FA773 (Cout[691], Cout[692], Cout[693], S[802], Cout[802]);
	Full_Adder FA774 (S[694], S[695], S[696], S[803], Cout[803]);
	Full_Adder FA775 (Cout[694], Cout[695], Cout[696], S[804], Cout[804]);
	Full_Adder FA776 (S[697], S[698], S[699], S[805], Cout[805]);
	Full_Adder FA777 (pp31[25], Cout[697], Cout[698], S[806], Cout[806]);
	Full_Adder FA778 (Cout[699], S[700], S[701], S[807], Cout[807]);
	Full_Adder FA779 (pp29[28], pp30[27], pp31[26], S[808], Cout[808]);
	Full_Adder FA780 (Cout[700], Cout[701], S[702], S[809], Cout[809]);
	Full_Adder FA781 (pp27[31], pp28[30], pp29[29], S[810], Cout[810]);
	Full_Adder FA782 (pp30[28], pp31[27], Cout[702], S[811], Cout[811]);
	Full_Adder FA783 (pp28[31], pp29[30], pp30[29], S[812], Cout[812]);
	Half_Adder HA30 (pp0[3], pp1[2], S[813], Cout[813]);
	Full_Adder FA784 (pp2[2], pp3[1], pp4[0], S[814], Cout[814]);
	Full_Adder FA785 (pp5[0], Cout[703], S[704], S[815], Cout[815]);
	Full_Adder FA786 (Cout[704], Cout[705], S[706], S[816], Cout[816]);
	Full_Adder FA787 (Cout[706], Cout[707], S[708], S[817], Cout[817]);
	Full_Adder FA788 (Cout[708], Cout[709], S[710], S[818], Cout[818]);
	Full_Adder FA789 (Cout[710], Cout[711], S[712], S[819], Cout[819]);
	Full_Adder FA790 (Cout[712], Cout[713], S[714], S[820], Cout[820]);
	Full_Adder FA791 (Cout[714], Cout[715], S[716], S[821], Cout[821]);
	Full_Adder FA792 (Cout[716], Cout[717], S[718], S[822], Cout[822]);
	Full_Adder FA793 (Cout[718], Cout[719], S[720], S[823], Cout[823]);
	Full_Adder FA794 (Cout[720], Cout[721], S[722], S[824], Cout[824]);
	Full_Adder FA795 (Cout[722], Cout[723], S[724], S[825], Cout[825]);
	Full_Adder FA796 (Cout[724], Cout[725], S[726], S[826], Cout[826]);
	Full_Adder FA797 (Cout[726], Cout[727], S[728], S[827], Cout[827]);
	Full_Adder FA798 (Cout[728], Cout[729], S[730], S[828], Cout[828]);
	Full_Adder FA799 (Cout[730], Cout[731], S[732], S[829], Cout[829]);
	Full_Adder FA800 (Cout[732], Cout[733], S[734], S[830], Cout[830]);
	Full_Adder FA801 (Cout[734], Cout[735], S[736], S[831], Cout[831]);
	Full_Adder FA802 (Cout[736], Cout[737], S[738], S[832], Cout[832]);
	Full_Adder FA803 (Cout[738], Cout[739], S[740], S[833], Cout[833]);
	Full_Adder FA804 (Cout[740], Cout[741], S[742], S[834], Cout[834]);
	Full_Adder FA805 (Cout[742], Cout[743], S[744], S[835], Cout[835]);
	Full_Adder FA806 (Cout[744], Cout[745], S[746], S[836], Cout[836]);
	Full_Adder FA807 (Cout[746], Cout[747], S[748], S[837], Cout[837]);
	Full_Adder FA808 (Cout[748], Cout[749], S[750], S[838], Cout[838]);
	Full_Adder FA809 (Cout[750], Cout[751], S[752], S[839], Cout[839]);
	Full_Adder FA810 (Cout[752], Cout[753], S[754], S[840], Cout[840]);
	Full_Adder FA811 (Cout[754], Cout[755], S[756], S[841], Cout[841]);
	Full_Adder FA812 (Cout[756], Cout[757], S[758], S[842], Cout[842]);
	Full_Adder FA813 (Cout[758], Cout[759], S[760], S[843], Cout[843]);
	Full_Adder FA814 (Cout[760], Cout[761], S[762], S[844], Cout[844]);
	Full_Adder FA815 (Cout[762], Cout[763], S[764], S[845], Cout[845]);
	Full_Adder FA816 (Cout[764], Cout[765], S[766], S[846], Cout[846]);
	Full_Adder FA817 (Cout[766], Cout[767], S[768], S[847], Cout[847]);
	Full_Adder FA818 (Cout[768], Cout[769], S[770], S[848], Cout[848]);
	Full_Adder FA819 (Cout[770], Cout[771], S[772], S[849], Cout[849]);
	Full_Adder FA820 (Cout[772], Cout[773], S[774], S[850], Cout[850]);
	Full_Adder FA821 (Cout[774], Cout[775], S[776], S[851], Cout[851]);
	Full_Adder FA822 (Cout[776], Cout[777], S[778], S[852], Cout[852]);
	Full_Adder FA823 (Cout[778], Cout[779], S[780], S[853], Cout[853]);
	Full_Adder FA824 (Cout[780], Cout[781], S[782], S[854], Cout[854]);
	Full_Adder FA825 (Cout[782], Cout[783], S[784], S[855], Cout[855]);
	Full_Adder FA826 (Cout[784], Cout[785], S[786], S[856], Cout[856]);
	Full_Adder FA827 (Cout[786], Cout[787], S[788], S[857], Cout[857]);
	Full_Adder FA828 (Cout[788], Cout[789], S[790], S[858], Cout[858]);
	Full_Adder FA829 (Cout[790], Cout[791], S[792], S[859], Cout[859]);
	Full_Adder FA830 (Cout[792], Cout[793], S[794], S[860], Cout[860]);
	Full_Adder FA831 (Cout[794], Cout[795], S[796], S[861], Cout[861]);
	Full_Adder FA832 (Cout[796], Cout[797], S[798], S[862], Cout[862]);
	Full_Adder FA833 (Cout[798], Cout[799], S[800], S[863], Cout[863]);
	Full_Adder FA834 (Cout[800], Cout[801], S[802], S[864], Cout[864]);
	Full_Adder FA835 (Cout[802], Cout[803], S[804], S[865], Cout[865]);
	Full_Adder FA836 (Cout[804], Cout[805], S[806], S[866], Cout[866]);
	Full_Adder FA837 (Cout[806], Cout[807], S[808], S[867], Cout[867]);
	Full_Adder FA838 (Cout[808], Cout[809], S[810], S[868], Cout[868]);
	Full_Adder FA839 (pp31[28], Cout[810], Cout[811], S[869], Cout[869]);
	Full_Adder FA840 (pp29[31], pp30[30], pp31[29], S[870], Cout[870]);
	Half_Adder HA31 (pp0[2], pp1[1], S[871], Cout[871]);
	Full_Adder FA841 (pp2[1], pp3[0], S[813], S[872], Cout[872]);
	Full_Adder FA842 (S[703], Cout[813], S[814], S[873], Cout[873]);
	Full_Adder FA843 (S[705], Cout[814], S[815], S[874], Cout[874]);
	Full_Adder FA844 (S[707], Cout[815], S[816], S[875], Cout[875]);
	Full_Adder FA845 (S[709], Cout[816], S[817], S[876], Cout[876]);
	Full_Adder FA846 (S[711], Cout[817], S[818], S[877], Cout[877]);
	Full_Adder FA847 (S[713], Cout[818], S[819], S[878], Cout[878]);
	Full_Adder FA848 (S[715], Cout[819], S[820], S[879], Cout[879]);
	Full_Adder FA849 (S[717], Cout[820], S[821], S[880], Cout[880]);
	Full_Adder FA850 (S[719], Cout[821], S[822], S[881], Cout[881]);
	Full_Adder FA851 (S[721], Cout[822], S[823], S[882], Cout[882]);
	Full_Adder FA852 (S[723], Cout[823], S[824], S[883], Cout[883]);
	Full_Adder FA853 (S[725], Cout[824], S[825], S[884], Cout[884]);
	Full_Adder FA854 (S[727], Cout[825], S[826], S[885], Cout[885]);
	Full_Adder FA855 (S[729], Cout[826], S[827], S[886], Cout[886]);
	Full_Adder FA856 (S[731], Cout[827], S[828], S[887], Cout[887]);
	Full_Adder FA857 (S[733], Cout[828], S[829], S[888], Cout[888]);
	Full_Adder FA858 (S[735], Cout[829], S[830], S[889], Cout[889]);
	Full_Adder FA859 (S[737], Cout[830], S[831], S[890], Cout[890]);
	Full_Adder FA860 (S[739], Cout[831], S[832], S[891], Cout[891]);
	Full_Adder FA861 (S[741], Cout[832], S[833], S[892], Cout[892]);
	Full_Adder FA862 (S[743], Cout[833], S[834], S[893], Cout[893]);
	Full_Adder FA863 (S[745], Cout[834], S[835], S[894], Cout[894]);
	Full_Adder FA864 (S[747], Cout[835], S[836], S[895], Cout[895]);
	Full_Adder FA865 (S[749], Cout[836], S[837], S[896], Cout[896]);
	Full_Adder FA866 (S[751], Cout[837], S[838], S[897], Cout[897]);
	Full_Adder FA867 (S[753], Cout[838], S[839], S[898], Cout[898]);
	Full_Adder FA868 (S[755], Cout[839], S[840], S[899], Cout[899]);
	Full_Adder FA869 (S[757], Cout[840], S[841], S[900], Cout[900]);
	Full_Adder FA870 (S[759], Cout[841], S[842], S[901], Cout[901]);
	Full_Adder FA871 (S[761], Cout[842], S[843], S[902], Cout[902]);
	Full_Adder FA872 (S[763], Cout[843], S[844], S[903], Cout[903]);
	Full_Adder FA873 (S[765], Cout[844], S[845], S[904], Cout[904]);
	Full_Adder FA874 (S[767], Cout[845], S[846], S[905], Cout[905]);
	Full_Adder FA875 (S[769], Cout[846], S[847], S[906], Cout[906]);
	Full_Adder FA876 (S[771], Cout[847], S[848], S[907], Cout[907]);
	Full_Adder FA877 (S[773], Cout[848], S[849], S[908], Cout[908]);
	Full_Adder FA878 (S[775], Cout[849], S[850], S[909], Cout[909]);
	Full_Adder FA879 (S[777], Cout[850], S[851], S[910], Cout[910]);
	Full_Adder FA880 (S[779], Cout[851], S[852], S[911], Cout[911]);
	Full_Adder FA881 (S[781], Cout[852], S[853], S[912], Cout[912]);
	Full_Adder FA882 (S[783], Cout[853], S[854], S[913], Cout[913]);
	Full_Adder FA883 (S[785], Cout[854], S[855], S[914], Cout[914]);
	Full_Adder FA884 (S[787], Cout[855], S[856], S[915], Cout[915]);
	Full_Adder FA885 (S[789], Cout[856], S[857], S[916], Cout[916]);
	Full_Adder FA886 (S[791], Cout[857], S[858], S[917], Cout[917]);
	Full_Adder FA887 (S[793], Cout[858], S[859], S[918], Cout[918]);
	Full_Adder FA888 (S[795], Cout[859], S[860], S[919], Cout[919]);
	Full_Adder FA889 (S[797], Cout[860], S[861], S[920], Cout[920]);
	Full_Adder FA890 (S[799], Cout[861], S[862], S[921], Cout[921]);
	Full_Adder FA891 (S[801], Cout[862], S[863], S[922], Cout[922]);
	Full_Adder FA892 (S[803], Cout[863], S[864], S[923], Cout[923]);
	Full_Adder FA893 (S[805], Cout[864], S[865], S[924], Cout[924]);
	Full_Adder FA894 (S[807], Cout[865], S[866], S[925], Cout[925]);
	Full_Adder FA895 (S[809], Cout[866], S[867], S[926], Cout[926]);
	Full_Adder FA896 (S[811], Cout[867], S[868], S[927], Cout[927]);
	Full_Adder FA897 (S[812], Cout[868], S[869], S[928], Cout[928]);
	Full_Adder FA898 (Cout[812], Cout[869], S[870], S[929], Cout[929]);
	Full_Adder FA899 (pp30[31], pp31[30], Cout[870], S[930], Cout[930]);
	Half_Adder HA32 (pp0[1], pp1[0], S[0], Cout[0]);
	Full_Adder FA900 (pp2[0], S[871], Cout[0], S[931], Cout[931]);
	Full_Adder FA901 (Cout[871], S[872], Cout[931], S[932], Cout[932]);
	Full_Adder FA902 (Cout[872], S[873], Cout[932], S[933], Cout[933]);
	Full_Adder FA903 (Cout[873], S[874], Cout[933], S[934], Cout[934]);
	Full_Adder FA904 (Cout[874], S[875], Cout[934], S[935], Cout[935]);
	Full_Adder FA905 (Cout[875], S[876], Cout[935], S[936], Cout[936]);
	Full_Adder FA906 (Cout[876], S[877], Cout[936], S[937], Cout[937]);
	Full_Adder FA907 (Cout[877], S[878], Cout[937], S[938], Cout[938]);
	Full_Adder FA908 (Cout[878], S[879], Cout[938], S[939], Cout[939]);
	Full_Adder FA909 (Cout[879], S[880], Cout[939], S[940], Cout[940]);
	Full_Adder FA910 (Cout[880], S[881], Cout[940], S[941], Cout[941]);
	Full_Adder FA911 (Cout[881], S[882], Cout[941], S[942], Cout[942]);
	Full_Adder FA912 (Cout[882], S[883], Cout[942], S[943], Cout[943]);
	Full_Adder FA913 (Cout[883], S[884], Cout[943], S[944], Cout[944]);
	Full_Adder FA914 (Cout[884], S[885], Cout[944], S[945], Cout[945]);
	Full_Adder FA915 (Cout[885], S[886], Cout[945], S[946], Cout[946]);
	Full_Adder FA916 (Cout[886], S[887], Cout[946], S[947], Cout[947]);
	Full_Adder FA917 (Cout[887], S[888], Cout[947], S[948], Cout[948]);
	Full_Adder FA918 (Cout[888], S[889], Cout[948], S[949], Cout[949]);
	Full_Adder FA919 (Cout[889], S[890], Cout[949], S[950], Cout[950]);
	Full_Adder FA920 (Cout[890], S[891], Cout[950], S[951], Cout[951]);
	Full_Adder FA921 (Cout[891], S[892], Cout[951], S[952], Cout[952]);
	Full_Adder FA922 (Cout[892], S[893], Cout[952], S[953], Cout[953]);
	Full_Adder FA923 (Cout[893], S[894], Cout[953], S[954], Cout[954]);
	Full_Adder FA924 (Cout[894], S[895], Cout[954], S[955], Cout[955]);
	Full_Adder FA925 (Cout[895], S[896], Cout[955], S[956], Cout[956]);
	Full_Adder FA926 (Cout[896], S[897], Cout[956], S[957], Cout[957]);
	Full_Adder FA927 (Cout[897], S[898], Cout[957], S[958], Cout[958]);
	Full_Adder FA928 (Cout[898], S[899], Cout[958], S[959], Cout[959]);
	Full_Adder FA929 (Cout[899], S[900], Cout[959], S[960], Cout[960]);
	Full_Adder FA930 (Cout[900], S[901], Cout[960], S[961], Cout[961]);
	Full_Adder FA931 (Cout[901], S[902], Cout[961], S[962], Cout[962]);
	Full_Adder FA932 (Cout[902], S[903], Cout[962], S[963], Cout[963]);
	Full_Adder FA933 (Cout[903], S[904], Cout[963], S[964], Cout[964]);
	Full_Adder FA934 (Cout[904], S[905], Cout[964], S[965], Cout[965]);
	Full_Adder FA935 (Cout[905], S[906], Cout[965], S[966], Cout[966]);
	Full_Adder FA936 (Cout[906], S[907], Cout[966], S[967], Cout[967]);
	Full_Adder FA937 (Cout[907], S[908], Cout[967], S[968], Cout[968]);
	Full_Adder FA938 (Cout[908], S[909], Cout[968], S[969], Cout[969]);
	Full_Adder FA939 (Cout[909], S[910], Cout[969], S[970], Cout[970]);
	Full_Adder FA940 (Cout[910], S[911], Cout[970], S[971], Cout[971]);
	Full_Adder FA941 (Cout[911], S[912], Cout[971], S[972], Cout[972]);
	Full_Adder FA942 (Cout[912], S[913], Cout[972], S[973], Cout[973]);
	Full_Adder FA943 (Cout[913], S[914], Cout[973], S[974], Cout[974]);
	Full_Adder FA944 (Cout[914], S[915], Cout[974], S[975], Cout[975]);
	Full_Adder FA945 (Cout[915], S[916], Cout[975], S[976], Cout[976]);
	Full_Adder FA946 (Cout[916], S[917], Cout[976], S[977], Cout[977]);
	Full_Adder FA947 (Cout[917], S[918], Cout[977], S[978], Cout[978]);
	Full_Adder FA948 (Cout[918], S[919], Cout[978], S[979], Cout[979]);
	Full_Adder FA949 (Cout[919], S[920], Cout[979], S[980], Cout[980]);
	Full_Adder FA950 (Cout[920], S[921], Cout[980], S[981], Cout[981]);
	Full_Adder FA951 (Cout[921], S[922], Cout[981], S[982], Cout[982]);
	Full_Adder FA952 (Cout[922], S[923], Cout[982], S[983], Cout[983]);
	Full_Adder FA953 (Cout[923], S[924], Cout[983], S[984], Cout[984]);
	Full_Adder FA954 (Cout[924], S[925], Cout[984], S[985], Cout[985]);
	Full_Adder FA955 (Cout[925], S[926], Cout[985], S[986], Cout[986]);
	Full_Adder FA956 (Cout[926], S[927], Cout[986], S[987], Cout[987]);
	Full_Adder FA957 (Cout[927], S[928], Cout[987], S[988], Cout[988]);
	Full_Adder FA958 (Cout[928], S[929], Cout[988], S[989], Cout[989]);
	Full_Adder FA959 (Cout[929], S[930], Cout[989], S[990], Cout[990]);
	Full_Adder FA960 (pp31[31], Cout[930], Cout[990], S[991], Cout[991]);

	assign product[63] = Cout[991];
	assign product[62] = S[991];
	assign product[61] = S[990];
	assign product[60] = S[989];
	assign product[59] = S[988];
	assign product[58] = S[987];
	assign product[57] = S[986];
	assign product[56] = S[985];
	assign product[55] = S[984];
	assign product[54] = S[983];
	assign product[53] = S[982];
	assign product[52] = S[981];
	assign product[51] = S[980];
	assign product[50] = S[979];
	assign product[49] = S[978];
	assign product[48] = S[977];
	assign product[47] = S[976];
	assign product[46] = S[975];
	assign product[45] = S[974];
	assign product[44] = S[973];
	assign product[43] = S[972];
	assign product[42] = S[971];
	assign product[41] = S[970];
	assign product[40] = S[969];
	assign product[39] = S[968];
	assign product[38] = S[967];
	assign product[37] = S[966];
	assign product[36] = S[965];
	assign product[35] = S[964];
	assign product[34] = S[963];
	assign product[33] = S[962];
	assign product[32] = S[961];
	assign product[31] = S[960];
	assign product[30] = S[959];
	assign product[29] = S[958];
	assign product[28] = S[957];
	assign product[27] = S[956];
	assign product[26] = S[955];
	assign product[25] = S[954];
	assign product[24] = S[953];
	assign product[23] = S[952];
	assign product[22] = S[951];
	assign product[21] = S[950];
	assign product[20] = S[949];
	assign product[19] = S[948];
	assign product[18] = S[947];
	assign product[17] = S[946];
	assign product[16] = S[945];
	assign product[15] = S[944];
	assign product[14] = S[943];
	assign product[13] = S[942];
	assign product[12] = S[941];
	assign product[11] = S[940];
	assign product[10] = S[939];
	assign product[9] = S[938];
	assign product[8] = S[937];
	assign product[7] = S[936];
	assign product[6] = S[935];
	assign product[5] = S[934];
	assign product[4] = S[933];
	assign product[3] = S[932];
	assign product[2] = S[931];
	assign product[1] = S[0];
	assign product[0] = pp0[0];
endmodule

module Half_Adder(input wire in1,
                  input wire in2,
				  output wire sum,
                  output wire cout);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(input wire in1,
                  input wire in2,
                  input wire cin,
				  output wire sum,
                  output wire cout);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule
