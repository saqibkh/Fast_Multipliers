module wallace_unsigned_multiplier_RCA_16(product, A, B);
    input [15:0] A, B;
    output [31:0] product;

wire [15:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;

assign P[0][0] = x[0] & y[0];
assign P[0][1] = x[0] & y[1];
assign P[0][2] = x[0] & y[2];
assign P[0][3] = x[0] & y[3];
assign P[0][4] = x[0] & y[4];
assign P[0][5] = x[0] & y[5];
assign P[0][6] = x[0] & y[6];
assign P[0][7] = x[0] & y[7];
assign P[0][8] = x[0] & y[8];
assign P[0][9] = x[0] & y[9];
assign P[0][10] = x[0] & y[10];
assign P[0][11] = x[0] & y[11];
assign P[0][12] = x[0] & y[12];
assign P[0][13] = x[0] & y[13];
assign P[0][14] = x[0] & y[14];
assign P[0][15] = x[0] & y[15];
assign P[1][0] = x[1] & y[0];
assign P[1][1] = x[1] & y[1];
assign P[1][2] = x[1] & y[2];
assign P[1][3] = x[1] & y[3];
assign P[1][4] = x[1] & y[4];
assign P[1][5] = x[1] & y[5];
assign P[1][6] = x[1] & y[6];
assign P[1][7] = x[1] & y[7];
assign P[1][8] = x[1] & y[8];
assign P[1][9] = x[1] & y[9];
assign P[1][10] = x[1] & y[10];
assign P[1][11] = x[1] & y[11];
assign P[1][12] = x[1] & y[12];
assign P[1][13] = x[1] & y[13];
assign P[1][14] = x[1] & y[14];
assign P[1][15] = x[1] & y[15];
assign P[2][0] = x[2] & y[0];
assign P[2][1] = x[2] & y[1];
assign P[2][2] = x[2] & y[2];
assign P[2][3] = x[2] & y[3];
assign P[2][4] = x[2] & y[4];
assign P[2][5] = x[2] & y[5];
assign P[2][6] = x[2] & y[6];
assign P[2][7] = x[2] & y[7];
assign P[2][8] = x[2] & y[8];
assign P[2][9] = x[2] & y[9];
assign P[2][10] = x[2] & y[10];
assign P[2][11] = x[2] & y[11];
assign P[2][12] = x[2] & y[12];
assign P[2][13] = x[2] & y[13];
assign P[2][14] = x[2] & y[14];
assign P[2][15] = x[2] & y[15];
assign P[3][0] = x[3] & y[0];
assign P[3][1] = x[3] & y[1];
assign P[3][2] = x[3] & y[2];
assign P[3][3] = x[3] & y[3];
assign P[3][4] = x[3] & y[4];
assign P[3][5] = x[3] & y[5];
assign P[3][6] = x[3] & y[6];
assign P[3][7] = x[3] & y[7];
assign P[3][8] = x[3] & y[8];
assign P[3][9] = x[3] & y[9];
assign P[3][10] = x[3] & y[10];
assign P[3][11] = x[3] & y[11];
assign P[3][12] = x[3] & y[12];
assign P[3][13] = x[3] & y[13];
assign P[3][14] = x[3] & y[14];
assign P[3][15] = x[3] & y[15];
assign P[4][0] = x[4] & y[0];
assign P[4][1] = x[4] & y[1];
assign P[4][2] = x[4] & y[2];
assign P[4][3] = x[4] & y[3];
assign P[4][4] = x[4] & y[4];
assign P[4][5] = x[4] & y[5];
assign P[4][6] = x[4] & y[6];
assign P[4][7] = x[4] & y[7];
assign P[4][8] = x[4] & y[8];
assign P[4][9] = x[4] & y[9];
assign P[4][10] = x[4] & y[10];
assign P[4][11] = x[4] & y[11];
assign P[4][12] = x[4] & y[12];
assign P[4][13] = x[4] & y[13];
assign P[4][14] = x[4] & y[14];
assign P[4][15] = x[4] & y[15];
assign P[5][0] = x[5] & y[0];
assign P[5][1] = x[5] & y[1];
assign P[5][2] = x[5] & y[2];
assign P[5][3] = x[5] & y[3];
assign P[5][4] = x[5] & y[4];
assign P[5][5] = x[5] & y[5];
assign P[5][6] = x[5] & y[6];
assign P[5][7] = x[5] & y[7];
assign P[5][8] = x[5] & y[8];
assign P[5][9] = x[5] & y[9];
assign P[5][10] = x[5] & y[10];
assign P[5][11] = x[5] & y[11];
assign P[5][12] = x[5] & y[12];
assign P[5][13] = x[5] & y[13];
assign P[5][14] = x[5] & y[14];
assign P[5][15] = x[5] & y[15];
assign P[6][0] = x[6] & y[0];
assign P[6][1] = x[6] & y[1];
assign P[6][2] = x[6] & y[2];
assign P[6][3] = x[6] & y[3];
assign P[6][4] = x[6] & y[4];
assign P[6][5] = x[6] & y[5];
assign P[6][6] = x[6] & y[6];
assign P[6][7] = x[6] & y[7];
assign P[6][8] = x[6] & y[8];
assign P[6][9] = x[6] & y[9];
assign P[6][10] = x[6] & y[10];
assign P[6][11] = x[6] & y[11];
assign P[6][12] = x[6] & y[12];
assign P[6][13] = x[6] & y[13];
assign P[6][14] = x[6] & y[14];
assign P[6][15] = x[6] & y[15];
assign P[7][0] = x[7] & y[0];
assign P[7][1] = x[7] & y[1];
assign P[7][2] = x[7] & y[2];
assign P[7][3] = x[7] & y[3];
assign P[7][4] = x[7] & y[4];
assign P[7][5] = x[7] & y[5];
assign P[7][6] = x[7] & y[6];
assign P[7][7] = x[7] & y[7];
assign P[7][8] = x[7] & y[8];
assign P[7][9] = x[7] & y[9];
assign P[7][10] = x[7] & y[10];
assign P[7][11] = x[7] & y[11];
assign P[7][12] = x[7] & y[12];
assign P[7][13] = x[7] & y[13];
assign P[7][14] = x[7] & y[14];
assign P[7][15] = x[7] & y[15];
assign P[8][0] = x[8] & y[0];
assign P[8][1] = x[8] & y[1];
assign P[8][2] = x[8] & y[2];
assign P[8][3] = x[8] & y[3];
assign P[8][4] = x[8] & y[4];
assign P[8][5] = x[8] & y[5];
assign P[8][6] = x[8] & y[6];
assign P[8][7] = x[8] & y[7];
assign P[8][8] = x[8] & y[8];
assign P[8][9] = x[8] & y[9];
assign P[8][10] = x[8] & y[10];
assign P[8][11] = x[8] & y[11];
assign P[8][12] = x[8] & y[12];
assign P[8][13] = x[8] & y[13];
assign P[8][14] = x[8] & y[14];
assign P[8][15] = x[8] & y[15];
assign P[9][0] = x[9] & y[0];
assign P[9][1] = x[9] & y[1];
assign P[9][2] = x[9] & y[2];
assign P[9][3] = x[9] & y[3];
assign P[9][4] = x[9] & y[4];
assign P[9][5] = x[9] & y[5];
assign P[9][6] = x[9] & y[6];
assign P[9][7] = x[9] & y[7];
assign P[9][8] = x[9] & y[8];
assign P[9][9] = x[9] & y[9];
assign P[9][10] = x[9] & y[10];
assign P[9][11] = x[9] & y[11];
assign P[9][12] = x[9] & y[12];
assign P[9][13] = x[9] & y[13];
assign P[9][14] = x[9] & y[14];
assign P[9][15] = x[9] & y[15];
assign P[10][0] = x[10] & y[0];
assign P[10][1] = x[10] & y[1];
assign P[10][2] = x[10] & y[2];
assign P[10][3] = x[10] & y[3];
assign P[10][4] = x[10] & y[4];
assign P[10][5] = x[10] & y[5];
assign P[10][6] = x[10] & y[6];
assign P[10][7] = x[10] & y[7];
assign P[10][8] = x[10] & y[8];
assign P[10][9] = x[10] & y[9];
assign P[10][10] = x[10] & y[10];
assign P[10][11] = x[10] & y[11];
assign P[10][12] = x[10] & y[12];
assign P[10][13] = x[10] & y[13];
assign P[10][14] = x[10] & y[14];
assign P[10][15] = x[10] & y[15];
assign P[11][0] = x[11] & y[0];
assign P[11][1] = x[11] & y[1];
assign P[11][2] = x[11] & y[2];
assign P[11][3] = x[11] & y[3];
assign P[11][4] = x[11] & y[4];
assign P[11][5] = x[11] & y[5];
assign P[11][6] = x[11] & y[6];
assign P[11][7] = x[11] & y[7];
assign P[11][8] = x[11] & y[8];
assign P[11][9] = x[11] & y[9];
assign P[11][10] = x[11] & y[10];
assign P[11][11] = x[11] & y[11];
assign P[11][12] = x[11] & y[12];
assign P[11][13] = x[11] & y[13];
assign P[11][14] = x[11] & y[14];
assign P[11][15] = x[11] & y[15];
assign P[12][0] = x[12] & y[0];
assign P[12][1] = x[12] & y[1];
assign P[12][2] = x[12] & y[2];
assign P[12][3] = x[12] & y[3];
assign P[12][4] = x[12] & y[4];
assign P[12][5] = x[12] & y[5];
assign P[12][6] = x[12] & y[6];
assign P[12][7] = x[12] & y[7];
assign P[12][8] = x[12] & y[8];
assign P[12][9] = x[12] & y[9];
assign P[12][10] = x[12] & y[10];
assign P[12][11] = x[12] & y[11];
assign P[12][12] = x[12] & y[12];
assign P[12][13] = x[12] & y[13];
assign P[12][14] = x[12] & y[14];
assign P[12][15] = x[12] & y[15];
assign P[13][0] = x[13] & y[0];
assign P[13][1] = x[13] & y[1];
assign P[13][2] = x[13] & y[2];
assign P[13][3] = x[13] & y[3];
assign P[13][4] = x[13] & y[4];
assign P[13][5] = x[13] & y[5];
assign P[13][6] = x[13] & y[6];
assign P[13][7] = x[13] & y[7];
assign P[13][8] = x[13] & y[8];
assign P[13][9] = x[13] & y[9];
assign P[13][10] = x[13] & y[10];
assign P[13][11] = x[13] & y[11];
assign P[13][12] = x[13] & y[12];
assign P[13][13] = x[13] & y[13];
assign P[13][14] = x[13] & y[14];
assign P[13][15] = x[13] & y[15];
assign P[14][0] = x[14] & y[0];
assign P[14][1] = x[14] & y[1];
assign P[14][2] = x[14] & y[2];
assign P[14][3] = x[14] & y[3];
assign P[14][4] = x[14] & y[4];
assign P[14][5] = x[14] & y[5];
assign P[14][6] = x[14] & y[6];
assign P[14][7] = x[14] & y[7];
assign P[14][8] = x[14] & y[8];
assign P[14][9] = x[14] & y[9];
assign P[14][10] = x[14] & y[10];
assign P[14][11] = x[14] & y[11];
assign P[14][12] = x[14] & y[12];
assign P[14][13] = x[14] & y[13];
assign P[14][14] = x[14] & y[14];
assign P[14][15] = x[14] & y[15];
assign P[15][0] = x[15] & y[0];
assign P[15][1] = x[15] & y[1];
assign P[15][2] = x[15] & y[2];
assign P[15][3] = x[15] & y[3];
assign P[15][4] = x[15] & y[4];
assign P[15][5] = x[15] & y[5];
assign P[15][6] = x[15] & y[6];
assign P[15][7] = x[15] & y[7];
assign P[15][8] = x[15] & y[8];
assign P[15][9] = x[15] & y[9];
assign P[15][10] = x[15] & y[10];
assign P[15][11] = x[15] & y[11];
assign P[15][12] = x[15] & y[12];
assign P[15][13] = x[15] & y[13];
assign P[15][14] = x[15] & y[14];
assign P[15][15] = x[15] & y[15];

wire [276:0] S;
wire [276:0] Cout;

Half_Adder HA1 (P[0][1], P[1][0], S[0], Cout[0]);
Full_Adder FA2 (P[0][2], P[1][1], P[2][0], S[1], Cout[1]);
Full_Adder FA3 (P[0][3], P[1][2], P[2][1], S[2], Cout[2]);
Full_Adder FA4 (P[0][4], P[1][3], P[2][2], S[3], Cout[3]);
Half_Adder HA5 (P[3][1], P[4][0], S[4], Cout[4]);
Full_Adder FA6 (P[0][5], P[1][4], P[2][3], S[5], Cout[5]);
Full_Adder FA7 (P[3][2], P[4][1], P[5][0], S[6], Cout[6]);
Full_Adder FA8 (P[0][6], P[1][5], P[2][4], S[7], Cout[7]);
Full_Adder FA9 (P[3][3], P[4][2], P[5][1], S[8], Cout[8]);
Full_Adder FA10 (P[0][7], P[1][6], P[2][5], S[9], Cout[9]);
Full_Adder FA11 (P[3][4], P[4][3], P[5][2], S[10], Cout[10]);
Half_Adder HA12 (P[6][1], P[7][0], S[11], Cout[11]);
Full_Adder FA13 (P[0][8], P[1][7], P[2][6], S[12], Cout[12]);
Full_Adder FA14 (P[3][5], P[4][4], P[5][3], S[13], Cout[13]);
Full_Adder FA15 (P[6][2], P[7][1], P[8][0], S[14], Cout[14]);
Full_Adder FA16 (P[0][9], P[1][8], P[2][7], S[15], Cout[15]);
Full_Adder FA17 (P[3][6], P[4][5], P[5][4], S[16], Cout[16]);
Full_Adder FA18 (P[6][3], P[7][2], P[8][1], S[17], Cout[17]);
Full_Adder FA19 (P[0][10], P[1][9], P[2][8], S[18], Cout[18]);
Full_Adder FA20 (P[3][7], P[4][6], P[5][5], S[19], Cout[19]);
Full_Adder FA21 (P[6][4], P[7][3], P[8][2], S[20], Cout[20]);
Half_Adder HA22 (P[9][1], P[10][0], S[21], Cout[21]);
Full_Adder FA23 (P[0][11], P[1][10], P[2][9], S[22], Cout[22]);
Full_Adder FA24 (P[3][8], P[4][7], P[5][6], S[23], Cout[23]);
Full_Adder FA25 (P[6][5], P[7][4], P[8][3], S[24], Cout[24]);
Full_Adder FA26 (P[9][2], P[10][1], P[11][0], S[25], Cout[25]);
Full_Adder FA27 (P[0][12], P[1][11], P[2][10], S[26], Cout[26]);
Full_Adder FA28 (P[3][9], P[4][8], P[5][7], S[27], Cout[27]);
Full_Adder FA29 (P[6][6], P[7][5], P[8][4], S[28], Cout[28]);
Full_Adder FA30 (P[9][3], P[10][2], P[11][1], S[29], Cout[29]);
Full_Adder FA31 (P[0][13], P[1][12], P[2][11], S[30], Cout[30]);
Full_Adder FA32 (P[3][10], P[4][9], P[5][8], S[31], Cout[31]);
Full_Adder FA33 (P[6][7], P[7][6], P[8][5], S[32], Cout[32]);
Full_Adder FA34 (P[9][4], P[10][3], P[11][2], S[33], Cout[33]);
Half_Adder HA35 (P[12][1], P[13][0], S[34], Cout[34]);
Full_Adder FA36 (P[0][14], P[1][13], P[2][12], S[35], Cout[35]);
Full_Adder FA37 (P[3][11], P[4][10], P[5][9], S[36], Cout[36]);
Full_Adder FA38 (P[6][8], P[7][7], P[8][6], S[37], Cout[37]);
Full_Adder FA39 (P[9][5], P[10][4], P[11][3], S[38], Cout[38]);
Full_Adder FA40 (P[12][2], P[13][1], P[14][0], S[39], Cout[39]);
Full_Adder FA41 (P[0][15], P[1][14], P[2][13], S[40], Cout[40]);
Full_Adder FA42 (P[3][12], P[4][11], P[5][10], S[41], Cout[41]);
Full_Adder FA43 (P[6][9], P[7][8], P[8][7], S[42], Cout[42]);
Full_Adder FA44 (P[9][6], P[10][5], P[11][4], S[43], Cout[43]);
Full_Adder FA45 (P[12][3], P[13][2], P[14][1], S[44], Cout[44]);
Full_Adder FA46 (P[1][15], P[2][14], P[3][13], S[45], Cout[45]);
Full_Adder FA47 (P[4][12], P[5][11], P[6][10], S[46], Cout[46]);
Full_Adder FA48 (P[7][9], P[8][8], P[9][7], S[47], Cout[47]);
Full_Adder FA49 (P[10][6], P[11][5], P[12][4], S[48], Cout[48]);
Half_Adder HA50 (P[13][3], P[14][2], S[49], Cout[49]);
Full_Adder FA51 (P[2][15], P[3][14], P[4][13], S[50], Cout[50]);
Full_Adder FA52 (P[5][12], P[6][11], P[7][10], S[51], Cout[51]);
Full_Adder FA53 (P[8][9], P[9][8], P[10][7], S[52], Cout[52]);
Full_Adder FA54 (P[11][6], P[12][5], P[13][4], S[53], Cout[53]);
Full_Adder FA55 (P[3][15], P[4][14], P[5][13], S[54], Cout[54]);
Full_Adder FA56 (P[6][12], P[7][11], P[8][10], S[55], Cout[55]);
Full_Adder FA57 (P[9][9], P[10][8], P[11][7], S[56], Cout[56]);
Full_Adder FA58 (P[12][6], P[13][5], P[14][4], S[57], Cout[57]);
Full_Adder FA59 (P[4][15], P[5][14], P[6][13], S[58], Cout[58]);
Full_Adder FA60 (P[7][12], P[8][11], P[9][10], S[59], Cout[59]);
Full_Adder FA61 (P[10][9], P[11][8], P[12][7], S[60], Cout[60]);
Half_Adder HA62 (P[13][6], P[14][5], S[61], Cout[61]);
Full_Adder FA63 (P[5][15], P[6][14], P[7][13], S[62], Cout[62]);
Full_Adder FA64 (P[8][12], P[9][11], P[10][10], S[63], Cout[63]);
Full_Adder FA65 (P[11][9], P[12][8], P[13][7], S[64], Cout[64]);
Full_Adder FA66 (P[6][15], P[7][14], P[8][13], S[65], Cout[65]);
Full_Adder FA67 (P[9][12], P[10][11], P[11][10], S[66], Cout[66]);
Full_Adder FA68 (P[12][9], P[13][8], P[14][7], S[67], Cout[67]);
Full_Adder FA69 (P[7][15], P[8][14], P[9][13], S[68], Cout[68]);
Full_Adder FA70 (P[10][12], P[11][11], P[12][10], S[69], Cout[69]);
Half_Adder HA71 (P[13][9], P[14][8], S[70], Cout[70]);
Full_Adder FA72 (P[8][15], P[9][14], P[10][13], S[71], Cout[71]);
Full_Adder FA73 (P[11][12], P[12][11], P[13][10], S[72], Cout[72]);
Full_Adder FA74 (P[9][15], P[10][14], P[11][13], S[73], Cout[73]);
Full_Adder FA75 (P[12][12], P[13][11], P[14][10], S[74], Cout[74]);
Full_Adder FA76 (P[10][15], P[11][14], P[12][13], S[75], Cout[75]);
Half_Adder HA77 (P[13][12], P[14][11], S[76], Cout[76]);
Full_Adder FA78 (P[11][15], P[12][14], P[13][13], S[77], Cout[77]);
Full_Adder FA79 (P[12][15], P[13][14], P[14][13], S[78], Cout[78]);
Half_Adder HA80 (P[13][15], P[14][14], S[79], Cout[79]);
Half_Adder HA81 (Cout[0], S[1], S[80], Cout[80]);
Full_Adder FA82 (P[3][0], Cout[1], S[2], S[81], Cout[81]);
Full_Adder FA83 (Cout[2], S[3], S[4], S[82], Cout[82]);
Full_Adder FA84 (Cout[3], Cout[4], S[5], S[83], Cout[83]);
Full_Adder FA85 (P[6][0], Cout[5], Cout[6], S[84], Cout[84]);
Half_Adder HA86 (S[7], S[8], S[85], Cout[85]);
Full_Adder FA87 (Cout[7], Cout[8], S[9], S[86], Cout[86]);
Half_Adder HA88 (S[10], S[11], S[87], Cout[87]);
Full_Adder FA89 (Cout[9], Cout[10], Cout[11], S[88], Cout[88]);
Full_Adder FA90 (S[12], S[13], S[14], S[89], Cout[89]);
Full_Adder FA91 (P[9][0], Cout[12], Cout[13], S[90], Cout[90]);
Full_Adder FA92 (Cout[14], S[15], S[16], S[91], Cout[91]);
Full_Adder FA93 (Cout[15], Cout[16], Cout[17], S[92], Cout[92]);
Full_Adder FA94 (S[18], S[19], S[20], S[93], Cout[93]);
Full_Adder FA95 (Cout[18], Cout[19], Cout[20], S[94], Cout[94]);
Full_Adder FA96 (Cout[21], S[22], S[23], S[95], Cout[95]);
Half_Adder HA97 (S[24], S[25], S[96], Cout[96]);
Full_Adder FA98 (P[12][0], Cout[22], Cout[23], S[97], Cout[97]);
Full_Adder FA99 (Cout[24], Cout[25], S[26], S[98], Cout[98]);
Full_Adder FA100 (S[27], S[28], S[29], S[99], Cout[99]);
Full_Adder FA101 (Cout[26], Cout[27], Cout[28], S[100], Cout[100]);
Full_Adder FA102 (Cout[29], S[30], S[31], S[101], Cout[101]);
Full_Adder FA103 (S[32], S[33], S[34], S[102], Cout[102]);
Full_Adder FA104 (Cout[30], Cout[31], Cout[32], S[103], Cout[103]);
Full_Adder FA105 (Cout[33], Cout[34], S[35], S[104], Cout[104]);
Full_Adder FA106 (S[36], S[37], S[38], S[105], Cout[105]);
Full_Adder FA107 (P[15][0], Cout[35], Cout[36], S[106], Cout[106]);
Full_Adder FA108 (Cout[37], Cout[38], Cout[39], S[107], Cout[107]);
Full_Adder FA109 (S[40], S[41], S[42], S[108], Cout[108]);
Full_Adder FA110 (P[15][1], Cout[40], Cout[41], S[109], Cout[109]);
Full_Adder FA111 (Cout[42], Cout[43], Cout[44], S[110], Cout[110]);
Full_Adder FA112 (S[45], S[46], S[47], S[111], Cout[111]);
Full_Adder FA113 (P[14][3], P[15][2], Cout[45], S[112], Cout[112]);
Full_Adder FA114 (Cout[46], Cout[47], Cout[48], S[113], Cout[113]);
Full_Adder FA115 (Cout[49], S[50], S[51], S[114], Cout[114]);
Full_Adder FA116 (P[15][3], Cout[50], Cout[51], S[115], Cout[115]);
Full_Adder FA117 (Cout[52], Cout[53], S[54], S[116], Cout[116]);
Full_Adder FA118 (P[15][4], Cout[54], Cout[55], S[117], Cout[117]);
Full_Adder FA119 (Cout[56], Cout[57], S[58], S[118], Cout[118]);
Full_Adder FA120 (P[14][6], P[15][5], Cout[58], S[119], Cout[119]);
Full_Adder FA121 (Cout[59], Cout[60], Cout[61], S[120], Cout[120]);
Full_Adder FA122 (P[15][6], Cout[62], Cout[63], S[121], Cout[121]);
Half_Adder HA123 (Cout[64], S[65], S[122], Cout[122]);
Full_Adder FA124 (P[15][7], Cout[65], Cout[66], S[123], Cout[123]);
Half_Adder HA125 (Cout[67], S[68], S[124], Cout[124]);
Full_Adder FA126 (P[14][9], P[15][8], Cout[68], S[125], Cout[125]);
Half_Adder HA127 (Cout[69], Cout[70], S[126], Cout[126]);
Full_Adder FA128 (P[15][9], Cout[71], Cout[72], S[127], Cout[127]);
Full_Adder FA129 (P[15][10], Cout[73], Cout[74], S[128], Cout[128]);
Full_Adder FA130 (P[14][12], P[15][11], Cout[75], S[129], Cout[129]);
Half_Adder HA131 (Cout[80], S[81], S[130], Cout[130]);
Half_Adder HA132 (Cout[81], S[82], S[131], Cout[131]);
Full_Adder FA133 (S[6], Cout[82], S[83], S[132], Cout[132]);
Full_Adder FA134 (Cout[83], S[84], S[85], S[133], Cout[133]);
Full_Adder FA135 (Cout[84], Cout[85], S[86], S[134], Cout[134]);
Full_Adder FA136 (Cout[86], Cout[87], S[88], S[135], Cout[135]);
Full_Adder FA137 (S[17], Cout[88], Cout[89], S[136], Cout[136]);
Half_Adder HA138 (S[90], S[91], S[137], Cout[137]);
Full_Adder FA139 (S[21], Cout[90], Cout[91], S[138], Cout[138]);
Half_Adder HA140 (S[92], S[93], S[139], Cout[139]);
Full_Adder FA141 (Cout[92], Cout[93], S[94], S[140], Cout[140]);
Half_Adder HA142 (S[95], S[96], S[141], Cout[141]);
Full_Adder FA143 (Cout[94], Cout[95], Cout[96], S[142], Cout[142]);
Full_Adder FA144 (S[97], S[98], S[99], S[143], Cout[143]);
Full_Adder FA145 (Cout[97], Cout[98], Cout[99], S[144], Cout[144]);
Full_Adder FA146 (S[100], S[101], S[102], S[145], Cout[145]);
Full_Adder FA147 (S[39], Cout[100], Cout[101], S[146], Cout[146]);
Full_Adder FA148 (Cout[102], S[103], S[104], S[147], Cout[147]);
Full_Adder FA149 (S[43], S[44], Cout[103], S[148], Cout[148]);
Full_Adder FA150 (Cout[104], Cout[105], S[106], S[149], Cout[149]);
Full_Adder FA151 (S[48], S[49], Cout[106], S[150], Cout[150]);
Full_Adder FA152 (Cout[107], Cout[108], S[109], S[151], Cout[151]);
Full_Adder FA153 (S[52], S[53], Cout[109], S[152], Cout[152]);
Full_Adder FA154 (Cout[110], Cout[111], S[112], S[153], Cout[153]);
Full_Adder FA155 (S[55], S[56], S[57], S[154], Cout[154]);
Full_Adder FA156 (Cout[112], Cout[113], Cout[114], S[155], Cout[155]);
Full_Adder FA157 (S[59], S[60], S[61], S[156], Cout[156]);
Half_Adder HA158 (Cout[115], Cout[116], S[157], Cout[157]);
Full_Adder FA159 (S[62], S[63], S[64], S[158], Cout[158]);
Half_Adder HA160 (Cout[117], Cout[118], S[159], Cout[159]);
Full_Adder FA161 (S[66], S[67], Cout[119], S[160], Cout[160]);
Full_Adder FA162 (S[69], S[70], Cout[121], S[161], Cout[161]);
Full_Adder FA163 (S[71], S[72], Cout[123], S[162], Cout[162]);
Full_Adder FA164 (S[73], S[74], Cout[125], S[163], Cout[163]);
Half_Adder HA165 (S[75], S[76], S[164], Cout[164]);
Half_Adder HA166 (Cout[76], S[77], S[165], Cout[165]);
Half_Adder HA167 (P[15][12], Cout[77], S[166], Cout[166]);
Half_Adder HA168 (Cout[130], S[131], S[167], Cout[167]);
Half_Adder HA169 (Cout[131], S[132], S[168], Cout[168]);
Half_Adder HA170 (Cout[132], S[133], S[169], Cout[169]);
Full_Adder FA171 (S[87], Cout[133], S[134], S[170], Cout[170]);
Full_Adder FA172 (S[89], Cout[134], S[135], S[171], Cout[171]);
Full_Adder FA173 (Cout[135], S[136], S[137], S[172], Cout[172]);
Full_Adder FA174 (Cout[136], Cout[137], S[138], S[173], Cout[173]);
Full_Adder FA175 (Cout[138], Cout[139], S[140], S[174], Cout[174]);
Full_Adder FA176 (Cout[140], Cout[141], S[142], S[175], Cout[175]);
Full_Adder FA177 (Cout[142], Cout[143], S[144], S[176], Cout[176]);
Full_Adder FA178 (S[105], Cout[144], Cout[145], S[177], Cout[177]);
Half_Adder HA179 (S[146], S[147], S[178], Cout[178]);
Full_Adder FA180 (S[107], S[108], Cout[146], S[179], Cout[179]);
Full_Adder FA181 (Cout[147], S[148], S[149], S[180], Cout[180]);
Full_Adder FA182 (S[110], S[111], Cout[148], S[181], Cout[181]);
Full_Adder FA183 (Cout[149], S[150], S[151], S[182], Cout[182]);
Full_Adder FA184 (S[113], S[114], Cout[150], S[183], Cout[183]);
Full_Adder FA185 (Cout[151], S[152], S[153], S[184], Cout[184]);
Full_Adder FA186 (S[115], S[116], Cout[152], S[185], Cout[185]);
Full_Adder FA187 (Cout[153], S[154], S[155], S[186], Cout[186]);
Full_Adder FA188 (S[117], S[118], Cout[154], S[187], Cout[187]);
Full_Adder FA189 (Cout[155], S[156], S[157], S[188], Cout[188]);
Full_Adder FA190 (S[119], S[120], Cout[156], S[189], Cout[189]);
Full_Adder FA191 (Cout[157], S[158], S[159], S[190], Cout[190]);
Full_Adder FA192 (Cout[120], S[121], S[122], S[191], Cout[191]);
Full_Adder FA193 (Cout[158], Cout[159], S[160], S[192], Cout[192]);
Full_Adder FA194 (Cout[122], S[123], S[124], S[193], Cout[193]);
Half_Adder HA195 (Cout[160], S[161], S[194], Cout[194]);
Full_Adder FA196 (Cout[124], S[125], S[126], S[195], Cout[195]);
Half_Adder HA197 (Cout[161], S[162], S[196], Cout[196]);
Full_Adder FA198 (Cout[126], S[127], Cout[162], S[197], Cout[197]);
Full_Adder FA199 (Cout[127], S[128], Cout[163], S[198], Cout[198]);
Full_Adder FA200 (Cout[128], S[129], Cout[164], S[199], Cout[199]);
Full_Adder FA201 (S[78], Cout[129], Cout[165], S[200], Cout[200]);
Full_Adder FA202 (P[15][13], Cout[78], S[79], S[201], Cout[201]);
Full_Adder FA203 (P[14][15], P[15][14], Cout[79], S[202], Cout[202]);
Half_Adder HA204 (Cout[167], S[168], S[203], Cout[203]);
Half_Adder HA205 (Cout[168], S[169], S[204], Cout[204]);
Half_Adder HA206 (Cout[169], S[170], S[205], Cout[205]);
Half_Adder HA207 (Cout[170], S[171], S[206], Cout[206]);
Half_Adder HA208 (Cout[171], S[172], S[207], Cout[207]);
Full_Adder FA209 (S[139], Cout[172], S[173], S[208], Cout[208]);
Full_Adder FA210 (S[141], Cout[173], S[174], S[209], Cout[209]);
Full_Adder FA211 (S[143], Cout[174], S[175], S[210], Cout[210]);
Full_Adder FA212 (S[145], Cout[175], S[176], S[211], Cout[211]);
Full_Adder FA213 (Cout[176], S[177], S[178], S[212], Cout[212]);
Full_Adder FA214 (Cout[177], Cout[178], S[179], S[213], Cout[213]);
Full_Adder FA215 (Cout[179], Cout[180], S[181], S[214], Cout[214]);
Full_Adder FA216 (Cout[181], Cout[182], S[183], S[215], Cout[215]);
Full_Adder FA217 (Cout[183], Cout[184], S[185], S[216], Cout[216]);
Full_Adder FA218 (Cout[185], Cout[186], S[187], S[217], Cout[217]);
Full_Adder FA219 (Cout[187], Cout[188], S[189], S[218], Cout[218]);
Full_Adder FA220 (Cout[189], Cout[190], S[191], S[219], Cout[219]);
Full_Adder FA221 (Cout[191], Cout[192], S[193], S[220], Cout[220]);
Full_Adder FA222 (Cout[193], Cout[194], S[195], S[221], Cout[221]);
Full_Adder FA223 (S[163], Cout[195], Cout[196], S[222], Cout[222]);
Half_Adder HA224 (S[164], Cout[197], S[223], Cout[223]);
Half_Adder HA225 (S[165], Cout[198], S[224], Cout[224]);
Half_Adder HA226 (S[166], Cout[199], S[225], Cout[225]);
Half_Adder HA227 (Cout[166], Cout[200], S[226], Cout[226]);
Half_Adder HA228 (Cout[203], S[204], S[227], Cout[227]);
Half_Adder HA229 (Cout[204], S[205], S[228], Cout[228]);
Half_Adder HA230 (Cout[205], S[206], S[229], Cout[229]);
Half_Adder HA231 (Cout[206], S[207], S[230], Cout[230]);
Half_Adder HA232 (Cout[207], S[208], S[231], Cout[231]);
Half_Adder HA233 (Cout[208], S[209], S[232], Cout[232]);
Half_Adder HA234 (Cout[209], S[210], S[233], Cout[233]);
Half_Adder HA235 (Cout[210], S[211], S[234], Cout[234]);
Half_Adder HA236 (Cout[211], S[212], S[235], Cout[235]);
Full_Adder FA237 (S[180], Cout[212], S[213], S[236], Cout[236]);
Full_Adder FA238 (S[182], Cout[213], S[214], S[237], Cout[237]);
Full_Adder FA239 (S[184], Cout[214], S[215], S[238], Cout[238]);
Full_Adder FA240 (S[186], Cout[215], S[216], S[239], Cout[239]);
Full_Adder FA241 (S[188], Cout[216], S[217], S[240], Cout[240]);
Full_Adder FA242 (S[190], Cout[217], S[218], S[241], Cout[241]);
Full_Adder FA243 (S[192], Cout[218], S[219], S[242], Cout[242]);
Full_Adder FA244 (S[194], Cout[219], S[220], S[243], Cout[243]);
Full_Adder FA245 (S[196], Cout[220], S[221], S[244], Cout[244]);
Full_Adder FA246 (S[197], Cout[221], S[222], S[245], Cout[245]);
Full_Adder FA247 (S[198], Cout[222], S[223], S[246], Cout[246]);
Full_Adder FA248 (S[199], Cout[223], S[224], S[247], Cout[247]);
Full_Adder FA249 (S[200], Cout[224], S[225], S[248], Cout[248]);
Full_Adder FA250 (S[201], Cout[225], S[226], S[249], Cout[249]);
Full_Adder FA251 (Cout[201], S[202], Cout[226], S[250], Cout[250]);
Half_Adder HA252 (P[15][15], Cout[202], S[251], Cout[251]);
Half_Adder HA253 (Cout[227], S[228], S[252], Cout[252]);
Full_Adder FA254 (Cout[228], S[229], Cout[252], S[253], Cout[253]);
Full_Adder FA255 (Cout[229], S[230], Cout[253], S[254], Cout[254]);
Full_Adder FA256 (Cout[230], S[231], Cout[254], S[255], Cout[255]);
Full_Adder FA257 (Cout[231], S[232], Cout[255], S[256], Cout[256]);
Full_Adder FA258 (Cout[232], S[233], Cout[256], S[257], Cout[257]);
Full_Adder FA259 (Cout[233], S[234], Cout[257], S[258], Cout[258]);
Full_Adder FA260 (Cout[234], S[235], Cout[258], S[259], Cout[259]);
Full_Adder FA261 (Cout[235], S[236], Cout[259], S[260], Cout[260]);
Full_Adder FA262 (Cout[236], S[237], Cout[260], S[261], Cout[261]);
Full_Adder FA263 (Cout[237], S[238], Cout[261], S[262], Cout[262]);
Full_Adder FA264 (Cout[238], S[239], Cout[262], S[263], Cout[263]);
Full_Adder FA265 (Cout[239], S[240], Cout[263], S[264], Cout[264]);
Full_Adder FA266 (Cout[240], S[241], Cout[264], S[265], Cout[265]);
Full_Adder FA267 (Cout[241], S[242], Cout[265], S[266], Cout[266]);
Full_Adder FA268 (Cout[242], S[243], Cout[266], S[267], Cout[267]);
Full_Adder FA269 (Cout[243], S[244], Cout[267], S[268], Cout[268]);
Full_Adder FA270 (Cout[244], S[245], Cout[268], S[269], Cout[269]);
Full_Adder FA271 (Cout[245], S[246], Cout[269], S[270], Cout[270]);
Full_Adder FA272 (Cout[246], S[247], Cout[270], S[271], Cout[271]);
Full_Adder FA273 (Cout[247], S[248], Cout[271], S[272], Cout[272]);
Full_Adder FA274 (Cout[248], S[249], Cout[272], S[273], Cout[273]);
Full_Adder FA275 (Cout[249], S[250], Cout[273], S[274], Cout[274]);
Full_Adder FA276 (Cout[250], S[251], Cout[274], S[275], Cout[275]);
Half_Adder HA277 (Cout[251], Cout[275], S[276], Cout[276]);

assign z[31] = S[276];
assign z[30] = S[275];
assign z[29] = S[274];
assign z[28] = S[273];
assign z[27] = S[272];
assign z[26] = S[271];
assign z[25] = S[270];
assign z[24] = S[269];
assign z[23] = S[268];
assign z[22] = S[267];
assign z[21] = S[266];
assign z[20] = S[265];
assign z[19] = S[264];
assign z[18] = S[263];
assign z[17] = S[262];
assign z[16] = S[261];
assign z[15] = S[260];
assign z[14] = S[259];
assign z[13] = S[258];
assign z[12] = S[257];
assign z[11] = S[256];
assign z[10] = S[255];
assign z[9] = S[254];
assign z[8] = S[253];
assign z[7] = S[252];
assign z[6] = S[227];
assign z[5] = S[203];
assign z[4] = S[167];
assign z[3] = S[130];
assign z[2] = S[80];
assign z[1] = S[0];
assign z[0] = P[0][0];

endmodule
