module dadda_unsigned_multiplier_CLA_16(product, A, B);
    input [15:0] A, B;
    output [31:0] product;

    wire [15:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;

	assign pp0[0] = A[0] & B[0];
	assign pp0[1] = A[0] & B[1];
	assign pp0[2] = A[0] & B[2];
	assign pp0[3] = A[0] & B[3];
	assign pp0[4] = A[0] & B[4];
	assign pp0[5] = A[0] & B[5];
	assign pp0[6] = A[0] & B[6];
	assign pp0[7] = A[0] & B[7];
	assign pp0[8] = A[0] & B[8];
	assign pp0[9] = A[0] & B[9];
	assign pp0[10] = A[0] & B[10];
	assign pp0[11] = A[0] & B[11];
	assign pp0[12] = A[0] & B[12];
	assign pp0[13] = A[0] & B[13];
	assign pp0[14] = A[0] & B[14];
	assign pp0[15] = A[0] & B[15];
	assign pp1[0] = A[1] & B[0];
	assign pp1[1] = A[1] & B[1];
	assign pp1[2] = A[1] & B[2];
	assign pp1[3] = A[1] & B[3];
	assign pp1[4] = A[1] & B[4];
	assign pp1[5] = A[1] & B[5];
	assign pp1[6] = A[1] & B[6];
	assign pp1[7] = A[1] & B[7];
	assign pp1[8] = A[1] & B[8];
	assign pp1[9] = A[1] & B[9];
	assign pp1[10] = A[1] & B[10];
	assign pp1[11] = A[1] & B[11];
	assign pp1[12] = A[1] & B[12];
	assign pp1[13] = A[1] & B[13];
	assign pp1[14] = A[1] & B[14];
	assign pp1[15] = A[1] & B[15];
	assign pp2[0] = A[2] & B[0];
	assign pp2[1] = A[2] & B[1];
	assign pp2[2] = A[2] & B[2];
	assign pp2[3] = A[2] & B[3];
	assign pp2[4] = A[2] & B[4];
	assign pp2[5] = A[2] & B[5];
	assign pp2[6] = A[2] & B[6];
	assign pp2[7] = A[2] & B[7];
	assign pp2[8] = A[2] & B[8];
	assign pp2[9] = A[2] & B[9];
	assign pp2[10] = A[2] & B[10];
	assign pp2[11] = A[2] & B[11];
	assign pp2[12] = A[2] & B[12];
	assign pp2[13] = A[2] & B[13];
	assign pp2[14] = A[2] & B[14];
	assign pp2[15] = A[2] & B[15];
	assign pp3[0] = A[3] & B[0];
	assign pp3[1] = A[3] & B[1];
	assign pp3[2] = A[3] & B[2];
	assign pp3[3] = A[3] & B[3];
	assign pp3[4] = A[3] & B[4];
	assign pp3[5] = A[3] & B[5];
	assign pp3[6] = A[3] & B[6];
	assign pp3[7] = A[3] & B[7];
	assign pp3[8] = A[3] & B[8];
	assign pp3[9] = A[3] & B[9];
	assign pp3[10] = A[3] & B[10];
	assign pp3[11] = A[3] & B[11];
	assign pp3[12] = A[3] & B[12];
	assign pp3[13] = A[3] & B[13];
	assign pp3[14] = A[3] & B[14];
	assign pp3[15] = A[3] & B[15];
	assign pp4[0] = A[4] & B[0];
	assign pp4[1] = A[4] & B[1];
	assign pp4[2] = A[4] & B[2];
	assign pp4[3] = A[4] & B[3];
	assign pp4[4] = A[4] & B[4];
	assign pp4[5] = A[4] & B[5];
	assign pp4[6] = A[4] & B[6];
	assign pp4[7] = A[4] & B[7];
	assign pp4[8] = A[4] & B[8];
	assign pp4[9] = A[4] & B[9];
	assign pp4[10] = A[4] & B[10];
	assign pp4[11] = A[4] & B[11];
	assign pp4[12] = A[4] & B[12];
	assign pp4[13] = A[4] & B[13];
	assign pp4[14] = A[4] & B[14];
	assign pp4[15] = A[4] & B[15];
	assign pp5[0] = A[5] & B[0];
	assign pp5[1] = A[5] & B[1];
	assign pp5[2] = A[5] & B[2];
	assign pp5[3] = A[5] & B[3];
	assign pp5[4] = A[5] & B[4];
	assign pp5[5] = A[5] & B[5];
	assign pp5[6] = A[5] & B[6];
	assign pp5[7] = A[5] & B[7];
	assign pp5[8] = A[5] & B[8];
	assign pp5[9] = A[5] & B[9];
	assign pp5[10] = A[5] & B[10];
	assign pp5[11] = A[5] & B[11];
	assign pp5[12] = A[5] & B[12];
	assign pp5[13] = A[5] & B[13];
	assign pp5[14] = A[5] & B[14];
	assign pp5[15] = A[5] & B[15];
	assign pp6[0] = A[6] & B[0];
	assign pp6[1] = A[6] & B[1];
	assign pp6[2] = A[6] & B[2];
	assign pp6[3] = A[6] & B[3];
	assign pp6[4] = A[6] & B[4];
	assign pp6[5] = A[6] & B[5];
	assign pp6[6] = A[6] & B[6];
	assign pp6[7] = A[6] & B[7];
	assign pp6[8] = A[6] & B[8];
	assign pp6[9] = A[6] & B[9];
	assign pp6[10] = A[6] & B[10];
	assign pp6[11] = A[6] & B[11];
	assign pp6[12] = A[6] & B[12];
	assign pp6[13] = A[6] & B[13];
	assign pp6[14] = A[6] & B[14];
	assign pp6[15] = A[6] & B[15];
	assign pp7[0] = A[7] & B[0];
	assign pp7[1] = A[7] & B[1];
	assign pp7[2] = A[7] & B[2];
	assign pp7[3] = A[7] & B[3];
	assign pp7[4] = A[7] & B[4];
	assign pp7[5] = A[7] & B[5];
	assign pp7[6] = A[7] & B[6];
	assign pp7[7] = A[7] & B[7];
	assign pp7[8] = A[7] & B[8];
	assign pp7[9] = A[7] & B[9];
	assign pp7[10] = A[7] & B[10];
	assign pp7[11] = A[7] & B[11];
	assign pp7[12] = A[7] & B[12];
	assign pp7[13] = A[7] & B[13];
	assign pp7[14] = A[7] & B[14];
	assign pp7[15] = A[7] & B[15];
	assign pp8[0] = A[8] & B[0];
	assign pp8[1] = A[8] & B[1];
	assign pp8[2] = A[8] & B[2];
	assign pp8[3] = A[8] & B[3];
	assign pp8[4] = A[8] & B[4];
	assign pp8[5] = A[8] & B[5];
	assign pp8[6] = A[8] & B[6];
	assign pp8[7] = A[8] & B[7];
	assign pp8[8] = A[8] & B[8];
	assign pp8[9] = A[8] & B[9];
	assign pp8[10] = A[8] & B[10];
	assign pp8[11] = A[8] & B[11];
	assign pp8[12] = A[8] & B[12];
	assign pp8[13] = A[8] & B[13];
	assign pp8[14] = A[8] & B[14];
	assign pp8[15] = A[8] & B[15];
	assign pp9[0] = A[9] & B[0];
	assign pp9[1] = A[9] & B[1];
	assign pp9[2] = A[9] & B[2];
	assign pp9[3] = A[9] & B[3];
	assign pp9[4] = A[9] & B[4];
	assign pp9[5] = A[9] & B[5];
	assign pp9[6] = A[9] & B[6];
	assign pp9[7] = A[9] & B[7];
	assign pp9[8] = A[9] & B[8];
	assign pp9[9] = A[9] & B[9];
	assign pp9[10] = A[9] & B[10];
	assign pp9[11] = A[9] & B[11];
	assign pp9[12] = A[9] & B[12];
	assign pp9[13] = A[9] & B[13];
	assign pp9[14] = A[9] & B[14];
	assign pp9[15] = A[9] & B[15];
	assign pp10[0] = A[10] & B[0];
	assign pp10[1] = A[10] & B[1];
	assign pp10[2] = A[10] & B[2];
	assign pp10[3] = A[10] & B[3];
	assign pp10[4] = A[10] & B[4];
	assign pp10[5] = A[10] & B[5];
	assign pp10[6] = A[10] & B[6];
	assign pp10[7] = A[10] & B[7];
	assign pp10[8] = A[10] & B[8];
	assign pp10[9] = A[10] & B[9];
	assign pp10[10] = A[10] & B[10];
	assign pp10[11] = A[10] & B[11];
	assign pp10[12] = A[10] & B[12];
	assign pp10[13] = A[10] & B[13];
	assign pp10[14] = A[10] & B[14];
	assign pp10[15] = A[10] & B[15];
	assign pp11[0] = A[11] & B[0];
	assign pp11[1] = A[11] & B[1];
	assign pp11[2] = A[11] & B[2];
	assign pp11[3] = A[11] & B[3];
	assign pp11[4] = A[11] & B[4];
	assign pp11[5] = A[11] & B[5];
	assign pp11[6] = A[11] & B[6];
	assign pp11[7] = A[11] & B[7];
	assign pp11[8] = A[11] & B[8];
	assign pp11[9] = A[11] & B[9];
	assign pp11[10] = A[11] & B[10];
	assign pp11[11] = A[11] & B[11];
	assign pp11[12] = A[11] & B[12];
	assign pp11[13] = A[11] & B[13];
	assign pp11[14] = A[11] & B[14];
	assign pp11[15] = A[11] & B[15];
	assign pp12[0] = A[12] & B[0];
	assign pp12[1] = A[12] & B[1];
	assign pp12[2] = A[12] & B[2];
	assign pp12[3] = A[12] & B[3];
	assign pp12[4] = A[12] & B[4];
	assign pp12[5] = A[12] & B[5];
	assign pp12[6] = A[12] & B[6];
	assign pp12[7] = A[12] & B[7];
	assign pp12[8] = A[12] & B[8];
	assign pp12[9] = A[12] & B[9];
	assign pp12[10] = A[12] & B[10];
	assign pp12[11] = A[12] & B[11];
	assign pp12[12] = A[12] & B[12];
	assign pp12[13] = A[12] & B[13];
	assign pp12[14] = A[12] & B[14];
	assign pp12[15] = A[12] & B[15];
	assign pp13[0] = A[13] & B[0];
	assign pp13[1] = A[13] & B[1];
	assign pp13[2] = A[13] & B[2];
	assign pp13[3] = A[13] & B[3];
	assign pp13[4] = A[13] & B[4];
	assign pp13[5] = A[13] & B[5];
	assign pp13[6] = A[13] & B[6];
	assign pp13[7] = A[13] & B[7];
	assign pp13[8] = A[13] & B[8];
	assign pp13[9] = A[13] & B[9];
	assign pp13[10] = A[13] & B[10];
	assign pp13[11] = A[13] & B[11];
	assign pp13[12] = A[13] & B[12];
	assign pp13[13] = A[13] & B[13];
	assign pp13[14] = A[13] & B[14];
	assign pp13[15] = A[13] & B[15];
	assign pp14[0] = A[14] & B[0];
	assign pp14[1] = A[14] & B[1];
	assign pp14[2] = A[14] & B[2];
	assign pp14[3] = A[14] & B[3];
	assign pp14[4] = A[14] & B[4];
	assign pp14[5] = A[14] & B[5];
	assign pp14[6] = A[14] & B[6];
	assign pp14[7] = A[14] & B[7];
	assign pp14[8] = A[14] & B[8];
	assign pp14[9] = A[14] & B[9];
	assign pp14[10] = A[14] & B[10];
	assign pp14[11] = A[14] & B[11];
	assign pp14[12] = A[14] & B[12];
	assign pp14[13] = A[14] & B[13];
	assign pp14[14] = A[14] & B[14];
	assign pp14[15] = A[14] & B[15];
	assign pp15[0] = A[15] & B[0];
	assign pp15[1] = A[15] & B[1];
	assign pp15[2] = A[15] & B[2];
	assign pp15[3] = A[15] & B[3];
	assign pp15[4] = A[15] & B[4];
	assign pp15[5] = A[15] & B[5];
	assign pp15[6] = A[15] & B[6];
	assign pp15[7] = A[15] & B[7];
	assign pp15[8] = A[15] & B[8];
	assign pp15[9] = A[15] & B[9];
	assign pp15[10] = A[15] & B[10];
	assign pp15[11] = A[15] & B[11];
	assign pp15[12] = A[15] & B[12];
	assign pp15[13] = A[15] & B[13];
	assign pp15[14] = A[15] & B[14];
	assign pp15[15] = A[15] & B[15];

	wire [240:0] S;
	wire [240:0] Cout;
	Half_Adder HA1 (pp0[13], pp1[12], S[1], Cout[1]);
	Full_Adder FA1 (pp0[14], pp1[13], pp2[12], S[2], Cout[2]);
	Half_Adder HA2 (pp3[11], pp4[10], S[3], Cout[3]);
	Full_Adder FA2 (pp0[15], pp1[14], pp2[13], S[4], Cout[4]);
	Full_Adder FA3 (pp3[12], pp4[11], pp5[10], S[5], Cout[5]);
	Half_Adder HA3 (pp6[9], pp7[8], S[6], Cout[6]);
	Full_Adder FA4 (pp1[15], pp2[14], pp3[13], S[7], Cout[7]);
	Full_Adder FA5 (pp4[12], pp5[11], pp6[10], S[8], Cout[8]);
	Half_Adder HA4 (pp7[9], pp8[8], S[9], Cout[9]);
	Full_Adder FA6 (pp2[15], pp3[14], pp4[13], S[10], Cout[10]);
	Full_Adder FA7 (pp5[12], pp6[11], pp7[10], S[11], Cout[11]);
	Full_Adder FA8 (pp3[15], pp4[14], pp5[13], S[12], Cout[12]);
	Half_Adder HA5 (pp0[9], pp1[8], S[13], Cout[13]);
	Full_Adder FA9 (pp0[10], pp1[9], pp2[8], S[14], Cout[14]);
	Half_Adder HA6 (pp3[7], pp4[6], S[15], Cout[15]);
	Full_Adder FA10 (pp0[11], pp1[10], pp2[9], S[16], Cout[16]);
	Full_Adder FA11 (pp3[8], pp4[7], pp5[6], S[17], Cout[17]);
	Half_Adder HA7 (pp6[5], pp7[4], S[18], Cout[18]);
	Full_Adder FA12 (pp0[12], pp1[11], pp2[10], S[19], Cout[19]);
	Full_Adder FA13 (pp3[9], pp4[8], pp5[7], S[20], Cout[20]);
	Full_Adder FA14 (pp6[6], pp7[5], pp8[4], S[21], Cout[21]);
	Half_Adder HA8 (pp9[3], pp10[2], S[22], Cout[22]);
	Full_Adder FA15 (pp2[11], pp3[10], pp4[9], S[23], Cout[23]);
	Full_Adder FA16 (pp5[8], pp6[7], pp7[6], S[24], Cout[24]);
	Full_Adder FA17 (pp8[5], pp9[4], pp10[3], S[25], Cout[25]);
	Full_Adder FA18 (pp11[2], pp12[1], pp13[0], S[26], Cout[26]);
	Full_Adder FA19 (pp5[9], pp6[8], pp7[7], S[27], Cout[27]);
	Full_Adder FA20 (pp8[6], pp9[5], pp10[4], S[28], Cout[28]);
	Full_Adder FA21 (pp11[3], pp12[2], pp13[1], S[29], Cout[29]);
	Full_Adder FA22 (pp14[0], Cout[1], S[2], S[30], Cout[30]);
	Full_Adder FA23 (pp8[7], pp9[6], pp10[5], S[31], Cout[31]);
	Full_Adder FA24 (pp11[4], pp12[3], pp13[2], S[32], Cout[32]);
	Full_Adder FA25 (pp14[1], pp15[0], Cout[2], S[33], Cout[33]);
	Full_Adder FA26 (Cout[3], S[4], S[5], S[34], Cout[34]);
	Full_Adder FA27 (pp9[7], pp10[6], pp11[5], S[35], Cout[35]);
	Full_Adder FA28 (pp12[4], pp13[3], pp14[2], S[36], Cout[36]);
	Full_Adder FA29 (pp15[1], Cout[4], Cout[5], S[37], Cout[37]);
	Full_Adder FA30 (Cout[6], S[7], S[8], S[38], Cout[38]);
	Full_Adder FA31 (pp8[9], pp9[8], pp10[7], S[39], Cout[39]);
	Full_Adder FA32 (pp11[6], pp12[5], pp13[4], S[40], Cout[40]);
	Full_Adder FA33 (pp14[3], pp15[2], Cout[7], S[41], Cout[41]);
	Full_Adder FA34 (Cout[8], Cout[9], S[10], S[42], Cout[42]);
	Full_Adder FA35 (pp6[12], pp7[11], pp8[10], S[43], Cout[43]);
	Full_Adder FA36 (pp9[9], pp10[8], pp11[7], S[44], Cout[44]);
	Full_Adder FA37 (pp12[6], pp13[5], pp14[4], S[45], Cout[45]);
	Full_Adder FA38 (pp15[3], Cout[10], Cout[11], S[46], Cout[46]);
	Full_Adder FA39 (pp4[15], pp5[14], pp6[13], S[47], Cout[47]);
	Full_Adder FA40 (pp7[12], pp8[11], pp9[10], S[48], Cout[48]);
	Full_Adder FA41 (pp10[9], pp11[8], pp12[7], S[49], Cout[49]);
	Full_Adder FA42 (pp13[6], pp14[5], pp15[4], S[50], Cout[50]);
	Full_Adder FA43 (pp5[15], pp6[14], pp7[13], S[51], Cout[51]);
	Full_Adder FA44 (pp8[12], pp9[11], pp10[10], S[52], Cout[52]);
	Full_Adder FA45 (pp11[9], pp12[8], pp13[7], S[53], Cout[53]);
	Full_Adder FA46 (pp6[15], pp7[14], pp8[13], S[54], Cout[54]);
	Full_Adder FA47 (pp9[12], pp10[11], pp11[10], S[55], Cout[55]);
	Full_Adder FA48 (pp7[15], pp8[14], pp9[13], S[56], Cout[56]);
	Half_Adder HA9 (pp0[6], pp1[5], S[57], Cout[57]);
	Full_Adder FA49 (pp0[7], pp1[6], pp2[5], S[58], Cout[58]);
	Half_Adder HA10 (pp3[4], pp4[3], S[59], Cout[59]);
	Full_Adder FA50 (pp0[8], pp1[7], pp2[6], S[60], Cout[60]);
	Full_Adder FA51 (pp3[5], pp4[4], pp5[3], S[61], Cout[61]);
	Half_Adder HA11 (pp6[2], pp7[1], S[62], Cout[62]);
	Full_Adder FA52 (pp2[7], pp3[6], pp4[5], S[63], Cout[63]);
	Full_Adder FA53 (pp5[4], pp6[3], pp7[2], S[64], Cout[64]);
	Full_Adder FA54 (pp8[1], pp9[0], S[13], S[65], Cout[65]);
	Full_Adder FA55 (pp5[5], pp6[4], pp7[3], S[66], Cout[66]);
	Full_Adder FA56 (pp8[2], pp9[1], pp10[0], S[67], Cout[67]);
	Full_Adder FA57 (Cout[13], S[14], S[15], S[68], Cout[68]);
	Full_Adder FA58 (pp8[3], pp9[2], pp10[1], S[69], Cout[69]);
	Full_Adder FA59 (pp11[0], Cout[14], Cout[15], S[70], Cout[70]);
	Full_Adder FA60 (S[16], S[17], S[18], S[71], Cout[71]);
	Full_Adder FA61 (pp11[1], pp12[0], Cout[16], S[72], Cout[72]);
	Full_Adder FA62 (Cout[17], Cout[18], S[19], S[73], Cout[73]);
	Full_Adder FA63 (S[20], S[21], S[22], S[74], Cout[74]);
	Full_Adder FA64 (S[1], Cout[19], Cout[20], S[75], Cout[75]);
	Full_Adder FA65 (Cout[21], Cout[22], S[23], S[76], Cout[76]);
	Full_Adder FA66 (S[24], S[25], S[26], S[77], Cout[77]);
	Full_Adder FA67 (S[3], Cout[23], Cout[24], S[78], Cout[78]);
	Full_Adder FA68 (Cout[25], Cout[26], S[27], S[79], Cout[79]);
	Full_Adder FA69 (S[28], S[29], S[30], S[80], Cout[80]);
	Full_Adder FA70 (S[6], Cout[27], Cout[28], S[81], Cout[81]);
	Full_Adder FA71 (Cout[29], Cout[30], S[31], S[82], Cout[82]);
	Full_Adder FA72 (S[32], S[33], S[34], S[83], Cout[83]);
	Full_Adder FA73 (S[9], Cout[31], Cout[32], S[84], Cout[84]);
	Full_Adder FA74 (Cout[33], Cout[34], S[35], S[85], Cout[85]);
	Full_Adder FA75 (S[36], S[37], S[38], S[86], Cout[86]);
	Full_Adder FA76 (S[11], Cout[35], Cout[36], S[87], Cout[87]);
	Full_Adder FA77 (Cout[37], Cout[38], S[39], S[88], Cout[88]);
	Full_Adder FA78 (S[40], S[41], S[42], S[89], Cout[89]);
	Full_Adder FA79 (S[12], Cout[39], Cout[40], S[90], Cout[90]);
	Full_Adder FA80 (Cout[41], Cout[42], S[43], S[91], Cout[91]);
	Full_Adder FA81 (S[44], S[45], S[46], S[92], Cout[92]);
	Full_Adder FA82 (Cout[12], Cout[43], Cout[44], S[93], Cout[93]);
	Full_Adder FA83 (Cout[45], Cout[46], S[47], S[94], Cout[94]);
	Full_Adder FA84 (S[48], S[49], S[50], S[95], Cout[95]);
	Full_Adder FA85 (pp14[6], pp15[5], Cout[47], S[96], Cout[96]);
	Full_Adder FA86 (Cout[48], Cout[49], Cout[50], S[97], Cout[97]);
	Full_Adder FA87 (S[51], S[52], S[53], S[98], Cout[98]);
	Full_Adder FA88 (pp12[9], pp13[8], pp14[7], S[99], Cout[99]);
	Full_Adder FA89 (pp15[6], Cout[51], Cout[52], S[100], Cout[100]);
	Full_Adder FA90 (Cout[53], S[54], S[55], S[101], Cout[101]);
	Full_Adder FA91 (pp10[12], pp11[11], pp12[10], S[102], Cout[102]);
	Full_Adder FA92 (pp13[9], pp14[8], pp15[7], S[103], Cout[103]);
	Full_Adder FA93 (Cout[54], Cout[55], S[56], S[104], Cout[104]);
	Full_Adder FA94 (pp8[15], pp9[14], pp10[13], S[105], Cout[105]);
	Full_Adder FA95 (pp11[12], pp12[11], pp13[10], S[106], Cout[106]);
	Full_Adder FA96 (pp14[9], pp15[8], Cout[56], S[107], Cout[107]);
	Full_Adder FA97 (pp9[15], pp10[14], pp11[13], S[108], Cout[108]);
	Full_Adder FA98 (pp12[12], pp13[11], pp14[10], S[109], Cout[109]);
	Full_Adder FA99 (pp10[15], pp11[14], pp12[13], S[110], Cout[110]);
	Half_Adder HA12 (pp0[4], pp1[3], S[111], Cout[111]);
	Full_Adder FA100 (pp0[5], pp1[4], pp2[3], S[112], Cout[112]);
	Half_Adder HA13 (pp3[2], pp4[1], S[113], Cout[113]);
	Full_Adder FA101 (pp2[4], pp3[3], pp4[2], S[114], Cout[114]);
	Full_Adder FA102 (pp5[1], pp6[0], S[57], S[115], Cout[115]);
	Full_Adder FA103 (pp5[2], pp6[1], pp7[0], S[116], Cout[116]);
	Full_Adder FA104 (Cout[57], S[58], S[59], S[117], Cout[117]);
	Full_Adder FA105 (pp8[0], Cout[58], Cout[59], S[118], Cout[118]);
	Full_Adder FA106 (S[60], S[61], S[62], S[119], Cout[119]);
	Full_Adder FA107 (Cout[60], Cout[61], Cout[62], S[120], Cout[120]);
	Full_Adder FA108 (S[63], S[64], S[65], S[121], Cout[121]);
	Full_Adder FA109 (Cout[63], Cout[64], Cout[65], S[122], Cout[122]);
	Full_Adder FA110 (S[66], S[67], S[68], S[123], Cout[123]);
	Full_Adder FA111 (Cout[66], Cout[67], Cout[68], S[124], Cout[124]);
	Full_Adder FA112 (S[69], S[70], S[71], S[125], Cout[125]);
	Full_Adder FA113 (Cout[69], Cout[70], Cout[71], S[126], Cout[126]);
	Full_Adder FA114 (S[72], S[73], S[74], S[127], Cout[127]);
	Full_Adder FA115 (Cout[72], Cout[73], Cout[74], S[128], Cout[128]);
	Full_Adder FA116 (S[75], S[76], S[77], S[129], Cout[129]);
	Full_Adder FA117 (Cout[75], Cout[76], Cout[77], S[130], Cout[130]);
	Full_Adder FA118 (S[78], S[79], S[80], S[131], Cout[131]);
	Full_Adder FA119 (Cout[78], Cout[79], Cout[80], S[132], Cout[132]);
	Full_Adder FA120 (S[81], S[82], S[83], S[133], Cout[133]);
	Full_Adder FA121 (Cout[81], Cout[82], Cout[83], S[134], Cout[134]);
	Full_Adder FA122 (S[84], S[85], S[86], S[135], Cout[135]);
	Full_Adder FA123 (Cout[84], Cout[85], Cout[86], S[136], Cout[136]);
	Full_Adder FA124 (S[87], S[88], S[89], S[137], Cout[137]);
	Full_Adder FA125 (Cout[87], Cout[88], Cout[89], S[138], Cout[138]);
	Full_Adder FA126 (S[90], S[91], S[92], S[139], Cout[139]);
	Full_Adder FA127 (Cout[90], Cout[91], Cout[92], S[140], Cout[140]);
	Full_Adder FA128 (S[93], S[94], S[95], S[141], Cout[141]);
	Full_Adder FA129 (Cout[93], Cout[94], Cout[95], S[142], Cout[142]);
	Full_Adder FA130 (S[96], S[97], S[98], S[143], Cout[143]);
	Full_Adder FA131 (Cout[96], Cout[97], Cout[98], S[144], Cout[144]);
	Full_Adder FA132 (S[99], S[100], S[101], S[145], Cout[145]);
	Full_Adder FA133 (Cout[99], Cout[100], Cout[101], S[146], Cout[146]);
	Full_Adder FA134 (S[102], S[103], S[104], S[147], Cout[147]);
	Full_Adder FA135 (Cout[102], Cout[103], Cout[104], S[148], Cout[148]);
	Full_Adder FA136 (S[105], S[106], S[107], S[149], Cout[149]);
	Full_Adder FA137 (pp15[9], Cout[105], Cout[106], S[150], Cout[150]);
	Full_Adder FA138 (Cout[107], S[108], S[109], S[151], Cout[151]);
	Full_Adder FA139 (pp13[12], pp14[11], pp15[10], S[152], Cout[152]);
	Full_Adder FA140 (Cout[108], Cout[109], S[110], S[153], Cout[153]);
	Full_Adder FA141 (pp11[15], pp12[14], pp13[13], S[154], Cout[154]);
	Full_Adder FA142 (pp14[12], pp15[11], Cout[110], S[155], Cout[155]);
	Full_Adder FA143 (pp12[15], pp13[14], pp14[13], S[156], Cout[156]);
	Half_Adder HA14 (pp0[3], pp1[2], S[157], Cout[157]);
	Full_Adder FA144 (pp2[2], pp3[1], pp4[0], S[158], Cout[158]);
	Full_Adder FA145 (pp5[0], Cout[111], S[112], S[159], Cout[159]);
	Full_Adder FA146 (Cout[112], Cout[113], S[114], S[160], Cout[160]);
	Full_Adder FA147 (Cout[114], Cout[115], S[116], S[161], Cout[161]);
	Full_Adder FA148 (Cout[116], Cout[117], S[118], S[162], Cout[162]);
	Full_Adder FA149 (Cout[118], Cout[119], S[120], S[163], Cout[163]);
	Full_Adder FA150 (Cout[120], Cout[121], S[122], S[164], Cout[164]);
	Full_Adder FA151 (Cout[122], Cout[123], S[124], S[165], Cout[165]);
	Full_Adder FA152 (Cout[124], Cout[125], S[126], S[166], Cout[166]);
	Full_Adder FA153 (Cout[126], Cout[127], S[128], S[167], Cout[167]);
	Full_Adder FA154 (Cout[128], Cout[129], S[130], S[168], Cout[168]);
	Full_Adder FA155 (Cout[130], Cout[131], S[132], S[169], Cout[169]);
	Full_Adder FA156 (Cout[132], Cout[133], S[134], S[170], Cout[170]);
	Full_Adder FA157 (Cout[134], Cout[135], S[136], S[171], Cout[171]);
	Full_Adder FA158 (Cout[136], Cout[137], S[138], S[172], Cout[172]);
	Full_Adder FA159 (Cout[138], Cout[139], S[140], S[173], Cout[173]);
	Full_Adder FA160 (Cout[140], Cout[141], S[142], S[174], Cout[174]);
	Full_Adder FA161 (Cout[142], Cout[143], S[144], S[175], Cout[175]);
	Full_Adder FA162 (Cout[144], Cout[145], S[146], S[176], Cout[176]);
	Full_Adder FA163 (Cout[146], Cout[147], S[148], S[177], Cout[177]);
	Full_Adder FA164 (Cout[148], Cout[149], S[150], S[178], Cout[178]);
	Full_Adder FA165 (Cout[150], Cout[151], S[152], S[179], Cout[179]);
	Full_Adder FA166 (Cout[152], Cout[153], S[154], S[180], Cout[180]);
	Full_Adder FA167 (pp15[12], Cout[154], Cout[155], S[181], Cout[181]);
	Full_Adder FA168 (pp13[15], pp14[14], pp15[13], S[182], Cout[182]);
	Half_Adder HA15 (pp0[2], pp1[1], S[183], Cout[183]);
	Full_Adder FA169 (pp2[1], pp3[0], S[157], S[184], Cout[184]);
	Full_Adder FA170 (S[111], Cout[157], S[158], S[185], Cout[185]);
	Full_Adder FA171 (S[113], Cout[158], S[159], S[186], Cout[186]);
	Full_Adder FA172 (S[115], Cout[159], S[160], S[187], Cout[187]);
	Full_Adder FA173 (S[117], Cout[160], S[161], S[188], Cout[188]);
	Full_Adder FA174 (S[119], Cout[161], S[162], S[189], Cout[189]);
	Full_Adder FA175 (S[121], Cout[162], S[163], S[190], Cout[190]);
	Full_Adder FA176 (S[123], Cout[163], S[164], S[191], Cout[191]);
	Full_Adder FA177 (S[125], Cout[164], S[165], S[192], Cout[192]);
	Full_Adder FA178 (S[127], Cout[165], S[166], S[193], Cout[193]);
	Full_Adder FA179 (S[129], Cout[166], S[167], S[194], Cout[194]);
	Full_Adder FA180 (S[131], Cout[167], S[168], S[195], Cout[195]);
	Full_Adder FA181 (S[133], Cout[168], S[169], S[196], Cout[196]);
	Full_Adder FA182 (S[135], Cout[169], S[170], S[197], Cout[197]);
	Full_Adder FA183 (S[137], Cout[170], S[171], S[198], Cout[198]);
	Full_Adder FA184 (S[139], Cout[171], S[172], S[199], Cout[199]);
	Full_Adder FA185 (S[141], Cout[172], S[173], S[200], Cout[200]);
	Full_Adder FA186 (S[143], Cout[173], S[174], S[201], Cout[201]);
	Full_Adder FA187 (S[145], Cout[174], S[175], S[202], Cout[202]);
	Full_Adder FA188 (S[147], Cout[175], S[176], S[203], Cout[203]);
	Full_Adder FA189 (S[149], Cout[176], S[177], S[204], Cout[204]);
	Full_Adder FA190 (S[151], Cout[177], S[178], S[205], Cout[205]);
	Full_Adder FA191 (S[153], Cout[178], S[179], S[206], Cout[206]);
	Full_Adder FA192 (S[155], Cout[179], S[180], S[207], Cout[207]);
	Full_Adder FA193 (S[156], Cout[180], S[181], S[208], Cout[208]);
	Full_Adder FA194 (Cout[156], Cout[181], S[182], S[209], Cout[209]);
	Full_Adder FA195 (pp14[15], pp15[14], Cout[182], S[210], Cout[210]);


    wire [29:0] G, P, C;
    assign G[0]  =  pp0[1]    & pp1[0];
    assign G[1]  =  pp2[0]    & S[183];
    assign G[2]  =  Cout[183] & S[184];
    assign G[3]  =  Cout[184] & S[185];
    assign G[4]  =  Cout[185] & S[186];
    assign G[5]  =  Cout[186] & S[187];
    assign G[6]  =  Cout[187] & S[188];
    assign G[7]  =  Cout[188] & S[189];
    assign G[8]  =  Cout[189] & S[190];
    assign G[9]  =  Cout[190] & S[191];
    assign G[10] =  Cout[191] & S[192];
    assign G[11] = Cout[192] & S[193];
    assign G[12] = Cout[193] & S[194];
    assign G[13] = Cout[194] & S[195];
    assign G[14] = Cout[195] & S[196];
    assign G[15] = Cout[196] & S[197];
    assign G[16] = Cout[197] & S[198];
    assign G[17] = Cout[198] & S[199];
    assign G[18] = Cout[199] & S[200];
    assign G[19] = Cout[200] & S[201];
    assign G[20] = Cout[201] & S[202];
    assign G[21] = Cout[202] & S[203];
    assign G[22] = Cout[203] & S[204];
    assign G[23] = Cout[204] & S[205];
    assign G[24] = Cout[205] & S[206];
    assign G[25] = Cout[206] & S[207];
    assign G[26] = Cout[207] & S[208];
    assign G[27] = Cout[208] & S[209];
    assign G[28] = Cout[209] & S[210];
    assign G[29] = pp15[15]  & Cout[210];
    assign P[0]  = pp0[1]    ^ pp1[0];
    assign P[1]  = pp2[0]    ^ S[183];
    assign P[2]  =  Cout[183] ^ S[184];
    assign P[3]  =  Cout[184] ^ S[185];
    assign P[4]  =  Cout[185] ^ S[186];
    assign P[5]  =  Cout[186] ^ S[187];
    assign P[6]  =  Cout[187] ^ S[188];
    assign P[7]  =  Cout[188] ^ S[189];
    assign P[8]  =  Cout[189] ^ S[190];
    assign P[9]  =  Cout[190] ^ S[191];
    assign P[10] =  Cout[191] ^ S[192];
    assign P[11] = Cout[192] ^ S[193];
    assign P[12] = Cout[193] ^ S[194];
    assign P[13] = Cout[194] ^ S[195];
    assign P[14] = Cout[195] ^ S[196];
    assign P[15] = Cout[196] ^ S[197];
    assign P[16] = Cout[197] ^ S[198];
    assign P[17] = Cout[198] ^ S[199];
    assign P[18] = Cout[199] ^ S[200];
    assign P[19] = Cout[200] ^ S[201];
    assign P[20] = Cout[201] ^ S[202];
    assign P[21] = Cout[202] ^ S[203];
    assign P[22] = Cout[203] ^ S[204];
    assign P[23] = Cout[204] ^ S[205];
    assign P[24] = Cout[205] ^ S[206];
    assign P[25] = Cout[206] ^ S[207];
    assign P[26] = Cout[207] ^ S[208];
    assign P[27] = Cout[208] ^ S[209];
    assign P[28] = Cout[209] ^ S[210];
    assign P[29] = pp15[15]  ^ Cout[210];

    assign C[0] = 0;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign product[31] = G[29] | (P[29] & C[29]);

    assign product[1]  = P[0];
    assign product[2]  = P[1]  ^ C[1];
    assign product[3]  = P[2]  ^ C[2];
    assign product[4]  = P[3]  ^ C[3];
    assign product[5]  = P[4]  ^ C[4];
    assign product[6]  = P[5]  ^ C[5];
    assign product[7]  = P[6]  ^ C[6];
    assign product[8]  = P[7]  ^ C[7];
    assign product[9]  = P[8]  ^ C[8];
    assign product[10] = P[9]  ^ C[9];
    assign product[11] = P[10] ^ C[10];
    assign product[12] = P[11] ^ C[11];
    assign product[13] = P[12] ^ C[12];
    assign product[14] = P[13] ^ C[13];
    assign product[15] = P[14] ^ C[14];
    assign product[16] = P[15] ^ C[15];
    assign product[17] = P[16] ^ C[16];
    assign product[18] = P[17] ^ C[17];
    assign product[19] = P[18] ^ C[18];
    assign product[20] = P[19] ^ C[19];
    assign product[21] = P[20] ^ C[20];
    assign product[22] = P[21] ^ C[21];
    assign product[23] = P[22] ^ C[22];
    assign product[24] = P[23] ^ C[23];
    assign product[25] = P[24] ^ C[24];
    assign product[26] = P[25] ^ C[25];
    assign product[27] = P[26] ^ C[26];
    assign product[28] = P[27] ^ C[27];
    assign product[29] = P[28] ^ C[28];
    assign product[30] = P[29] ^ C[29];


    assign product[0] = pp0[0];

	
endmodule

module Half_Adder(input wire in1,
                  input wire in2,
				  output wire sum,
                  output wire cout);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(input wire in1,
                  input wire in2,
                  input wire cin,
				  output wire sum,
                  output wire cout);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule
