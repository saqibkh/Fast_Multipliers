module multiplier_16bits_version14(product, A, B);

    output [31:0] product;
    input [15:0] A, B;

    wire [15:0] pp0;
    wire [15:0] pp1;
    wire [15:0] pp2;
    wire [15:0] pp3;
    wire [15:0] pp4;
    wire [15:0] pp5;
    wire [15:0] pp6;
    wire [15:0] pp7;
    wire [15:0] pp8;
    wire [15:0] pp9;
    wire [15:0] pp10;
    wire [15:0] pp11;
    wire [15:0] pp12;
    wire [15:0] pp13;
    wire [15:0] pp14;
    wire [15:0] pp15;


    assign pp0 = A[0] ? B: 16'b0000000000000000;
    assign pp1 = A[1] ? B: 16'b0000000000000000;
    assign pp2 = A[2] ? B: 16'b0000000000000000;
    assign pp3 = A[3] ? B: 16'b0000000000000000;
    assign pp4 = A[4] ? B: 16'b0000000000000000;
    assign pp5 = A[5] ? B: 16'b0000000000000000;
    assign pp6 = A[6] ? B: 16'b0000000000000000;
    assign pp7 = A[7] ? B: 16'b0000000000000000;
    assign pp8 = A[8] ? B: 16'b0000000000000000;
    assign pp9 = A[9] ? B: 16'b0000000000000000;
    assign pp10 = A[10] ? B: 16'b0000000000000000;
    assign pp11 = A[11] ? B: 16'b0000000000000000;
    assign pp12 = A[12] ? B: 16'b0000000000000000;
    assign pp13 = A[13] ? B: 16'b0000000000000000;
    assign pp14 = A[14] ? B: 16'b0000000000000000;
    assign pp15 = A[15] ? B: 16'b0000000000000000;


    /*Stage 1*/
    wire[0:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[11]};
    assign in1_2 = {pp1[10]};
    Half_Adder HA_1(s1, c1, in1_1, in1_2);
    wire[0:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp1[11]};
    assign in2_2 = {pp2[10]};
    Full_Adder FA_2(s2, c2, in2_1, in2_2, pp0[12]);
    wire[0:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp3[9]};
    assign in3_2 = {pp4[8]};
    Half_Adder HA_3(s3, c3, in3_1, in3_2);
    wire[0:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp1[12]};
    assign in4_2 = {pp2[11]};
    Full_Adder FA_4(s4, c4, in4_1, in4_2, pp0[13]);
    wire[0:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp4[9]};
    assign in5_2 = {pp5[8]};
    Full_Adder FA_5(s5, c5, in5_1, in5_2, pp3[10]);
    wire[0:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp6[7]};
    assign in6_2 = {pp7[6]};
    Half_Adder HA_6(s6, c6, in6_1, in6_2);
    wire[0:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp1[13]};
    assign in7_2 = {pp2[12]};
    Full_Adder FA_7(s7, c7, in7_1, in7_2, pp0[14]);
    wire[0:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp4[10]};
    assign in8_2 = {pp5[9]};
    Full_Adder FA_8(s8, c8, in8_1, in8_2, pp3[11]);
    wire[0:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp7[7]};
    assign in9_2 = {pp8[6]};
    Full_Adder FA_9(s9, c9, in9_1, in9_2, pp6[8]);
    wire[0:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp9[5]};
    assign in10_2 = {pp10[4]};
    Half_Adder HA_10(s10, c10, in10_1, in10_2);
    wire[0:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp1[14]};
    assign in11_2 = {pp2[13]};
    Full_Adder FA_11(s11, c11, in11_1, in11_2, pp0[15]);
    wire[0:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp4[11]};
    assign in12_2 = {pp5[10]};
    Full_Adder FA_12(s12, c12, in12_1, in12_2, pp3[12]);
    wire[0:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp7[8]};
    assign in13_2 = {pp8[7]};
    Full_Adder FA_13(s13, c13, in13_1, in13_2, pp6[9]);
    wire[0:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp10[5]};
    assign in14_2 = {pp11[4]};
    Full_Adder FA_14(s14, c14, in14_1, in14_2, pp9[6]);
    wire[0:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp12[3]};
    assign in15_2 = {pp13[2]};
    Half_Adder HA_15(s15, c15, in15_1, in15_2);
    wire[0:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp2[14]};
    assign in16_2 = {pp3[13]};
    Full_Adder FA_16(s16, c16, in16_1, in16_2, pp1[15]);
    wire[0:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp5[11]};
    assign in17_2 = {pp6[10]};
    Full_Adder FA_17(s17, c17, in17_1, in17_2, pp4[12]);
    wire[0:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp8[8]};
    assign in18_2 = {pp9[7]};
    Full_Adder FA_18(s18, c18, in18_1, in18_2, pp7[9]);
    wire[0:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp11[5]};
    assign in19_2 = {pp12[4]};
    Full_Adder FA_19(s19, c19, in19_1, in19_2, pp10[6]);
    wire[0:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp13[3]};
    assign in20_2 = {pp14[2]};
    Half_Adder HA_20(s20, c20, in20_1, in20_2);
    wire[0:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp3[14]};
    assign in21_2 = {pp4[13]};
    Full_Adder FA_21(s21, c21, in21_1, in21_2, pp2[15]);
    wire[0:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp6[11]};
    assign in22_2 = {pp7[10]};
    Full_Adder FA_22(s22, c22, in22_1, in22_2, pp5[12]);
    wire[0:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp9[8]};
    assign in23_2 = {pp10[7]};
    Full_Adder FA_23(s23, c23, in23_1, in23_2, pp8[9]);
    wire[0:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp12[5]};
    assign in24_2 = {pp13[4]};
    Full_Adder FA_24(s24, c24, in24_1, in24_2, pp11[6]);
    wire[0:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp4[14]};
    assign in25_2 = {pp5[13]};
    Full_Adder FA_25(s25, c25, in25_1, in25_2, pp3[15]);
    wire[0:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp7[11]};
    assign in26_2 = {pp8[10]};
    Full_Adder FA_26(s26, c26, in26_1, in26_2, pp6[12]);
    wire[0:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp10[8]};
    assign in27_2 = {pp11[7]};
    Full_Adder FA_27(s27, c27, in27_1, in27_2, pp9[9]);
    wire[0:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp5[14]};
    assign in28_2 = {pp6[13]};
    Full_Adder FA_28(s28, c28, in28_1, in28_2, pp4[15]);
    wire[0:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp8[11]};
    assign in29_2 = {pp9[10]};
    Full_Adder FA_29(s29, c29, in29_1, in29_2, pp7[12]);
    wire[0:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp6[14]};
    assign in30_2 = {pp7[13]};
    Full_Adder FA_30(s30, c30, in30_1, in30_2, pp5[15]);

    /*Stage 2*/
    wire[0:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp0[8]};
    assign in31_2 = {pp1[7]};
    Half_Adder HA_31(s31, c31, in31_1, in31_2);
    wire[0:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp1[8]};
    assign in32_2 = {pp2[7]};
    Full_Adder FA_32(s32, c32, in32_1, in32_2, pp0[9]);
    wire[0:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp3[6]};
    assign in33_2 = {pp4[5]};
    Half_Adder HA_33(s33, c33, in33_1, in33_2);
    wire[0:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp1[9]};
    assign in34_2 = {pp2[8]};
    Full_Adder FA_34(s34, c34, in34_1, in34_2, pp0[10]);
    wire[0:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp4[6]};
    assign in35_2 = {pp5[5]};
    Full_Adder FA_35(s35, c35, in35_1, in35_2, pp3[7]);
    wire[0:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp6[4]};
    assign in36_2 = {pp7[3]};
    Half_Adder HA_36(s36, c36, in36_1, in36_2);
    wire[0:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp3[8]};
    assign in37_2 = {pp4[7]};
    Full_Adder FA_37(s37, c37, in37_1, in37_2, pp2[9]);
    wire[0:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp6[5]};
    assign in38_2 = {pp7[4]};
    Full_Adder FA_38(s38, c38, in38_1, in38_2, pp5[6]);
    wire[0:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp9[2]};
    assign in39_2 = {pp10[1]};
    Full_Adder FA_39(s39, c39, in39_1, in39_2, pp8[3]);
    wire[0:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp6[6]};
    assign in40_2 = {pp7[5]};
    Full_Adder FA_40(s40, c40, in40_1, in40_2, pp5[7]);
    wire[0:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp9[3]};
    assign in41_2 = {pp10[2]};
    Full_Adder FA_41(s41, c41, in41_1, in41_2, pp8[4]);
    wire[0:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp12[0]};
    assign in42_2 = {c1};
    Full_Adder FA_42(s42, c42, in42_1, in42_2, pp11[1]);
    wire[0:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp9[4]};
    assign in43_2 = {pp10[3]};
    Full_Adder FA_43(s43, c43, in43_1, in43_2, pp8[5]);
    wire[0:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp12[1]};
    assign in44_2 = {pp13[0]};
    Full_Adder FA_44(s44, c44, in44_1, in44_2, pp11[2]);
    wire[0:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {c3};
    assign in45_2 = {s4[0]};
    Full_Adder FA_45(s45, c45, in45_1, in45_2, c2);
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp12[2]};
    assign in46_2 = {pp13[1]};
    Full_Adder FA_46(s46, c46, in46_1, in46_2, pp11[3]);
    wire[0:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {c4};
    assign in47_2 = {c5};
    Full_Adder FA_47(s47, c47, in47_1, in47_2, pp14[0]);
    wire[0:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {s7[0]};
    assign in48_2 = {s8[0]};
    Full_Adder FA_48(s48, c48, in48_1, in48_2, c6);
    wire[0:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp15[0]};
    assign in49_2 = {c7};
    Full_Adder FA_49(s49, c49, in49_1, in49_2, pp14[1]);
    wire[0:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {c9};
    assign in50_2 = {c10};
    Full_Adder FA_50(s50, c50, in50_1, in50_2, c8);
    wire[0:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {s12[0]};
    assign in51_2 = {s13[0]};
    Full_Adder FA_51(s51, c51, in51_1, in51_2, s11[0]);
    wire[0:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {c11};
    assign in52_2 = {c12};
    Full_Adder FA_52(s52, c52, in52_1, in52_2, pp15[1]);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {c14};
    assign in53_2 = {c15};
    Full_Adder FA_53(s53, c53, in53_1, in53_2, c13);
    wire[0:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {s17[0]};
    assign in54_2 = {s18[0]};
    Full_Adder FA_54(s54, c54, in54_1, in54_2, s16[0]);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp15[2]};
    assign in55_2 = {c16};
    Full_Adder FA_55(s55, c55, in55_1, in55_2, pp14[3]);
    wire[0:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {c18};
    assign in56_2 = {c19};
    Full_Adder FA_56(s56, c56, in56_1, in56_2, c17);
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {s21[0]};
    assign in57_2 = {s22[0]};
    Full_Adder FA_57(s57, c57, in57_1, in57_2, c20);
    wire[0:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp13[5]};
    assign in58_2 = {pp14[4]};
    Full_Adder FA_58(s58, c58, in58_1, in58_2, pp12[6]);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {c21};
    assign in59_2 = {c22};
    Full_Adder FA_59(s59, c59, in59_1, in59_2, pp15[3]);
    wire[0:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {c24};
    assign in60_2 = {s25[0]};
    Full_Adder FA_60(s60, c60, in60_1, in60_2, c23);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp11[8]};
    assign in61_2 = {pp12[7]};
    Full_Adder FA_61(s61, c61, in61_1, in61_2, pp10[9]);
    wire[0:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp14[5]};
    assign in62_2 = {pp15[4]};
    Full_Adder FA_62(s62, c62, in62_1, in62_2, pp13[6]);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {c26};
    assign in63_2 = {c27};
    Full_Adder FA_63(s63, c63, in63_1, in63_2, c25);
    wire[0:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp9[11]};
    assign in64_2 = {pp10[10]};
    Full_Adder FA_64(s64, c64, in64_1, in64_2, pp8[12]);
    wire[0:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp12[8]};
    assign in65_2 = {pp13[7]};
    Full_Adder FA_65(s65, c65, in65_1, in65_2, pp11[9]);
    wire[0:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp15[5]};
    assign in66_2 = {c28};
    Full_Adder FA_66(s66, c66, in66_1, in66_2, pp14[6]);
    wire[0:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp7[14]};
    assign in67_2 = {pp8[13]};
    Full_Adder FA_67(s67, c67, in67_1, in67_2, pp6[15]);
    wire[0:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp10[11]};
    assign in68_2 = {pp11[10]};
    Full_Adder FA_68(s68, c68, in68_1, in68_2, pp9[12]);
    wire[0:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp13[8]};
    assign in69_2 = {pp14[7]};
    Full_Adder FA_69(s69, c69, in69_1, in69_2, pp12[9]);
    wire[0:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp8[14]};
    assign in70_2 = {pp9[13]};
    Full_Adder FA_70(s70, c70, in70_1, in70_2, pp7[15]);
    wire[0:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp11[11]};
    assign in71_2 = {pp12[10]};
    Full_Adder FA_71(s71, c71, in71_1, in71_2, pp10[12]);
    wire[0:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp9[14]};
    assign in72_2 = {pp10[13]};
    Full_Adder FA_72(s72, c72, in72_1, in72_2, pp8[15]);

    /*Stage 3*/
    wire[0:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp0[6]};
    assign in73_2 = {pp1[5]};
    Half_Adder HA_73(s73, c73, in73_1, in73_2);
    wire[0:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp1[6]};
    assign in74_2 = {pp2[5]};
    Full_Adder FA_74(s74, c74, in74_1, in74_2, pp0[7]);
    wire[0:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp3[4]};
    assign in75_2 = {pp4[3]};
    Half_Adder HA_75(s75, c75, in75_1, in75_2);
    wire[0:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp3[5]};
    assign in76_2 = {pp4[4]};
    Full_Adder FA_76(s76, c76, in76_1, in76_2, pp2[6]);
    wire[0:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp6[2]};
    assign in77_2 = {pp7[1]};
    Full_Adder FA_77(s77, c77, in77_1, in77_2, pp5[3]);
    wire[0:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp6[3]};
    assign in78_2 = {pp7[2]};
    Full_Adder FA_78(s78, c78, in78_1, in78_2, pp5[4]);
    wire[0:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp9[0]};
    assign in79_2 = {c31};
    Full_Adder FA_79(s79, c79, in79_1, in79_2, pp8[1]);
    wire[0:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp9[1]};
    assign in80_2 = {pp10[0]};
    Full_Adder FA_80(s80, c80, in80_1, in80_2, pp8[2]);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {c33};
    assign in81_2 = {s34[0]};
    Full_Adder FA_81(s81, c81, in81_1, in81_2, c32);
    wire[0:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {s1[0]};
    assign in82_2 = {c34};
    Full_Adder FA_82(s82, c82, in82_1, in82_2, pp11[0]);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {c36};
    assign in83_2 = {s37[0]};
    Full_Adder FA_83(s83, c83, in83_1, in83_2, c35);
    wire[0:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {s3[0]};
    assign in84_2 = {c37};
    Full_Adder FA_84(s84, c84, in84_1, in84_2, s2[0]);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {c39};
    assign in85_2 = {s40[0]};
    Full_Adder FA_85(s85, c85, in85_1, in85_2, c38);
    wire[0:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {s6[0]};
    assign in86_2 = {c40};
    Full_Adder FA_86(s86, c86, in86_1, in86_2, s5[0]);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {c42};
    assign in87_2 = {s43[0]};
    Full_Adder FA_87(s87, c87, in87_1, in87_2, c41);
    wire[0:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {s10[0]};
    assign in88_2 = {c43};
    Full_Adder FA_88(s88, c88, in88_1, in88_2, s9[0]);
    wire[0:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {c45};
    assign in89_2 = {s46[0]};
    Full_Adder FA_89(s89, c89, in89_1, in89_2, c44);
    wire[0:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {s15[0]};
    assign in90_2 = {c46};
    Full_Adder FA_90(s90, c90, in90_1, in90_2, s14[0]);
    wire[0:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {c48};
    assign in91_2 = {s49[0]};
    Full_Adder FA_91(s91, c91, in91_1, in91_2, c47);
    wire[0:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {s20[0]};
    assign in92_2 = {c49};
    Full_Adder FA_92(s92, c92, in92_1, in92_2, s19[0]);
    wire[0:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {c51};
    assign in93_2 = {s52[0]};
    Full_Adder FA_93(s93, c93, in93_1, in93_2, c50);
    wire[0:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {s24[0]};
    assign in94_2 = {c52};
    Full_Adder FA_94(s94, c94, in94_1, in94_2, s23[0]);
    wire[0:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {c54};
    assign in95_2 = {s55[0]};
    Full_Adder FA_95(s95, c95, in95_1, in95_2, c53);
    wire[0:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {s27[0]};
    assign in96_2 = {c55};
    Full_Adder FA_96(s96, c96, in96_1, in96_2, s26[0]);
    wire[0:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {c57};
    assign in97_2 = {s58[0]};
    Full_Adder FA_97(s97, c97, in97_1, in97_2, c56);
    wire[0:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {s29[0]};
    assign in98_2 = {c58};
    Full_Adder FA_98(s98, c98, in98_1, in98_2, s28[0]);
    wire[0:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {c60};
    assign in99_2 = {s61[0]};
    Full_Adder FA_99(s99, c99, in99_1, in99_2, c59);
    wire[0:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {s30[0]};
    assign in100_2 = {c61};
    Full_Adder FA_100(s100, c100, in100_1, in100_2, c29);
    wire[0:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {c63};
    assign in101_2 = {s64[0]};
    Full_Adder FA_101(s101, c101, in101_1, in101_2, c62);
    wire[0:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {c30};
    assign in102_2 = {c64};
    Full_Adder FA_102(s102, c102, in102_1, in102_2, pp15[6]);
    wire[0:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {c66};
    assign in103_2 = {s67[0]};
    Full_Adder FA_103(s103, c103, in103_1, in103_2, c65);
    wire[0:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp14[8]};
    assign in104_2 = {pp15[7]};
    Full_Adder FA_104(s104, c104, in104_1, in104_2, pp13[9]);
    wire[0:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {c68};
    assign in105_2 = {c69};
    Full_Adder FA_105(s105, c105, in105_1, in105_2, c67);
    wire[0:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp12[11]};
    assign in106_2 = {pp13[10]};
    Full_Adder FA_106(s106, c106, in106_1, in106_2, pp11[12]);
    wire[0:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp15[8]};
    assign in107_2 = {c70};
    Full_Adder FA_107(s107, c107, in107_1, in107_2, pp14[9]);
    wire[0:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp10[14]};
    assign in108_2 = {pp11[13]};
    Full_Adder FA_108(s108, c108, in108_1, in108_2, pp9[15]);
    wire[0:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp13[11]};
    assign in109_2 = {pp14[10]};
    Full_Adder FA_109(s109, c109, in109_1, in109_2, pp12[12]);
    wire[0:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp11[14]};
    assign in110_2 = {pp12[13]};
    Full_Adder FA_110(s110, c110, in110_1, in110_2, pp10[15]);

    /*Stage 4*/
    wire[0:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp0[4]};
    assign in111_2 = {pp1[3]};
    Half_Adder HA_111(s111, c111, in111_1, in111_2);
    wire[0:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp1[4]};
    assign in112_2 = {pp2[3]};
    Full_Adder FA_112(s112, c112, in112_1, in112_2, pp0[5]);
    wire[0:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp3[2]};
    assign in113_2 = {pp4[1]};
    Half_Adder HA_113(s113, c113, in113_1, in113_2);
    wire[0:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp3[3]};
    assign in114_2 = {pp4[2]};
    Full_Adder FA_114(s114, c114, in114_1, in114_2, pp2[4]);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp6[0]};
    assign in115_2 = {s73[0]};
    Full_Adder FA_115(s115, c115, in115_1, in115_2, pp5[1]);
    wire[0:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp6[1]};
    assign in116_2 = {pp7[0]};
    Full_Adder FA_116(s116, c116, in116_1, in116_2, pp5[2]);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {s74[0]};
    assign in117_2 = {s75[0]};
    Full_Adder FA_117(s117, c117, in117_1, in117_2, c73);
    wire[0:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {s31[0]};
    assign in118_2 = {c74};
    Full_Adder FA_118(s118, c118, in118_1, in118_2, pp8[0]);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {s76[0]};
    assign in119_2 = {s77[0]};
    Full_Adder FA_119(s119, c119, in119_1, in119_2, c75);
    wire[0:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {s33[0]};
    assign in120_2 = {c76};
    Full_Adder FA_120(s120, c120, in120_1, in120_2, s32[0]);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {s78[0]};
    assign in121_2 = {s79[0]};
    Full_Adder FA_121(s121, c121, in121_1, in121_2, c77);
    wire[0:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {s36[0]};
    assign in122_2 = {c78};
    Full_Adder FA_122(s122, c122, in122_1, in122_2, s35[0]);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {s80[0]};
    assign in123_2 = {s81[0]};
    Full_Adder FA_123(s123, c123, in123_1, in123_2, c79);
    wire[0:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {s39[0]};
    assign in124_2 = {c80};
    Full_Adder FA_124(s124, c124, in124_1, in124_2, s38[0]);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {s82[0]};
    assign in125_2 = {s83[0]};
    Full_Adder FA_125(s125, c125, in125_1, in125_2, c81);
    wire[0:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {s42[0]};
    assign in126_2 = {c82};
    Full_Adder FA_126(s126, c126, in126_1, in126_2, s41[0]);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {s84[0]};
    assign in127_2 = {s85[0]};
    Full_Adder FA_127(s127, c127, in127_1, in127_2, c83);
    wire[0:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {s45[0]};
    assign in128_2 = {c84};
    Full_Adder FA_128(s128, c128, in128_1, in128_2, s44[0]);
    wire[0:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {s86[0]};
    assign in129_2 = {s87[0]};
    Full_Adder FA_129(s129, c129, in129_1, in129_2, c85);
    wire[0:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {s48[0]};
    assign in130_2 = {c86};
    Full_Adder FA_130(s130, c130, in130_1, in130_2, s47[0]);
    wire[0:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {s88[0]};
    assign in131_2 = {s89[0]};
    Full_Adder FA_131(s131, c131, in131_1, in131_2, c87);
    wire[0:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {s51[0]};
    assign in132_2 = {c88};
    Full_Adder FA_132(s132, c132, in132_1, in132_2, s50[0]);
    wire[0:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {s90[0]};
    assign in133_2 = {s91[0]};
    Full_Adder FA_133(s133, c133, in133_1, in133_2, c89);
    wire[0:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {s54[0]};
    assign in134_2 = {c90};
    Full_Adder FA_134(s134, c134, in134_1, in134_2, s53[0]);
    wire[0:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {s92[0]};
    assign in135_2 = {s93[0]};
    Full_Adder FA_135(s135, c135, in135_1, in135_2, c91);
    wire[0:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {s57[0]};
    assign in136_2 = {c92};
    Full_Adder FA_136(s136, c136, in136_1, in136_2, s56[0]);
    wire[0:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {s94[0]};
    assign in137_2 = {s95[0]};
    Full_Adder FA_137(s137, c137, in137_1, in137_2, c93);
    wire[0:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {s60[0]};
    assign in138_2 = {c94};
    Full_Adder FA_138(s138, c138, in138_1, in138_2, s59[0]);
    wire[0:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {s96[0]};
    assign in139_2 = {s97[0]};
    Full_Adder FA_139(s139, c139, in139_1, in139_2, c95);
    wire[0:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {s63[0]};
    assign in140_2 = {c96};
    Full_Adder FA_140(s140, c140, in140_1, in140_2, s62[0]);
    wire[0:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {s98[0]};
    assign in141_2 = {s99[0]};
    Full_Adder FA_141(s141, c141, in141_1, in141_2, c97);
    wire[0:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {s66[0]};
    assign in142_2 = {c98};
    Full_Adder FA_142(s142, c142, in142_1, in142_2, s65[0]);
    wire[0:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {s100[0]};
    assign in143_2 = {s101[0]};
    Full_Adder FA_143(s143, c143, in143_1, in143_2, c99);
    wire[0:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {s69[0]};
    assign in144_2 = {c100};
    Full_Adder FA_144(s144, c144, in144_1, in144_2, s68[0]);
    wire[0:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {s102[0]};
    assign in145_2 = {s103[0]};
    Full_Adder FA_145(s145, c145, in145_1, in145_2, c101);
    wire[0:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {s71[0]};
    assign in146_2 = {c102};
    Full_Adder FA_146(s146, c146, in146_1, in146_2, s70[0]);
    wire[0:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {s104[0]};
    assign in147_2 = {s105[0]};
    Full_Adder FA_147(s147, c147, in147_1, in147_2, c103);
    wire[0:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {s72[0]};
    assign in148_2 = {c104};
    Full_Adder FA_148(s148, c148, in148_1, in148_2, c71);
    wire[0:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {s106[0]};
    assign in149_2 = {s107[0]};
    Full_Adder FA_149(s149, c149, in149_1, in149_2, c105);
    wire[0:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {c72};
    assign in150_2 = {c106};
    Full_Adder FA_150(s150, c150, in150_1, in150_2, pp15[9]);
    wire[0:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {s108[0]};
    assign in151_2 = {s109[0]};
    Full_Adder FA_151(s151, c151, in151_1, in151_2, c107);
    wire[0:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp14[11]};
    assign in152_2 = {pp15[10]};
    Full_Adder FA_152(s152, c152, in152_1, in152_2, pp13[12]);
    wire[0:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {c109};
    assign in153_2 = {s110[0]};
    Full_Adder FA_153(s153, c153, in153_1, in153_2, c108);
    wire[0:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp12[14]};
    assign in154_2 = {pp13[13]};
    Full_Adder FA_154(s154, c154, in154_1, in154_2, pp11[15]);
    wire[0:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp15[11]};
    assign in155_2 = {c110};
    Full_Adder FA_155(s155, c155, in155_1, in155_2, pp14[12]);
    wire[0:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp13[14]};
    assign in156_2 = {pp14[13]};
    Full_Adder FA_156(s156, c156, in156_1, in156_2, pp12[15]);

    /*Stage 5*/
    wire[0:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp0[3]};
    assign in157_2 = {pp1[2]};
    Half_Adder HA_157(s157, c157, in157_1, in157_2);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp3[1]};
    assign in158_2 = {pp4[0]};
    Full_Adder FA_158(s158, c158, in158_1, in158_2, pp2[2]);
    wire[0:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {c111};
    assign in159_2 = {s112[0]};
    Full_Adder FA_159(s159, c159, in159_1, in159_2, pp5[0]);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {c113};
    assign in160_2 = {s114[0]};
    Full_Adder FA_160(s160, c160, in160_1, in160_2, c112);
    wire[0:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {c115};
    assign in161_2 = {s116[0]};
    Full_Adder FA_161(s161, c161, in161_1, in161_2, c114);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {c117};
    assign in162_2 = {s118[0]};
    Full_Adder FA_162(s162, c162, in162_1, in162_2, c116);
    wire[0:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {c119};
    assign in163_2 = {s120[0]};
    Full_Adder FA_163(s163, c163, in163_1, in163_2, c118);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {c121};
    assign in164_2 = {s122[0]};
    Full_Adder FA_164(s164, c164, in164_1, in164_2, c120);
    wire[0:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {c123};
    assign in165_2 = {s124[0]};
    Full_Adder FA_165(s165, c165, in165_1, in165_2, c122);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {c125};
    assign in166_2 = {s126[0]};
    Full_Adder FA_166(s166, c166, in166_1, in166_2, c124);
    wire[0:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {c127};
    assign in167_2 = {s128[0]};
    Full_Adder FA_167(s167, c167, in167_1, in167_2, c126);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {c129};
    assign in168_2 = {s130[0]};
    Full_Adder FA_168(s168, c168, in168_1, in168_2, c128);
    wire[0:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {c131};
    assign in169_2 = {s132[0]};
    Full_Adder FA_169(s169, c169, in169_1, in169_2, c130);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {c133};
    assign in170_2 = {s134[0]};
    Full_Adder FA_170(s170, c170, in170_1, in170_2, c132);
    wire[0:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {c135};
    assign in171_2 = {s136[0]};
    Full_Adder FA_171(s171, c171, in171_1, in171_2, c134);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {c137};
    assign in172_2 = {s138[0]};
    Full_Adder FA_172(s172, c172, in172_1, in172_2, c136);
    wire[0:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {c139};
    assign in173_2 = {s140[0]};
    Full_Adder FA_173(s173, c173, in173_1, in173_2, c138);
    wire[0:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {c141};
    assign in174_2 = {s142[0]};
    Full_Adder FA_174(s174, c174, in174_1, in174_2, c140);
    wire[0:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {c143};
    assign in175_2 = {s144[0]};
    Full_Adder FA_175(s175, c175, in175_1, in175_2, c142);
    wire[0:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {c145};
    assign in176_2 = {s146[0]};
    Full_Adder FA_176(s176, c176, in176_1, in176_2, c144);
    wire[0:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {c147};
    assign in177_2 = {s148[0]};
    Full_Adder FA_177(s177, c177, in177_1, in177_2, c146);
    wire[0:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {c149};
    assign in178_2 = {s150[0]};
    Full_Adder FA_178(s178, c178, in178_1, in178_2, c148);
    wire[0:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {c151};
    assign in179_2 = {s152[0]};
    Full_Adder FA_179(s179, c179, in179_1, in179_2, c150);
    wire[0:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {c153};
    assign in180_2 = {s154[0]};
    Full_Adder FA_180(s180, c180, in180_1, in180_2, c152);
    wire[0:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {c154};
    assign in181_2 = {c155};
    Full_Adder FA_181(s181, c181, in181_1, in181_2, pp15[12]);
    wire[0:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp14[14]};
    assign in182_2 = {pp15[13]};
    Full_Adder FA_182(s182, c182, in182_1, in182_2, pp13[15]);

    /*Stage 6*/
    wire[0:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp0[2]};
    assign in183_2 = {pp1[1]};
    Half_Adder HA_183(s183, c183, in183_1, in183_2);
    wire[0:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp3[0]};
    assign in184_2 = {s157[0]};
    Full_Adder FA_184(s184, c184, in184_1, in184_2, pp2[1]);
    wire[0:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {c157};
    assign in185_2 = {s158[0]};
    Full_Adder FA_185(s185, c185, in185_1, in185_2, s111[0]);
    wire[0:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {c158};
    assign in186_2 = {s159[0]};
    Full_Adder FA_186(s186, c186, in186_1, in186_2, s113[0]);
    wire[0:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {c159};
    assign in187_2 = {s160[0]};
    Full_Adder FA_187(s187, c187, in187_1, in187_2, s115[0]);
    wire[0:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {c160};
    assign in188_2 = {s161[0]};
    Full_Adder FA_188(s188, c188, in188_1, in188_2, s117[0]);
    wire[0:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {c161};
    assign in189_2 = {s162[0]};
    Full_Adder FA_189(s189, c189, in189_1, in189_2, s119[0]);
    wire[0:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {c162};
    assign in190_2 = {s163[0]};
    Full_Adder FA_190(s190, c190, in190_1, in190_2, s121[0]);
    wire[0:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {c163};
    assign in191_2 = {s164[0]};
    Full_Adder FA_191(s191, c191, in191_1, in191_2, s123[0]);
    wire[0:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {c164};
    assign in192_2 = {s165[0]};
    Full_Adder FA_192(s192, c192, in192_1, in192_2, s125[0]);
    wire[0:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {c165};
    assign in193_2 = {s166[0]};
    Full_Adder FA_193(s193, c193, in193_1, in193_2, s127[0]);
    wire[0:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {c166};
    assign in194_2 = {s167[0]};
    Full_Adder FA_194(s194, c194, in194_1, in194_2, s129[0]);
    wire[0:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {c167};
    assign in195_2 = {s168[0]};
    Full_Adder FA_195(s195, c195, in195_1, in195_2, s131[0]);
    wire[0:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {c168};
    assign in196_2 = {s169[0]};
    Full_Adder FA_196(s196, c196, in196_1, in196_2, s133[0]);
    wire[0:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {c169};
    assign in197_2 = {s170[0]};
    Full_Adder FA_197(s197, c197, in197_1, in197_2, s135[0]);
    wire[0:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {c170};
    assign in198_2 = {s171[0]};
    Full_Adder FA_198(s198, c198, in198_1, in198_2, s137[0]);
    wire[0:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {c171};
    assign in199_2 = {s172[0]};
    Full_Adder FA_199(s199, c199, in199_1, in199_2, s139[0]);
    wire[0:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {c172};
    assign in200_2 = {s173[0]};
    Full_Adder FA_200(s200, c200, in200_1, in200_2, s141[0]);
    wire[0:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {c173};
    assign in201_2 = {s174[0]};
    Full_Adder FA_201(s201, c201, in201_1, in201_2, s143[0]);
    wire[0:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {c174};
    assign in202_2 = {s175[0]};
    Full_Adder FA_202(s202, c202, in202_1, in202_2, s145[0]);
    wire[0:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {c175};
    assign in203_2 = {s176[0]};
    Full_Adder FA_203(s203, c203, in203_1, in203_2, s147[0]);
    wire[0:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {c176};
    assign in204_2 = {s177[0]};
    Full_Adder FA_204(s204, c204, in204_1, in204_2, s149[0]);
    wire[0:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {c177};
    assign in205_2 = {s178[0]};
    Full_Adder FA_205(s205, c205, in205_1, in205_2, s151[0]);
    wire[0:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {c178};
    assign in206_2 = {s179[0]};
    Full_Adder FA_206(s206, c206, in206_1, in206_2, s153[0]);
    wire[0:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {c179};
    assign in207_2 = {s180[0]};
    Full_Adder FA_207(s207, c207, in207_1, in207_2, s155[0]);
    wire[0:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {c180};
    assign in208_2 = {s181[0]};
    Full_Adder FA_208(s208, c208, in208_1, in208_2, s156[0]);
    wire[0:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {c181};
    assign in209_2 = {s182[0]};
    Full_Adder FA_209(s209, c209, in209_1, in209_2, c156);
    wire[0:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {pp15[14]};
    assign in210_2 = {c182};
    Full_Adder FA_210(s210, c210, in210_1, in210_2, pp14[15]);


    /*Final Stage 6*/
    wire[29:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],c183,c184,c185,c186,c187,c188,c189,c190,c191,c192,c193,c194,c195,c196,c197,c198,c199,c200,c201,c202,c203,c204,c205,c206,c207,c208,c209,pp15[15]};
    assign in_2 = {pp1[0],s183[0],s184[0],s185[0],s186[0],s187[0],s188[0],s189[0],s190[0],s191[0],s192[0],s193[0],s194[0],s195[0],s196[0],s197[0],s198[0],s199[0],s200[0],s201[0],s202[0],s203[0],s204[0],s205[0],s206[0],s207[0],s208[0],s209[0],s210[0],c210};
    CLA_30(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = c;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule


module CLA_30(output [29:0] sum, output cout, input [29:0] in1, input [29:0] in2);

    wire[29:0] G;
    wire[29:0] C;
    wire[29:0] P;

    assign G[0] = in1[29] & in2[29];
    assign P[0] = in1[29] ^ in2[29];
    assign G[1] = in1[28] & in2[28];
    assign P[1] = in1[28] ^ in2[28];
    assign G[2] = in1[27] & in2[27];
    assign P[2] = in1[27] ^ in2[27];
    assign G[3] = in1[26] & in2[26];
    assign P[3] = in1[26] ^ in2[26];
    assign G[4] = in1[25] & in2[25];
    assign P[4] = in1[25] ^ in2[25];
    assign G[5] = in1[24] & in2[24];
    assign P[5] = in1[24] ^ in2[24];
    assign G[6] = in1[23] & in2[23];
    assign P[6] = in1[23] ^ in2[23];
    assign G[7] = in1[22] & in2[22];
    assign P[7] = in1[22] ^ in2[22];
    assign G[8] = in1[21] & in2[21];
    assign P[8] = in1[21] ^ in2[21];
    assign G[9] = in1[20] & in2[20];
    assign P[9] = in1[20] ^ in2[20];
    assign G[10] = in1[19] & in2[19];
    assign P[10] = in1[19] ^ in2[19];
    assign G[11] = in1[18] & in2[18];
    assign P[11] = in1[18] ^ in2[18];
    assign G[12] = in1[17] & in2[17];
    assign P[12] = in1[17] ^ in2[17];
    assign G[13] = in1[16] & in2[16];
    assign P[13] = in1[16] ^ in2[16];
    assign G[14] = in1[15] & in2[15];
    assign P[14] = in1[15] ^ in2[15];
    assign G[15] = in1[14] & in2[14];
    assign P[15] = in1[14] ^ in2[14];
    assign G[16] = in1[13] & in2[13];
    assign P[16] = in1[13] ^ in2[13];
    assign G[17] = in1[12] & in2[12];
    assign P[17] = in1[12] ^ in2[12];
    assign G[18] = in1[11] & in2[11];
    assign P[18] = in1[11] ^ in2[11];
    assign G[19] = in1[10] & in2[10];
    assign P[19] = in1[10] ^ in2[10];
    assign G[20] = in1[9] & in2[9];
    assign P[20] = in1[9] ^ in2[9];
    assign G[21] = in1[8] & in2[8];
    assign P[21] = in1[8] ^ in2[8];
    assign G[22] = in1[7] & in2[7];
    assign P[22] = in1[7] ^ in2[7];
    assign G[23] = in1[6] & in2[6];
    assign P[23] = in1[6] ^ in2[6];
    assign G[24] = in1[5] & in2[5];
    assign P[24] = in1[5] ^ in2[5];
    assign G[25] = in1[4] & in2[4];
    assign P[25] = in1[4] ^ in2[4];
    assign G[26] = in1[3] & in2[3];
    assign P[26] = in1[3] ^ in2[3];
    assign G[27] = in1[2] & in2[2];
    assign P[27] = in1[2] ^ in2[2];
    assign G[28] = in1[1] & in2[1];
    assign P[28] = in1[1] ^ in2[1];
    assign G[29] = in1[0] & in2[0];
    assign P[29] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign cout = G[29] | (P[29] & C[29]);
    assign sum = P ^ C;
endmodule

