module multiplier_64bits_version14(product, A, B);

    output [127:0] product;
    input [63:0] A, B;

    wire [63:0] pp0;
    wire [63:0] pp1;
    wire [63:0] pp2;
    wire [63:0] pp3;
    wire [63:0] pp4;
    wire [63:0] pp5;
    wire [63:0] pp6;
    wire [63:0] pp7;
    wire [63:0] pp8;
    wire [63:0] pp9;
    wire [63:0] pp10;
    wire [63:0] pp11;
    wire [63:0] pp12;
    wire [63:0] pp13;
    wire [63:0] pp14;
    wire [63:0] pp15;
    wire [63:0] pp16;
    wire [63:0] pp17;
    wire [63:0] pp18;
    wire [63:0] pp19;
    wire [63:0] pp20;
    wire [63:0] pp21;
    wire [63:0] pp22;
    wire [63:0] pp23;
    wire [63:0] pp24;
    wire [63:0] pp25;
    wire [63:0] pp26;
    wire [63:0] pp27;
    wire [63:0] pp28;
    wire [63:0] pp29;
    wire [63:0] pp30;
    wire [63:0] pp31;
    wire [63:0] pp32;
    wire [63:0] pp33;
    wire [63:0] pp34;
    wire [63:0] pp35;
    wire [63:0] pp36;
    wire [63:0] pp37;
    wire [63:0] pp38;
    wire [63:0] pp39;
    wire [63:0] pp40;
    wire [63:0] pp41;
    wire [63:0] pp42;
    wire [63:0] pp43;
    wire [63:0] pp44;
    wire [63:0] pp45;
    wire [63:0] pp46;
    wire [63:0] pp47;
    wire [63:0] pp48;
    wire [63:0] pp49;
    wire [63:0] pp50;
    wire [63:0] pp51;
    wire [63:0] pp52;
    wire [63:0] pp53;
    wire [63:0] pp54;
    wire [63:0] pp55;
    wire [63:0] pp56;
    wire [63:0] pp57;
    wire [63:0] pp58;
    wire [63:0] pp59;
    wire [63:0] pp60;
    wire [63:0] pp61;
    wire [63:0] pp62;
    wire [63:0] pp63;


    assign pp0 = A[0] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[0:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[43]};
    assign in1_2 = {pp1[42]};
    Half_Adder HA_1(s1, c1, in1_1, in1_2);
    wire[0:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp1[43]};
    assign in2_2 = {pp2[42]};
    Full_Adder FA_2(s2, c2, in2_1, in2_2, pp0[44]);
    wire[0:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp3[41]};
    assign in3_2 = {pp4[40]};
    Half_Adder HA_3(s3, c3, in3_1, in3_2);
    wire[0:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp1[44]};
    assign in4_2 = {pp2[43]};
    Full_Adder FA_4(s4, c4, in4_1, in4_2, pp0[45]);
    wire[0:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp4[41]};
    assign in5_2 = {pp5[40]};
    Full_Adder FA_5(s5, c5, in5_1, in5_2, pp3[42]);
    wire[0:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp6[39]};
    assign in6_2 = {pp7[38]};
    Half_Adder HA_6(s6, c6, in6_1, in6_2);
    wire[0:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp1[45]};
    assign in7_2 = {pp2[44]};
    Full_Adder FA_7(s7, c7, in7_1, in7_2, pp0[46]);
    wire[0:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp4[42]};
    assign in8_2 = {pp5[41]};
    Full_Adder FA_8(s8, c8, in8_1, in8_2, pp3[43]);
    wire[0:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp7[39]};
    assign in9_2 = {pp8[38]};
    Full_Adder FA_9(s9, c9, in9_1, in9_2, pp6[40]);
    wire[0:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp9[37]};
    assign in10_2 = {pp10[36]};
    Half_Adder HA_10(s10, c10, in10_1, in10_2);
    wire[0:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp1[46]};
    assign in11_2 = {pp2[45]};
    Full_Adder FA_11(s11, c11, in11_1, in11_2, pp0[47]);
    wire[0:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp4[43]};
    assign in12_2 = {pp5[42]};
    Full_Adder FA_12(s12, c12, in12_1, in12_2, pp3[44]);
    wire[0:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp7[40]};
    assign in13_2 = {pp8[39]};
    Full_Adder FA_13(s13, c13, in13_1, in13_2, pp6[41]);
    wire[0:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp10[37]};
    assign in14_2 = {pp11[36]};
    Full_Adder FA_14(s14, c14, in14_1, in14_2, pp9[38]);
    wire[0:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp12[35]};
    assign in15_2 = {pp13[34]};
    Half_Adder HA_15(s15, c15, in15_1, in15_2);
    wire[0:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp1[47]};
    assign in16_2 = {pp2[46]};
    Full_Adder FA_16(s16, c16, in16_1, in16_2, pp0[48]);
    wire[0:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp4[44]};
    assign in17_2 = {pp5[43]};
    Full_Adder FA_17(s17, c17, in17_1, in17_2, pp3[45]);
    wire[0:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp7[41]};
    assign in18_2 = {pp8[40]};
    Full_Adder FA_18(s18, c18, in18_1, in18_2, pp6[42]);
    wire[0:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp10[38]};
    assign in19_2 = {pp11[37]};
    Full_Adder FA_19(s19, c19, in19_1, in19_2, pp9[39]);
    wire[0:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp13[35]};
    assign in20_2 = {pp14[34]};
    Full_Adder FA_20(s20, c20, in20_1, in20_2, pp12[36]);
    wire[0:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp15[33]};
    assign in21_2 = {pp16[32]};
    Half_Adder HA_21(s21, c21, in21_1, in21_2);
    wire[0:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp1[48]};
    assign in22_2 = {pp2[47]};
    Full_Adder FA_22(s22, c22, in22_1, in22_2, pp0[49]);
    wire[0:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp4[45]};
    assign in23_2 = {pp5[44]};
    Full_Adder FA_23(s23, c23, in23_1, in23_2, pp3[46]);
    wire[0:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp7[42]};
    assign in24_2 = {pp8[41]};
    Full_Adder FA_24(s24, c24, in24_1, in24_2, pp6[43]);
    wire[0:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp10[39]};
    assign in25_2 = {pp11[38]};
    Full_Adder FA_25(s25, c25, in25_1, in25_2, pp9[40]);
    wire[0:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp13[36]};
    assign in26_2 = {pp14[35]};
    Full_Adder FA_26(s26, c26, in26_1, in26_2, pp12[37]);
    wire[0:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp16[33]};
    assign in27_2 = {pp17[32]};
    Full_Adder FA_27(s27, c27, in27_1, in27_2, pp15[34]);
    wire[0:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp18[31]};
    assign in28_2 = {pp19[30]};
    Half_Adder HA_28(s28, c28, in28_1, in28_2);
    wire[0:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp1[49]};
    assign in29_2 = {pp2[48]};
    Full_Adder FA_29(s29, c29, in29_1, in29_2, pp0[50]);
    wire[0:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp4[46]};
    assign in30_2 = {pp5[45]};
    Full_Adder FA_30(s30, c30, in30_1, in30_2, pp3[47]);
    wire[0:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp7[43]};
    assign in31_2 = {pp8[42]};
    Full_Adder FA_31(s31, c31, in31_1, in31_2, pp6[44]);
    wire[0:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp10[40]};
    assign in32_2 = {pp11[39]};
    Full_Adder FA_32(s32, c32, in32_1, in32_2, pp9[41]);
    wire[0:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp13[37]};
    assign in33_2 = {pp14[36]};
    Full_Adder FA_33(s33, c33, in33_1, in33_2, pp12[38]);
    wire[0:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp16[34]};
    assign in34_2 = {pp17[33]};
    Full_Adder FA_34(s34, c34, in34_1, in34_2, pp15[35]);
    wire[0:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp19[31]};
    assign in35_2 = {pp20[30]};
    Full_Adder FA_35(s35, c35, in35_1, in35_2, pp18[32]);
    wire[0:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp21[29]};
    assign in36_2 = {pp22[28]};
    Half_Adder HA_36(s36, c36, in36_1, in36_2);
    wire[0:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp1[50]};
    assign in37_2 = {pp2[49]};
    Full_Adder FA_37(s37, c37, in37_1, in37_2, pp0[51]);
    wire[0:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp4[47]};
    assign in38_2 = {pp5[46]};
    Full_Adder FA_38(s38, c38, in38_1, in38_2, pp3[48]);
    wire[0:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp7[44]};
    assign in39_2 = {pp8[43]};
    Full_Adder FA_39(s39, c39, in39_1, in39_2, pp6[45]);
    wire[0:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp10[41]};
    assign in40_2 = {pp11[40]};
    Full_Adder FA_40(s40, c40, in40_1, in40_2, pp9[42]);
    wire[0:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp13[38]};
    assign in41_2 = {pp14[37]};
    Full_Adder FA_41(s41, c41, in41_1, in41_2, pp12[39]);
    wire[0:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp16[35]};
    assign in42_2 = {pp17[34]};
    Full_Adder FA_42(s42, c42, in42_1, in42_2, pp15[36]);
    wire[0:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp19[32]};
    assign in43_2 = {pp20[31]};
    Full_Adder FA_43(s43, c43, in43_1, in43_2, pp18[33]);
    wire[0:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[29]};
    assign in44_2 = {pp23[28]};
    Full_Adder FA_44(s44, c44, in44_1, in44_2, pp21[30]);
    wire[0:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[27]};
    assign in45_2 = {pp25[26]};
    Half_Adder HA_45(s45, c45, in45_1, in45_2);
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp1[51]};
    assign in46_2 = {pp2[50]};
    Full_Adder FA_46(s46, c46, in46_1, in46_2, pp0[52]);
    wire[0:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp4[48]};
    assign in47_2 = {pp5[47]};
    Full_Adder FA_47(s47, c47, in47_1, in47_2, pp3[49]);
    wire[0:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp7[45]};
    assign in48_2 = {pp8[44]};
    Full_Adder FA_48(s48, c48, in48_1, in48_2, pp6[46]);
    wire[0:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp10[42]};
    assign in49_2 = {pp11[41]};
    Full_Adder FA_49(s49, c49, in49_1, in49_2, pp9[43]);
    wire[0:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp13[39]};
    assign in50_2 = {pp14[38]};
    Full_Adder FA_50(s50, c50, in50_1, in50_2, pp12[40]);
    wire[0:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp16[36]};
    assign in51_2 = {pp17[35]};
    Full_Adder FA_51(s51, c51, in51_1, in51_2, pp15[37]);
    wire[0:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp19[33]};
    assign in52_2 = {pp20[32]};
    Full_Adder FA_52(s52, c52, in52_1, in52_2, pp18[34]);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp22[30]};
    assign in53_2 = {pp23[29]};
    Full_Adder FA_53(s53, c53, in53_1, in53_2, pp21[31]);
    wire[0:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp25[27]};
    assign in54_2 = {pp26[26]};
    Full_Adder FA_54(s54, c54, in54_1, in54_2, pp24[28]);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp27[25]};
    assign in55_2 = {pp28[24]};
    Half_Adder HA_55(s55, c55, in55_1, in55_2);
    wire[0:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp1[52]};
    assign in56_2 = {pp2[51]};
    Full_Adder FA_56(s56, c56, in56_1, in56_2, pp0[53]);
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp4[49]};
    assign in57_2 = {pp5[48]};
    Full_Adder FA_57(s57, c57, in57_1, in57_2, pp3[50]);
    wire[0:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp7[46]};
    assign in58_2 = {pp8[45]};
    Full_Adder FA_58(s58, c58, in58_1, in58_2, pp6[47]);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp10[43]};
    assign in59_2 = {pp11[42]};
    Full_Adder FA_59(s59, c59, in59_1, in59_2, pp9[44]);
    wire[0:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp13[40]};
    assign in60_2 = {pp14[39]};
    Full_Adder FA_60(s60, c60, in60_1, in60_2, pp12[41]);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp16[37]};
    assign in61_2 = {pp17[36]};
    Full_Adder FA_61(s61, c61, in61_1, in61_2, pp15[38]);
    wire[0:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp19[34]};
    assign in62_2 = {pp20[33]};
    Full_Adder FA_62(s62, c62, in62_1, in62_2, pp18[35]);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp22[31]};
    assign in63_2 = {pp23[30]};
    Full_Adder FA_63(s63, c63, in63_1, in63_2, pp21[32]);
    wire[0:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp25[28]};
    assign in64_2 = {pp26[27]};
    Full_Adder FA_64(s64, c64, in64_1, in64_2, pp24[29]);
    wire[0:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp28[25]};
    assign in65_2 = {pp29[24]};
    Full_Adder FA_65(s65, c65, in65_1, in65_2, pp27[26]);
    wire[0:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp30[23]};
    assign in66_2 = {pp31[22]};
    Half_Adder HA_66(s66, c66, in66_1, in66_2);
    wire[0:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp1[53]};
    assign in67_2 = {pp2[52]};
    Full_Adder FA_67(s67, c67, in67_1, in67_2, pp0[54]);
    wire[0:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp4[50]};
    assign in68_2 = {pp5[49]};
    Full_Adder FA_68(s68, c68, in68_1, in68_2, pp3[51]);
    wire[0:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp7[47]};
    assign in69_2 = {pp8[46]};
    Full_Adder FA_69(s69, c69, in69_1, in69_2, pp6[48]);
    wire[0:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp10[44]};
    assign in70_2 = {pp11[43]};
    Full_Adder FA_70(s70, c70, in70_1, in70_2, pp9[45]);
    wire[0:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp13[41]};
    assign in71_2 = {pp14[40]};
    Full_Adder FA_71(s71, c71, in71_1, in71_2, pp12[42]);
    wire[0:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp16[38]};
    assign in72_2 = {pp17[37]};
    Full_Adder FA_72(s72, c72, in72_1, in72_2, pp15[39]);
    wire[0:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp19[35]};
    assign in73_2 = {pp20[34]};
    Full_Adder FA_73(s73, c73, in73_1, in73_2, pp18[36]);
    wire[0:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp22[32]};
    assign in74_2 = {pp23[31]};
    Full_Adder FA_74(s74, c74, in74_1, in74_2, pp21[33]);
    wire[0:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp25[29]};
    assign in75_2 = {pp26[28]};
    Full_Adder FA_75(s75, c75, in75_1, in75_2, pp24[30]);
    wire[0:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp28[26]};
    assign in76_2 = {pp29[25]};
    Full_Adder FA_76(s76, c76, in76_1, in76_2, pp27[27]);
    wire[0:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp31[23]};
    assign in77_2 = {pp32[22]};
    Full_Adder FA_77(s77, c77, in77_1, in77_2, pp30[24]);
    wire[0:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp33[21]};
    assign in78_2 = {pp34[20]};
    Half_Adder HA_78(s78, c78, in78_1, in78_2);
    wire[0:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp1[54]};
    assign in79_2 = {pp2[53]};
    Full_Adder FA_79(s79, c79, in79_1, in79_2, pp0[55]);
    wire[0:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp4[51]};
    assign in80_2 = {pp5[50]};
    Full_Adder FA_80(s80, c80, in80_1, in80_2, pp3[52]);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp7[48]};
    assign in81_2 = {pp8[47]};
    Full_Adder FA_81(s81, c81, in81_1, in81_2, pp6[49]);
    wire[0:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp10[45]};
    assign in82_2 = {pp11[44]};
    Full_Adder FA_82(s82, c82, in82_1, in82_2, pp9[46]);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp13[42]};
    assign in83_2 = {pp14[41]};
    Full_Adder FA_83(s83, c83, in83_1, in83_2, pp12[43]);
    wire[0:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp16[39]};
    assign in84_2 = {pp17[38]};
    Full_Adder FA_84(s84, c84, in84_1, in84_2, pp15[40]);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp19[36]};
    assign in85_2 = {pp20[35]};
    Full_Adder FA_85(s85, c85, in85_1, in85_2, pp18[37]);
    wire[0:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp22[33]};
    assign in86_2 = {pp23[32]};
    Full_Adder FA_86(s86, c86, in86_1, in86_2, pp21[34]);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp25[30]};
    assign in87_2 = {pp26[29]};
    Full_Adder FA_87(s87, c87, in87_1, in87_2, pp24[31]);
    wire[0:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp28[27]};
    assign in88_2 = {pp29[26]};
    Full_Adder FA_88(s88, c88, in88_1, in88_2, pp27[28]);
    wire[0:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp31[24]};
    assign in89_2 = {pp32[23]};
    Full_Adder FA_89(s89, c89, in89_1, in89_2, pp30[25]);
    wire[0:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp34[21]};
    assign in90_2 = {pp35[20]};
    Full_Adder FA_90(s90, c90, in90_1, in90_2, pp33[22]);
    wire[0:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp36[19]};
    assign in91_2 = {pp37[18]};
    Half_Adder HA_91(s91, c91, in91_1, in91_2);
    wire[0:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp1[55]};
    assign in92_2 = {pp2[54]};
    Full_Adder FA_92(s92, c92, in92_1, in92_2, pp0[56]);
    wire[0:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp4[52]};
    assign in93_2 = {pp5[51]};
    Full_Adder FA_93(s93, c93, in93_1, in93_2, pp3[53]);
    wire[0:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp7[49]};
    assign in94_2 = {pp8[48]};
    Full_Adder FA_94(s94, c94, in94_1, in94_2, pp6[50]);
    wire[0:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp10[46]};
    assign in95_2 = {pp11[45]};
    Full_Adder FA_95(s95, c95, in95_1, in95_2, pp9[47]);
    wire[0:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp13[43]};
    assign in96_2 = {pp14[42]};
    Full_Adder FA_96(s96, c96, in96_1, in96_2, pp12[44]);
    wire[0:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp16[40]};
    assign in97_2 = {pp17[39]};
    Full_Adder FA_97(s97, c97, in97_1, in97_2, pp15[41]);
    wire[0:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp19[37]};
    assign in98_2 = {pp20[36]};
    Full_Adder FA_98(s98, c98, in98_1, in98_2, pp18[38]);
    wire[0:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp22[34]};
    assign in99_2 = {pp23[33]};
    Full_Adder FA_99(s99, c99, in99_1, in99_2, pp21[35]);
    wire[0:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp25[31]};
    assign in100_2 = {pp26[30]};
    Full_Adder FA_100(s100, c100, in100_1, in100_2, pp24[32]);
    wire[0:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp28[28]};
    assign in101_2 = {pp29[27]};
    Full_Adder FA_101(s101, c101, in101_1, in101_2, pp27[29]);
    wire[0:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp31[25]};
    assign in102_2 = {pp32[24]};
    Full_Adder FA_102(s102, c102, in102_1, in102_2, pp30[26]);
    wire[0:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp34[22]};
    assign in103_2 = {pp35[21]};
    Full_Adder FA_103(s103, c103, in103_1, in103_2, pp33[23]);
    wire[0:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp37[19]};
    assign in104_2 = {pp38[18]};
    Full_Adder FA_104(s104, c104, in104_1, in104_2, pp36[20]);
    wire[0:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp39[17]};
    assign in105_2 = {pp40[16]};
    Half_Adder HA_105(s105, c105, in105_1, in105_2);
    wire[0:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp1[56]};
    assign in106_2 = {pp2[55]};
    Full_Adder FA_106(s106, c106, in106_1, in106_2, pp0[57]);
    wire[0:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp4[53]};
    assign in107_2 = {pp5[52]};
    Full_Adder FA_107(s107, c107, in107_1, in107_2, pp3[54]);
    wire[0:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp7[50]};
    assign in108_2 = {pp8[49]};
    Full_Adder FA_108(s108, c108, in108_1, in108_2, pp6[51]);
    wire[0:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp10[47]};
    assign in109_2 = {pp11[46]};
    Full_Adder FA_109(s109, c109, in109_1, in109_2, pp9[48]);
    wire[0:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp13[44]};
    assign in110_2 = {pp14[43]};
    Full_Adder FA_110(s110, c110, in110_1, in110_2, pp12[45]);
    wire[0:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp16[41]};
    assign in111_2 = {pp17[40]};
    Full_Adder FA_111(s111, c111, in111_1, in111_2, pp15[42]);
    wire[0:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp19[38]};
    assign in112_2 = {pp20[37]};
    Full_Adder FA_112(s112, c112, in112_1, in112_2, pp18[39]);
    wire[0:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp22[35]};
    assign in113_2 = {pp23[34]};
    Full_Adder FA_113(s113, c113, in113_1, in113_2, pp21[36]);
    wire[0:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp25[32]};
    assign in114_2 = {pp26[31]};
    Full_Adder FA_114(s114, c114, in114_1, in114_2, pp24[33]);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp28[29]};
    assign in115_2 = {pp29[28]};
    Full_Adder FA_115(s115, c115, in115_1, in115_2, pp27[30]);
    wire[0:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp31[26]};
    assign in116_2 = {pp32[25]};
    Full_Adder FA_116(s116, c116, in116_1, in116_2, pp30[27]);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp34[23]};
    assign in117_2 = {pp35[22]};
    Full_Adder FA_117(s117, c117, in117_1, in117_2, pp33[24]);
    wire[0:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp37[20]};
    assign in118_2 = {pp38[19]};
    Full_Adder FA_118(s118, c118, in118_1, in118_2, pp36[21]);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp40[17]};
    assign in119_2 = {pp41[16]};
    Full_Adder FA_119(s119, c119, in119_1, in119_2, pp39[18]);
    wire[0:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {pp42[15]};
    assign in120_2 = {pp43[14]};
    Half_Adder HA_120(s120, c120, in120_1, in120_2);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp1[57]};
    assign in121_2 = {pp2[56]};
    Full_Adder FA_121(s121, c121, in121_1, in121_2, pp0[58]);
    wire[0:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp4[54]};
    assign in122_2 = {pp5[53]};
    Full_Adder FA_122(s122, c122, in122_1, in122_2, pp3[55]);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp7[51]};
    assign in123_2 = {pp8[50]};
    Full_Adder FA_123(s123, c123, in123_1, in123_2, pp6[52]);
    wire[0:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp10[48]};
    assign in124_2 = {pp11[47]};
    Full_Adder FA_124(s124, c124, in124_1, in124_2, pp9[49]);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp13[45]};
    assign in125_2 = {pp14[44]};
    Full_Adder FA_125(s125, c125, in125_1, in125_2, pp12[46]);
    wire[0:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp16[42]};
    assign in126_2 = {pp17[41]};
    Full_Adder FA_126(s126, c126, in126_1, in126_2, pp15[43]);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {pp19[39]};
    assign in127_2 = {pp20[38]};
    Full_Adder FA_127(s127, c127, in127_1, in127_2, pp18[40]);
    wire[0:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {pp22[36]};
    assign in128_2 = {pp23[35]};
    Full_Adder FA_128(s128, c128, in128_1, in128_2, pp21[37]);
    wire[0:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp25[33]};
    assign in129_2 = {pp26[32]};
    Full_Adder FA_129(s129, c129, in129_1, in129_2, pp24[34]);
    wire[0:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp28[30]};
    assign in130_2 = {pp29[29]};
    Full_Adder FA_130(s130, c130, in130_1, in130_2, pp27[31]);
    wire[0:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp31[27]};
    assign in131_2 = {pp32[26]};
    Full_Adder FA_131(s131, c131, in131_1, in131_2, pp30[28]);
    wire[0:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp34[24]};
    assign in132_2 = {pp35[23]};
    Full_Adder FA_132(s132, c132, in132_1, in132_2, pp33[25]);
    wire[0:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp37[21]};
    assign in133_2 = {pp38[20]};
    Full_Adder FA_133(s133, c133, in133_1, in133_2, pp36[22]);
    wire[0:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp40[18]};
    assign in134_2 = {pp41[17]};
    Full_Adder FA_134(s134, c134, in134_1, in134_2, pp39[19]);
    wire[0:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp43[15]};
    assign in135_2 = {pp44[14]};
    Full_Adder FA_135(s135, c135, in135_1, in135_2, pp42[16]);
    wire[0:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp45[13]};
    assign in136_2 = {pp46[12]};
    Half_Adder HA_136(s136, c136, in136_1, in136_2);
    wire[0:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp1[58]};
    assign in137_2 = {pp2[57]};
    Full_Adder FA_137(s137, c137, in137_1, in137_2, pp0[59]);
    wire[0:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp4[55]};
    assign in138_2 = {pp5[54]};
    Full_Adder FA_138(s138, c138, in138_1, in138_2, pp3[56]);
    wire[0:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp7[52]};
    assign in139_2 = {pp8[51]};
    Full_Adder FA_139(s139, c139, in139_1, in139_2, pp6[53]);
    wire[0:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp10[49]};
    assign in140_2 = {pp11[48]};
    Full_Adder FA_140(s140, c140, in140_1, in140_2, pp9[50]);
    wire[0:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp13[46]};
    assign in141_2 = {pp14[45]};
    Full_Adder FA_141(s141, c141, in141_1, in141_2, pp12[47]);
    wire[0:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp16[43]};
    assign in142_2 = {pp17[42]};
    Full_Adder FA_142(s142, c142, in142_1, in142_2, pp15[44]);
    wire[0:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp19[40]};
    assign in143_2 = {pp20[39]};
    Full_Adder FA_143(s143, c143, in143_1, in143_2, pp18[41]);
    wire[0:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp22[37]};
    assign in144_2 = {pp23[36]};
    Full_Adder FA_144(s144, c144, in144_1, in144_2, pp21[38]);
    wire[0:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp25[34]};
    assign in145_2 = {pp26[33]};
    Full_Adder FA_145(s145, c145, in145_1, in145_2, pp24[35]);
    wire[0:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp28[31]};
    assign in146_2 = {pp29[30]};
    Full_Adder FA_146(s146, c146, in146_1, in146_2, pp27[32]);
    wire[0:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp31[28]};
    assign in147_2 = {pp32[27]};
    Full_Adder FA_147(s147, c147, in147_1, in147_2, pp30[29]);
    wire[0:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp34[25]};
    assign in148_2 = {pp35[24]};
    Full_Adder FA_148(s148, c148, in148_1, in148_2, pp33[26]);
    wire[0:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp37[22]};
    assign in149_2 = {pp38[21]};
    Full_Adder FA_149(s149, c149, in149_1, in149_2, pp36[23]);
    wire[0:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp40[19]};
    assign in150_2 = {pp41[18]};
    Full_Adder FA_150(s150, c150, in150_1, in150_2, pp39[20]);
    wire[0:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp43[16]};
    assign in151_2 = {pp44[15]};
    Full_Adder FA_151(s151, c151, in151_1, in151_2, pp42[17]);
    wire[0:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp46[13]};
    assign in152_2 = {pp47[12]};
    Full_Adder FA_152(s152, c152, in152_1, in152_2, pp45[14]);
    wire[0:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp48[11]};
    assign in153_2 = {pp49[10]};
    Half_Adder HA_153(s153, c153, in153_1, in153_2);
    wire[0:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp1[59]};
    assign in154_2 = {pp2[58]};
    Full_Adder FA_154(s154, c154, in154_1, in154_2, pp0[60]);
    wire[0:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp4[56]};
    assign in155_2 = {pp5[55]};
    Full_Adder FA_155(s155, c155, in155_1, in155_2, pp3[57]);
    wire[0:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp7[53]};
    assign in156_2 = {pp8[52]};
    Full_Adder FA_156(s156, c156, in156_1, in156_2, pp6[54]);
    wire[0:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp10[50]};
    assign in157_2 = {pp11[49]};
    Full_Adder FA_157(s157, c157, in157_1, in157_2, pp9[51]);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp13[47]};
    assign in158_2 = {pp14[46]};
    Full_Adder FA_158(s158, c158, in158_1, in158_2, pp12[48]);
    wire[0:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp16[44]};
    assign in159_2 = {pp17[43]};
    Full_Adder FA_159(s159, c159, in159_1, in159_2, pp15[45]);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp19[41]};
    assign in160_2 = {pp20[40]};
    Full_Adder FA_160(s160, c160, in160_1, in160_2, pp18[42]);
    wire[0:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp22[38]};
    assign in161_2 = {pp23[37]};
    Full_Adder FA_161(s161, c161, in161_1, in161_2, pp21[39]);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp25[35]};
    assign in162_2 = {pp26[34]};
    Full_Adder FA_162(s162, c162, in162_1, in162_2, pp24[36]);
    wire[0:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp28[32]};
    assign in163_2 = {pp29[31]};
    Full_Adder FA_163(s163, c163, in163_1, in163_2, pp27[33]);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp31[29]};
    assign in164_2 = {pp32[28]};
    Full_Adder FA_164(s164, c164, in164_1, in164_2, pp30[30]);
    wire[0:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {pp34[26]};
    assign in165_2 = {pp35[25]};
    Full_Adder FA_165(s165, c165, in165_1, in165_2, pp33[27]);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {pp37[23]};
    assign in166_2 = {pp38[22]};
    Full_Adder FA_166(s166, c166, in166_1, in166_2, pp36[24]);
    wire[0:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {pp40[20]};
    assign in167_2 = {pp41[19]};
    Full_Adder FA_167(s167, c167, in167_1, in167_2, pp39[21]);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {pp43[17]};
    assign in168_2 = {pp44[16]};
    Full_Adder FA_168(s168, c168, in168_1, in168_2, pp42[18]);
    wire[0:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {pp46[14]};
    assign in169_2 = {pp47[13]};
    Full_Adder FA_169(s169, c169, in169_1, in169_2, pp45[15]);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {pp49[11]};
    assign in170_2 = {pp50[10]};
    Full_Adder FA_170(s170, c170, in170_1, in170_2, pp48[12]);
    wire[0:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {pp51[9]};
    assign in171_2 = {pp52[8]};
    Half_Adder HA_171(s171, c171, in171_1, in171_2);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {pp1[60]};
    assign in172_2 = {pp2[59]};
    Full_Adder FA_172(s172, c172, in172_1, in172_2, pp0[61]);
    wire[0:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {pp4[57]};
    assign in173_2 = {pp5[56]};
    Full_Adder FA_173(s173, c173, in173_1, in173_2, pp3[58]);
    wire[0:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp7[54]};
    assign in174_2 = {pp8[53]};
    Full_Adder FA_174(s174, c174, in174_1, in174_2, pp6[55]);
    wire[0:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp10[51]};
    assign in175_2 = {pp11[50]};
    Full_Adder FA_175(s175, c175, in175_1, in175_2, pp9[52]);
    wire[0:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp13[48]};
    assign in176_2 = {pp14[47]};
    Full_Adder FA_176(s176, c176, in176_1, in176_2, pp12[49]);
    wire[0:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp16[45]};
    assign in177_2 = {pp17[44]};
    Full_Adder FA_177(s177, c177, in177_1, in177_2, pp15[46]);
    wire[0:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {pp19[42]};
    assign in178_2 = {pp20[41]};
    Full_Adder FA_178(s178, c178, in178_1, in178_2, pp18[43]);
    wire[0:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {pp22[39]};
    assign in179_2 = {pp23[38]};
    Full_Adder FA_179(s179, c179, in179_1, in179_2, pp21[40]);
    wire[0:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {pp25[36]};
    assign in180_2 = {pp26[35]};
    Full_Adder FA_180(s180, c180, in180_1, in180_2, pp24[37]);
    wire[0:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp28[33]};
    assign in181_2 = {pp29[32]};
    Full_Adder FA_181(s181, c181, in181_1, in181_2, pp27[34]);
    wire[0:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp31[30]};
    assign in182_2 = {pp32[29]};
    Full_Adder FA_182(s182, c182, in182_1, in182_2, pp30[31]);
    wire[0:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp34[27]};
    assign in183_2 = {pp35[26]};
    Full_Adder FA_183(s183, c183, in183_1, in183_2, pp33[28]);
    wire[0:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp37[24]};
    assign in184_2 = {pp38[23]};
    Full_Adder FA_184(s184, c184, in184_1, in184_2, pp36[25]);
    wire[0:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {pp40[21]};
    assign in185_2 = {pp41[20]};
    Full_Adder FA_185(s185, c185, in185_1, in185_2, pp39[22]);
    wire[0:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {pp43[18]};
    assign in186_2 = {pp44[17]};
    Full_Adder FA_186(s186, c186, in186_1, in186_2, pp42[19]);
    wire[0:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {pp46[15]};
    assign in187_2 = {pp47[14]};
    Full_Adder FA_187(s187, c187, in187_1, in187_2, pp45[16]);
    wire[0:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp49[12]};
    assign in188_2 = {pp50[11]};
    Full_Adder FA_188(s188, c188, in188_1, in188_2, pp48[13]);
    wire[0:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp52[9]};
    assign in189_2 = {pp53[8]};
    Full_Adder FA_189(s189, c189, in189_1, in189_2, pp51[10]);
    wire[0:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {pp54[7]};
    assign in190_2 = {pp55[6]};
    Half_Adder HA_190(s190, c190, in190_1, in190_2);
    wire[0:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {pp1[61]};
    assign in191_2 = {pp2[60]};
    Full_Adder FA_191(s191, c191, in191_1, in191_2, pp0[62]);
    wire[0:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {pp4[58]};
    assign in192_2 = {pp5[57]};
    Full_Adder FA_192(s192, c192, in192_1, in192_2, pp3[59]);
    wire[0:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {pp7[55]};
    assign in193_2 = {pp8[54]};
    Full_Adder FA_193(s193, c193, in193_1, in193_2, pp6[56]);
    wire[0:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {pp10[52]};
    assign in194_2 = {pp11[51]};
    Full_Adder FA_194(s194, c194, in194_1, in194_2, pp9[53]);
    wire[0:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp13[49]};
    assign in195_2 = {pp14[48]};
    Full_Adder FA_195(s195, c195, in195_1, in195_2, pp12[50]);
    wire[0:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp16[46]};
    assign in196_2 = {pp17[45]};
    Full_Adder FA_196(s196, c196, in196_1, in196_2, pp15[47]);
    wire[0:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {pp19[43]};
    assign in197_2 = {pp20[42]};
    Full_Adder FA_197(s197, c197, in197_1, in197_2, pp18[44]);
    wire[0:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {pp22[40]};
    assign in198_2 = {pp23[39]};
    Full_Adder FA_198(s198, c198, in198_1, in198_2, pp21[41]);
    wire[0:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {pp25[37]};
    assign in199_2 = {pp26[36]};
    Full_Adder FA_199(s199, c199, in199_1, in199_2, pp24[38]);
    wire[0:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {pp28[34]};
    assign in200_2 = {pp29[33]};
    Full_Adder FA_200(s200, c200, in200_1, in200_2, pp27[35]);
    wire[0:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {pp31[31]};
    assign in201_2 = {pp32[30]};
    Full_Adder FA_201(s201, c201, in201_1, in201_2, pp30[32]);
    wire[0:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp34[28]};
    assign in202_2 = {pp35[27]};
    Full_Adder FA_202(s202, c202, in202_1, in202_2, pp33[29]);
    wire[0:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {pp37[25]};
    assign in203_2 = {pp38[24]};
    Full_Adder FA_203(s203, c203, in203_1, in203_2, pp36[26]);
    wire[0:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {pp40[22]};
    assign in204_2 = {pp41[21]};
    Full_Adder FA_204(s204, c204, in204_1, in204_2, pp39[23]);
    wire[0:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {pp43[19]};
    assign in205_2 = {pp44[18]};
    Full_Adder FA_205(s205, c205, in205_1, in205_2, pp42[20]);
    wire[0:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {pp46[16]};
    assign in206_2 = {pp47[15]};
    Full_Adder FA_206(s206, c206, in206_1, in206_2, pp45[17]);
    wire[0:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {pp49[13]};
    assign in207_2 = {pp50[12]};
    Full_Adder FA_207(s207, c207, in207_1, in207_2, pp48[14]);
    wire[0:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {pp52[10]};
    assign in208_2 = {pp53[9]};
    Full_Adder FA_208(s208, c208, in208_1, in208_2, pp51[11]);
    wire[0:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {pp55[7]};
    assign in209_2 = {pp56[6]};
    Full_Adder FA_209(s209, c209, in209_1, in209_2, pp54[8]);
    wire[0:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {pp57[5]};
    assign in210_2 = {pp58[4]};
    Half_Adder HA_210(s210, c210, in210_1, in210_2);
    wire[0:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {pp1[62]};
    assign in211_2 = {pp2[61]};
    Full_Adder FA_211(s211, c211, in211_1, in211_2, pp0[63]);
    wire[0:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {pp4[59]};
    assign in212_2 = {pp5[58]};
    Full_Adder FA_212(s212, c212, in212_1, in212_2, pp3[60]);
    wire[0:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {pp7[56]};
    assign in213_2 = {pp8[55]};
    Full_Adder FA_213(s213, c213, in213_1, in213_2, pp6[57]);
    wire[0:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {pp10[53]};
    assign in214_2 = {pp11[52]};
    Full_Adder FA_214(s214, c214, in214_1, in214_2, pp9[54]);
    wire[0:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {pp13[50]};
    assign in215_2 = {pp14[49]};
    Full_Adder FA_215(s215, c215, in215_1, in215_2, pp12[51]);
    wire[0:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {pp16[47]};
    assign in216_2 = {pp17[46]};
    Full_Adder FA_216(s216, c216, in216_1, in216_2, pp15[48]);
    wire[0:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {pp19[44]};
    assign in217_2 = {pp20[43]};
    Full_Adder FA_217(s217, c217, in217_1, in217_2, pp18[45]);
    wire[0:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {pp22[41]};
    assign in218_2 = {pp23[40]};
    Full_Adder FA_218(s218, c218, in218_1, in218_2, pp21[42]);
    wire[0:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {pp25[38]};
    assign in219_2 = {pp26[37]};
    Full_Adder FA_219(s219, c219, in219_1, in219_2, pp24[39]);
    wire[0:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {pp28[35]};
    assign in220_2 = {pp29[34]};
    Full_Adder FA_220(s220, c220, in220_1, in220_2, pp27[36]);
    wire[0:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {pp31[32]};
    assign in221_2 = {pp32[31]};
    Full_Adder FA_221(s221, c221, in221_1, in221_2, pp30[33]);
    wire[0:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {pp34[29]};
    assign in222_2 = {pp35[28]};
    Full_Adder FA_222(s222, c222, in222_1, in222_2, pp33[30]);
    wire[0:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {pp37[26]};
    assign in223_2 = {pp38[25]};
    Full_Adder FA_223(s223, c223, in223_1, in223_2, pp36[27]);
    wire[0:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {pp40[23]};
    assign in224_2 = {pp41[22]};
    Full_Adder FA_224(s224, c224, in224_1, in224_2, pp39[24]);
    wire[0:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {pp43[20]};
    assign in225_2 = {pp44[19]};
    Full_Adder FA_225(s225, c225, in225_1, in225_2, pp42[21]);
    wire[0:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {pp46[17]};
    assign in226_2 = {pp47[16]};
    Full_Adder FA_226(s226, c226, in226_1, in226_2, pp45[18]);
    wire[0:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {pp49[14]};
    assign in227_2 = {pp50[13]};
    Full_Adder FA_227(s227, c227, in227_1, in227_2, pp48[15]);
    wire[0:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {pp52[11]};
    assign in228_2 = {pp53[10]};
    Full_Adder FA_228(s228, c228, in228_1, in228_2, pp51[12]);
    wire[0:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {pp55[8]};
    assign in229_2 = {pp56[7]};
    Full_Adder FA_229(s229, c229, in229_1, in229_2, pp54[9]);
    wire[0:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp58[5]};
    assign in230_2 = {pp59[4]};
    Full_Adder FA_230(s230, c230, in230_1, in230_2, pp57[6]);
    wire[0:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp60[3]};
    assign in231_2 = {pp61[2]};
    Half_Adder HA_231(s231, c231, in231_1, in231_2);
    wire[0:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {pp2[62]};
    assign in232_2 = {pp3[61]};
    Full_Adder FA_232(s232, c232, in232_1, in232_2, pp1[63]);
    wire[0:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {pp5[59]};
    assign in233_2 = {pp6[58]};
    Full_Adder FA_233(s233, c233, in233_1, in233_2, pp4[60]);
    wire[0:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {pp8[56]};
    assign in234_2 = {pp9[55]};
    Full_Adder FA_234(s234, c234, in234_1, in234_2, pp7[57]);
    wire[0:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {pp11[53]};
    assign in235_2 = {pp12[52]};
    Full_Adder FA_235(s235, c235, in235_1, in235_2, pp10[54]);
    wire[0:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {pp14[50]};
    assign in236_2 = {pp15[49]};
    Full_Adder FA_236(s236, c236, in236_1, in236_2, pp13[51]);
    wire[0:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {pp17[47]};
    assign in237_2 = {pp18[46]};
    Full_Adder FA_237(s237, c237, in237_1, in237_2, pp16[48]);
    wire[0:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {pp20[44]};
    assign in238_2 = {pp21[43]};
    Full_Adder FA_238(s238, c238, in238_1, in238_2, pp19[45]);
    wire[0:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {pp23[41]};
    assign in239_2 = {pp24[40]};
    Full_Adder FA_239(s239, c239, in239_1, in239_2, pp22[42]);
    wire[0:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {pp26[38]};
    assign in240_2 = {pp27[37]};
    Full_Adder FA_240(s240, c240, in240_1, in240_2, pp25[39]);
    wire[0:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {pp29[35]};
    assign in241_2 = {pp30[34]};
    Full_Adder FA_241(s241, c241, in241_1, in241_2, pp28[36]);
    wire[0:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {pp32[32]};
    assign in242_2 = {pp33[31]};
    Full_Adder FA_242(s242, c242, in242_1, in242_2, pp31[33]);
    wire[0:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {pp35[29]};
    assign in243_2 = {pp36[28]};
    Full_Adder FA_243(s243, c243, in243_1, in243_2, pp34[30]);
    wire[0:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp38[26]};
    assign in244_2 = {pp39[25]};
    Full_Adder FA_244(s244, c244, in244_1, in244_2, pp37[27]);
    wire[0:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {pp41[23]};
    assign in245_2 = {pp42[22]};
    Full_Adder FA_245(s245, c245, in245_1, in245_2, pp40[24]);
    wire[0:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {pp44[20]};
    assign in246_2 = {pp45[19]};
    Full_Adder FA_246(s246, c246, in246_1, in246_2, pp43[21]);
    wire[0:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {pp47[17]};
    assign in247_2 = {pp48[16]};
    Full_Adder FA_247(s247, c247, in247_1, in247_2, pp46[18]);
    wire[0:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {pp50[14]};
    assign in248_2 = {pp51[13]};
    Full_Adder FA_248(s248, c248, in248_1, in248_2, pp49[15]);
    wire[0:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {pp53[11]};
    assign in249_2 = {pp54[10]};
    Full_Adder FA_249(s249, c249, in249_1, in249_2, pp52[12]);
    wire[0:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {pp56[8]};
    assign in250_2 = {pp57[7]};
    Full_Adder FA_250(s250, c250, in250_1, in250_2, pp55[9]);
    wire[0:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp59[5]};
    assign in251_2 = {pp60[4]};
    Full_Adder FA_251(s251, c251, in251_1, in251_2, pp58[6]);
    wire[0:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp61[3]};
    assign in252_2 = {pp62[2]};
    Half_Adder HA_252(s252, c252, in252_1, in252_2);
    wire[0:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp3[62]};
    assign in253_2 = {pp4[61]};
    Full_Adder FA_253(s253, c253, in253_1, in253_2, pp2[63]);
    wire[0:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp6[59]};
    assign in254_2 = {pp7[58]};
    Full_Adder FA_254(s254, c254, in254_1, in254_2, pp5[60]);
    wire[0:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {pp9[56]};
    assign in255_2 = {pp10[55]};
    Full_Adder FA_255(s255, c255, in255_1, in255_2, pp8[57]);
    wire[0:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {pp12[53]};
    assign in256_2 = {pp13[52]};
    Full_Adder FA_256(s256, c256, in256_1, in256_2, pp11[54]);
    wire[0:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {pp15[50]};
    assign in257_2 = {pp16[49]};
    Full_Adder FA_257(s257, c257, in257_1, in257_2, pp14[51]);
    wire[0:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {pp18[47]};
    assign in258_2 = {pp19[46]};
    Full_Adder FA_258(s258, c258, in258_1, in258_2, pp17[48]);
    wire[0:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {pp21[44]};
    assign in259_2 = {pp22[43]};
    Full_Adder FA_259(s259, c259, in259_1, in259_2, pp20[45]);
    wire[0:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {pp24[41]};
    assign in260_2 = {pp25[40]};
    Full_Adder FA_260(s260, c260, in260_1, in260_2, pp23[42]);
    wire[0:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {pp27[38]};
    assign in261_2 = {pp28[37]};
    Full_Adder FA_261(s261, c261, in261_1, in261_2, pp26[39]);
    wire[0:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {pp30[35]};
    assign in262_2 = {pp31[34]};
    Full_Adder FA_262(s262, c262, in262_1, in262_2, pp29[36]);
    wire[0:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {pp33[32]};
    assign in263_2 = {pp34[31]};
    Full_Adder FA_263(s263, c263, in263_1, in263_2, pp32[33]);
    wire[0:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {pp36[29]};
    assign in264_2 = {pp37[28]};
    Full_Adder FA_264(s264, c264, in264_1, in264_2, pp35[30]);
    wire[0:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {pp39[26]};
    assign in265_2 = {pp40[25]};
    Full_Adder FA_265(s265, c265, in265_1, in265_2, pp38[27]);
    wire[0:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {pp42[23]};
    assign in266_2 = {pp43[22]};
    Full_Adder FA_266(s266, c266, in266_1, in266_2, pp41[24]);
    wire[0:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {pp45[20]};
    assign in267_2 = {pp46[19]};
    Full_Adder FA_267(s267, c267, in267_1, in267_2, pp44[21]);
    wire[0:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {pp48[17]};
    assign in268_2 = {pp49[16]};
    Full_Adder FA_268(s268, c268, in268_1, in268_2, pp47[18]);
    wire[0:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {pp51[14]};
    assign in269_2 = {pp52[13]};
    Full_Adder FA_269(s269, c269, in269_1, in269_2, pp50[15]);
    wire[0:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {pp54[11]};
    assign in270_2 = {pp55[10]};
    Full_Adder FA_270(s270, c270, in270_1, in270_2, pp53[12]);
    wire[0:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {pp57[8]};
    assign in271_2 = {pp58[7]};
    Full_Adder FA_271(s271, c271, in271_1, in271_2, pp56[9]);
    wire[0:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {pp60[5]};
    assign in272_2 = {pp61[4]};
    Full_Adder FA_272(s272, c272, in272_1, in272_2, pp59[6]);
    wire[0:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {pp4[62]};
    assign in273_2 = {pp5[61]};
    Full_Adder FA_273(s273, c273, in273_1, in273_2, pp3[63]);
    wire[0:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {pp7[59]};
    assign in274_2 = {pp8[58]};
    Full_Adder FA_274(s274, c274, in274_1, in274_2, pp6[60]);
    wire[0:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp10[56]};
    assign in275_2 = {pp11[55]};
    Full_Adder FA_275(s275, c275, in275_1, in275_2, pp9[57]);
    wire[0:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {pp13[53]};
    assign in276_2 = {pp14[52]};
    Full_Adder FA_276(s276, c276, in276_1, in276_2, pp12[54]);
    wire[0:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {pp16[50]};
    assign in277_2 = {pp17[49]};
    Full_Adder FA_277(s277, c277, in277_1, in277_2, pp15[51]);
    wire[0:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {pp19[47]};
    assign in278_2 = {pp20[46]};
    Full_Adder FA_278(s278, c278, in278_1, in278_2, pp18[48]);
    wire[0:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {pp22[44]};
    assign in279_2 = {pp23[43]};
    Full_Adder FA_279(s279, c279, in279_1, in279_2, pp21[45]);
    wire[0:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {pp25[41]};
    assign in280_2 = {pp26[40]};
    Full_Adder FA_280(s280, c280, in280_1, in280_2, pp24[42]);
    wire[0:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {pp28[38]};
    assign in281_2 = {pp29[37]};
    Full_Adder FA_281(s281, c281, in281_1, in281_2, pp27[39]);
    wire[0:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {pp31[35]};
    assign in282_2 = {pp32[34]};
    Full_Adder FA_282(s282, c282, in282_1, in282_2, pp30[36]);
    wire[0:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {pp34[32]};
    assign in283_2 = {pp35[31]};
    Full_Adder FA_283(s283, c283, in283_1, in283_2, pp33[33]);
    wire[0:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {pp37[29]};
    assign in284_2 = {pp38[28]};
    Full_Adder FA_284(s284, c284, in284_1, in284_2, pp36[30]);
    wire[0:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {pp40[26]};
    assign in285_2 = {pp41[25]};
    Full_Adder FA_285(s285, c285, in285_1, in285_2, pp39[27]);
    wire[0:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {pp43[23]};
    assign in286_2 = {pp44[22]};
    Full_Adder FA_286(s286, c286, in286_1, in286_2, pp42[24]);
    wire[0:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {pp46[20]};
    assign in287_2 = {pp47[19]};
    Full_Adder FA_287(s287, c287, in287_1, in287_2, pp45[21]);
    wire[0:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {pp49[17]};
    assign in288_2 = {pp50[16]};
    Full_Adder FA_288(s288, c288, in288_1, in288_2, pp48[18]);
    wire[0:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {pp52[14]};
    assign in289_2 = {pp53[13]};
    Full_Adder FA_289(s289, c289, in289_1, in289_2, pp51[15]);
    wire[0:0] s290, in290_1, in290_2;
    wire c290;
    assign in290_1 = {pp55[11]};
    assign in290_2 = {pp56[10]};
    Full_Adder FA_290(s290, c290, in290_1, in290_2, pp54[12]);
    wire[0:0] s291, in291_1, in291_2;
    wire c291;
    assign in291_1 = {pp58[8]};
    assign in291_2 = {pp59[7]};
    Full_Adder FA_291(s291, c291, in291_1, in291_2, pp57[9]);
    wire[0:0] s292, in292_1, in292_2;
    wire c292;
    assign in292_1 = {pp5[62]};
    assign in292_2 = {pp6[61]};
    Full_Adder FA_292(s292, c292, in292_1, in292_2, pp4[63]);
    wire[0:0] s293, in293_1, in293_2;
    wire c293;
    assign in293_1 = {pp8[59]};
    assign in293_2 = {pp9[58]};
    Full_Adder FA_293(s293, c293, in293_1, in293_2, pp7[60]);
    wire[0:0] s294, in294_1, in294_2;
    wire c294;
    assign in294_1 = {pp11[56]};
    assign in294_2 = {pp12[55]};
    Full_Adder FA_294(s294, c294, in294_1, in294_2, pp10[57]);
    wire[0:0] s295, in295_1, in295_2;
    wire c295;
    assign in295_1 = {pp14[53]};
    assign in295_2 = {pp15[52]};
    Full_Adder FA_295(s295, c295, in295_1, in295_2, pp13[54]);
    wire[0:0] s296, in296_1, in296_2;
    wire c296;
    assign in296_1 = {pp17[50]};
    assign in296_2 = {pp18[49]};
    Full_Adder FA_296(s296, c296, in296_1, in296_2, pp16[51]);
    wire[0:0] s297, in297_1, in297_2;
    wire c297;
    assign in297_1 = {pp20[47]};
    assign in297_2 = {pp21[46]};
    Full_Adder FA_297(s297, c297, in297_1, in297_2, pp19[48]);
    wire[0:0] s298, in298_1, in298_2;
    wire c298;
    assign in298_1 = {pp23[44]};
    assign in298_2 = {pp24[43]};
    Full_Adder FA_298(s298, c298, in298_1, in298_2, pp22[45]);
    wire[0:0] s299, in299_1, in299_2;
    wire c299;
    assign in299_1 = {pp26[41]};
    assign in299_2 = {pp27[40]};
    Full_Adder FA_299(s299, c299, in299_1, in299_2, pp25[42]);
    wire[0:0] s300, in300_1, in300_2;
    wire c300;
    assign in300_1 = {pp29[38]};
    assign in300_2 = {pp30[37]};
    Full_Adder FA_300(s300, c300, in300_1, in300_2, pp28[39]);
    wire[0:0] s301, in301_1, in301_2;
    wire c301;
    assign in301_1 = {pp32[35]};
    assign in301_2 = {pp33[34]};
    Full_Adder FA_301(s301, c301, in301_1, in301_2, pp31[36]);
    wire[0:0] s302, in302_1, in302_2;
    wire c302;
    assign in302_1 = {pp35[32]};
    assign in302_2 = {pp36[31]};
    Full_Adder FA_302(s302, c302, in302_1, in302_2, pp34[33]);
    wire[0:0] s303, in303_1, in303_2;
    wire c303;
    assign in303_1 = {pp38[29]};
    assign in303_2 = {pp39[28]};
    Full_Adder FA_303(s303, c303, in303_1, in303_2, pp37[30]);
    wire[0:0] s304, in304_1, in304_2;
    wire c304;
    assign in304_1 = {pp41[26]};
    assign in304_2 = {pp42[25]};
    Full_Adder FA_304(s304, c304, in304_1, in304_2, pp40[27]);
    wire[0:0] s305, in305_1, in305_2;
    wire c305;
    assign in305_1 = {pp44[23]};
    assign in305_2 = {pp45[22]};
    Full_Adder FA_305(s305, c305, in305_1, in305_2, pp43[24]);
    wire[0:0] s306, in306_1, in306_2;
    wire c306;
    assign in306_1 = {pp47[20]};
    assign in306_2 = {pp48[19]};
    Full_Adder FA_306(s306, c306, in306_1, in306_2, pp46[21]);
    wire[0:0] s307, in307_1, in307_2;
    wire c307;
    assign in307_1 = {pp50[17]};
    assign in307_2 = {pp51[16]};
    Full_Adder FA_307(s307, c307, in307_1, in307_2, pp49[18]);
    wire[0:0] s308, in308_1, in308_2;
    wire c308;
    assign in308_1 = {pp53[14]};
    assign in308_2 = {pp54[13]};
    Full_Adder FA_308(s308, c308, in308_1, in308_2, pp52[15]);
    wire[0:0] s309, in309_1, in309_2;
    wire c309;
    assign in309_1 = {pp56[11]};
    assign in309_2 = {pp57[10]};
    Full_Adder FA_309(s309, c309, in309_1, in309_2, pp55[12]);
    wire[0:0] s310, in310_1, in310_2;
    wire c310;
    assign in310_1 = {pp6[62]};
    assign in310_2 = {pp7[61]};
    Full_Adder FA_310(s310, c310, in310_1, in310_2, pp5[63]);
    wire[0:0] s311, in311_1, in311_2;
    wire c311;
    assign in311_1 = {pp9[59]};
    assign in311_2 = {pp10[58]};
    Full_Adder FA_311(s311, c311, in311_1, in311_2, pp8[60]);
    wire[0:0] s312, in312_1, in312_2;
    wire c312;
    assign in312_1 = {pp12[56]};
    assign in312_2 = {pp13[55]};
    Full_Adder FA_312(s312, c312, in312_1, in312_2, pp11[57]);
    wire[0:0] s313, in313_1, in313_2;
    wire c313;
    assign in313_1 = {pp15[53]};
    assign in313_2 = {pp16[52]};
    Full_Adder FA_313(s313, c313, in313_1, in313_2, pp14[54]);
    wire[0:0] s314, in314_1, in314_2;
    wire c314;
    assign in314_1 = {pp18[50]};
    assign in314_2 = {pp19[49]};
    Full_Adder FA_314(s314, c314, in314_1, in314_2, pp17[51]);
    wire[0:0] s315, in315_1, in315_2;
    wire c315;
    assign in315_1 = {pp21[47]};
    assign in315_2 = {pp22[46]};
    Full_Adder FA_315(s315, c315, in315_1, in315_2, pp20[48]);
    wire[0:0] s316, in316_1, in316_2;
    wire c316;
    assign in316_1 = {pp24[44]};
    assign in316_2 = {pp25[43]};
    Full_Adder FA_316(s316, c316, in316_1, in316_2, pp23[45]);
    wire[0:0] s317, in317_1, in317_2;
    wire c317;
    assign in317_1 = {pp27[41]};
    assign in317_2 = {pp28[40]};
    Full_Adder FA_317(s317, c317, in317_1, in317_2, pp26[42]);
    wire[0:0] s318, in318_1, in318_2;
    wire c318;
    assign in318_1 = {pp30[38]};
    assign in318_2 = {pp31[37]};
    Full_Adder FA_318(s318, c318, in318_1, in318_2, pp29[39]);
    wire[0:0] s319, in319_1, in319_2;
    wire c319;
    assign in319_1 = {pp33[35]};
    assign in319_2 = {pp34[34]};
    Full_Adder FA_319(s319, c319, in319_1, in319_2, pp32[36]);
    wire[0:0] s320, in320_1, in320_2;
    wire c320;
    assign in320_1 = {pp36[32]};
    assign in320_2 = {pp37[31]};
    Full_Adder FA_320(s320, c320, in320_1, in320_2, pp35[33]);
    wire[0:0] s321, in321_1, in321_2;
    wire c321;
    assign in321_1 = {pp39[29]};
    assign in321_2 = {pp40[28]};
    Full_Adder FA_321(s321, c321, in321_1, in321_2, pp38[30]);
    wire[0:0] s322, in322_1, in322_2;
    wire c322;
    assign in322_1 = {pp42[26]};
    assign in322_2 = {pp43[25]};
    Full_Adder FA_322(s322, c322, in322_1, in322_2, pp41[27]);
    wire[0:0] s323, in323_1, in323_2;
    wire c323;
    assign in323_1 = {pp45[23]};
    assign in323_2 = {pp46[22]};
    Full_Adder FA_323(s323, c323, in323_1, in323_2, pp44[24]);
    wire[0:0] s324, in324_1, in324_2;
    wire c324;
    assign in324_1 = {pp48[20]};
    assign in324_2 = {pp49[19]};
    Full_Adder FA_324(s324, c324, in324_1, in324_2, pp47[21]);
    wire[0:0] s325, in325_1, in325_2;
    wire c325;
    assign in325_1 = {pp51[17]};
    assign in325_2 = {pp52[16]};
    Full_Adder FA_325(s325, c325, in325_1, in325_2, pp50[18]);
    wire[0:0] s326, in326_1, in326_2;
    wire c326;
    assign in326_1 = {pp54[14]};
    assign in326_2 = {pp55[13]};
    Full_Adder FA_326(s326, c326, in326_1, in326_2, pp53[15]);
    wire[0:0] s327, in327_1, in327_2;
    wire c327;
    assign in327_1 = {pp7[62]};
    assign in327_2 = {pp8[61]};
    Full_Adder FA_327(s327, c327, in327_1, in327_2, pp6[63]);
    wire[0:0] s328, in328_1, in328_2;
    wire c328;
    assign in328_1 = {pp10[59]};
    assign in328_2 = {pp11[58]};
    Full_Adder FA_328(s328, c328, in328_1, in328_2, pp9[60]);
    wire[0:0] s329, in329_1, in329_2;
    wire c329;
    assign in329_1 = {pp13[56]};
    assign in329_2 = {pp14[55]};
    Full_Adder FA_329(s329, c329, in329_1, in329_2, pp12[57]);
    wire[0:0] s330, in330_1, in330_2;
    wire c330;
    assign in330_1 = {pp16[53]};
    assign in330_2 = {pp17[52]};
    Full_Adder FA_330(s330, c330, in330_1, in330_2, pp15[54]);
    wire[0:0] s331, in331_1, in331_2;
    wire c331;
    assign in331_1 = {pp19[50]};
    assign in331_2 = {pp20[49]};
    Full_Adder FA_331(s331, c331, in331_1, in331_2, pp18[51]);
    wire[0:0] s332, in332_1, in332_2;
    wire c332;
    assign in332_1 = {pp22[47]};
    assign in332_2 = {pp23[46]};
    Full_Adder FA_332(s332, c332, in332_1, in332_2, pp21[48]);
    wire[0:0] s333, in333_1, in333_2;
    wire c333;
    assign in333_1 = {pp25[44]};
    assign in333_2 = {pp26[43]};
    Full_Adder FA_333(s333, c333, in333_1, in333_2, pp24[45]);
    wire[0:0] s334, in334_1, in334_2;
    wire c334;
    assign in334_1 = {pp28[41]};
    assign in334_2 = {pp29[40]};
    Full_Adder FA_334(s334, c334, in334_1, in334_2, pp27[42]);
    wire[0:0] s335, in335_1, in335_2;
    wire c335;
    assign in335_1 = {pp31[38]};
    assign in335_2 = {pp32[37]};
    Full_Adder FA_335(s335, c335, in335_1, in335_2, pp30[39]);
    wire[0:0] s336, in336_1, in336_2;
    wire c336;
    assign in336_1 = {pp34[35]};
    assign in336_2 = {pp35[34]};
    Full_Adder FA_336(s336, c336, in336_1, in336_2, pp33[36]);
    wire[0:0] s337, in337_1, in337_2;
    wire c337;
    assign in337_1 = {pp37[32]};
    assign in337_2 = {pp38[31]};
    Full_Adder FA_337(s337, c337, in337_1, in337_2, pp36[33]);
    wire[0:0] s338, in338_1, in338_2;
    wire c338;
    assign in338_1 = {pp40[29]};
    assign in338_2 = {pp41[28]};
    Full_Adder FA_338(s338, c338, in338_1, in338_2, pp39[30]);
    wire[0:0] s339, in339_1, in339_2;
    wire c339;
    assign in339_1 = {pp43[26]};
    assign in339_2 = {pp44[25]};
    Full_Adder FA_339(s339, c339, in339_1, in339_2, pp42[27]);
    wire[0:0] s340, in340_1, in340_2;
    wire c340;
    assign in340_1 = {pp46[23]};
    assign in340_2 = {pp47[22]};
    Full_Adder FA_340(s340, c340, in340_1, in340_2, pp45[24]);
    wire[0:0] s341, in341_1, in341_2;
    wire c341;
    assign in341_1 = {pp49[20]};
    assign in341_2 = {pp50[19]};
    Full_Adder FA_341(s341, c341, in341_1, in341_2, pp48[21]);
    wire[0:0] s342, in342_1, in342_2;
    wire c342;
    assign in342_1 = {pp52[17]};
    assign in342_2 = {pp53[16]};
    Full_Adder FA_342(s342, c342, in342_1, in342_2, pp51[18]);
    wire[0:0] s343, in343_1, in343_2;
    wire c343;
    assign in343_1 = {pp8[62]};
    assign in343_2 = {pp9[61]};
    Full_Adder FA_343(s343, c343, in343_1, in343_2, pp7[63]);
    wire[0:0] s344, in344_1, in344_2;
    wire c344;
    assign in344_1 = {pp11[59]};
    assign in344_2 = {pp12[58]};
    Full_Adder FA_344(s344, c344, in344_1, in344_2, pp10[60]);
    wire[0:0] s345, in345_1, in345_2;
    wire c345;
    assign in345_1 = {pp14[56]};
    assign in345_2 = {pp15[55]};
    Full_Adder FA_345(s345, c345, in345_1, in345_2, pp13[57]);
    wire[0:0] s346, in346_1, in346_2;
    wire c346;
    assign in346_1 = {pp17[53]};
    assign in346_2 = {pp18[52]};
    Full_Adder FA_346(s346, c346, in346_1, in346_2, pp16[54]);
    wire[0:0] s347, in347_1, in347_2;
    wire c347;
    assign in347_1 = {pp20[50]};
    assign in347_2 = {pp21[49]};
    Full_Adder FA_347(s347, c347, in347_1, in347_2, pp19[51]);
    wire[0:0] s348, in348_1, in348_2;
    wire c348;
    assign in348_1 = {pp23[47]};
    assign in348_2 = {pp24[46]};
    Full_Adder FA_348(s348, c348, in348_1, in348_2, pp22[48]);
    wire[0:0] s349, in349_1, in349_2;
    wire c349;
    assign in349_1 = {pp26[44]};
    assign in349_2 = {pp27[43]};
    Full_Adder FA_349(s349, c349, in349_1, in349_2, pp25[45]);
    wire[0:0] s350, in350_1, in350_2;
    wire c350;
    assign in350_1 = {pp29[41]};
    assign in350_2 = {pp30[40]};
    Full_Adder FA_350(s350, c350, in350_1, in350_2, pp28[42]);
    wire[0:0] s351, in351_1, in351_2;
    wire c351;
    assign in351_1 = {pp32[38]};
    assign in351_2 = {pp33[37]};
    Full_Adder FA_351(s351, c351, in351_1, in351_2, pp31[39]);
    wire[0:0] s352, in352_1, in352_2;
    wire c352;
    assign in352_1 = {pp35[35]};
    assign in352_2 = {pp36[34]};
    Full_Adder FA_352(s352, c352, in352_1, in352_2, pp34[36]);
    wire[0:0] s353, in353_1, in353_2;
    wire c353;
    assign in353_1 = {pp38[32]};
    assign in353_2 = {pp39[31]};
    Full_Adder FA_353(s353, c353, in353_1, in353_2, pp37[33]);
    wire[0:0] s354, in354_1, in354_2;
    wire c354;
    assign in354_1 = {pp41[29]};
    assign in354_2 = {pp42[28]};
    Full_Adder FA_354(s354, c354, in354_1, in354_2, pp40[30]);
    wire[0:0] s355, in355_1, in355_2;
    wire c355;
    assign in355_1 = {pp44[26]};
    assign in355_2 = {pp45[25]};
    Full_Adder FA_355(s355, c355, in355_1, in355_2, pp43[27]);
    wire[0:0] s356, in356_1, in356_2;
    wire c356;
    assign in356_1 = {pp47[23]};
    assign in356_2 = {pp48[22]};
    Full_Adder FA_356(s356, c356, in356_1, in356_2, pp46[24]);
    wire[0:0] s357, in357_1, in357_2;
    wire c357;
    assign in357_1 = {pp50[20]};
    assign in357_2 = {pp51[19]};
    Full_Adder FA_357(s357, c357, in357_1, in357_2, pp49[21]);
    wire[0:0] s358, in358_1, in358_2;
    wire c358;
    assign in358_1 = {pp9[62]};
    assign in358_2 = {pp10[61]};
    Full_Adder FA_358(s358, c358, in358_1, in358_2, pp8[63]);
    wire[0:0] s359, in359_1, in359_2;
    wire c359;
    assign in359_1 = {pp12[59]};
    assign in359_2 = {pp13[58]};
    Full_Adder FA_359(s359, c359, in359_1, in359_2, pp11[60]);
    wire[0:0] s360, in360_1, in360_2;
    wire c360;
    assign in360_1 = {pp15[56]};
    assign in360_2 = {pp16[55]};
    Full_Adder FA_360(s360, c360, in360_1, in360_2, pp14[57]);
    wire[0:0] s361, in361_1, in361_2;
    wire c361;
    assign in361_1 = {pp18[53]};
    assign in361_2 = {pp19[52]};
    Full_Adder FA_361(s361, c361, in361_1, in361_2, pp17[54]);
    wire[0:0] s362, in362_1, in362_2;
    wire c362;
    assign in362_1 = {pp21[50]};
    assign in362_2 = {pp22[49]};
    Full_Adder FA_362(s362, c362, in362_1, in362_2, pp20[51]);
    wire[0:0] s363, in363_1, in363_2;
    wire c363;
    assign in363_1 = {pp24[47]};
    assign in363_2 = {pp25[46]};
    Full_Adder FA_363(s363, c363, in363_1, in363_2, pp23[48]);
    wire[0:0] s364, in364_1, in364_2;
    wire c364;
    assign in364_1 = {pp27[44]};
    assign in364_2 = {pp28[43]};
    Full_Adder FA_364(s364, c364, in364_1, in364_2, pp26[45]);
    wire[0:0] s365, in365_1, in365_2;
    wire c365;
    assign in365_1 = {pp30[41]};
    assign in365_2 = {pp31[40]};
    Full_Adder FA_365(s365, c365, in365_1, in365_2, pp29[42]);
    wire[0:0] s366, in366_1, in366_2;
    wire c366;
    assign in366_1 = {pp33[38]};
    assign in366_2 = {pp34[37]};
    Full_Adder FA_366(s366, c366, in366_1, in366_2, pp32[39]);
    wire[0:0] s367, in367_1, in367_2;
    wire c367;
    assign in367_1 = {pp36[35]};
    assign in367_2 = {pp37[34]};
    Full_Adder FA_367(s367, c367, in367_1, in367_2, pp35[36]);
    wire[0:0] s368, in368_1, in368_2;
    wire c368;
    assign in368_1 = {pp39[32]};
    assign in368_2 = {pp40[31]};
    Full_Adder FA_368(s368, c368, in368_1, in368_2, pp38[33]);
    wire[0:0] s369, in369_1, in369_2;
    wire c369;
    assign in369_1 = {pp42[29]};
    assign in369_2 = {pp43[28]};
    Full_Adder FA_369(s369, c369, in369_1, in369_2, pp41[30]);
    wire[0:0] s370, in370_1, in370_2;
    wire c370;
    assign in370_1 = {pp45[26]};
    assign in370_2 = {pp46[25]};
    Full_Adder FA_370(s370, c370, in370_1, in370_2, pp44[27]);
    wire[0:0] s371, in371_1, in371_2;
    wire c371;
    assign in371_1 = {pp48[23]};
    assign in371_2 = {pp49[22]};
    Full_Adder FA_371(s371, c371, in371_1, in371_2, pp47[24]);
    wire[0:0] s372, in372_1, in372_2;
    wire c372;
    assign in372_1 = {pp10[62]};
    assign in372_2 = {pp11[61]};
    Full_Adder FA_372(s372, c372, in372_1, in372_2, pp9[63]);
    wire[0:0] s373, in373_1, in373_2;
    wire c373;
    assign in373_1 = {pp13[59]};
    assign in373_2 = {pp14[58]};
    Full_Adder FA_373(s373, c373, in373_1, in373_2, pp12[60]);
    wire[0:0] s374, in374_1, in374_2;
    wire c374;
    assign in374_1 = {pp16[56]};
    assign in374_2 = {pp17[55]};
    Full_Adder FA_374(s374, c374, in374_1, in374_2, pp15[57]);
    wire[0:0] s375, in375_1, in375_2;
    wire c375;
    assign in375_1 = {pp19[53]};
    assign in375_2 = {pp20[52]};
    Full_Adder FA_375(s375, c375, in375_1, in375_2, pp18[54]);
    wire[0:0] s376, in376_1, in376_2;
    wire c376;
    assign in376_1 = {pp22[50]};
    assign in376_2 = {pp23[49]};
    Full_Adder FA_376(s376, c376, in376_1, in376_2, pp21[51]);
    wire[0:0] s377, in377_1, in377_2;
    wire c377;
    assign in377_1 = {pp25[47]};
    assign in377_2 = {pp26[46]};
    Full_Adder FA_377(s377, c377, in377_1, in377_2, pp24[48]);
    wire[0:0] s378, in378_1, in378_2;
    wire c378;
    assign in378_1 = {pp28[44]};
    assign in378_2 = {pp29[43]};
    Full_Adder FA_378(s378, c378, in378_1, in378_2, pp27[45]);
    wire[0:0] s379, in379_1, in379_2;
    wire c379;
    assign in379_1 = {pp31[41]};
    assign in379_2 = {pp32[40]};
    Full_Adder FA_379(s379, c379, in379_1, in379_2, pp30[42]);
    wire[0:0] s380, in380_1, in380_2;
    wire c380;
    assign in380_1 = {pp34[38]};
    assign in380_2 = {pp35[37]};
    Full_Adder FA_380(s380, c380, in380_1, in380_2, pp33[39]);
    wire[0:0] s381, in381_1, in381_2;
    wire c381;
    assign in381_1 = {pp37[35]};
    assign in381_2 = {pp38[34]};
    Full_Adder FA_381(s381, c381, in381_1, in381_2, pp36[36]);
    wire[0:0] s382, in382_1, in382_2;
    wire c382;
    assign in382_1 = {pp40[32]};
    assign in382_2 = {pp41[31]};
    Full_Adder FA_382(s382, c382, in382_1, in382_2, pp39[33]);
    wire[0:0] s383, in383_1, in383_2;
    wire c383;
    assign in383_1 = {pp43[29]};
    assign in383_2 = {pp44[28]};
    Full_Adder FA_383(s383, c383, in383_1, in383_2, pp42[30]);
    wire[0:0] s384, in384_1, in384_2;
    wire c384;
    assign in384_1 = {pp46[26]};
    assign in384_2 = {pp47[25]};
    Full_Adder FA_384(s384, c384, in384_1, in384_2, pp45[27]);
    wire[0:0] s385, in385_1, in385_2;
    wire c385;
    assign in385_1 = {pp11[62]};
    assign in385_2 = {pp12[61]};
    Full_Adder FA_385(s385, c385, in385_1, in385_2, pp10[63]);
    wire[0:0] s386, in386_1, in386_2;
    wire c386;
    assign in386_1 = {pp14[59]};
    assign in386_2 = {pp15[58]};
    Full_Adder FA_386(s386, c386, in386_1, in386_2, pp13[60]);
    wire[0:0] s387, in387_1, in387_2;
    wire c387;
    assign in387_1 = {pp17[56]};
    assign in387_2 = {pp18[55]};
    Full_Adder FA_387(s387, c387, in387_1, in387_2, pp16[57]);
    wire[0:0] s388, in388_1, in388_2;
    wire c388;
    assign in388_1 = {pp20[53]};
    assign in388_2 = {pp21[52]};
    Full_Adder FA_388(s388, c388, in388_1, in388_2, pp19[54]);
    wire[0:0] s389, in389_1, in389_2;
    wire c389;
    assign in389_1 = {pp23[50]};
    assign in389_2 = {pp24[49]};
    Full_Adder FA_389(s389, c389, in389_1, in389_2, pp22[51]);
    wire[0:0] s390, in390_1, in390_2;
    wire c390;
    assign in390_1 = {pp26[47]};
    assign in390_2 = {pp27[46]};
    Full_Adder FA_390(s390, c390, in390_1, in390_2, pp25[48]);
    wire[0:0] s391, in391_1, in391_2;
    wire c391;
    assign in391_1 = {pp29[44]};
    assign in391_2 = {pp30[43]};
    Full_Adder FA_391(s391, c391, in391_1, in391_2, pp28[45]);
    wire[0:0] s392, in392_1, in392_2;
    wire c392;
    assign in392_1 = {pp32[41]};
    assign in392_2 = {pp33[40]};
    Full_Adder FA_392(s392, c392, in392_1, in392_2, pp31[42]);
    wire[0:0] s393, in393_1, in393_2;
    wire c393;
    assign in393_1 = {pp35[38]};
    assign in393_2 = {pp36[37]};
    Full_Adder FA_393(s393, c393, in393_1, in393_2, pp34[39]);
    wire[0:0] s394, in394_1, in394_2;
    wire c394;
    assign in394_1 = {pp38[35]};
    assign in394_2 = {pp39[34]};
    Full_Adder FA_394(s394, c394, in394_1, in394_2, pp37[36]);
    wire[0:0] s395, in395_1, in395_2;
    wire c395;
    assign in395_1 = {pp41[32]};
    assign in395_2 = {pp42[31]};
    Full_Adder FA_395(s395, c395, in395_1, in395_2, pp40[33]);
    wire[0:0] s396, in396_1, in396_2;
    wire c396;
    assign in396_1 = {pp44[29]};
    assign in396_2 = {pp45[28]};
    Full_Adder FA_396(s396, c396, in396_1, in396_2, pp43[30]);
    wire[0:0] s397, in397_1, in397_2;
    wire c397;
    assign in397_1 = {pp12[62]};
    assign in397_2 = {pp13[61]};
    Full_Adder FA_397(s397, c397, in397_1, in397_2, pp11[63]);
    wire[0:0] s398, in398_1, in398_2;
    wire c398;
    assign in398_1 = {pp15[59]};
    assign in398_2 = {pp16[58]};
    Full_Adder FA_398(s398, c398, in398_1, in398_2, pp14[60]);
    wire[0:0] s399, in399_1, in399_2;
    wire c399;
    assign in399_1 = {pp18[56]};
    assign in399_2 = {pp19[55]};
    Full_Adder FA_399(s399, c399, in399_1, in399_2, pp17[57]);
    wire[0:0] s400, in400_1, in400_2;
    wire c400;
    assign in400_1 = {pp21[53]};
    assign in400_2 = {pp22[52]};
    Full_Adder FA_400(s400, c400, in400_1, in400_2, pp20[54]);
    wire[0:0] s401, in401_1, in401_2;
    wire c401;
    assign in401_1 = {pp24[50]};
    assign in401_2 = {pp25[49]};
    Full_Adder FA_401(s401, c401, in401_1, in401_2, pp23[51]);
    wire[0:0] s402, in402_1, in402_2;
    wire c402;
    assign in402_1 = {pp27[47]};
    assign in402_2 = {pp28[46]};
    Full_Adder FA_402(s402, c402, in402_1, in402_2, pp26[48]);
    wire[0:0] s403, in403_1, in403_2;
    wire c403;
    assign in403_1 = {pp30[44]};
    assign in403_2 = {pp31[43]};
    Full_Adder FA_403(s403, c403, in403_1, in403_2, pp29[45]);
    wire[0:0] s404, in404_1, in404_2;
    wire c404;
    assign in404_1 = {pp33[41]};
    assign in404_2 = {pp34[40]};
    Full_Adder FA_404(s404, c404, in404_1, in404_2, pp32[42]);
    wire[0:0] s405, in405_1, in405_2;
    wire c405;
    assign in405_1 = {pp36[38]};
    assign in405_2 = {pp37[37]};
    Full_Adder FA_405(s405, c405, in405_1, in405_2, pp35[39]);
    wire[0:0] s406, in406_1, in406_2;
    wire c406;
    assign in406_1 = {pp39[35]};
    assign in406_2 = {pp40[34]};
    Full_Adder FA_406(s406, c406, in406_1, in406_2, pp38[36]);
    wire[0:0] s407, in407_1, in407_2;
    wire c407;
    assign in407_1 = {pp42[32]};
    assign in407_2 = {pp43[31]};
    Full_Adder FA_407(s407, c407, in407_1, in407_2, pp41[33]);
    wire[0:0] s408, in408_1, in408_2;
    wire c408;
    assign in408_1 = {pp13[62]};
    assign in408_2 = {pp14[61]};
    Full_Adder FA_408(s408, c408, in408_1, in408_2, pp12[63]);
    wire[0:0] s409, in409_1, in409_2;
    wire c409;
    assign in409_1 = {pp16[59]};
    assign in409_2 = {pp17[58]};
    Full_Adder FA_409(s409, c409, in409_1, in409_2, pp15[60]);
    wire[0:0] s410, in410_1, in410_2;
    wire c410;
    assign in410_1 = {pp19[56]};
    assign in410_2 = {pp20[55]};
    Full_Adder FA_410(s410, c410, in410_1, in410_2, pp18[57]);
    wire[0:0] s411, in411_1, in411_2;
    wire c411;
    assign in411_1 = {pp22[53]};
    assign in411_2 = {pp23[52]};
    Full_Adder FA_411(s411, c411, in411_1, in411_2, pp21[54]);
    wire[0:0] s412, in412_1, in412_2;
    wire c412;
    assign in412_1 = {pp25[50]};
    assign in412_2 = {pp26[49]};
    Full_Adder FA_412(s412, c412, in412_1, in412_2, pp24[51]);
    wire[0:0] s413, in413_1, in413_2;
    wire c413;
    assign in413_1 = {pp28[47]};
    assign in413_2 = {pp29[46]};
    Full_Adder FA_413(s413, c413, in413_1, in413_2, pp27[48]);
    wire[0:0] s414, in414_1, in414_2;
    wire c414;
    assign in414_1 = {pp31[44]};
    assign in414_2 = {pp32[43]};
    Full_Adder FA_414(s414, c414, in414_1, in414_2, pp30[45]);
    wire[0:0] s415, in415_1, in415_2;
    wire c415;
    assign in415_1 = {pp34[41]};
    assign in415_2 = {pp35[40]};
    Full_Adder FA_415(s415, c415, in415_1, in415_2, pp33[42]);
    wire[0:0] s416, in416_1, in416_2;
    wire c416;
    assign in416_1 = {pp37[38]};
    assign in416_2 = {pp38[37]};
    Full_Adder FA_416(s416, c416, in416_1, in416_2, pp36[39]);
    wire[0:0] s417, in417_1, in417_2;
    wire c417;
    assign in417_1 = {pp40[35]};
    assign in417_2 = {pp41[34]};
    Full_Adder FA_417(s417, c417, in417_1, in417_2, pp39[36]);
    wire[0:0] s418, in418_1, in418_2;
    wire c418;
    assign in418_1 = {pp14[62]};
    assign in418_2 = {pp15[61]};
    Full_Adder FA_418(s418, c418, in418_1, in418_2, pp13[63]);
    wire[0:0] s419, in419_1, in419_2;
    wire c419;
    assign in419_1 = {pp17[59]};
    assign in419_2 = {pp18[58]};
    Full_Adder FA_419(s419, c419, in419_1, in419_2, pp16[60]);
    wire[0:0] s420, in420_1, in420_2;
    wire c420;
    assign in420_1 = {pp20[56]};
    assign in420_2 = {pp21[55]};
    Full_Adder FA_420(s420, c420, in420_1, in420_2, pp19[57]);
    wire[0:0] s421, in421_1, in421_2;
    wire c421;
    assign in421_1 = {pp23[53]};
    assign in421_2 = {pp24[52]};
    Full_Adder FA_421(s421, c421, in421_1, in421_2, pp22[54]);
    wire[0:0] s422, in422_1, in422_2;
    wire c422;
    assign in422_1 = {pp26[50]};
    assign in422_2 = {pp27[49]};
    Full_Adder FA_422(s422, c422, in422_1, in422_2, pp25[51]);
    wire[0:0] s423, in423_1, in423_2;
    wire c423;
    assign in423_1 = {pp29[47]};
    assign in423_2 = {pp30[46]};
    Full_Adder FA_423(s423, c423, in423_1, in423_2, pp28[48]);
    wire[0:0] s424, in424_1, in424_2;
    wire c424;
    assign in424_1 = {pp32[44]};
    assign in424_2 = {pp33[43]};
    Full_Adder FA_424(s424, c424, in424_1, in424_2, pp31[45]);
    wire[0:0] s425, in425_1, in425_2;
    wire c425;
    assign in425_1 = {pp35[41]};
    assign in425_2 = {pp36[40]};
    Full_Adder FA_425(s425, c425, in425_1, in425_2, pp34[42]);
    wire[0:0] s426, in426_1, in426_2;
    wire c426;
    assign in426_1 = {pp38[38]};
    assign in426_2 = {pp39[37]};
    Full_Adder FA_426(s426, c426, in426_1, in426_2, pp37[39]);
    wire[0:0] s427, in427_1, in427_2;
    wire c427;
    assign in427_1 = {pp15[62]};
    assign in427_2 = {pp16[61]};
    Full_Adder FA_427(s427, c427, in427_1, in427_2, pp14[63]);
    wire[0:0] s428, in428_1, in428_2;
    wire c428;
    assign in428_1 = {pp18[59]};
    assign in428_2 = {pp19[58]};
    Full_Adder FA_428(s428, c428, in428_1, in428_2, pp17[60]);
    wire[0:0] s429, in429_1, in429_2;
    wire c429;
    assign in429_1 = {pp21[56]};
    assign in429_2 = {pp22[55]};
    Full_Adder FA_429(s429, c429, in429_1, in429_2, pp20[57]);
    wire[0:0] s430, in430_1, in430_2;
    wire c430;
    assign in430_1 = {pp24[53]};
    assign in430_2 = {pp25[52]};
    Full_Adder FA_430(s430, c430, in430_1, in430_2, pp23[54]);
    wire[0:0] s431, in431_1, in431_2;
    wire c431;
    assign in431_1 = {pp27[50]};
    assign in431_2 = {pp28[49]};
    Full_Adder FA_431(s431, c431, in431_1, in431_2, pp26[51]);
    wire[0:0] s432, in432_1, in432_2;
    wire c432;
    assign in432_1 = {pp30[47]};
    assign in432_2 = {pp31[46]};
    Full_Adder FA_432(s432, c432, in432_1, in432_2, pp29[48]);
    wire[0:0] s433, in433_1, in433_2;
    wire c433;
    assign in433_1 = {pp33[44]};
    assign in433_2 = {pp34[43]};
    Full_Adder FA_433(s433, c433, in433_1, in433_2, pp32[45]);
    wire[0:0] s434, in434_1, in434_2;
    wire c434;
    assign in434_1 = {pp36[41]};
    assign in434_2 = {pp37[40]};
    Full_Adder FA_434(s434, c434, in434_1, in434_2, pp35[42]);
    wire[0:0] s435, in435_1, in435_2;
    wire c435;
    assign in435_1 = {pp16[62]};
    assign in435_2 = {pp17[61]};
    Full_Adder FA_435(s435, c435, in435_1, in435_2, pp15[63]);
    wire[0:0] s436, in436_1, in436_2;
    wire c436;
    assign in436_1 = {pp19[59]};
    assign in436_2 = {pp20[58]};
    Full_Adder FA_436(s436, c436, in436_1, in436_2, pp18[60]);
    wire[0:0] s437, in437_1, in437_2;
    wire c437;
    assign in437_1 = {pp22[56]};
    assign in437_2 = {pp23[55]};
    Full_Adder FA_437(s437, c437, in437_1, in437_2, pp21[57]);
    wire[0:0] s438, in438_1, in438_2;
    wire c438;
    assign in438_1 = {pp25[53]};
    assign in438_2 = {pp26[52]};
    Full_Adder FA_438(s438, c438, in438_1, in438_2, pp24[54]);
    wire[0:0] s439, in439_1, in439_2;
    wire c439;
    assign in439_1 = {pp28[50]};
    assign in439_2 = {pp29[49]};
    Full_Adder FA_439(s439, c439, in439_1, in439_2, pp27[51]);
    wire[0:0] s440, in440_1, in440_2;
    wire c440;
    assign in440_1 = {pp31[47]};
    assign in440_2 = {pp32[46]};
    Full_Adder FA_440(s440, c440, in440_1, in440_2, pp30[48]);
    wire[0:0] s441, in441_1, in441_2;
    wire c441;
    assign in441_1 = {pp34[44]};
    assign in441_2 = {pp35[43]};
    Full_Adder FA_441(s441, c441, in441_1, in441_2, pp33[45]);
    wire[0:0] s442, in442_1, in442_2;
    wire c442;
    assign in442_1 = {pp17[62]};
    assign in442_2 = {pp18[61]};
    Full_Adder FA_442(s442, c442, in442_1, in442_2, pp16[63]);
    wire[0:0] s443, in443_1, in443_2;
    wire c443;
    assign in443_1 = {pp20[59]};
    assign in443_2 = {pp21[58]};
    Full_Adder FA_443(s443, c443, in443_1, in443_2, pp19[60]);
    wire[0:0] s444, in444_1, in444_2;
    wire c444;
    assign in444_1 = {pp23[56]};
    assign in444_2 = {pp24[55]};
    Full_Adder FA_444(s444, c444, in444_1, in444_2, pp22[57]);
    wire[0:0] s445, in445_1, in445_2;
    wire c445;
    assign in445_1 = {pp26[53]};
    assign in445_2 = {pp27[52]};
    Full_Adder FA_445(s445, c445, in445_1, in445_2, pp25[54]);
    wire[0:0] s446, in446_1, in446_2;
    wire c446;
    assign in446_1 = {pp29[50]};
    assign in446_2 = {pp30[49]};
    Full_Adder FA_446(s446, c446, in446_1, in446_2, pp28[51]);
    wire[0:0] s447, in447_1, in447_2;
    wire c447;
    assign in447_1 = {pp32[47]};
    assign in447_2 = {pp33[46]};
    Full_Adder FA_447(s447, c447, in447_1, in447_2, pp31[48]);
    wire[0:0] s448, in448_1, in448_2;
    wire c448;
    assign in448_1 = {pp18[62]};
    assign in448_2 = {pp19[61]};
    Full_Adder FA_448(s448, c448, in448_1, in448_2, pp17[63]);
    wire[0:0] s449, in449_1, in449_2;
    wire c449;
    assign in449_1 = {pp21[59]};
    assign in449_2 = {pp22[58]};
    Full_Adder FA_449(s449, c449, in449_1, in449_2, pp20[60]);
    wire[0:0] s450, in450_1, in450_2;
    wire c450;
    assign in450_1 = {pp24[56]};
    assign in450_2 = {pp25[55]};
    Full_Adder FA_450(s450, c450, in450_1, in450_2, pp23[57]);
    wire[0:0] s451, in451_1, in451_2;
    wire c451;
    assign in451_1 = {pp27[53]};
    assign in451_2 = {pp28[52]};
    Full_Adder FA_451(s451, c451, in451_1, in451_2, pp26[54]);
    wire[0:0] s452, in452_1, in452_2;
    wire c452;
    assign in452_1 = {pp30[50]};
    assign in452_2 = {pp31[49]};
    Full_Adder FA_452(s452, c452, in452_1, in452_2, pp29[51]);
    wire[0:0] s453, in453_1, in453_2;
    wire c453;
    assign in453_1 = {pp19[62]};
    assign in453_2 = {pp20[61]};
    Full_Adder FA_453(s453, c453, in453_1, in453_2, pp18[63]);
    wire[0:0] s454, in454_1, in454_2;
    wire c454;
    assign in454_1 = {pp22[59]};
    assign in454_2 = {pp23[58]};
    Full_Adder FA_454(s454, c454, in454_1, in454_2, pp21[60]);
    wire[0:0] s455, in455_1, in455_2;
    wire c455;
    assign in455_1 = {pp25[56]};
    assign in455_2 = {pp26[55]};
    Full_Adder FA_455(s455, c455, in455_1, in455_2, pp24[57]);
    wire[0:0] s456, in456_1, in456_2;
    wire c456;
    assign in456_1 = {pp28[53]};
    assign in456_2 = {pp29[52]};
    Full_Adder FA_456(s456, c456, in456_1, in456_2, pp27[54]);
    wire[0:0] s457, in457_1, in457_2;
    wire c457;
    assign in457_1 = {pp20[62]};
    assign in457_2 = {pp21[61]};
    Full_Adder FA_457(s457, c457, in457_1, in457_2, pp19[63]);
    wire[0:0] s458, in458_1, in458_2;
    wire c458;
    assign in458_1 = {pp23[59]};
    assign in458_2 = {pp24[58]};
    Full_Adder FA_458(s458, c458, in458_1, in458_2, pp22[60]);
    wire[0:0] s459, in459_1, in459_2;
    wire c459;
    assign in459_1 = {pp26[56]};
    assign in459_2 = {pp27[55]};
    Full_Adder FA_459(s459, c459, in459_1, in459_2, pp25[57]);
    wire[0:0] s460, in460_1, in460_2;
    wire c460;
    assign in460_1 = {pp21[62]};
    assign in460_2 = {pp22[61]};
    Full_Adder FA_460(s460, c460, in460_1, in460_2, pp20[63]);
    wire[0:0] s461, in461_1, in461_2;
    wire c461;
    assign in461_1 = {pp24[59]};
    assign in461_2 = {pp25[58]};
    Full_Adder FA_461(s461, c461, in461_1, in461_2, pp23[60]);
    wire[0:0] s462, in462_1, in462_2;
    wire c462;
    assign in462_1 = {pp22[62]};
    assign in462_2 = {pp23[61]};
    Full_Adder FA_462(s462, c462, in462_1, in462_2, pp21[63]);

    /*Stage 2*/
    wire[0:0] s463, in463_1, in463_2;
    wire c463;
    assign in463_1 = {pp0[29]};
    assign in463_2 = {pp1[28]};
    Half_Adder HA_463(s463, c463, in463_1, in463_2);
    wire[0:0] s464, in464_1, in464_2;
    wire c464;
    assign in464_1 = {pp1[29]};
    assign in464_2 = {pp2[28]};
    Full_Adder FA_464(s464, c464, in464_1, in464_2, pp0[30]);
    wire[0:0] s465, in465_1, in465_2;
    wire c465;
    assign in465_1 = {pp3[27]};
    assign in465_2 = {pp4[26]};
    Half_Adder HA_465(s465, c465, in465_1, in465_2);
    wire[0:0] s466, in466_1, in466_2;
    wire c466;
    assign in466_1 = {pp1[30]};
    assign in466_2 = {pp2[29]};
    Full_Adder FA_466(s466, c466, in466_1, in466_2, pp0[31]);
    wire[0:0] s467, in467_1, in467_2;
    wire c467;
    assign in467_1 = {pp4[27]};
    assign in467_2 = {pp5[26]};
    Full_Adder FA_467(s467, c467, in467_1, in467_2, pp3[28]);
    wire[0:0] s468, in468_1, in468_2;
    wire c468;
    assign in468_1 = {pp6[25]};
    assign in468_2 = {pp7[24]};
    Half_Adder HA_468(s468, c468, in468_1, in468_2);
    wire[0:0] s469, in469_1, in469_2;
    wire c469;
    assign in469_1 = {pp1[31]};
    assign in469_2 = {pp2[30]};
    Full_Adder FA_469(s469, c469, in469_1, in469_2, pp0[32]);
    wire[0:0] s470, in470_1, in470_2;
    wire c470;
    assign in470_1 = {pp4[28]};
    assign in470_2 = {pp5[27]};
    Full_Adder FA_470(s470, c470, in470_1, in470_2, pp3[29]);
    wire[0:0] s471, in471_1, in471_2;
    wire c471;
    assign in471_1 = {pp7[25]};
    assign in471_2 = {pp8[24]};
    Full_Adder FA_471(s471, c471, in471_1, in471_2, pp6[26]);
    wire[0:0] s472, in472_1, in472_2;
    wire c472;
    assign in472_1 = {pp9[23]};
    assign in472_2 = {pp10[22]};
    Half_Adder HA_472(s472, c472, in472_1, in472_2);
    wire[0:0] s473, in473_1, in473_2;
    wire c473;
    assign in473_1 = {pp1[32]};
    assign in473_2 = {pp2[31]};
    Full_Adder FA_473(s473, c473, in473_1, in473_2, pp0[33]);
    wire[0:0] s474, in474_1, in474_2;
    wire c474;
    assign in474_1 = {pp4[29]};
    assign in474_2 = {pp5[28]};
    Full_Adder FA_474(s474, c474, in474_1, in474_2, pp3[30]);
    wire[0:0] s475, in475_1, in475_2;
    wire c475;
    assign in475_1 = {pp7[26]};
    assign in475_2 = {pp8[25]};
    Full_Adder FA_475(s475, c475, in475_1, in475_2, pp6[27]);
    wire[0:0] s476, in476_1, in476_2;
    wire c476;
    assign in476_1 = {pp10[23]};
    assign in476_2 = {pp11[22]};
    Full_Adder FA_476(s476, c476, in476_1, in476_2, pp9[24]);
    wire[0:0] s477, in477_1, in477_2;
    wire c477;
    assign in477_1 = {pp12[21]};
    assign in477_2 = {pp13[20]};
    Half_Adder HA_477(s477, c477, in477_1, in477_2);
    wire[0:0] s478, in478_1, in478_2;
    wire c478;
    assign in478_1 = {pp1[33]};
    assign in478_2 = {pp2[32]};
    Full_Adder FA_478(s478, c478, in478_1, in478_2, pp0[34]);
    wire[0:0] s479, in479_1, in479_2;
    wire c479;
    assign in479_1 = {pp4[30]};
    assign in479_2 = {pp5[29]};
    Full_Adder FA_479(s479, c479, in479_1, in479_2, pp3[31]);
    wire[0:0] s480, in480_1, in480_2;
    wire c480;
    assign in480_1 = {pp7[27]};
    assign in480_2 = {pp8[26]};
    Full_Adder FA_480(s480, c480, in480_1, in480_2, pp6[28]);
    wire[0:0] s481, in481_1, in481_2;
    wire c481;
    assign in481_1 = {pp10[24]};
    assign in481_2 = {pp11[23]};
    Full_Adder FA_481(s481, c481, in481_1, in481_2, pp9[25]);
    wire[0:0] s482, in482_1, in482_2;
    wire c482;
    assign in482_1 = {pp13[21]};
    assign in482_2 = {pp14[20]};
    Full_Adder FA_482(s482, c482, in482_1, in482_2, pp12[22]);
    wire[0:0] s483, in483_1, in483_2;
    wire c483;
    assign in483_1 = {pp15[19]};
    assign in483_2 = {pp16[18]};
    Half_Adder HA_483(s483, c483, in483_1, in483_2);
    wire[0:0] s484, in484_1, in484_2;
    wire c484;
    assign in484_1 = {pp1[34]};
    assign in484_2 = {pp2[33]};
    Full_Adder FA_484(s484, c484, in484_1, in484_2, pp0[35]);
    wire[0:0] s485, in485_1, in485_2;
    wire c485;
    assign in485_1 = {pp4[31]};
    assign in485_2 = {pp5[30]};
    Full_Adder FA_485(s485, c485, in485_1, in485_2, pp3[32]);
    wire[0:0] s486, in486_1, in486_2;
    wire c486;
    assign in486_1 = {pp7[28]};
    assign in486_2 = {pp8[27]};
    Full_Adder FA_486(s486, c486, in486_1, in486_2, pp6[29]);
    wire[0:0] s487, in487_1, in487_2;
    wire c487;
    assign in487_1 = {pp10[25]};
    assign in487_2 = {pp11[24]};
    Full_Adder FA_487(s487, c487, in487_1, in487_2, pp9[26]);
    wire[0:0] s488, in488_1, in488_2;
    wire c488;
    assign in488_1 = {pp13[22]};
    assign in488_2 = {pp14[21]};
    Full_Adder FA_488(s488, c488, in488_1, in488_2, pp12[23]);
    wire[0:0] s489, in489_1, in489_2;
    wire c489;
    assign in489_1 = {pp16[19]};
    assign in489_2 = {pp17[18]};
    Full_Adder FA_489(s489, c489, in489_1, in489_2, pp15[20]);
    wire[0:0] s490, in490_1, in490_2;
    wire c490;
    assign in490_1 = {pp18[17]};
    assign in490_2 = {pp19[16]};
    Half_Adder HA_490(s490, c490, in490_1, in490_2);
    wire[0:0] s491, in491_1, in491_2;
    wire c491;
    assign in491_1 = {pp1[35]};
    assign in491_2 = {pp2[34]};
    Full_Adder FA_491(s491, c491, in491_1, in491_2, pp0[36]);
    wire[0:0] s492, in492_1, in492_2;
    wire c492;
    assign in492_1 = {pp4[32]};
    assign in492_2 = {pp5[31]};
    Full_Adder FA_492(s492, c492, in492_1, in492_2, pp3[33]);
    wire[0:0] s493, in493_1, in493_2;
    wire c493;
    assign in493_1 = {pp7[29]};
    assign in493_2 = {pp8[28]};
    Full_Adder FA_493(s493, c493, in493_1, in493_2, pp6[30]);
    wire[0:0] s494, in494_1, in494_2;
    wire c494;
    assign in494_1 = {pp10[26]};
    assign in494_2 = {pp11[25]};
    Full_Adder FA_494(s494, c494, in494_1, in494_2, pp9[27]);
    wire[0:0] s495, in495_1, in495_2;
    wire c495;
    assign in495_1 = {pp13[23]};
    assign in495_2 = {pp14[22]};
    Full_Adder FA_495(s495, c495, in495_1, in495_2, pp12[24]);
    wire[0:0] s496, in496_1, in496_2;
    wire c496;
    assign in496_1 = {pp16[20]};
    assign in496_2 = {pp17[19]};
    Full_Adder FA_496(s496, c496, in496_1, in496_2, pp15[21]);
    wire[0:0] s497, in497_1, in497_2;
    wire c497;
    assign in497_1 = {pp19[17]};
    assign in497_2 = {pp20[16]};
    Full_Adder FA_497(s497, c497, in497_1, in497_2, pp18[18]);
    wire[0:0] s498, in498_1, in498_2;
    wire c498;
    assign in498_1 = {pp21[15]};
    assign in498_2 = {pp22[14]};
    Half_Adder HA_498(s498, c498, in498_1, in498_2);
    wire[0:0] s499, in499_1, in499_2;
    wire c499;
    assign in499_1 = {pp1[36]};
    assign in499_2 = {pp2[35]};
    Full_Adder FA_499(s499, c499, in499_1, in499_2, pp0[37]);
    wire[0:0] s500, in500_1, in500_2;
    wire c500;
    assign in500_1 = {pp4[33]};
    assign in500_2 = {pp5[32]};
    Full_Adder FA_500(s500, c500, in500_1, in500_2, pp3[34]);
    wire[0:0] s501, in501_1, in501_2;
    wire c501;
    assign in501_1 = {pp7[30]};
    assign in501_2 = {pp8[29]};
    Full_Adder FA_501(s501, c501, in501_1, in501_2, pp6[31]);
    wire[0:0] s502, in502_1, in502_2;
    wire c502;
    assign in502_1 = {pp10[27]};
    assign in502_2 = {pp11[26]};
    Full_Adder FA_502(s502, c502, in502_1, in502_2, pp9[28]);
    wire[0:0] s503, in503_1, in503_2;
    wire c503;
    assign in503_1 = {pp13[24]};
    assign in503_2 = {pp14[23]};
    Full_Adder FA_503(s503, c503, in503_1, in503_2, pp12[25]);
    wire[0:0] s504, in504_1, in504_2;
    wire c504;
    assign in504_1 = {pp16[21]};
    assign in504_2 = {pp17[20]};
    Full_Adder FA_504(s504, c504, in504_1, in504_2, pp15[22]);
    wire[0:0] s505, in505_1, in505_2;
    wire c505;
    assign in505_1 = {pp19[18]};
    assign in505_2 = {pp20[17]};
    Full_Adder FA_505(s505, c505, in505_1, in505_2, pp18[19]);
    wire[0:0] s506, in506_1, in506_2;
    wire c506;
    assign in506_1 = {pp22[15]};
    assign in506_2 = {pp23[14]};
    Full_Adder FA_506(s506, c506, in506_1, in506_2, pp21[16]);
    wire[0:0] s507, in507_1, in507_2;
    wire c507;
    assign in507_1 = {pp24[13]};
    assign in507_2 = {pp25[12]};
    Half_Adder HA_507(s507, c507, in507_1, in507_2);
    wire[0:0] s508, in508_1, in508_2;
    wire c508;
    assign in508_1 = {pp1[37]};
    assign in508_2 = {pp2[36]};
    Full_Adder FA_508(s508, c508, in508_1, in508_2, pp0[38]);
    wire[0:0] s509, in509_1, in509_2;
    wire c509;
    assign in509_1 = {pp4[34]};
    assign in509_2 = {pp5[33]};
    Full_Adder FA_509(s509, c509, in509_1, in509_2, pp3[35]);
    wire[0:0] s510, in510_1, in510_2;
    wire c510;
    assign in510_1 = {pp7[31]};
    assign in510_2 = {pp8[30]};
    Full_Adder FA_510(s510, c510, in510_1, in510_2, pp6[32]);
    wire[0:0] s511, in511_1, in511_2;
    wire c511;
    assign in511_1 = {pp10[28]};
    assign in511_2 = {pp11[27]};
    Full_Adder FA_511(s511, c511, in511_1, in511_2, pp9[29]);
    wire[0:0] s512, in512_1, in512_2;
    wire c512;
    assign in512_1 = {pp13[25]};
    assign in512_2 = {pp14[24]};
    Full_Adder FA_512(s512, c512, in512_1, in512_2, pp12[26]);
    wire[0:0] s513, in513_1, in513_2;
    wire c513;
    assign in513_1 = {pp16[22]};
    assign in513_2 = {pp17[21]};
    Full_Adder FA_513(s513, c513, in513_1, in513_2, pp15[23]);
    wire[0:0] s514, in514_1, in514_2;
    wire c514;
    assign in514_1 = {pp19[19]};
    assign in514_2 = {pp20[18]};
    Full_Adder FA_514(s514, c514, in514_1, in514_2, pp18[20]);
    wire[0:0] s515, in515_1, in515_2;
    wire c515;
    assign in515_1 = {pp22[16]};
    assign in515_2 = {pp23[15]};
    Full_Adder FA_515(s515, c515, in515_1, in515_2, pp21[17]);
    wire[0:0] s516, in516_1, in516_2;
    wire c516;
    assign in516_1 = {pp25[13]};
    assign in516_2 = {pp26[12]};
    Full_Adder FA_516(s516, c516, in516_1, in516_2, pp24[14]);
    wire[0:0] s517, in517_1, in517_2;
    wire c517;
    assign in517_1 = {pp27[11]};
    assign in517_2 = {pp28[10]};
    Half_Adder HA_517(s517, c517, in517_1, in517_2);
    wire[0:0] s518, in518_1, in518_2;
    wire c518;
    assign in518_1 = {pp1[38]};
    assign in518_2 = {pp2[37]};
    Full_Adder FA_518(s518, c518, in518_1, in518_2, pp0[39]);
    wire[0:0] s519, in519_1, in519_2;
    wire c519;
    assign in519_1 = {pp4[35]};
    assign in519_2 = {pp5[34]};
    Full_Adder FA_519(s519, c519, in519_1, in519_2, pp3[36]);
    wire[0:0] s520, in520_1, in520_2;
    wire c520;
    assign in520_1 = {pp7[32]};
    assign in520_2 = {pp8[31]};
    Full_Adder FA_520(s520, c520, in520_1, in520_2, pp6[33]);
    wire[0:0] s521, in521_1, in521_2;
    wire c521;
    assign in521_1 = {pp10[29]};
    assign in521_2 = {pp11[28]};
    Full_Adder FA_521(s521, c521, in521_1, in521_2, pp9[30]);
    wire[0:0] s522, in522_1, in522_2;
    wire c522;
    assign in522_1 = {pp13[26]};
    assign in522_2 = {pp14[25]};
    Full_Adder FA_522(s522, c522, in522_1, in522_2, pp12[27]);
    wire[0:0] s523, in523_1, in523_2;
    wire c523;
    assign in523_1 = {pp16[23]};
    assign in523_2 = {pp17[22]};
    Full_Adder FA_523(s523, c523, in523_1, in523_2, pp15[24]);
    wire[0:0] s524, in524_1, in524_2;
    wire c524;
    assign in524_1 = {pp19[20]};
    assign in524_2 = {pp20[19]};
    Full_Adder FA_524(s524, c524, in524_1, in524_2, pp18[21]);
    wire[0:0] s525, in525_1, in525_2;
    wire c525;
    assign in525_1 = {pp22[17]};
    assign in525_2 = {pp23[16]};
    Full_Adder FA_525(s525, c525, in525_1, in525_2, pp21[18]);
    wire[0:0] s526, in526_1, in526_2;
    wire c526;
    assign in526_1 = {pp25[14]};
    assign in526_2 = {pp26[13]};
    Full_Adder FA_526(s526, c526, in526_1, in526_2, pp24[15]);
    wire[0:0] s527, in527_1, in527_2;
    wire c527;
    assign in527_1 = {pp28[11]};
    assign in527_2 = {pp29[10]};
    Full_Adder FA_527(s527, c527, in527_1, in527_2, pp27[12]);
    wire[0:0] s528, in528_1, in528_2;
    wire c528;
    assign in528_1 = {pp30[9]};
    assign in528_2 = {pp31[8]};
    Half_Adder HA_528(s528, c528, in528_1, in528_2);
    wire[0:0] s529, in529_1, in529_2;
    wire c529;
    assign in529_1 = {pp1[39]};
    assign in529_2 = {pp2[38]};
    Full_Adder FA_529(s529, c529, in529_1, in529_2, pp0[40]);
    wire[0:0] s530, in530_1, in530_2;
    wire c530;
    assign in530_1 = {pp4[36]};
    assign in530_2 = {pp5[35]};
    Full_Adder FA_530(s530, c530, in530_1, in530_2, pp3[37]);
    wire[0:0] s531, in531_1, in531_2;
    wire c531;
    assign in531_1 = {pp7[33]};
    assign in531_2 = {pp8[32]};
    Full_Adder FA_531(s531, c531, in531_1, in531_2, pp6[34]);
    wire[0:0] s532, in532_1, in532_2;
    wire c532;
    assign in532_1 = {pp10[30]};
    assign in532_2 = {pp11[29]};
    Full_Adder FA_532(s532, c532, in532_1, in532_2, pp9[31]);
    wire[0:0] s533, in533_1, in533_2;
    wire c533;
    assign in533_1 = {pp13[27]};
    assign in533_2 = {pp14[26]};
    Full_Adder FA_533(s533, c533, in533_1, in533_2, pp12[28]);
    wire[0:0] s534, in534_1, in534_2;
    wire c534;
    assign in534_1 = {pp16[24]};
    assign in534_2 = {pp17[23]};
    Full_Adder FA_534(s534, c534, in534_1, in534_2, pp15[25]);
    wire[0:0] s535, in535_1, in535_2;
    wire c535;
    assign in535_1 = {pp19[21]};
    assign in535_2 = {pp20[20]};
    Full_Adder FA_535(s535, c535, in535_1, in535_2, pp18[22]);
    wire[0:0] s536, in536_1, in536_2;
    wire c536;
    assign in536_1 = {pp22[18]};
    assign in536_2 = {pp23[17]};
    Full_Adder FA_536(s536, c536, in536_1, in536_2, pp21[19]);
    wire[0:0] s537, in537_1, in537_2;
    wire c537;
    assign in537_1 = {pp25[15]};
    assign in537_2 = {pp26[14]};
    Full_Adder FA_537(s537, c537, in537_1, in537_2, pp24[16]);
    wire[0:0] s538, in538_1, in538_2;
    wire c538;
    assign in538_1 = {pp28[12]};
    assign in538_2 = {pp29[11]};
    Full_Adder FA_538(s538, c538, in538_1, in538_2, pp27[13]);
    wire[0:0] s539, in539_1, in539_2;
    wire c539;
    assign in539_1 = {pp31[9]};
    assign in539_2 = {pp32[8]};
    Full_Adder FA_539(s539, c539, in539_1, in539_2, pp30[10]);
    wire[0:0] s540, in540_1, in540_2;
    wire c540;
    assign in540_1 = {pp33[7]};
    assign in540_2 = {pp34[6]};
    Half_Adder HA_540(s540, c540, in540_1, in540_2);
    wire[0:0] s541, in541_1, in541_2;
    wire c541;
    assign in541_1 = {pp1[40]};
    assign in541_2 = {pp2[39]};
    Full_Adder FA_541(s541, c541, in541_1, in541_2, pp0[41]);
    wire[0:0] s542, in542_1, in542_2;
    wire c542;
    assign in542_1 = {pp4[37]};
    assign in542_2 = {pp5[36]};
    Full_Adder FA_542(s542, c542, in542_1, in542_2, pp3[38]);
    wire[0:0] s543, in543_1, in543_2;
    wire c543;
    assign in543_1 = {pp7[34]};
    assign in543_2 = {pp8[33]};
    Full_Adder FA_543(s543, c543, in543_1, in543_2, pp6[35]);
    wire[0:0] s544, in544_1, in544_2;
    wire c544;
    assign in544_1 = {pp10[31]};
    assign in544_2 = {pp11[30]};
    Full_Adder FA_544(s544, c544, in544_1, in544_2, pp9[32]);
    wire[0:0] s545, in545_1, in545_2;
    wire c545;
    assign in545_1 = {pp13[28]};
    assign in545_2 = {pp14[27]};
    Full_Adder FA_545(s545, c545, in545_1, in545_2, pp12[29]);
    wire[0:0] s546, in546_1, in546_2;
    wire c546;
    assign in546_1 = {pp16[25]};
    assign in546_2 = {pp17[24]};
    Full_Adder FA_546(s546, c546, in546_1, in546_2, pp15[26]);
    wire[0:0] s547, in547_1, in547_2;
    wire c547;
    assign in547_1 = {pp19[22]};
    assign in547_2 = {pp20[21]};
    Full_Adder FA_547(s547, c547, in547_1, in547_2, pp18[23]);
    wire[0:0] s548, in548_1, in548_2;
    wire c548;
    assign in548_1 = {pp22[19]};
    assign in548_2 = {pp23[18]};
    Full_Adder FA_548(s548, c548, in548_1, in548_2, pp21[20]);
    wire[0:0] s549, in549_1, in549_2;
    wire c549;
    assign in549_1 = {pp25[16]};
    assign in549_2 = {pp26[15]};
    Full_Adder FA_549(s549, c549, in549_1, in549_2, pp24[17]);
    wire[0:0] s550, in550_1, in550_2;
    wire c550;
    assign in550_1 = {pp28[13]};
    assign in550_2 = {pp29[12]};
    Full_Adder FA_550(s550, c550, in550_1, in550_2, pp27[14]);
    wire[0:0] s551, in551_1, in551_2;
    wire c551;
    assign in551_1 = {pp31[10]};
    assign in551_2 = {pp32[9]};
    Full_Adder FA_551(s551, c551, in551_1, in551_2, pp30[11]);
    wire[0:0] s552, in552_1, in552_2;
    wire c552;
    assign in552_1 = {pp34[7]};
    assign in552_2 = {pp35[6]};
    Full_Adder FA_552(s552, c552, in552_1, in552_2, pp33[8]);
    wire[0:0] s553, in553_1, in553_2;
    wire c553;
    assign in553_1 = {pp36[5]};
    assign in553_2 = {pp37[4]};
    Half_Adder HA_553(s553, c553, in553_1, in553_2);
    wire[0:0] s554, in554_1, in554_2;
    wire c554;
    assign in554_1 = {pp1[41]};
    assign in554_2 = {pp2[40]};
    Full_Adder FA_554(s554, c554, in554_1, in554_2, pp0[42]);
    wire[0:0] s555, in555_1, in555_2;
    wire c555;
    assign in555_1 = {pp4[38]};
    assign in555_2 = {pp5[37]};
    Full_Adder FA_555(s555, c555, in555_1, in555_2, pp3[39]);
    wire[0:0] s556, in556_1, in556_2;
    wire c556;
    assign in556_1 = {pp7[35]};
    assign in556_2 = {pp8[34]};
    Full_Adder FA_556(s556, c556, in556_1, in556_2, pp6[36]);
    wire[0:0] s557, in557_1, in557_2;
    wire c557;
    assign in557_1 = {pp10[32]};
    assign in557_2 = {pp11[31]};
    Full_Adder FA_557(s557, c557, in557_1, in557_2, pp9[33]);
    wire[0:0] s558, in558_1, in558_2;
    wire c558;
    assign in558_1 = {pp13[29]};
    assign in558_2 = {pp14[28]};
    Full_Adder FA_558(s558, c558, in558_1, in558_2, pp12[30]);
    wire[0:0] s559, in559_1, in559_2;
    wire c559;
    assign in559_1 = {pp16[26]};
    assign in559_2 = {pp17[25]};
    Full_Adder FA_559(s559, c559, in559_1, in559_2, pp15[27]);
    wire[0:0] s560, in560_1, in560_2;
    wire c560;
    assign in560_1 = {pp19[23]};
    assign in560_2 = {pp20[22]};
    Full_Adder FA_560(s560, c560, in560_1, in560_2, pp18[24]);
    wire[0:0] s561, in561_1, in561_2;
    wire c561;
    assign in561_1 = {pp22[20]};
    assign in561_2 = {pp23[19]};
    Full_Adder FA_561(s561, c561, in561_1, in561_2, pp21[21]);
    wire[0:0] s562, in562_1, in562_2;
    wire c562;
    assign in562_1 = {pp25[17]};
    assign in562_2 = {pp26[16]};
    Full_Adder FA_562(s562, c562, in562_1, in562_2, pp24[18]);
    wire[0:0] s563, in563_1, in563_2;
    wire c563;
    assign in563_1 = {pp28[14]};
    assign in563_2 = {pp29[13]};
    Full_Adder FA_563(s563, c563, in563_1, in563_2, pp27[15]);
    wire[0:0] s564, in564_1, in564_2;
    wire c564;
    assign in564_1 = {pp31[11]};
    assign in564_2 = {pp32[10]};
    Full_Adder FA_564(s564, c564, in564_1, in564_2, pp30[12]);
    wire[0:0] s565, in565_1, in565_2;
    wire c565;
    assign in565_1 = {pp34[8]};
    assign in565_2 = {pp35[7]};
    Full_Adder FA_565(s565, c565, in565_1, in565_2, pp33[9]);
    wire[0:0] s566, in566_1, in566_2;
    wire c566;
    assign in566_1 = {pp37[5]};
    assign in566_2 = {pp38[4]};
    Full_Adder FA_566(s566, c566, in566_1, in566_2, pp36[6]);
    wire[0:0] s567, in567_1, in567_2;
    wire c567;
    assign in567_1 = {pp39[3]};
    assign in567_2 = {pp40[2]};
    Half_Adder HA_567(s567, c567, in567_1, in567_2);
    wire[0:0] s568, in568_1, in568_2;
    wire c568;
    assign in568_1 = {pp3[40]};
    assign in568_2 = {pp4[39]};
    Full_Adder FA_568(s568, c568, in568_1, in568_2, pp2[41]);
    wire[0:0] s569, in569_1, in569_2;
    wire c569;
    assign in569_1 = {pp6[37]};
    assign in569_2 = {pp7[36]};
    Full_Adder FA_569(s569, c569, in569_1, in569_2, pp5[38]);
    wire[0:0] s570, in570_1, in570_2;
    wire c570;
    assign in570_1 = {pp9[34]};
    assign in570_2 = {pp10[33]};
    Full_Adder FA_570(s570, c570, in570_1, in570_2, pp8[35]);
    wire[0:0] s571, in571_1, in571_2;
    wire c571;
    assign in571_1 = {pp12[31]};
    assign in571_2 = {pp13[30]};
    Full_Adder FA_571(s571, c571, in571_1, in571_2, pp11[32]);
    wire[0:0] s572, in572_1, in572_2;
    wire c572;
    assign in572_1 = {pp15[28]};
    assign in572_2 = {pp16[27]};
    Full_Adder FA_572(s572, c572, in572_1, in572_2, pp14[29]);
    wire[0:0] s573, in573_1, in573_2;
    wire c573;
    assign in573_1 = {pp18[25]};
    assign in573_2 = {pp19[24]};
    Full_Adder FA_573(s573, c573, in573_1, in573_2, pp17[26]);
    wire[0:0] s574, in574_1, in574_2;
    wire c574;
    assign in574_1 = {pp21[22]};
    assign in574_2 = {pp22[21]};
    Full_Adder FA_574(s574, c574, in574_1, in574_2, pp20[23]);
    wire[0:0] s575, in575_1, in575_2;
    wire c575;
    assign in575_1 = {pp24[19]};
    assign in575_2 = {pp25[18]};
    Full_Adder FA_575(s575, c575, in575_1, in575_2, pp23[20]);
    wire[0:0] s576, in576_1, in576_2;
    wire c576;
    assign in576_1 = {pp27[16]};
    assign in576_2 = {pp28[15]};
    Full_Adder FA_576(s576, c576, in576_1, in576_2, pp26[17]);
    wire[0:0] s577, in577_1, in577_2;
    wire c577;
    assign in577_1 = {pp30[13]};
    assign in577_2 = {pp31[12]};
    Full_Adder FA_577(s577, c577, in577_1, in577_2, pp29[14]);
    wire[0:0] s578, in578_1, in578_2;
    wire c578;
    assign in578_1 = {pp33[10]};
    assign in578_2 = {pp34[9]};
    Full_Adder FA_578(s578, c578, in578_1, in578_2, pp32[11]);
    wire[0:0] s579, in579_1, in579_2;
    wire c579;
    assign in579_1 = {pp36[7]};
    assign in579_2 = {pp37[6]};
    Full_Adder FA_579(s579, c579, in579_1, in579_2, pp35[8]);
    wire[0:0] s580, in580_1, in580_2;
    wire c580;
    assign in580_1 = {pp39[4]};
    assign in580_2 = {pp40[3]};
    Full_Adder FA_580(s580, c580, in580_1, in580_2, pp38[5]);
    wire[0:0] s581, in581_1, in581_2;
    wire c581;
    assign in581_1 = {pp42[1]};
    assign in581_2 = {pp43[0]};
    Full_Adder FA_581(s581, c581, in581_1, in581_2, pp41[2]);
    wire[0:0] s582, in582_1, in582_2;
    wire c582;
    assign in582_1 = {pp6[38]};
    assign in582_2 = {pp7[37]};
    Full_Adder FA_582(s582, c582, in582_1, in582_2, pp5[39]);
    wire[0:0] s583, in583_1, in583_2;
    wire c583;
    assign in583_1 = {pp9[35]};
    assign in583_2 = {pp10[34]};
    Full_Adder FA_583(s583, c583, in583_1, in583_2, pp8[36]);
    wire[0:0] s584, in584_1, in584_2;
    wire c584;
    assign in584_1 = {pp12[32]};
    assign in584_2 = {pp13[31]};
    Full_Adder FA_584(s584, c584, in584_1, in584_2, pp11[33]);
    wire[0:0] s585, in585_1, in585_2;
    wire c585;
    assign in585_1 = {pp15[29]};
    assign in585_2 = {pp16[28]};
    Full_Adder FA_585(s585, c585, in585_1, in585_2, pp14[30]);
    wire[0:0] s586, in586_1, in586_2;
    wire c586;
    assign in586_1 = {pp18[26]};
    assign in586_2 = {pp19[25]};
    Full_Adder FA_586(s586, c586, in586_1, in586_2, pp17[27]);
    wire[0:0] s587, in587_1, in587_2;
    wire c587;
    assign in587_1 = {pp21[23]};
    assign in587_2 = {pp22[22]};
    Full_Adder FA_587(s587, c587, in587_1, in587_2, pp20[24]);
    wire[0:0] s588, in588_1, in588_2;
    wire c588;
    assign in588_1 = {pp24[20]};
    assign in588_2 = {pp25[19]};
    Full_Adder FA_588(s588, c588, in588_1, in588_2, pp23[21]);
    wire[0:0] s589, in589_1, in589_2;
    wire c589;
    assign in589_1 = {pp27[17]};
    assign in589_2 = {pp28[16]};
    Full_Adder FA_589(s589, c589, in589_1, in589_2, pp26[18]);
    wire[0:0] s590, in590_1, in590_2;
    wire c590;
    assign in590_1 = {pp30[14]};
    assign in590_2 = {pp31[13]};
    Full_Adder FA_590(s590, c590, in590_1, in590_2, pp29[15]);
    wire[0:0] s591, in591_1, in591_2;
    wire c591;
    assign in591_1 = {pp33[11]};
    assign in591_2 = {pp34[10]};
    Full_Adder FA_591(s591, c591, in591_1, in591_2, pp32[12]);
    wire[0:0] s592, in592_1, in592_2;
    wire c592;
    assign in592_1 = {pp36[8]};
    assign in592_2 = {pp37[7]};
    Full_Adder FA_592(s592, c592, in592_1, in592_2, pp35[9]);
    wire[0:0] s593, in593_1, in593_2;
    wire c593;
    assign in593_1 = {pp39[5]};
    assign in593_2 = {pp40[4]};
    Full_Adder FA_593(s593, c593, in593_1, in593_2, pp38[6]);
    wire[0:0] s594, in594_1, in594_2;
    wire c594;
    assign in594_1 = {pp42[2]};
    assign in594_2 = {pp43[1]};
    Full_Adder FA_594(s594, c594, in594_1, in594_2, pp41[3]);
    wire[0:0] s595, in595_1, in595_2;
    wire c595;
    assign in595_1 = {c1};
    assign in595_2 = {s2[0]};
    Full_Adder FA_595(s595, c595, in595_1, in595_2, pp44[0]);
    wire[0:0] s596, in596_1, in596_2;
    wire c596;
    assign in596_1 = {pp9[36]};
    assign in596_2 = {pp10[35]};
    Full_Adder FA_596(s596, c596, in596_1, in596_2, pp8[37]);
    wire[0:0] s597, in597_1, in597_2;
    wire c597;
    assign in597_1 = {pp12[33]};
    assign in597_2 = {pp13[32]};
    Full_Adder FA_597(s597, c597, in597_1, in597_2, pp11[34]);
    wire[0:0] s598, in598_1, in598_2;
    wire c598;
    assign in598_1 = {pp15[30]};
    assign in598_2 = {pp16[29]};
    Full_Adder FA_598(s598, c598, in598_1, in598_2, pp14[31]);
    wire[0:0] s599, in599_1, in599_2;
    wire c599;
    assign in599_1 = {pp18[27]};
    assign in599_2 = {pp19[26]};
    Full_Adder FA_599(s599, c599, in599_1, in599_2, pp17[28]);
    wire[0:0] s600, in600_1, in600_2;
    wire c600;
    assign in600_1 = {pp21[24]};
    assign in600_2 = {pp22[23]};
    Full_Adder FA_600(s600, c600, in600_1, in600_2, pp20[25]);
    wire[0:0] s601, in601_1, in601_2;
    wire c601;
    assign in601_1 = {pp24[21]};
    assign in601_2 = {pp25[20]};
    Full_Adder FA_601(s601, c601, in601_1, in601_2, pp23[22]);
    wire[0:0] s602, in602_1, in602_2;
    wire c602;
    assign in602_1 = {pp27[18]};
    assign in602_2 = {pp28[17]};
    Full_Adder FA_602(s602, c602, in602_1, in602_2, pp26[19]);
    wire[0:0] s603, in603_1, in603_2;
    wire c603;
    assign in603_1 = {pp30[15]};
    assign in603_2 = {pp31[14]};
    Full_Adder FA_603(s603, c603, in603_1, in603_2, pp29[16]);
    wire[0:0] s604, in604_1, in604_2;
    wire c604;
    assign in604_1 = {pp33[12]};
    assign in604_2 = {pp34[11]};
    Full_Adder FA_604(s604, c604, in604_1, in604_2, pp32[13]);
    wire[0:0] s605, in605_1, in605_2;
    wire c605;
    assign in605_1 = {pp36[9]};
    assign in605_2 = {pp37[8]};
    Full_Adder FA_605(s605, c605, in605_1, in605_2, pp35[10]);
    wire[0:0] s606, in606_1, in606_2;
    wire c606;
    assign in606_1 = {pp39[6]};
    assign in606_2 = {pp40[5]};
    Full_Adder FA_606(s606, c606, in606_1, in606_2, pp38[7]);
    wire[0:0] s607, in607_1, in607_2;
    wire c607;
    assign in607_1 = {pp42[3]};
    assign in607_2 = {pp43[2]};
    Full_Adder FA_607(s607, c607, in607_1, in607_2, pp41[4]);
    wire[0:0] s608, in608_1, in608_2;
    wire c608;
    assign in608_1 = {pp45[0]};
    assign in608_2 = {c2};
    Full_Adder FA_608(s608, c608, in608_1, in608_2, pp44[1]);
    wire[0:0] s609, in609_1, in609_2;
    wire c609;
    assign in609_1 = {s4[0]};
    assign in609_2 = {s5[0]};
    Full_Adder FA_609(s609, c609, in609_1, in609_2, c3);
    wire[0:0] s610, in610_1, in610_2;
    wire c610;
    assign in610_1 = {pp12[34]};
    assign in610_2 = {pp13[33]};
    Full_Adder FA_610(s610, c610, in610_1, in610_2, pp11[35]);
    wire[0:0] s611, in611_1, in611_2;
    wire c611;
    assign in611_1 = {pp15[31]};
    assign in611_2 = {pp16[30]};
    Full_Adder FA_611(s611, c611, in611_1, in611_2, pp14[32]);
    wire[0:0] s612, in612_1, in612_2;
    wire c612;
    assign in612_1 = {pp18[28]};
    assign in612_2 = {pp19[27]};
    Full_Adder FA_612(s612, c612, in612_1, in612_2, pp17[29]);
    wire[0:0] s613, in613_1, in613_2;
    wire c613;
    assign in613_1 = {pp21[25]};
    assign in613_2 = {pp22[24]};
    Full_Adder FA_613(s613, c613, in613_1, in613_2, pp20[26]);
    wire[0:0] s614, in614_1, in614_2;
    wire c614;
    assign in614_1 = {pp24[22]};
    assign in614_2 = {pp25[21]};
    Full_Adder FA_614(s614, c614, in614_1, in614_2, pp23[23]);
    wire[0:0] s615, in615_1, in615_2;
    wire c615;
    assign in615_1 = {pp27[19]};
    assign in615_2 = {pp28[18]};
    Full_Adder FA_615(s615, c615, in615_1, in615_2, pp26[20]);
    wire[0:0] s616, in616_1, in616_2;
    wire c616;
    assign in616_1 = {pp30[16]};
    assign in616_2 = {pp31[15]};
    Full_Adder FA_616(s616, c616, in616_1, in616_2, pp29[17]);
    wire[0:0] s617, in617_1, in617_2;
    wire c617;
    assign in617_1 = {pp33[13]};
    assign in617_2 = {pp34[12]};
    Full_Adder FA_617(s617, c617, in617_1, in617_2, pp32[14]);
    wire[0:0] s618, in618_1, in618_2;
    wire c618;
    assign in618_1 = {pp36[10]};
    assign in618_2 = {pp37[9]};
    Full_Adder FA_618(s618, c618, in618_1, in618_2, pp35[11]);
    wire[0:0] s619, in619_1, in619_2;
    wire c619;
    assign in619_1 = {pp39[7]};
    assign in619_2 = {pp40[6]};
    Full_Adder FA_619(s619, c619, in619_1, in619_2, pp38[8]);
    wire[0:0] s620, in620_1, in620_2;
    wire c620;
    assign in620_1 = {pp42[4]};
    assign in620_2 = {pp43[3]};
    Full_Adder FA_620(s620, c620, in620_1, in620_2, pp41[5]);
    wire[0:0] s621, in621_1, in621_2;
    wire c621;
    assign in621_1 = {pp45[1]};
    assign in621_2 = {pp46[0]};
    Full_Adder FA_621(s621, c621, in621_1, in621_2, pp44[2]);
    wire[0:0] s622, in622_1, in622_2;
    wire c622;
    assign in622_1 = {c5};
    assign in622_2 = {c6};
    Full_Adder FA_622(s622, c622, in622_1, in622_2, c4);
    wire[0:0] s623, in623_1, in623_2;
    wire c623;
    assign in623_1 = {s8[0]};
    assign in623_2 = {s9[0]};
    Full_Adder FA_623(s623, c623, in623_1, in623_2, s7[0]);
    wire[0:0] s624, in624_1, in624_2;
    wire c624;
    assign in624_1 = {pp15[32]};
    assign in624_2 = {pp16[31]};
    Full_Adder FA_624(s624, c624, in624_1, in624_2, pp14[33]);
    wire[0:0] s625, in625_1, in625_2;
    wire c625;
    assign in625_1 = {pp18[29]};
    assign in625_2 = {pp19[28]};
    Full_Adder FA_625(s625, c625, in625_1, in625_2, pp17[30]);
    wire[0:0] s626, in626_1, in626_2;
    wire c626;
    assign in626_1 = {pp21[26]};
    assign in626_2 = {pp22[25]};
    Full_Adder FA_626(s626, c626, in626_1, in626_2, pp20[27]);
    wire[0:0] s627, in627_1, in627_2;
    wire c627;
    assign in627_1 = {pp24[23]};
    assign in627_2 = {pp25[22]};
    Full_Adder FA_627(s627, c627, in627_1, in627_2, pp23[24]);
    wire[0:0] s628, in628_1, in628_2;
    wire c628;
    assign in628_1 = {pp27[20]};
    assign in628_2 = {pp28[19]};
    Full_Adder FA_628(s628, c628, in628_1, in628_2, pp26[21]);
    wire[0:0] s629, in629_1, in629_2;
    wire c629;
    assign in629_1 = {pp30[17]};
    assign in629_2 = {pp31[16]};
    Full_Adder FA_629(s629, c629, in629_1, in629_2, pp29[18]);
    wire[0:0] s630, in630_1, in630_2;
    wire c630;
    assign in630_1 = {pp33[14]};
    assign in630_2 = {pp34[13]};
    Full_Adder FA_630(s630, c630, in630_1, in630_2, pp32[15]);
    wire[0:0] s631, in631_1, in631_2;
    wire c631;
    assign in631_1 = {pp36[11]};
    assign in631_2 = {pp37[10]};
    Full_Adder FA_631(s631, c631, in631_1, in631_2, pp35[12]);
    wire[0:0] s632, in632_1, in632_2;
    wire c632;
    assign in632_1 = {pp39[8]};
    assign in632_2 = {pp40[7]};
    Full_Adder FA_632(s632, c632, in632_1, in632_2, pp38[9]);
    wire[0:0] s633, in633_1, in633_2;
    wire c633;
    assign in633_1 = {pp42[5]};
    assign in633_2 = {pp43[4]};
    Full_Adder FA_633(s633, c633, in633_1, in633_2, pp41[6]);
    wire[0:0] s634, in634_1, in634_2;
    wire c634;
    assign in634_1 = {pp45[2]};
    assign in634_2 = {pp46[1]};
    Full_Adder FA_634(s634, c634, in634_1, in634_2, pp44[3]);
    wire[0:0] s635, in635_1, in635_2;
    wire c635;
    assign in635_1 = {c7};
    assign in635_2 = {c8};
    Full_Adder FA_635(s635, c635, in635_1, in635_2, pp47[0]);
    wire[0:0] s636, in636_1, in636_2;
    wire c636;
    assign in636_1 = {c10};
    assign in636_2 = {s11[0]};
    Full_Adder FA_636(s636, c636, in636_1, in636_2, c9);
    wire[0:0] s637, in637_1, in637_2;
    wire c637;
    assign in637_1 = {s13[0]};
    assign in637_2 = {s14[0]};
    Full_Adder FA_637(s637, c637, in637_1, in637_2, s12[0]);
    wire[0:0] s638, in638_1, in638_2;
    wire c638;
    assign in638_1 = {pp18[30]};
    assign in638_2 = {pp19[29]};
    Full_Adder FA_638(s638, c638, in638_1, in638_2, pp17[31]);
    wire[0:0] s639, in639_1, in639_2;
    wire c639;
    assign in639_1 = {pp21[27]};
    assign in639_2 = {pp22[26]};
    Full_Adder FA_639(s639, c639, in639_1, in639_2, pp20[28]);
    wire[0:0] s640, in640_1, in640_2;
    wire c640;
    assign in640_1 = {pp24[24]};
    assign in640_2 = {pp25[23]};
    Full_Adder FA_640(s640, c640, in640_1, in640_2, pp23[25]);
    wire[0:0] s641, in641_1, in641_2;
    wire c641;
    assign in641_1 = {pp27[21]};
    assign in641_2 = {pp28[20]};
    Full_Adder FA_641(s641, c641, in641_1, in641_2, pp26[22]);
    wire[0:0] s642, in642_1, in642_2;
    wire c642;
    assign in642_1 = {pp30[18]};
    assign in642_2 = {pp31[17]};
    Full_Adder FA_642(s642, c642, in642_1, in642_2, pp29[19]);
    wire[0:0] s643, in643_1, in643_2;
    wire c643;
    assign in643_1 = {pp33[15]};
    assign in643_2 = {pp34[14]};
    Full_Adder FA_643(s643, c643, in643_1, in643_2, pp32[16]);
    wire[0:0] s644, in644_1, in644_2;
    wire c644;
    assign in644_1 = {pp36[12]};
    assign in644_2 = {pp37[11]};
    Full_Adder FA_644(s644, c644, in644_1, in644_2, pp35[13]);
    wire[0:0] s645, in645_1, in645_2;
    wire c645;
    assign in645_1 = {pp39[9]};
    assign in645_2 = {pp40[8]};
    Full_Adder FA_645(s645, c645, in645_1, in645_2, pp38[10]);
    wire[0:0] s646, in646_1, in646_2;
    wire c646;
    assign in646_1 = {pp42[6]};
    assign in646_2 = {pp43[5]};
    Full_Adder FA_646(s646, c646, in646_1, in646_2, pp41[7]);
    wire[0:0] s647, in647_1, in647_2;
    wire c647;
    assign in647_1 = {pp45[3]};
    assign in647_2 = {pp46[2]};
    Full_Adder FA_647(s647, c647, in647_1, in647_2, pp44[4]);
    wire[0:0] s648, in648_1, in648_2;
    wire c648;
    assign in648_1 = {pp48[0]};
    assign in648_2 = {c11};
    Full_Adder FA_648(s648, c648, in648_1, in648_2, pp47[1]);
    wire[0:0] s649, in649_1, in649_2;
    wire c649;
    assign in649_1 = {c13};
    assign in649_2 = {c14};
    Full_Adder FA_649(s649, c649, in649_1, in649_2, c12);
    wire[0:0] s650, in650_1, in650_2;
    wire c650;
    assign in650_1 = {s16[0]};
    assign in650_2 = {s17[0]};
    Full_Adder FA_650(s650, c650, in650_1, in650_2, c15);
    wire[0:0] s651, in651_1, in651_2;
    wire c651;
    assign in651_1 = {s19[0]};
    assign in651_2 = {s20[0]};
    Full_Adder FA_651(s651, c651, in651_1, in651_2, s18[0]);
    wire[0:0] s652, in652_1, in652_2;
    wire c652;
    assign in652_1 = {pp21[28]};
    assign in652_2 = {pp22[27]};
    Full_Adder FA_652(s652, c652, in652_1, in652_2, pp20[29]);
    wire[0:0] s653, in653_1, in653_2;
    wire c653;
    assign in653_1 = {pp24[25]};
    assign in653_2 = {pp25[24]};
    Full_Adder FA_653(s653, c653, in653_1, in653_2, pp23[26]);
    wire[0:0] s654, in654_1, in654_2;
    wire c654;
    assign in654_1 = {pp27[22]};
    assign in654_2 = {pp28[21]};
    Full_Adder FA_654(s654, c654, in654_1, in654_2, pp26[23]);
    wire[0:0] s655, in655_1, in655_2;
    wire c655;
    assign in655_1 = {pp30[19]};
    assign in655_2 = {pp31[18]};
    Full_Adder FA_655(s655, c655, in655_1, in655_2, pp29[20]);
    wire[0:0] s656, in656_1, in656_2;
    wire c656;
    assign in656_1 = {pp33[16]};
    assign in656_2 = {pp34[15]};
    Full_Adder FA_656(s656, c656, in656_1, in656_2, pp32[17]);
    wire[0:0] s657, in657_1, in657_2;
    wire c657;
    assign in657_1 = {pp36[13]};
    assign in657_2 = {pp37[12]};
    Full_Adder FA_657(s657, c657, in657_1, in657_2, pp35[14]);
    wire[0:0] s658, in658_1, in658_2;
    wire c658;
    assign in658_1 = {pp39[10]};
    assign in658_2 = {pp40[9]};
    Full_Adder FA_658(s658, c658, in658_1, in658_2, pp38[11]);
    wire[0:0] s659, in659_1, in659_2;
    wire c659;
    assign in659_1 = {pp42[7]};
    assign in659_2 = {pp43[6]};
    Full_Adder FA_659(s659, c659, in659_1, in659_2, pp41[8]);
    wire[0:0] s660, in660_1, in660_2;
    wire c660;
    assign in660_1 = {pp45[4]};
    assign in660_2 = {pp46[3]};
    Full_Adder FA_660(s660, c660, in660_1, in660_2, pp44[5]);
    wire[0:0] s661, in661_1, in661_2;
    wire c661;
    assign in661_1 = {pp48[1]};
    assign in661_2 = {pp49[0]};
    Full_Adder FA_661(s661, c661, in661_1, in661_2, pp47[2]);
    wire[0:0] s662, in662_1, in662_2;
    wire c662;
    assign in662_1 = {c17};
    assign in662_2 = {c18};
    Full_Adder FA_662(s662, c662, in662_1, in662_2, c16);
    wire[0:0] s663, in663_1, in663_2;
    wire c663;
    assign in663_1 = {c20};
    assign in663_2 = {c21};
    Full_Adder FA_663(s663, c663, in663_1, in663_2, c19);
    wire[0:0] s664, in664_1, in664_2;
    wire c664;
    assign in664_1 = {s23[0]};
    assign in664_2 = {s24[0]};
    Full_Adder FA_664(s664, c664, in664_1, in664_2, s22[0]);
    wire[0:0] s665, in665_1, in665_2;
    wire c665;
    assign in665_1 = {s26[0]};
    assign in665_2 = {s27[0]};
    Full_Adder FA_665(s665, c665, in665_1, in665_2, s25[0]);
    wire[0:0] s666, in666_1, in666_2;
    wire c666;
    assign in666_1 = {pp24[26]};
    assign in666_2 = {pp25[25]};
    Full_Adder FA_666(s666, c666, in666_1, in666_2, pp23[27]);
    wire[0:0] s667, in667_1, in667_2;
    wire c667;
    assign in667_1 = {pp27[23]};
    assign in667_2 = {pp28[22]};
    Full_Adder FA_667(s667, c667, in667_1, in667_2, pp26[24]);
    wire[0:0] s668, in668_1, in668_2;
    wire c668;
    assign in668_1 = {pp30[20]};
    assign in668_2 = {pp31[19]};
    Full_Adder FA_668(s668, c668, in668_1, in668_2, pp29[21]);
    wire[0:0] s669, in669_1, in669_2;
    wire c669;
    assign in669_1 = {pp33[17]};
    assign in669_2 = {pp34[16]};
    Full_Adder FA_669(s669, c669, in669_1, in669_2, pp32[18]);
    wire[0:0] s670, in670_1, in670_2;
    wire c670;
    assign in670_1 = {pp36[14]};
    assign in670_2 = {pp37[13]};
    Full_Adder FA_670(s670, c670, in670_1, in670_2, pp35[15]);
    wire[0:0] s671, in671_1, in671_2;
    wire c671;
    assign in671_1 = {pp39[11]};
    assign in671_2 = {pp40[10]};
    Full_Adder FA_671(s671, c671, in671_1, in671_2, pp38[12]);
    wire[0:0] s672, in672_1, in672_2;
    wire c672;
    assign in672_1 = {pp42[8]};
    assign in672_2 = {pp43[7]};
    Full_Adder FA_672(s672, c672, in672_1, in672_2, pp41[9]);
    wire[0:0] s673, in673_1, in673_2;
    wire c673;
    assign in673_1 = {pp45[5]};
    assign in673_2 = {pp46[4]};
    Full_Adder FA_673(s673, c673, in673_1, in673_2, pp44[6]);
    wire[0:0] s674, in674_1, in674_2;
    wire c674;
    assign in674_1 = {pp48[2]};
    assign in674_2 = {pp49[1]};
    Full_Adder FA_674(s674, c674, in674_1, in674_2, pp47[3]);
    wire[0:0] s675, in675_1, in675_2;
    wire c675;
    assign in675_1 = {c22};
    assign in675_2 = {c23};
    Full_Adder FA_675(s675, c675, in675_1, in675_2, pp50[0]);
    wire[0:0] s676, in676_1, in676_2;
    wire c676;
    assign in676_1 = {c25};
    assign in676_2 = {c26};
    Full_Adder FA_676(s676, c676, in676_1, in676_2, c24);
    wire[0:0] s677, in677_1, in677_2;
    wire c677;
    assign in677_1 = {c28};
    assign in677_2 = {s29[0]};
    Full_Adder FA_677(s677, c677, in677_1, in677_2, c27);
    wire[0:0] s678, in678_1, in678_2;
    wire c678;
    assign in678_1 = {s31[0]};
    assign in678_2 = {s32[0]};
    Full_Adder FA_678(s678, c678, in678_1, in678_2, s30[0]);
    wire[0:0] s679, in679_1, in679_2;
    wire c679;
    assign in679_1 = {s34[0]};
    assign in679_2 = {s35[0]};
    Full_Adder FA_679(s679, c679, in679_1, in679_2, s33[0]);
    wire[0:0] s680, in680_1, in680_2;
    wire c680;
    assign in680_1 = {pp27[24]};
    assign in680_2 = {pp28[23]};
    Full_Adder FA_680(s680, c680, in680_1, in680_2, pp26[25]);
    wire[0:0] s681, in681_1, in681_2;
    wire c681;
    assign in681_1 = {pp30[21]};
    assign in681_2 = {pp31[20]};
    Full_Adder FA_681(s681, c681, in681_1, in681_2, pp29[22]);
    wire[0:0] s682, in682_1, in682_2;
    wire c682;
    assign in682_1 = {pp33[18]};
    assign in682_2 = {pp34[17]};
    Full_Adder FA_682(s682, c682, in682_1, in682_2, pp32[19]);
    wire[0:0] s683, in683_1, in683_2;
    wire c683;
    assign in683_1 = {pp36[15]};
    assign in683_2 = {pp37[14]};
    Full_Adder FA_683(s683, c683, in683_1, in683_2, pp35[16]);
    wire[0:0] s684, in684_1, in684_2;
    wire c684;
    assign in684_1 = {pp39[12]};
    assign in684_2 = {pp40[11]};
    Full_Adder FA_684(s684, c684, in684_1, in684_2, pp38[13]);
    wire[0:0] s685, in685_1, in685_2;
    wire c685;
    assign in685_1 = {pp42[9]};
    assign in685_2 = {pp43[8]};
    Full_Adder FA_685(s685, c685, in685_1, in685_2, pp41[10]);
    wire[0:0] s686, in686_1, in686_2;
    wire c686;
    assign in686_1 = {pp45[6]};
    assign in686_2 = {pp46[5]};
    Full_Adder FA_686(s686, c686, in686_1, in686_2, pp44[7]);
    wire[0:0] s687, in687_1, in687_2;
    wire c687;
    assign in687_1 = {pp48[3]};
    assign in687_2 = {pp49[2]};
    Full_Adder FA_687(s687, c687, in687_1, in687_2, pp47[4]);
    wire[0:0] s688, in688_1, in688_2;
    wire c688;
    assign in688_1 = {pp51[0]};
    assign in688_2 = {c29};
    Full_Adder FA_688(s688, c688, in688_1, in688_2, pp50[1]);
    wire[0:0] s689, in689_1, in689_2;
    wire c689;
    assign in689_1 = {c31};
    assign in689_2 = {c32};
    Full_Adder FA_689(s689, c689, in689_1, in689_2, c30);
    wire[0:0] s690, in690_1, in690_2;
    wire c690;
    assign in690_1 = {c34};
    assign in690_2 = {c35};
    Full_Adder FA_690(s690, c690, in690_1, in690_2, c33);
    wire[0:0] s691, in691_1, in691_2;
    wire c691;
    assign in691_1 = {s37[0]};
    assign in691_2 = {s38[0]};
    Full_Adder FA_691(s691, c691, in691_1, in691_2, c36);
    wire[0:0] s692, in692_1, in692_2;
    wire c692;
    assign in692_1 = {s40[0]};
    assign in692_2 = {s41[0]};
    Full_Adder FA_692(s692, c692, in692_1, in692_2, s39[0]);
    wire[0:0] s693, in693_1, in693_2;
    wire c693;
    assign in693_1 = {s43[0]};
    assign in693_2 = {s44[0]};
    Full_Adder FA_693(s693, c693, in693_1, in693_2, s42[0]);
    wire[0:0] s694, in694_1, in694_2;
    wire c694;
    assign in694_1 = {pp30[22]};
    assign in694_2 = {pp31[21]};
    Full_Adder FA_694(s694, c694, in694_1, in694_2, pp29[23]);
    wire[0:0] s695, in695_1, in695_2;
    wire c695;
    assign in695_1 = {pp33[19]};
    assign in695_2 = {pp34[18]};
    Full_Adder FA_695(s695, c695, in695_1, in695_2, pp32[20]);
    wire[0:0] s696, in696_1, in696_2;
    wire c696;
    assign in696_1 = {pp36[16]};
    assign in696_2 = {pp37[15]};
    Full_Adder FA_696(s696, c696, in696_1, in696_2, pp35[17]);
    wire[0:0] s697, in697_1, in697_2;
    wire c697;
    assign in697_1 = {pp39[13]};
    assign in697_2 = {pp40[12]};
    Full_Adder FA_697(s697, c697, in697_1, in697_2, pp38[14]);
    wire[0:0] s698, in698_1, in698_2;
    wire c698;
    assign in698_1 = {pp42[10]};
    assign in698_2 = {pp43[9]};
    Full_Adder FA_698(s698, c698, in698_1, in698_2, pp41[11]);
    wire[0:0] s699, in699_1, in699_2;
    wire c699;
    assign in699_1 = {pp45[7]};
    assign in699_2 = {pp46[6]};
    Full_Adder FA_699(s699, c699, in699_1, in699_2, pp44[8]);
    wire[0:0] s700, in700_1, in700_2;
    wire c700;
    assign in700_1 = {pp48[4]};
    assign in700_2 = {pp49[3]};
    Full_Adder FA_700(s700, c700, in700_1, in700_2, pp47[5]);
    wire[0:0] s701, in701_1, in701_2;
    wire c701;
    assign in701_1 = {pp51[1]};
    assign in701_2 = {pp52[0]};
    Full_Adder FA_701(s701, c701, in701_1, in701_2, pp50[2]);
    wire[0:0] s702, in702_1, in702_2;
    wire c702;
    assign in702_1 = {c38};
    assign in702_2 = {c39};
    Full_Adder FA_702(s702, c702, in702_1, in702_2, c37);
    wire[0:0] s703, in703_1, in703_2;
    wire c703;
    assign in703_1 = {c41};
    assign in703_2 = {c42};
    Full_Adder FA_703(s703, c703, in703_1, in703_2, c40);
    wire[0:0] s704, in704_1, in704_2;
    wire c704;
    assign in704_1 = {c44};
    assign in704_2 = {c45};
    Full_Adder FA_704(s704, c704, in704_1, in704_2, c43);
    wire[0:0] s705, in705_1, in705_2;
    wire c705;
    assign in705_1 = {s47[0]};
    assign in705_2 = {s48[0]};
    Full_Adder FA_705(s705, c705, in705_1, in705_2, s46[0]);
    wire[0:0] s706, in706_1, in706_2;
    wire c706;
    assign in706_1 = {s50[0]};
    assign in706_2 = {s51[0]};
    Full_Adder FA_706(s706, c706, in706_1, in706_2, s49[0]);
    wire[0:0] s707, in707_1, in707_2;
    wire c707;
    assign in707_1 = {s53[0]};
    assign in707_2 = {s54[0]};
    Full_Adder FA_707(s707, c707, in707_1, in707_2, s52[0]);
    wire[0:0] s708, in708_1, in708_2;
    wire c708;
    assign in708_1 = {pp33[20]};
    assign in708_2 = {pp34[19]};
    Full_Adder FA_708(s708, c708, in708_1, in708_2, pp32[21]);
    wire[0:0] s709, in709_1, in709_2;
    wire c709;
    assign in709_1 = {pp36[17]};
    assign in709_2 = {pp37[16]};
    Full_Adder FA_709(s709, c709, in709_1, in709_2, pp35[18]);
    wire[0:0] s710, in710_1, in710_2;
    wire c710;
    assign in710_1 = {pp39[14]};
    assign in710_2 = {pp40[13]};
    Full_Adder FA_710(s710, c710, in710_1, in710_2, pp38[15]);
    wire[0:0] s711, in711_1, in711_2;
    wire c711;
    assign in711_1 = {pp42[11]};
    assign in711_2 = {pp43[10]};
    Full_Adder FA_711(s711, c711, in711_1, in711_2, pp41[12]);
    wire[0:0] s712, in712_1, in712_2;
    wire c712;
    assign in712_1 = {pp45[8]};
    assign in712_2 = {pp46[7]};
    Full_Adder FA_712(s712, c712, in712_1, in712_2, pp44[9]);
    wire[0:0] s713, in713_1, in713_2;
    wire c713;
    assign in713_1 = {pp48[5]};
    assign in713_2 = {pp49[4]};
    Full_Adder FA_713(s713, c713, in713_1, in713_2, pp47[6]);
    wire[0:0] s714, in714_1, in714_2;
    wire c714;
    assign in714_1 = {pp51[2]};
    assign in714_2 = {pp52[1]};
    Full_Adder FA_714(s714, c714, in714_1, in714_2, pp50[3]);
    wire[0:0] s715, in715_1, in715_2;
    wire c715;
    assign in715_1 = {c46};
    assign in715_2 = {c47};
    Full_Adder FA_715(s715, c715, in715_1, in715_2, pp53[0]);
    wire[0:0] s716, in716_1, in716_2;
    wire c716;
    assign in716_1 = {c49};
    assign in716_2 = {c50};
    Full_Adder FA_716(s716, c716, in716_1, in716_2, c48);
    wire[0:0] s717, in717_1, in717_2;
    wire c717;
    assign in717_1 = {c52};
    assign in717_2 = {c53};
    Full_Adder FA_717(s717, c717, in717_1, in717_2, c51);
    wire[0:0] s718, in718_1, in718_2;
    wire c718;
    assign in718_1 = {c55};
    assign in718_2 = {s56[0]};
    Full_Adder FA_718(s718, c718, in718_1, in718_2, c54);
    wire[0:0] s719, in719_1, in719_2;
    wire c719;
    assign in719_1 = {s58[0]};
    assign in719_2 = {s59[0]};
    Full_Adder FA_719(s719, c719, in719_1, in719_2, s57[0]);
    wire[0:0] s720, in720_1, in720_2;
    wire c720;
    assign in720_1 = {s61[0]};
    assign in720_2 = {s62[0]};
    Full_Adder FA_720(s720, c720, in720_1, in720_2, s60[0]);
    wire[0:0] s721, in721_1, in721_2;
    wire c721;
    assign in721_1 = {s64[0]};
    assign in721_2 = {s65[0]};
    Full_Adder FA_721(s721, c721, in721_1, in721_2, s63[0]);
    wire[0:0] s722, in722_1, in722_2;
    wire c722;
    assign in722_1 = {pp36[18]};
    assign in722_2 = {pp37[17]};
    Full_Adder FA_722(s722, c722, in722_1, in722_2, pp35[19]);
    wire[0:0] s723, in723_1, in723_2;
    wire c723;
    assign in723_1 = {pp39[15]};
    assign in723_2 = {pp40[14]};
    Full_Adder FA_723(s723, c723, in723_1, in723_2, pp38[16]);
    wire[0:0] s724, in724_1, in724_2;
    wire c724;
    assign in724_1 = {pp42[12]};
    assign in724_2 = {pp43[11]};
    Full_Adder FA_724(s724, c724, in724_1, in724_2, pp41[13]);
    wire[0:0] s725, in725_1, in725_2;
    wire c725;
    assign in725_1 = {pp45[9]};
    assign in725_2 = {pp46[8]};
    Full_Adder FA_725(s725, c725, in725_1, in725_2, pp44[10]);
    wire[0:0] s726, in726_1, in726_2;
    wire c726;
    assign in726_1 = {pp48[6]};
    assign in726_2 = {pp49[5]};
    Full_Adder FA_726(s726, c726, in726_1, in726_2, pp47[7]);
    wire[0:0] s727, in727_1, in727_2;
    wire c727;
    assign in727_1 = {pp51[3]};
    assign in727_2 = {pp52[2]};
    Full_Adder FA_727(s727, c727, in727_1, in727_2, pp50[4]);
    wire[0:0] s728, in728_1, in728_2;
    wire c728;
    assign in728_1 = {pp54[0]};
    assign in728_2 = {c56};
    Full_Adder FA_728(s728, c728, in728_1, in728_2, pp53[1]);
    wire[0:0] s729, in729_1, in729_2;
    wire c729;
    assign in729_1 = {c58};
    assign in729_2 = {c59};
    Full_Adder FA_729(s729, c729, in729_1, in729_2, c57);
    wire[0:0] s730, in730_1, in730_2;
    wire c730;
    assign in730_1 = {c61};
    assign in730_2 = {c62};
    Full_Adder FA_730(s730, c730, in730_1, in730_2, c60);
    wire[0:0] s731, in731_1, in731_2;
    wire c731;
    assign in731_1 = {c64};
    assign in731_2 = {c65};
    Full_Adder FA_731(s731, c731, in731_1, in731_2, c63);
    wire[0:0] s732, in732_1, in732_2;
    wire c732;
    assign in732_1 = {s67[0]};
    assign in732_2 = {s68[0]};
    Full_Adder FA_732(s732, c732, in732_1, in732_2, c66);
    wire[0:0] s733, in733_1, in733_2;
    wire c733;
    assign in733_1 = {s70[0]};
    assign in733_2 = {s71[0]};
    Full_Adder FA_733(s733, c733, in733_1, in733_2, s69[0]);
    wire[0:0] s734, in734_1, in734_2;
    wire c734;
    assign in734_1 = {s73[0]};
    assign in734_2 = {s74[0]};
    Full_Adder FA_734(s734, c734, in734_1, in734_2, s72[0]);
    wire[0:0] s735, in735_1, in735_2;
    wire c735;
    assign in735_1 = {s76[0]};
    assign in735_2 = {s77[0]};
    Full_Adder FA_735(s735, c735, in735_1, in735_2, s75[0]);
    wire[0:0] s736, in736_1, in736_2;
    wire c736;
    assign in736_1 = {pp39[16]};
    assign in736_2 = {pp40[15]};
    Full_Adder FA_736(s736, c736, in736_1, in736_2, pp38[17]);
    wire[0:0] s737, in737_1, in737_2;
    wire c737;
    assign in737_1 = {pp42[13]};
    assign in737_2 = {pp43[12]};
    Full_Adder FA_737(s737, c737, in737_1, in737_2, pp41[14]);
    wire[0:0] s738, in738_1, in738_2;
    wire c738;
    assign in738_1 = {pp45[10]};
    assign in738_2 = {pp46[9]};
    Full_Adder FA_738(s738, c738, in738_1, in738_2, pp44[11]);
    wire[0:0] s739, in739_1, in739_2;
    wire c739;
    assign in739_1 = {pp48[7]};
    assign in739_2 = {pp49[6]};
    Full_Adder FA_739(s739, c739, in739_1, in739_2, pp47[8]);
    wire[0:0] s740, in740_1, in740_2;
    wire c740;
    assign in740_1 = {pp51[4]};
    assign in740_2 = {pp52[3]};
    Full_Adder FA_740(s740, c740, in740_1, in740_2, pp50[5]);
    wire[0:0] s741, in741_1, in741_2;
    wire c741;
    assign in741_1 = {pp54[1]};
    assign in741_2 = {pp55[0]};
    Full_Adder FA_741(s741, c741, in741_1, in741_2, pp53[2]);
    wire[0:0] s742, in742_1, in742_2;
    wire c742;
    assign in742_1 = {c68};
    assign in742_2 = {c69};
    Full_Adder FA_742(s742, c742, in742_1, in742_2, c67);
    wire[0:0] s743, in743_1, in743_2;
    wire c743;
    assign in743_1 = {c71};
    assign in743_2 = {c72};
    Full_Adder FA_743(s743, c743, in743_1, in743_2, c70);
    wire[0:0] s744, in744_1, in744_2;
    wire c744;
    assign in744_1 = {c74};
    assign in744_2 = {c75};
    Full_Adder FA_744(s744, c744, in744_1, in744_2, c73);
    wire[0:0] s745, in745_1, in745_2;
    wire c745;
    assign in745_1 = {c77};
    assign in745_2 = {c78};
    Full_Adder FA_745(s745, c745, in745_1, in745_2, c76);
    wire[0:0] s746, in746_1, in746_2;
    wire c746;
    assign in746_1 = {s80[0]};
    assign in746_2 = {s81[0]};
    Full_Adder FA_746(s746, c746, in746_1, in746_2, s79[0]);
    wire[0:0] s747, in747_1, in747_2;
    wire c747;
    assign in747_1 = {s83[0]};
    assign in747_2 = {s84[0]};
    Full_Adder FA_747(s747, c747, in747_1, in747_2, s82[0]);
    wire[0:0] s748, in748_1, in748_2;
    wire c748;
    assign in748_1 = {s86[0]};
    assign in748_2 = {s87[0]};
    Full_Adder FA_748(s748, c748, in748_1, in748_2, s85[0]);
    wire[0:0] s749, in749_1, in749_2;
    wire c749;
    assign in749_1 = {s89[0]};
    assign in749_2 = {s90[0]};
    Full_Adder FA_749(s749, c749, in749_1, in749_2, s88[0]);
    wire[0:0] s750, in750_1, in750_2;
    wire c750;
    assign in750_1 = {pp42[14]};
    assign in750_2 = {pp43[13]};
    Full_Adder FA_750(s750, c750, in750_1, in750_2, pp41[15]);
    wire[0:0] s751, in751_1, in751_2;
    wire c751;
    assign in751_1 = {pp45[11]};
    assign in751_2 = {pp46[10]};
    Full_Adder FA_751(s751, c751, in751_1, in751_2, pp44[12]);
    wire[0:0] s752, in752_1, in752_2;
    wire c752;
    assign in752_1 = {pp48[8]};
    assign in752_2 = {pp49[7]};
    Full_Adder FA_752(s752, c752, in752_1, in752_2, pp47[9]);
    wire[0:0] s753, in753_1, in753_2;
    wire c753;
    assign in753_1 = {pp51[5]};
    assign in753_2 = {pp52[4]};
    Full_Adder FA_753(s753, c753, in753_1, in753_2, pp50[6]);
    wire[0:0] s754, in754_1, in754_2;
    wire c754;
    assign in754_1 = {pp54[2]};
    assign in754_2 = {pp55[1]};
    Full_Adder FA_754(s754, c754, in754_1, in754_2, pp53[3]);
    wire[0:0] s755, in755_1, in755_2;
    wire c755;
    assign in755_1 = {c79};
    assign in755_2 = {c80};
    Full_Adder FA_755(s755, c755, in755_1, in755_2, pp56[0]);
    wire[0:0] s756, in756_1, in756_2;
    wire c756;
    assign in756_1 = {c82};
    assign in756_2 = {c83};
    Full_Adder FA_756(s756, c756, in756_1, in756_2, c81);
    wire[0:0] s757, in757_1, in757_2;
    wire c757;
    assign in757_1 = {c85};
    assign in757_2 = {c86};
    Full_Adder FA_757(s757, c757, in757_1, in757_2, c84);
    wire[0:0] s758, in758_1, in758_2;
    wire c758;
    assign in758_1 = {c88};
    assign in758_2 = {c89};
    Full_Adder FA_758(s758, c758, in758_1, in758_2, c87);
    wire[0:0] s759, in759_1, in759_2;
    wire c759;
    assign in759_1 = {c91};
    assign in759_2 = {s92[0]};
    Full_Adder FA_759(s759, c759, in759_1, in759_2, c90);
    wire[0:0] s760, in760_1, in760_2;
    wire c760;
    assign in760_1 = {s94[0]};
    assign in760_2 = {s95[0]};
    Full_Adder FA_760(s760, c760, in760_1, in760_2, s93[0]);
    wire[0:0] s761, in761_1, in761_2;
    wire c761;
    assign in761_1 = {s97[0]};
    assign in761_2 = {s98[0]};
    Full_Adder FA_761(s761, c761, in761_1, in761_2, s96[0]);
    wire[0:0] s762, in762_1, in762_2;
    wire c762;
    assign in762_1 = {s100[0]};
    assign in762_2 = {s101[0]};
    Full_Adder FA_762(s762, c762, in762_1, in762_2, s99[0]);
    wire[0:0] s763, in763_1, in763_2;
    wire c763;
    assign in763_1 = {s103[0]};
    assign in763_2 = {s104[0]};
    Full_Adder FA_763(s763, c763, in763_1, in763_2, s102[0]);
    wire[0:0] s764, in764_1, in764_2;
    wire c764;
    assign in764_1 = {pp45[12]};
    assign in764_2 = {pp46[11]};
    Full_Adder FA_764(s764, c764, in764_1, in764_2, pp44[13]);
    wire[0:0] s765, in765_1, in765_2;
    wire c765;
    assign in765_1 = {pp48[9]};
    assign in765_2 = {pp49[8]};
    Full_Adder FA_765(s765, c765, in765_1, in765_2, pp47[10]);
    wire[0:0] s766, in766_1, in766_2;
    wire c766;
    assign in766_1 = {pp51[6]};
    assign in766_2 = {pp52[5]};
    Full_Adder FA_766(s766, c766, in766_1, in766_2, pp50[7]);
    wire[0:0] s767, in767_1, in767_2;
    wire c767;
    assign in767_1 = {pp54[3]};
    assign in767_2 = {pp55[2]};
    Full_Adder FA_767(s767, c767, in767_1, in767_2, pp53[4]);
    wire[0:0] s768, in768_1, in768_2;
    wire c768;
    assign in768_1 = {pp57[0]};
    assign in768_2 = {c92};
    Full_Adder FA_768(s768, c768, in768_1, in768_2, pp56[1]);
    wire[0:0] s769, in769_1, in769_2;
    wire c769;
    assign in769_1 = {c94};
    assign in769_2 = {c95};
    Full_Adder FA_769(s769, c769, in769_1, in769_2, c93);
    wire[0:0] s770, in770_1, in770_2;
    wire c770;
    assign in770_1 = {c97};
    assign in770_2 = {c98};
    Full_Adder FA_770(s770, c770, in770_1, in770_2, c96);
    wire[0:0] s771, in771_1, in771_2;
    wire c771;
    assign in771_1 = {c100};
    assign in771_2 = {c101};
    Full_Adder FA_771(s771, c771, in771_1, in771_2, c99);
    wire[0:0] s772, in772_1, in772_2;
    wire c772;
    assign in772_1 = {c103};
    assign in772_2 = {c104};
    Full_Adder FA_772(s772, c772, in772_1, in772_2, c102);
    wire[0:0] s773, in773_1, in773_2;
    wire c773;
    assign in773_1 = {s106[0]};
    assign in773_2 = {s107[0]};
    Full_Adder FA_773(s773, c773, in773_1, in773_2, c105);
    wire[0:0] s774, in774_1, in774_2;
    wire c774;
    assign in774_1 = {s109[0]};
    assign in774_2 = {s110[0]};
    Full_Adder FA_774(s774, c774, in774_1, in774_2, s108[0]);
    wire[0:0] s775, in775_1, in775_2;
    wire c775;
    assign in775_1 = {s112[0]};
    assign in775_2 = {s113[0]};
    Full_Adder FA_775(s775, c775, in775_1, in775_2, s111[0]);
    wire[0:0] s776, in776_1, in776_2;
    wire c776;
    assign in776_1 = {s115[0]};
    assign in776_2 = {s116[0]};
    Full_Adder FA_776(s776, c776, in776_1, in776_2, s114[0]);
    wire[0:0] s777, in777_1, in777_2;
    wire c777;
    assign in777_1 = {s118[0]};
    assign in777_2 = {s119[0]};
    Full_Adder FA_777(s777, c777, in777_1, in777_2, s117[0]);
    wire[0:0] s778, in778_1, in778_2;
    wire c778;
    assign in778_1 = {pp48[10]};
    assign in778_2 = {pp49[9]};
    Full_Adder FA_778(s778, c778, in778_1, in778_2, pp47[11]);
    wire[0:0] s779, in779_1, in779_2;
    wire c779;
    assign in779_1 = {pp51[7]};
    assign in779_2 = {pp52[6]};
    Full_Adder FA_779(s779, c779, in779_1, in779_2, pp50[8]);
    wire[0:0] s780, in780_1, in780_2;
    wire c780;
    assign in780_1 = {pp54[4]};
    assign in780_2 = {pp55[3]};
    Full_Adder FA_780(s780, c780, in780_1, in780_2, pp53[5]);
    wire[0:0] s781, in781_1, in781_2;
    wire c781;
    assign in781_1 = {pp57[1]};
    assign in781_2 = {pp58[0]};
    Full_Adder FA_781(s781, c781, in781_1, in781_2, pp56[2]);
    wire[0:0] s782, in782_1, in782_2;
    wire c782;
    assign in782_1 = {c107};
    assign in782_2 = {c108};
    Full_Adder FA_782(s782, c782, in782_1, in782_2, c106);
    wire[0:0] s783, in783_1, in783_2;
    wire c783;
    assign in783_1 = {c110};
    assign in783_2 = {c111};
    Full_Adder FA_783(s783, c783, in783_1, in783_2, c109);
    wire[0:0] s784, in784_1, in784_2;
    wire c784;
    assign in784_1 = {c113};
    assign in784_2 = {c114};
    Full_Adder FA_784(s784, c784, in784_1, in784_2, c112);
    wire[0:0] s785, in785_1, in785_2;
    wire c785;
    assign in785_1 = {c116};
    assign in785_2 = {c117};
    Full_Adder FA_785(s785, c785, in785_1, in785_2, c115);
    wire[0:0] s786, in786_1, in786_2;
    wire c786;
    assign in786_1 = {c119};
    assign in786_2 = {c120};
    Full_Adder FA_786(s786, c786, in786_1, in786_2, c118);
    wire[0:0] s787, in787_1, in787_2;
    wire c787;
    assign in787_1 = {s122[0]};
    assign in787_2 = {s123[0]};
    Full_Adder FA_787(s787, c787, in787_1, in787_2, s121[0]);
    wire[0:0] s788, in788_1, in788_2;
    wire c788;
    assign in788_1 = {s125[0]};
    assign in788_2 = {s126[0]};
    Full_Adder FA_788(s788, c788, in788_1, in788_2, s124[0]);
    wire[0:0] s789, in789_1, in789_2;
    wire c789;
    assign in789_1 = {s128[0]};
    assign in789_2 = {s129[0]};
    Full_Adder FA_789(s789, c789, in789_1, in789_2, s127[0]);
    wire[0:0] s790, in790_1, in790_2;
    wire c790;
    assign in790_1 = {s131[0]};
    assign in790_2 = {s132[0]};
    Full_Adder FA_790(s790, c790, in790_1, in790_2, s130[0]);
    wire[0:0] s791, in791_1, in791_2;
    wire c791;
    assign in791_1 = {s134[0]};
    assign in791_2 = {s135[0]};
    Full_Adder FA_791(s791, c791, in791_1, in791_2, s133[0]);
    wire[0:0] s792, in792_1, in792_2;
    wire c792;
    assign in792_1 = {pp51[8]};
    assign in792_2 = {pp52[7]};
    Full_Adder FA_792(s792, c792, in792_1, in792_2, pp50[9]);
    wire[0:0] s793, in793_1, in793_2;
    wire c793;
    assign in793_1 = {pp54[5]};
    assign in793_2 = {pp55[4]};
    Full_Adder FA_793(s793, c793, in793_1, in793_2, pp53[6]);
    wire[0:0] s794, in794_1, in794_2;
    wire c794;
    assign in794_1 = {pp57[2]};
    assign in794_2 = {pp58[1]};
    Full_Adder FA_794(s794, c794, in794_1, in794_2, pp56[3]);
    wire[0:0] s795, in795_1, in795_2;
    wire c795;
    assign in795_1 = {c121};
    assign in795_2 = {c122};
    Full_Adder FA_795(s795, c795, in795_1, in795_2, pp59[0]);
    wire[0:0] s796, in796_1, in796_2;
    wire c796;
    assign in796_1 = {c124};
    assign in796_2 = {c125};
    Full_Adder FA_796(s796, c796, in796_1, in796_2, c123);
    wire[0:0] s797, in797_1, in797_2;
    wire c797;
    assign in797_1 = {c127};
    assign in797_2 = {c128};
    Full_Adder FA_797(s797, c797, in797_1, in797_2, c126);
    wire[0:0] s798, in798_1, in798_2;
    wire c798;
    assign in798_1 = {c130};
    assign in798_2 = {c131};
    Full_Adder FA_798(s798, c798, in798_1, in798_2, c129);
    wire[0:0] s799, in799_1, in799_2;
    wire c799;
    assign in799_1 = {c133};
    assign in799_2 = {c134};
    Full_Adder FA_799(s799, c799, in799_1, in799_2, c132);
    wire[0:0] s800, in800_1, in800_2;
    wire c800;
    assign in800_1 = {c136};
    assign in800_2 = {s137[0]};
    Full_Adder FA_800(s800, c800, in800_1, in800_2, c135);
    wire[0:0] s801, in801_1, in801_2;
    wire c801;
    assign in801_1 = {s139[0]};
    assign in801_2 = {s140[0]};
    Full_Adder FA_801(s801, c801, in801_1, in801_2, s138[0]);
    wire[0:0] s802, in802_1, in802_2;
    wire c802;
    assign in802_1 = {s142[0]};
    assign in802_2 = {s143[0]};
    Full_Adder FA_802(s802, c802, in802_1, in802_2, s141[0]);
    wire[0:0] s803, in803_1, in803_2;
    wire c803;
    assign in803_1 = {s145[0]};
    assign in803_2 = {s146[0]};
    Full_Adder FA_803(s803, c803, in803_1, in803_2, s144[0]);
    wire[0:0] s804, in804_1, in804_2;
    wire c804;
    assign in804_1 = {s148[0]};
    assign in804_2 = {s149[0]};
    Full_Adder FA_804(s804, c804, in804_1, in804_2, s147[0]);
    wire[0:0] s805, in805_1, in805_2;
    wire c805;
    assign in805_1 = {s151[0]};
    assign in805_2 = {s152[0]};
    Full_Adder FA_805(s805, c805, in805_1, in805_2, s150[0]);
    wire[0:0] s806, in806_1, in806_2;
    wire c806;
    assign in806_1 = {pp54[6]};
    assign in806_2 = {pp55[5]};
    Full_Adder FA_806(s806, c806, in806_1, in806_2, pp53[7]);
    wire[0:0] s807, in807_1, in807_2;
    wire c807;
    assign in807_1 = {pp57[3]};
    assign in807_2 = {pp58[2]};
    Full_Adder FA_807(s807, c807, in807_1, in807_2, pp56[4]);
    wire[0:0] s808, in808_1, in808_2;
    wire c808;
    assign in808_1 = {pp60[0]};
    assign in808_2 = {c137};
    Full_Adder FA_808(s808, c808, in808_1, in808_2, pp59[1]);
    wire[0:0] s809, in809_1, in809_2;
    wire c809;
    assign in809_1 = {c139};
    assign in809_2 = {c140};
    Full_Adder FA_809(s809, c809, in809_1, in809_2, c138);
    wire[0:0] s810, in810_1, in810_2;
    wire c810;
    assign in810_1 = {c142};
    assign in810_2 = {c143};
    Full_Adder FA_810(s810, c810, in810_1, in810_2, c141);
    wire[0:0] s811, in811_1, in811_2;
    wire c811;
    assign in811_1 = {c145};
    assign in811_2 = {c146};
    Full_Adder FA_811(s811, c811, in811_1, in811_2, c144);
    wire[0:0] s812, in812_1, in812_2;
    wire c812;
    assign in812_1 = {c148};
    assign in812_2 = {c149};
    Full_Adder FA_812(s812, c812, in812_1, in812_2, c147);
    wire[0:0] s813, in813_1, in813_2;
    wire c813;
    assign in813_1 = {c151};
    assign in813_2 = {c152};
    Full_Adder FA_813(s813, c813, in813_1, in813_2, c150);
    wire[0:0] s814, in814_1, in814_2;
    wire c814;
    assign in814_1 = {s154[0]};
    assign in814_2 = {s155[0]};
    Full_Adder FA_814(s814, c814, in814_1, in814_2, c153);
    wire[0:0] s815, in815_1, in815_2;
    wire c815;
    assign in815_1 = {s157[0]};
    assign in815_2 = {s158[0]};
    Full_Adder FA_815(s815, c815, in815_1, in815_2, s156[0]);
    wire[0:0] s816, in816_1, in816_2;
    wire c816;
    assign in816_1 = {s160[0]};
    assign in816_2 = {s161[0]};
    Full_Adder FA_816(s816, c816, in816_1, in816_2, s159[0]);
    wire[0:0] s817, in817_1, in817_2;
    wire c817;
    assign in817_1 = {s163[0]};
    assign in817_2 = {s164[0]};
    Full_Adder FA_817(s817, c817, in817_1, in817_2, s162[0]);
    wire[0:0] s818, in818_1, in818_2;
    wire c818;
    assign in818_1 = {s166[0]};
    assign in818_2 = {s167[0]};
    Full_Adder FA_818(s818, c818, in818_1, in818_2, s165[0]);
    wire[0:0] s819, in819_1, in819_2;
    wire c819;
    assign in819_1 = {s169[0]};
    assign in819_2 = {s170[0]};
    Full_Adder FA_819(s819, c819, in819_1, in819_2, s168[0]);
    wire[0:0] s820, in820_1, in820_2;
    wire c820;
    assign in820_1 = {pp57[4]};
    assign in820_2 = {pp58[3]};
    Full_Adder FA_820(s820, c820, in820_1, in820_2, pp56[5]);
    wire[0:0] s821, in821_1, in821_2;
    wire c821;
    assign in821_1 = {pp60[1]};
    assign in821_2 = {pp61[0]};
    Full_Adder FA_821(s821, c821, in821_1, in821_2, pp59[2]);
    wire[0:0] s822, in822_1, in822_2;
    wire c822;
    assign in822_1 = {c155};
    assign in822_2 = {c156};
    Full_Adder FA_822(s822, c822, in822_1, in822_2, c154);
    wire[0:0] s823, in823_1, in823_2;
    wire c823;
    assign in823_1 = {c158};
    assign in823_2 = {c159};
    Full_Adder FA_823(s823, c823, in823_1, in823_2, c157);
    wire[0:0] s824, in824_1, in824_2;
    wire c824;
    assign in824_1 = {c161};
    assign in824_2 = {c162};
    Full_Adder FA_824(s824, c824, in824_1, in824_2, c160);
    wire[0:0] s825, in825_1, in825_2;
    wire c825;
    assign in825_1 = {c164};
    assign in825_2 = {c165};
    Full_Adder FA_825(s825, c825, in825_1, in825_2, c163);
    wire[0:0] s826, in826_1, in826_2;
    wire c826;
    assign in826_1 = {c167};
    assign in826_2 = {c168};
    Full_Adder FA_826(s826, c826, in826_1, in826_2, c166);
    wire[0:0] s827, in827_1, in827_2;
    wire c827;
    assign in827_1 = {c170};
    assign in827_2 = {c171};
    Full_Adder FA_827(s827, c827, in827_1, in827_2, c169);
    wire[0:0] s828, in828_1, in828_2;
    wire c828;
    assign in828_1 = {s173[0]};
    assign in828_2 = {s174[0]};
    Full_Adder FA_828(s828, c828, in828_1, in828_2, s172[0]);
    wire[0:0] s829, in829_1, in829_2;
    wire c829;
    assign in829_1 = {s176[0]};
    assign in829_2 = {s177[0]};
    Full_Adder FA_829(s829, c829, in829_1, in829_2, s175[0]);
    wire[0:0] s830, in830_1, in830_2;
    wire c830;
    assign in830_1 = {s179[0]};
    assign in830_2 = {s180[0]};
    Full_Adder FA_830(s830, c830, in830_1, in830_2, s178[0]);
    wire[0:0] s831, in831_1, in831_2;
    wire c831;
    assign in831_1 = {s182[0]};
    assign in831_2 = {s183[0]};
    Full_Adder FA_831(s831, c831, in831_1, in831_2, s181[0]);
    wire[0:0] s832, in832_1, in832_2;
    wire c832;
    assign in832_1 = {s185[0]};
    assign in832_2 = {s186[0]};
    Full_Adder FA_832(s832, c832, in832_1, in832_2, s184[0]);
    wire[0:0] s833, in833_1, in833_2;
    wire c833;
    assign in833_1 = {s188[0]};
    assign in833_2 = {s189[0]};
    Full_Adder FA_833(s833, c833, in833_1, in833_2, s187[0]);
    wire[0:0] s834, in834_1, in834_2;
    wire c834;
    assign in834_1 = {pp60[2]};
    assign in834_2 = {pp61[1]};
    Full_Adder FA_834(s834, c834, in834_1, in834_2, pp59[3]);
    wire[0:0] s835, in835_1, in835_2;
    wire c835;
    assign in835_1 = {c172};
    assign in835_2 = {c173};
    Full_Adder FA_835(s835, c835, in835_1, in835_2, pp62[0]);
    wire[0:0] s836, in836_1, in836_2;
    wire c836;
    assign in836_1 = {c175};
    assign in836_2 = {c176};
    Full_Adder FA_836(s836, c836, in836_1, in836_2, c174);
    wire[0:0] s837, in837_1, in837_2;
    wire c837;
    assign in837_1 = {c178};
    assign in837_2 = {c179};
    Full_Adder FA_837(s837, c837, in837_1, in837_2, c177);
    wire[0:0] s838, in838_1, in838_2;
    wire c838;
    assign in838_1 = {c181};
    assign in838_2 = {c182};
    Full_Adder FA_838(s838, c838, in838_1, in838_2, c180);
    wire[0:0] s839, in839_1, in839_2;
    wire c839;
    assign in839_1 = {c184};
    assign in839_2 = {c185};
    Full_Adder FA_839(s839, c839, in839_1, in839_2, c183);
    wire[0:0] s840, in840_1, in840_2;
    wire c840;
    assign in840_1 = {c187};
    assign in840_2 = {c188};
    Full_Adder FA_840(s840, c840, in840_1, in840_2, c186);
    wire[0:0] s841, in841_1, in841_2;
    wire c841;
    assign in841_1 = {c190};
    assign in841_2 = {s191[0]};
    Full_Adder FA_841(s841, c841, in841_1, in841_2, c189);
    wire[0:0] s842, in842_1, in842_2;
    wire c842;
    assign in842_1 = {s193[0]};
    assign in842_2 = {s194[0]};
    Full_Adder FA_842(s842, c842, in842_1, in842_2, s192[0]);
    wire[0:0] s843, in843_1, in843_2;
    wire c843;
    assign in843_1 = {s196[0]};
    assign in843_2 = {s197[0]};
    Full_Adder FA_843(s843, c843, in843_1, in843_2, s195[0]);
    wire[0:0] s844, in844_1, in844_2;
    wire c844;
    assign in844_1 = {s199[0]};
    assign in844_2 = {s200[0]};
    Full_Adder FA_844(s844, c844, in844_1, in844_2, s198[0]);
    wire[0:0] s845, in845_1, in845_2;
    wire c845;
    assign in845_1 = {s202[0]};
    assign in845_2 = {s203[0]};
    Full_Adder FA_845(s845, c845, in845_1, in845_2, s201[0]);
    wire[0:0] s846, in846_1, in846_2;
    wire c846;
    assign in846_1 = {s205[0]};
    assign in846_2 = {s206[0]};
    Full_Adder FA_846(s846, c846, in846_1, in846_2, s204[0]);
    wire[0:0] s847, in847_1, in847_2;
    wire c847;
    assign in847_1 = {s208[0]};
    assign in847_2 = {s209[0]};
    Full_Adder FA_847(s847, c847, in847_1, in847_2, s207[0]);
    wire[0:0] s848, in848_1, in848_2;
    wire c848;
    assign in848_1 = {pp63[0]};
    assign in848_2 = {c191};
    Full_Adder FA_848(s848, c848, in848_1, in848_2, pp62[1]);
    wire[0:0] s849, in849_1, in849_2;
    wire c849;
    assign in849_1 = {c193};
    assign in849_2 = {c194};
    Full_Adder FA_849(s849, c849, in849_1, in849_2, c192);
    wire[0:0] s850, in850_1, in850_2;
    wire c850;
    assign in850_1 = {c196};
    assign in850_2 = {c197};
    Full_Adder FA_850(s850, c850, in850_1, in850_2, c195);
    wire[0:0] s851, in851_1, in851_2;
    wire c851;
    assign in851_1 = {c199};
    assign in851_2 = {c200};
    Full_Adder FA_851(s851, c851, in851_1, in851_2, c198);
    wire[0:0] s852, in852_1, in852_2;
    wire c852;
    assign in852_1 = {c202};
    assign in852_2 = {c203};
    Full_Adder FA_852(s852, c852, in852_1, in852_2, c201);
    wire[0:0] s853, in853_1, in853_2;
    wire c853;
    assign in853_1 = {c205};
    assign in853_2 = {c206};
    Full_Adder FA_853(s853, c853, in853_1, in853_2, c204);
    wire[0:0] s854, in854_1, in854_2;
    wire c854;
    assign in854_1 = {c208};
    assign in854_2 = {c209};
    Full_Adder FA_854(s854, c854, in854_1, in854_2, c207);
    wire[0:0] s855, in855_1, in855_2;
    wire c855;
    assign in855_1 = {s211[0]};
    assign in855_2 = {s212[0]};
    Full_Adder FA_855(s855, c855, in855_1, in855_2, c210);
    wire[0:0] s856, in856_1, in856_2;
    wire c856;
    assign in856_1 = {s214[0]};
    assign in856_2 = {s215[0]};
    Full_Adder FA_856(s856, c856, in856_1, in856_2, s213[0]);
    wire[0:0] s857, in857_1, in857_2;
    wire c857;
    assign in857_1 = {s217[0]};
    assign in857_2 = {s218[0]};
    Full_Adder FA_857(s857, c857, in857_1, in857_2, s216[0]);
    wire[0:0] s858, in858_1, in858_2;
    wire c858;
    assign in858_1 = {s220[0]};
    assign in858_2 = {s221[0]};
    Full_Adder FA_858(s858, c858, in858_1, in858_2, s219[0]);
    wire[0:0] s859, in859_1, in859_2;
    wire c859;
    assign in859_1 = {s223[0]};
    assign in859_2 = {s224[0]};
    Full_Adder FA_859(s859, c859, in859_1, in859_2, s222[0]);
    wire[0:0] s860, in860_1, in860_2;
    wire c860;
    assign in860_1 = {s226[0]};
    assign in860_2 = {s227[0]};
    Full_Adder FA_860(s860, c860, in860_1, in860_2, s225[0]);
    wire[0:0] s861, in861_1, in861_2;
    wire c861;
    assign in861_1 = {s229[0]};
    assign in861_2 = {s230[0]};
    Full_Adder FA_861(s861, c861, in861_1, in861_2, s228[0]);
    wire[0:0] s862, in862_1, in862_2;
    wire c862;
    assign in862_1 = {c211};
    assign in862_2 = {c212};
    Full_Adder FA_862(s862, c862, in862_1, in862_2, pp63[1]);
    wire[0:0] s863, in863_1, in863_2;
    wire c863;
    assign in863_1 = {c214};
    assign in863_2 = {c215};
    Full_Adder FA_863(s863, c863, in863_1, in863_2, c213);
    wire[0:0] s864, in864_1, in864_2;
    wire c864;
    assign in864_1 = {c217};
    assign in864_2 = {c218};
    Full_Adder FA_864(s864, c864, in864_1, in864_2, c216);
    wire[0:0] s865, in865_1, in865_2;
    wire c865;
    assign in865_1 = {c220};
    assign in865_2 = {c221};
    Full_Adder FA_865(s865, c865, in865_1, in865_2, c219);
    wire[0:0] s866, in866_1, in866_2;
    wire c866;
    assign in866_1 = {c223};
    assign in866_2 = {c224};
    Full_Adder FA_866(s866, c866, in866_1, in866_2, c222);
    wire[0:0] s867, in867_1, in867_2;
    wire c867;
    assign in867_1 = {c226};
    assign in867_2 = {c227};
    Full_Adder FA_867(s867, c867, in867_1, in867_2, c225);
    wire[0:0] s868, in868_1, in868_2;
    wire c868;
    assign in868_1 = {c229};
    assign in868_2 = {c230};
    Full_Adder FA_868(s868, c868, in868_1, in868_2, c228);
    wire[0:0] s869, in869_1, in869_2;
    wire c869;
    assign in869_1 = {s232[0]};
    assign in869_2 = {s233[0]};
    Full_Adder FA_869(s869, c869, in869_1, in869_2, c231);
    wire[0:0] s870, in870_1, in870_2;
    wire c870;
    assign in870_1 = {s235[0]};
    assign in870_2 = {s236[0]};
    Full_Adder FA_870(s870, c870, in870_1, in870_2, s234[0]);
    wire[0:0] s871, in871_1, in871_2;
    wire c871;
    assign in871_1 = {s238[0]};
    assign in871_2 = {s239[0]};
    Full_Adder FA_871(s871, c871, in871_1, in871_2, s237[0]);
    wire[0:0] s872, in872_1, in872_2;
    wire c872;
    assign in872_1 = {s241[0]};
    assign in872_2 = {s242[0]};
    Full_Adder FA_872(s872, c872, in872_1, in872_2, s240[0]);
    wire[0:0] s873, in873_1, in873_2;
    wire c873;
    assign in873_1 = {s244[0]};
    assign in873_2 = {s245[0]};
    Full_Adder FA_873(s873, c873, in873_1, in873_2, s243[0]);
    wire[0:0] s874, in874_1, in874_2;
    wire c874;
    assign in874_1 = {s247[0]};
    assign in874_2 = {s248[0]};
    Full_Adder FA_874(s874, c874, in874_1, in874_2, s246[0]);
    wire[0:0] s875, in875_1, in875_2;
    wire c875;
    assign in875_1 = {s250[0]};
    assign in875_2 = {s251[0]};
    Full_Adder FA_875(s875, c875, in875_1, in875_2, s249[0]);
    wire[0:0] s876, in876_1, in876_2;
    wire c876;
    assign in876_1 = {pp63[2]};
    assign in876_2 = {c232};
    Full_Adder FA_876(s876, c876, in876_1, in876_2, pp62[3]);
    wire[0:0] s877, in877_1, in877_2;
    wire c877;
    assign in877_1 = {c234};
    assign in877_2 = {c235};
    Full_Adder FA_877(s877, c877, in877_1, in877_2, c233);
    wire[0:0] s878, in878_1, in878_2;
    wire c878;
    assign in878_1 = {c237};
    assign in878_2 = {c238};
    Full_Adder FA_878(s878, c878, in878_1, in878_2, c236);
    wire[0:0] s879, in879_1, in879_2;
    wire c879;
    assign in879_1 = {c240};
    assign in879_2 = {c241};
    Full_Adder FA_879(s879, c879, in879_1, in879_2, c239);
    wire[0:0] s880, in880_1, in880_2;
    wire c880;
    assign in880_1 = {c243};
    assign in880_2 = {c244};
    Full_Adder FA_880(s880, c880, in880_1, in880_2, c242);
    wire[0:0] s881, in881_1, in881_2;
    wire c881;
    assign in881_1 = {c246};
    assign in881_2 = {c247};
    Full_Adder FA_881(s881, c881, in881_1, in881_2, c245);
    wire[0:0] s882, in882_1, in882_2;
    wire c882;
    assign in882_1 = {c249};
    assign in882_2 = {c250};
    Full_Adder FA_882(s882, c882, in882_1, in882_2, c248);
    wire[0:0] s883, in883_1, in883_2;
    wire c883;
    assign in883_1 = {c252};
    assign in883_2 = {s253[0]};
    Full_Adder FA_883(s883, c883, in883_1, in883_2, c251);
    wire[0:0] s884, in884_1, in884_2;
    wire c884;
    assign in884_1 = {s255[0]};
    assign in884_2 = {s256[0]};
    Full_Adder FA_884(s884, c884, in884_1, in884_2, s254[0]);
    wire[0:0] s885, in885_1, in885_2;
    wire c885;
    assign in885_1 = {s258[0]};
    assign in885_2 = {s259[0]};
    Full_Adder FA_885(s885, c885, in885_1, in885_2, s257[0]);
    wire[0:0] s886, in886_1, in886_2;
    wire c886;
    assign in886_1 = {s261[0]};
    assign in886_2 = {s262[0]};
    Full_Adder FA_886(s886, c886, in886_1, in886_2, s260[0]);
    wire[0:0] s887, in887_1, in887_2;
    wire c887;
    assign in887_1 = {s264[0]};
    assign in887_2 = {s265[0]};
    Full_Adder FA_887(s887, c887, in887_1, in887_2, s263[0]);
    wire[0:0] s888, in888_1, in888_2;
    wire c888;
    assign in888_1 = {s267[0]};
    assign in888_2 = {s268[0]};
    Full_Adder FA_888(s888, c888, in888_1, in888_2, s266[0]);
    wire[0:0] s889, in889_1, in889_2;
    wire c889;
    assign in889_1 = {s270[0]};
    assign in889_2 = {s271[0]};
    Full_Adder FA_889(s889, c889, in889_1, in889_2, s269[0]);
    wire[0:0] s890, in890_1, in890_2;
    wire c890;
    assign in890_1 = {pp61[5]};
    assign in890_2 = {pp62[4]};
    Full_Adder FA_890(s890, c890, in890_1, in890_2, pp60[6]);
    wire[0:0] s891, in891_1, in891_2;
    wire c891;
    assign in891_1 = {c253};
    assign in891_2 = {c254};
    Full_Adder FA_891(s891, c891, in891_1, in891_2, pp63[3]);
    wire[0:0] s892, in892_1, in892_2;
    wire c892;
    assign in892_1 = {c256};
    assign in892_2 = {c257};
    Full_Adder FA_892(s892, c892, in892_1, in892_2, c255);
    wire[0:0] s893, in893_1, in893_2;
    wire c893;
    assign in893_1 = {c259};
    assign in893_2 = {c260};
    Full_Adder FA_893(s893, c893, in893_1, in893_2, c258);
    wire[0:0] s894, in894_1, in894_2;
    wire c894;
    assign in894_1 = {c262};
    assign in894_2 = {c263};
    Full_Adder FA_894(s894, c894, in894_1, in894_2, c261);
    wire[0:0] s895, in895_1, in895_2;
    wire c895;
    assign in895_1 = {c265};
    assign in895_2 = {c266};
    Full_Adder FA_895(s895, c895, in895_1, in895_2, c264);
    wire[0:0] s896, in896_1, in896_2;
    wire c896;
    assign in896_1 = {c268};
    assign in896_2 = {c269};
    Full_Adder FA_896(s896, c896, in896_1, in896_2, c267);
    wire[0:0] s897, in897_1, in897_2;
    wire c897;
    assign in897_1 = {c271};
    assign in897_2 = {c272};
    Full_Adder FA_897(s897, c897, in897_1, in897_2, c270);
    wire[0:0] s898, in898_1, in898_2;
    wire c898;
    assign in898_1 = {s274[0]};
    assign in898_2 = {s275[0]};
    Full_Adder FA_898(s898, c898, in898_1, in898_2, s273[0]);
    wire[0:0] s899, in899_1, in899_2;
    wire c899;
    assign in899_1 = {s277[0]};
    assign in899_2 = {s278[0]};
    Full_Adder FA_899(s899, c899, in899_1, in899_2, s276[0]);
    wire[0:0] s900, in900_1, in900_2;
    wire c900;
    assign in900_1 = {s280[0]};
    assign in900_2 = {s281[0]};
    Full_Adder FA_900(s900, c900, in900_1, in900_2, s279[0]);
    wire[0:0] s901, in901_1, in901_2;
    wire c901;
    assign in901_1 = {s283[0]};
    assign in901_2 = {s284[0]};
    Full_Adder FA_901(s901, c901, in901_1, in901_2, s282[0]);
    wire[0:0] s902, in902_1, in902_2;
    wire c902;
    assign in902_1 = {s286[0]};
    assign in902_2 = {s287[0]};
    Full_Adder FA_902(s902, c902, in902_1, in902_2, s285[0]);
    wire[0:0] s903, in903_1, in903_2;
    wire c903;
    assign in903_1 = {s289[0]};
    assign in903_2 = {s290[0]};
    Full_Adder FA_903(s903, c903, in903_1, in903_2, s288[0]);
    wire[0:0] s904, in904_1, in904_2;
    wire c904;
    assign in904_1 = {pp59[8]};
    assign in904_2 = {pp60[7]};
    Full_Adder FA_904(s904, c904, in904_1, in904_2, pp58[9]);
    wire[0:0] s905, in905_1, in905_2;
    wire c905;
    assign in905_1 = {pp62[5]};
    assign in905_2 = {pp63[4]};
    Full_Adder FA_905(s905, c905, in905_1, in905_2, pp61[6]);
    wire[0:0] s906, in906_1, in906_2;
    wire c906;
    assign in906_1 = {c274};
    assign in906_2 = {c275};
    Full_Adder FA_906(s906, c906, in906_1, in906_2, c273);
    wire[0:0] s907, in907_1, in907_2;
    wire c907;
    assign in907_1 = {c277};
    assign in907_2 = {c278};
    Full_Adder FA_907(s907, c907, in907_1, in907_2, c276);
    wire[0:0] s908, in908_1, in908_2;
    wire c908;
    assign in908_1 = {c280};
    assign in908_2 = {c281};
    Full_Adder FA_908(s908, c908, in908_1, in908_2, c279);
    wire[0:0] s909, in909_1, in909_2;
    wire c909;
    assign in909_1 = {c283};
    assign in909_2 = {c284};
    Full_Adder FA_909(s909, c909, in909_1, in909_2, c282);
    wire[0:0] s910, in910_1, in910_2;
    wire c910;
    assign in910_1 = {c286};
    assign in910_2 = {c287};
    Full_Adder FA_910(s910, c910, in910_1, in910_2, c285);
    wire[0:0] s911, in911_1, in911_2;
    wire c911;
    assign in911_1 = {c289};
    assign in911_2 = {c290};
    Full_Adder FA_911(s911, c911, in911_1, in911_2, c288);
    wire[0:0] s912, in912_1, in912_2;
    wire c912;
    assign in912_1 = {s292[0]};
    assign in912_2 = {s293[0]};
    Full_Adder FA_912(s912, c912, in912_1, in912_2, c291);
    wire[0:0] s913, in913_1, in913_2;
    wire c913;
    assign in913_1 = {s295[0]};
    assign in913_2 = {s296[0]};
    Full_Adder FA_913(s913, c913, in913_1, in913_2, s294[0]);
    wire[0:0] s914, in914_1, in914_2;
    wire c914;
    assign in914_1 = {s298[0]};
    assign in914_2 = {s299[0]};
    Full_Adder FA_914(s914, c914, in914_1, in914_2, s297[0]);
    wire[0:0] s915, in915_1, in915_2;
    wire c915;
    assign in915_1 = {s301[0]};
    assign in915_2 = {s302[0]};
    Full_Adder FA_915(s915, c915, in915_1, in915_2, s300[0]);
    wire[0:0] s916, in916_1, in916_2;
    wire c916;
    assign in916_1 = {s304[0]};
    assign in916_2 = {s305[0]};
    Full_Adder FA_916(s916, c916, in916_1, in916_2, s303[0]);
    wire[0:0] s917, in917_1, in917_2;
    wire c917;
    assign in917_1 = {s307[0]};
    assign in917_2 = {s308[0]};
    Full_Adder FA_917(s917, c917, in917_1, in917_2, s306[0]);
    wire[0:0] s918, in918_1, in918_2;
    wire c918;
    assign in918_1 = {pp57[11]};
    assign in918_2 = {pp58[10]};
    Full_Adder FA_918(s918, c918, in918_1, in918_2, pp56[12]);
    wire[0:0] s919, in919_1, in919_2;
    wire c919;
    assign in919_1 = {pp60[8]};
    assign in919_2 = {pp61[7]};
    Full_Adder FA_919(s919, c919, in919_1, in919_2, pp59[9]);
    wire[0:0] s920, in920_1, in920_2;
    wire c920;
    assign in920_1 = {pp63[5]};
    assign in920_2 = {c292};
    Full_Adder FA_920(s920, c920, in920_1, in920_2, pp62[6]);
    wire[0:0] s921, in921_1, in921_2;
    wire c921;
    assign in921_1 = {c294};
    assign in921_2 = {c295};
    Full_Adder FA_921(s921, c921, in921_1, in921_2, c293);
    wire[0:0] s922, in922_1, in922_2;
    wire c922;
    assign in922_1 = {c297};
    assign in922_2 = {c298};
    Full_Adder FA_922(s922, c922, in922_1, in922_2, c296);
    wire[0:0] s923, in923_1, in923_2;
    wire c923;
    assign in923_1 = {c300};
    assign in923_2 = {c301};
    Full_Adder FA_923(s923, c923, in923_1, in923_2, c299);
    wire[0:0] s924, in924_1, in924_2;
    wire c924;
    assign in924_1 = {c303};
    assign in924_2 = {c304};
    Full_Adder FA_924(s924, c924, in924_1, in924_2, c302);
    wire[0:0] s925, in925_1, in925_2;
    wire c925;
    assign in925_1 = {c306};
    assign in925_2 = {c307};
    Full_Adder FA_925(s925, c925, in925_1, in925_2, c305);
    wire[0:0] s926, in926_1, in926_2;
    wire c926;
    assign in926_1 = {c309};
    assign in926_2 = {s310[0]};
    Full_Adder FA_926(s926, c926, in926_1, in926_2, c308);
    wire[0:0] s927, in927_1, in927_2;
    wire c927;
    assign in927_1 = {s312[0]};
    assign in927_2 = {s313[0]};
    Full_Adder FA_927(s927, c927, in927_1, in927_2, s311[0]);
    wire[0:0] s928, in928_1, in928_2;
    wire c928;
    assign in928_1 = {s315[0]};
    assign in928_2 = {s316[0]};
    Full_Adder FA_928(s928, c928, in928_1, in928_2, s314[0]);
    wire[0:0] s929, in929_1, in929_2;
    wire c929;
    assign in929_1 = {s318[0]};
    assign in929_2 = {s319[0]};
    Full_Adder FA_929(s929, c929, in929_1, in929_2, s317[0]);
    wire[0:0] s930, in930_1, in930_2;
    wire c930;
    assign in930_1 = {s321[0]};
    assign in930_2 = {s322[0]};
    Full_Adder FA_930(s930, c930, in930_1, in930_2, s320[0]);
    wire[0:0] s931, in931_1, in931_2;
    wire c931;
    assign in931_1 = {s324[0]};
    assign in931_2 = {s325[0]};
    Full_Adder FA_931(s931, c931, in931_1, in931_2, s323[0]);
    wire[0:0] s932, in932_1, in932_2;
    wire c932;
    assign in932_1 = {pp55[14]};
    assign in932_2 = {pp56[13]};
    Full_Adder FA_932(s932, c932, in932_1, in932_2, pp54[15]);
    wire[0:0] s933, in933_1, in933_2;
    wire c933;
    assign in933_1 = {pp58[11]};
    assign in933_2 = {pp59[10]};
    Full_Adder FA_933(s933, c933, in933_1, in933_2, pp57[12]);
    wire[0:0] s934, in934_1, in934_2;
    wire c934;
    assign in934_1 = {pp61[8]};
    assign in934_2 = {pp62[7]};
    Full_Adder FA_934(s934, c934, in934_1, in934_2, pp60[9]);
    wire[0:0] s935, in935_1, in935_2;
    wire c935;
    assign in935_1 = {c310};
    assign in935_2 = {c311};
    Full_Adder FA_935(s935, c935, in935_1, in935_2, pp63[6]);
    wire[0:0] s936, in936_1, in936_2;
    wire c936;
    assign in936_1 = {c313};
    assign in936_2 = {c314};
    Full_Adder FA_936(s936, c936, in936_1, in936_2, c312);
    wire[0:0] s937, in937_1, in937_2;
    wire c937;
    assign in937_1 = {c316};
    assign in937_2 = {c317};
    Full_Adder FA_937(s937, c937, in937_1, in937_2, c315);
    wire[0:0] s938, in938_1, in938_2;
    wire c938;
    assign in938_1 = {c319};
    assign in938_2 = {c320};
    Full_Adder FA_938(s938, c938, in938_1, in938_2, c318);
    wire[0:0] s939, in939_1, in939_2;
    wire c939;
    assign in939_1 = {c322};
    assign in939_2 = {c323};
    Full_Adder FA_939(s939, c939, in939_1, in939_2, c321);
    wire[0:0] s940, in940_1, in940_2;
    wire c940;
    assign in940_1 = {c325};
    assign in940_2 = {c326};
    Full_Adder FA_940(s940, c940, in940_1, in940_2, c324);
    wire[0:0] s941, in941_1, in941_2;
    wire c941;
    assign in941_1 = {s328[0]};
    assign in941_2 = {s329[0]};
    Full_Adder FA_941(s941, c941, in941_1, in941_2, s327[0]);
    wire[0:0] s942, in942_1, in942_2;
    wire c942;
    assign in942_1 = {s331[0]};
    assign in942_2 = {s332[0]};
    Full_Adder FA_942(s942, c942, in942_1, in942_2, s330[0]);
    wire[0:0] s943, in943_1, in943_2;
    wire c943;
    assign in943_1 = {s334[0]};
    assign in943_2 = {s335[0]};
    Full_Adder FA_943(s943, c943, in943_1, in943_2, s333[0]);
    wire[0:0] s944, in944_1, in944_2;
    wire c944;
    assign in944_1 = {s337[0]};
    assign in944_2 = {s338[0]};
    Full_Adder FA_944(s944, c944, in944_1, in944_2, s336[0]);
    wire[0:0] s945, in945_1, in945_2;
    wire c945;
    assign in945_1 = {s340[0]};
    assign in945_2 = {s341[0]};
    Full_Adder FA_945(s945, c945, in945_1, in945_2, s339[0]);
    wire[0:0] s946, in946_1, in946_2;
    wire c946;
    assign in946_1 = {pp53[17]};
    assign in946_2 = {pp54[16]};
    Full_Adder FA_946(s946, c946, in946_1, in946_2, pp52[18]);
    wire[0:0] s947, in947_1, in947_2;
    wire c947;
    assign in947_1 = {pp56[14]};
    assign in947_2 = {pp57[13]};
    Full_Adder FA_947(s947, c947, in947_1, in947_2, pp55[15]);
    wire[0:0] s948, in948_1, in948_2;
    wire c948;
    assign in948_1 = {pp59[11]};
    assign in948_2 = {pp60[10]};
    Full_Adder FA_948(s948, c948, in948_1, in948_2, pp58[12]);
    wire[0:0] s949, in949_1, in949_2;
    wire c949;
    assign in949_1 = {pp62[8]};
    assign in949_2 = {pp63[7]};
    Full_Adder FA_949(s949, c949, in949_1, in949_2, pp61[9]);
    wire[0:0] s950, in950_1, in950_2;
    wire c950;
    assign in950_1 = {c328};
    assign in950_2 = {c329};
    Full_Adder FA_950(s950, c950, in950_1, in950_2, c327);
    wire[0:0] s951, in951_1, in951_2;
    wire c951;
    assign in951_1 = {c331};
    assign in951_2 = {c332};
    Full_Adder FA_951(s951, c951, in951_1, in951_2, c330);
    wire[0:0] s952, in952_1, in952_2;
    wire c952;
    assign in952_1 = {c334};
    assign in952_2 = {c335};
    Full_Adder FA_952(s952, c952, in952_1, in952_2, c333);
    wire[0:0] s953, in953_1, in953_2;
    wire c953;
    assign in953_1 = {c337};
    assign in953_2 = {c338};
    Full_Adder FA_953(s953, c953, in953_1, in953_2, c336);
    wire[0:0] s954, in954_1, in954_2;
    wire c954;
    assign in954_1 = {c340};
    assign in954_2 = {c341};
    Full_Adder FA_954(s954, c954, in954_1, in954_2, c339);
    wire[0:0] s955, in955_1, in955_2;
    wire c955;
    assign in955_1 = {s343[0]};
    assign in955_2 = {s344[0]};
    Full_Adder FA_955(s955, c955, in955_1, in955_2, c342);
    wire[0:0] s956, in956_1, in956_2;
    wire c956;
    assign in956_1 = {s346[0]};
    assign in956_2 = {s347[0]};
    Full_Adder FA_956(s956, c956, in956_1, in956_2, s345[0]);
    wire[0:0] s957, in957_1, in957_2;
    wire c957;
    assign in957_1 = {s349[0]};
    assign in957_2 = {s350[0]};
    Full_Adder FA_957(s957, c957, in957_1, in957_2, s348[0]);
    wire[0:0] s958, in958_1, in958_2;
    wire c958;
    assign in958_1 = {s352[0]};
    assign in958_2 = {s353[0]};
    Full_Adder FA_958(s958, c958, in958_1, in958_2, s351[0]);
    wire[0:0] s959, in959_1, in959_2;
    wire c959;
    assign in959_1 = {s355[0]};
    assign in959_2 = {s356[0]};
    Full_Adder FA_959(s959, c959, in959_1, in959_2, s354[0]);
    wire[0:0] s960, in960_1, in960_2;
    wire c960;
    assign in960_1 = {pp51[20]};
    assign in960_2 = {pp52[19]};
    Full_Adder FA_960(s960, c960, in960_1, in960_2, pp50[21]);
    wire[0:0] s961, in961_1, in961_2;
    wire c961;
    assign in961_1 = {pp54[17]};
    assign in961_2 = {pp55[16]};
    Full_Adder FA_961(s961, c961, in961_1, in961_2, pp53[18]);
    wire[0:0] s962, in962_1, in962_2;
    wire c962;
    assign in962_1 = {pp57[14]};
    assign in962_2 = {pp58[13]};
    Full_Adder FA_962(s962, c962, in962_1, in962_2, pp56[15]);
    wire[0:0] s963, in963_1, in963_2;
    wire c963;
    assign in963_1 = {pp60[11]};
    assign in963_2 = {pp61[10]};
    Full_Adder FA_963(s963, c963, in963_1, in963_2, pp59[12]);
    wire[0:0] s964, in964_1, in964_2;
    wire c964;
    assign in964_1 = {pp63[8]};
    assign in964_2 = {c343};
    Full_Adder FA_964(s964, c964, in964_1, in964_2, pp62[9]);
    wire[0:0] s965, in965_1, in965_2;
    wire c965;
    assign in965_1 = {c345};
    assign in965_2 = {c346};
    Full_Adder FA_965(s965, c965, in965_1, in965_2, c344);
    wire[0:0] s966, in966_1, in966_2;
    wire c966;
    assign in966_1 = {c348};
    assign in966_2 = {c349};
    Full_Adder FA_966(s966, c966, in966_1, in966_2, c347);
    wire[0:0] s967, in967_1, in967_2;
    wire c967;
    assign in967_1 = {c351};
    assign in967_2 = {c352};
    Full_Adder FA_967(s967, c967, in967_1, in967_2, c350);
    wire[0:0] s968, in968_1, in968_2;
    wire c968;
    assign in968_1 = {c354};
    assign in968_2 = {c355};
    Full_Adder FA_968(s968, c968, in968_1, in968_2, c353);
    wire[0:0] s969, in969_1, in969_2;
    wire c969;
    assign in969_1 = {c357};
    assign in969_2 = {s358[0]};
    Full_Adder FA_969(s969, c969, in969_1, in969_2, c356);
    wire[0:0] s970, in970_1, in970_2;
    wire c970;
    assign in970_1 = {s360[0]};
    assign in970_2 = {s361[0]};
    Full_Adder FA_970(s970, c970, in970_1, in970_2, s359[0]);
    wire[0:0] s971, in971_1, in971_2;
    wire c971;
    assign in971_1 = {s363[0]};
    assign in971_2 = {s364[0]};
    Full_Adder FA_971(s971, c971, in971_1, in971_2, s362[0]);
    wire[0:0] s972, in972_1, in972_2;
    wire c972;
    assign in972_1 = {s366[0]};
    assign in972_2 = {s367[0]};
    Full_Adder FA_972(s972, c972, in972_1, in972_2, s365[0]);
    wire[0:0] s973, in973_1, in973_2;
    wire c973;
    assign in973_1 = {s369[0]};
    assign in973_2 = {s370[0]};
    Full_Adder FA_973(s973, c973, in973_1, in973_2, s368[0]);
    wire[0:0] s974, in974_1, in974_2;
    wire c974;
    assign in974_1 = {pp49[23]};
    assign in974_2 = {pp50[22]};
    Full_Adder FA_974(s974, c974, in974_1, in974_2, pp48[24]);
    wire[0:0] s975, in975_1, in975_2;
    wire c975;
    assign in975_1 = {pp52[20]};
    assign in975_2 = {pp53[19]};
    Full_Adder FA_975(s975, c975, in975_1, in975_2, pp51[21]);
    wire[0:0] s976, in976_1, in976_2;
    wire c976;
    assign in976_1 = {pp55[17]};
    assign in976_2 = {pp56[16]};
    Full_Adder FA_976(s976, c976, in976_1, in976_2, pp54[18]);
    wire[0:0] s977, in977_1, in977_2;
    wire c977;
    assign in977_1 = {pp58[14]};
    assign in977_2 = {pp59[13]};
    Full_Adder FA_977(s977, c977, in977_1, in977_2, pp57[15]);
    wire[0:0] s978, in978_1, in978_2;
    wire c978;
    assign in978_1 = {pp61[11]};
    assign in978_2 = {pp62[10]};
    Full_Adder FA_978(s978, c978, in978_1, in978_2, pp60[12]);
    wire[0:0] s979, in979_1, in979_2;
    wire c979;
    assign in979_1 = {c358};
    assign in979_2 = {c359};
    Full_Adder FA_979(s979, c979, in979_1, in979_2, pp63[9]);
    wire[0:0] s980, in980_1, in980_2;
    wire c980;
    assign in980_1 = {c361};
    assign in980_2 = {c362};
    Full_Adder FA_980(s980, c980, in980_1, in980_2, c360);
    wire[0:0] s981, in981_1, in981_2;
    wire c981;
    assign in981_1 = {c364};
    assign in981_2 = {c365};
    Full_Adder FA_981(s981, c981, in981_1, in981_2, c363);
    wire[0:0] s982, in982_1, in982_2;
    wire c982;
    assign in982_1 = {c367};
    assign in982_2 = {c368};
    Full_Adder FA_982(s982, c982, in982_1, in982_2, c366);
    wire[0:0] s983, in983_1, in983_2;
    wire c983;
    assign in983_1 = {c370};
    assign in983_2 = {c371};
    Full_Adder FA_983(s983, c983, in983_1, in983_2, c369);
    wire[0:0] s984, in984_1, in984_2;
    wire c984;
    assign in984_1 = {s373[0]};
    assign in984_2 = {s374[0]};
    Full_Adder FA_984(s984, c984, in984_1, in984_2, s372[0]);
    wire[0:0] s985, in985_1, in985_2;
    wire c985;
    assign in985_1 = {s376[0]};
    assign in985_2 = {s377[0]};
    Full_Adder FA_985(s985, c985, in985_1, in985_2, s375[0]);
    wire[0:0] s986, in986_1, in986_2;
    wire c986;
    assign in986_1 = {s379[0]};
    assign in986_2 = {s380[0]};
    Full_Adder FA_986(s986, c986, in986_1, in986_2, s378[0]);
    wire[0:0] s987, in987_1, in987_2;
    wire c987;
    assign in987_1 = {s382[0]};
    assign in987_2 = {s383[0]};
    Full_Adder FA_987(s987, c987, in987_1, in987_2, s381[0]);
    wire[0:0] s988, in988_1, in988_2;
    wire c988;
    assign in988_1 = {pp47[26]};
    assign in988_2 = {pp48[25]};
    Full_Adder FA_988(s988, c988, in988_1, in988_2, pp46[27]);
    wire[0:0] s989, in989_1, in989_2;
    wire c989;
    assign in989_1 = {pp50[23]};
    assign in989_2 = {pp51[22]};
    Full_Adder FA_989(s989, c989, in989_1, in989_2, pp49[24]);
    wire[0:0] s990, in990_1, in990_2;
    wire c990;
    assign in990_1 = {pp53[20]};
    assign in990_2 = {pp54[19]};
    Full_Adder FA_990(s990, c990, in990_1, in990_2, pp52[21]);
    wire[0:0] s991, in991_1, in991_2;
    wire c991;
    assign in991_1 = {pp56[17]};
    assign in991_2 = {pp57[16]};
    Full_Adder FA_991(s991, c991, in991_1, in991_2, pp55[18]);
    wire[0:0] s992, in992_1, in992_2;
    wire c992;
    assign in992_1 = {pp59[14]};
    assign in992_2 = {pp60[13]};
    Full_Adder FA_992(s992, c992, in992_1, in992_2, pp58[15]);
    wire[0:0] s993, in993_1, in993_2;
    wire c993;
    assign in993_1 = {pp62[11]};
    assign in993_2 = {pp63[10]};
    Full_Adder FA_993(s993, c993, in993_1, in993_2, pp61[12]);
    wire[0:0] s994, in994_1, in994_2;
    wire c994;
    assign in994_1 = {c373};
    assign in994_2 = {c374};
    Full_Adder FA_994(s994, c994, in994_1, in994_2, c372);
    wire[0:0] s995, in995_1, in995_2;
    wire c995;
    assign in995_1 = {c376};
    assign in995_2 = {c377};
    Full_Adder FA_995(s995, c995, in995_1, in995_2, c375);
    wire[0:0] s996, in996_1, in996_2;
    wire c996;
    assign in996_1 = {c379};
    assign in996_2 = {c380};
    Full_Adder FA_996(s996, c996, in996_1, in996_2, c378);
    wire[0:0] s997, in997_1, in997_2;
    wire c997;
    assign in997_1 = {c382};
    assign in997_2 = {c383};
    Full_Adder FA_997(s997, c997, in997_1, in997_2, c381);
    wire[0:0] s998, in998_1, in998_2;
    wire c998;
    assign in998_1 = {s385[0]};
    assign in998_2 = {s386[0]};
    Full_Adder FA_998(s998, c998, in998_1, in998_2, c384);
    wire[0:0] s999, in999_1, in999_2;
    wire c999;
    assign in999_1 = {s388[0]};
    assign in999_2 = {s389[0]};
    Full_Adder FA_999(s999, c999, in999_1, in999_2, s387[0]);
    wire[0:0] s1000, in1000_1, in1000_2;
    wire c1000;
    assign in1000_1 = {s391[0]};
    assign in1000_2 = {s392[0]};
    Full_Adder FA_1000(s1000, c1000, in1000_1, in1000_2, s390[0]);
    wire[0:0] s1001, in1001_1, in1001_2;
    wire c1001;
    assign in1001_1 = {s394[0]};
    assign in1001_2 = {s395[0]};
    Full_Adder FA_1001(s1001, c1001, in1001_1, in1001_2, s393[0]);
    wire[0:0] s1002, in1002_1, in1002_2;
    wire c1002;
    assign in1002_1 = {pp45[29]};
    assign in1002_2 = {pp46[28]};
    Full_Adder FA_1002(s1002, c1002, in1002_1, in1002_2, pp44[30]);
    wire[0:0] s1003, in1003_1, in1003_2;
    wire c1003;
    assign in1003_1 = {pp48[26]};
    assign in1003_2 = {pp49[25]};
    Full_Adder FA_1003(s1003, c1003, in1003_1, in1003_2, pp47[27]);
    wire[0:0] s1004, in1004_1, in1004_2;
    wire c1004;
    assign in1004_1 = {pp51[23]};
    assign in1004_2 = {pp52[22]};
    Full_Adder FA_1004(s1004, c1004, in1004_1, in1004_2, pp50[24]);
    wire[0:0] s1005, in1005_1, in1005_2;
    wire c1005;
    assign in1005_1 = {pp54[20]};
    assign in1005_2 = {pp55[19]};
    Full_Adder FA_1005(s1005, c1005, in1005_1, in1005_2, pp53[21]);
    wire[0:0] s1006, in1006_1, in1006_2;
    wire c1006;
    assign in1006_1 = {pp57[17]};
    assign in1006_2 = {pp58[16]};
    Full_Adder FA_1006(s1006, c1006, in1006_1, in1006_2, pp56[18]);
    wire[0:0] s1007, in1007_1, in1007_2;
    wire c1007;
    assign in1007_1 = {pp60[14]};
    assign in1007_2 = {pp61[13]};
    Full_Adder FA_1007(s1007, c1007, in1007_1, in1007_2, pp59[15]);
    wire[0:0] s1008, in1008_1, in1008_2;
    wire c1008;
    assign in1008_1 = {pp63[11]};
    assign in1008_2 = {c385};
    Full_Adder FA_1008(s1008, c1008, in1008_1, in1008_2, pp62[12]);
    wire[0:0] s1009, in1009_1, in1009_2;
    wire c1009;
    assign in1009_1 = {c387};
    assign in1009_2 = {c388};
    Full_Adder FA_1009(s1009, c1009, in1009_1, in1009_2, c386);
    wire[0:0] s1010, in1010_1, in1010_2;
    wire c1010;
    assign in1010_1 = {c390};
    assign in1010_2 = {c391};
    Full_Adder FA_1010(s1010, c1010, in1010_1, in1010_2, c389);
    wire[0:0] s1011, in1011_1, in1011_2;
    wire c1011;
    assign in1011_1 = {c393};
    assign in1011_2 = {c394};
    Full_Adder FA_1011(s1011, c1011, in1011_1, in1011_2, c392);
    wire[0:0] s1012, in1012_1, in1012_2;
    wire c1012;
    assign in1012_1 = {c396};
    assign in1012_2 = {s397[0]};
    Full_Adder FA_1012(s1012, c1012, in1012_1, in1012_2, c395);
    wire[0:0] s1013, in1013_1, in1013_2;
    wire c1013;
    assign in1013_1 = {s399[0]};
    assign in1013_2 = {s400[0]};
    Full_Adder FA_1013(s1013, c1013, in1013_1, in1013_2, s398[0]);
    wire[0:0] s1014, in1014_1, in1014_2;
    wire c1014;
    assign in1014_1 = {s402[0]};
    assign in1014_2 = {s403[0]};
    Full_Adder FA_1014(s1014, c1014, in1014_1, in1014_2, s401[0]);
    wire[0:0] s1015, in1015_1, in1015_2;
    wire c1015;
    assign in1015_1 = {s405[0]};
    assign in1015_2 = {s406[0]};
    Full_Adder FA_1015(s1015, c1015, in1015_1, in1015_2, s404[0]);
    wire[0:0] s1016, in1016_1, in1016_2;
    wire c1016;
    assign in1016_1 = {pp43[32]};
    assign in1016_2 = {pp44[31]};
    Full_Adder FA_1016(s1016, c1016, in1016_1, in1016_2, pp42[33]);
    wire[0:0] s1017, in1017_1, in1017_2;
    wire c1017;
    assign in1017_1 = {pp46[29]};
    assign in1017_2 = {pp47[28]};
    Full_Adder FA_1017(s1017, c1017, in1017_1, in1017_2, pp45[30]);
    wire[0:0] s1018, in1018_1, in1018_2;
    wire c1018;
    assign in1018_1 = {pp49[26]};
    assign in1018_2 = {pp50[25]};
    Full_Adder FA_1018(s1018, c1018, in1018_1, in1018_2, pp48[27]);
    wire[0:0] s1019, in1019_1, in1019_2;
    wire c1019;
    assign in1019_1 = {pp52[23]};
    assign in1019_2 = {pp53[22]};
    Full_Adder FA_1019(s1019, c1019, in1019_1, in1019_2, pp51[24]);
    wire[0:0] s1020, in1020_1, in1020_2;
    wire c1020;
    assign in1020_1 = {pp55[20]};
    assign in1020_2 = {pp56[19]};
    Full_Adder FA_1020(s1020, c1020, in1020_1, in1020_2, pp54[21]);
    wire[0:0] s1021, in1021_1, in1021_2;
    wire c1021;
    assign in1021_1 = {pp58[17]};
    assign in1021_2 = {pp59[16]};
    Full_Adder FA_1021(s1021, c1021, in1021_1, in1021_2, pp57[18]);
    wire[0:0] s1022, in1022_1, in1022_2;
    wire c1022;
    assign in1022_1 = {pp61[14]};
    assign in1022_2 = {pp62[13]};
    Full_Adder FA_1022(s1022, c1022, in1022_1, in1022_2, pp60[15]);
    wire[0:0] s1023, in1023_1, in1023_2;
    wire c1023;
    assign in1023_1 = {c397};
    assign in1023_2 = {c398};
    Full_Adder FA_1023(s1023, c1023, in1023_1, in1023_2, pp63[12]);
    wire[0:0] s1024, in1024_1, in1024_2;
    wire c1024;
    assign in1024_1 = {c400};
    assign in1024_2 = {c401};
    Full_Adder FA_1024(s1024, c1024, in1024_1, in1024_2, c399);
    wire[0:0] s1025, in1025_1, in1025_2;
    wire c1025;
    assign in1025_1 = {c403};
    assign in1025_2 = {c404};
    Full_Adder FA_1025(s1025, c1025, in1025_1, in1025_2, c402);
    wire[0:0] s1026, in1026_1, in1026_2;
    wire c1026;
    assign in1026_1 = {c406};
    assign in1026_2 = {c407};
    Full_Adder FA_1026(s1026, c1026, in1026_1, in1026_2, c405);
    wire[0:0] s1027, in1027_1, in1027_2;
    wire c1027;
    assign in1027_1 = {s409[0]};
    assign in1027_2 = {s410[0]};
    Full_Adder FA_1027(s1027, c1027, in1027_1, in1027_2, s408[0]);
    wire[0:0] s1028, in1028_1, in1028_2;
    wire c1028;
    assign in1028_1 = {s412[0]};
    assign in1028_2 = {s413[0]};
    Full_Adder FA_1028(s1028, c1028, in1028_1, in1028_2, s411[0]);
    wire[0:0] s1029, in1029_1, in1029_2;
    wire c1029;
    assign in1029_1 = {s415[0]};
    assign in1029_2 = {s416[0]};
    Full_Adder FA_1029(s1029, c1029, in1029_1, in1029_2, s414[0]);
    wire[0:0] s1030, in1030_1, in1030_2;
    wire c1030;
    assign in1030_1 = {pp41[35]};
    assign in1030_2 = {pp42[34]};
    Full_Adder FA_1030(s1030, c1030, in1030_1, in1030_2, pp40[36]);
    wire[0:0] s1031, in1031_1, in1031_2;
    wire c1031;
    assign in1031_1 = {pp44[32]};
    assign in1031_2 = {pp45[31]};
    Full_Adder FA_1031(s1031, c1031, in1031_1, in1031_2, pp43[33]);
    wire[0:0] s1032, in1032_1, in1032_2;
    wire c1032;
    assign in1032_1 = {pp47[29]};
    assign in1032_2 = {pp48[28]};
    Full_Adder FA_1032(s1032, c1032, in1032_1, in1032_2, pp46[30]);
    wire[0:0] s1033, in1033_1, in1033_2;
    wire c1033;
    assign in1033_1 = {pp50[26]};
    assign in1033_2 = {pp51[25]};
    Full_Adder FA_1033(s1033, c1033, in1033_1, in1033_2, pp49[27]);
    wire[0:0] s1034, in1034_1, in1034_2;
    wire c1034;
    assign in1034_1 = {pp53[23]};
    assign in1034_2 = {pp54[22]};
    Full_Adder FA_1034(s1034, c1034, in1034_1, in1034_2, pp52[24]);
    wire[0:0] s1035, in1035_1, in1035_2;
    wire c1035;
    assign in1035_1 = {pp56[20]};
    assign in1035_2 = {pp57[19]};
    Full_Adder FA_1035(s1035, c1035, in1035_1, in1035_2, pp55[21]);
    wire[0:0] s1036, in1036_1, in1036_2;
    wire c1036;
    assign in1036_1 = {pp59[17]};
    assign in1036_2 = {pp60[16]};
    Full_Adder FA_1036(s1036, c1036, in1036_1, in1036_2, pp58[18]);
    wire[0:0] s1037, in1037_1, in1037_2;
    wire c1037;
    assign in1037_1 = {pp62[14]};
    assign in1037_2 = {pp63[13]};
    Full_Adder FA_1037(s1037, c1037, in1037_1, in1037_2, pp61[15]);
    wire[0:0] s1038, in1038_1, in1038_2;
    wire c1038;
    assign in1038_1 = {c409};
    assign in1038_2 = {c410};
    Full_Adder FA_1038(s1038, c1038, in1038_1, in1038_2, c408);
    wire[0:0] s1039, in1039_1, in1039_2;
    wire c1039;
    assign in1039_1 = {c412};
    assign in1039_2 = {c413};
    Full_Adder FA_1039(s1039, c1039, in1039_1, in1039_2, c411);
    wire[0:0] s1040, in1040_1, in1040_2;
    wire c1040;
    assign in1040_1 = {c415};
    assign in1040_2 = {c416};
    Full_Adder FA_1040(s1040, c1040, in1040_1, in1040_2, c414);
    wire[0:0] s1041, in1041_1, in1041_2;
    wire c1041;
    assign in1041_1 = {s418[0]};
    assign in1041_2 = {s419[0]};
    Full_Adder FA_1041(s1041, c1041, in1041_1, in1041_2, c417);
    wire[0:0] s1042, in1042_1, in1042_2;
    wire c1042;
    assign in1042_1 = {s421[0]};
    assign in1042_2 = {s422[0]};
    Full_Adder FA_1042(s1042, c1042, in1042_1, in1042_2, s420[0]);
    wire[0:0] s1043, in1043_1, in1043_2;
    wire c1043;
    assign in1043_1 = {s424[0]};
    assign in1043_2 = {s425[0]};
    Full_Adder FA_1043(s1043, c1043, in1043_1, in1043_2, s423[0]);
    wire[0:0] s1044, in1044_1, in1044_2;
    wire c1044;
    assign in1044_1 = {pp39[38]};
    assign in1044_2 = {pp40[37]};
    Full_Adder FA_1044(s1044, c1044, in1044_1, in1044_2, pp38[39]);
    wire[0:0] s1045, in1045_1, in1045_2;
    wire c1045;
    assign in1045_1 = {pp42[35]};
    assign in1045_2 = {pp43[34]};
    Full_Adder FA_1045(s1045, c1045, in1045_1, in1045_2, pp41[36]);
    wire[0:0] s1046, in1046_1, in1046_2;
    wire c1046;
    assign in1046_1 = {pp45[32]};
    assign in1046_2 = {pp46[31]};
    Full_Adder FA_1046(s1046, c1046, in1046_1, in1046_2, pp44[33]);
    wire[0:0] s1047, in1047_1, in1047_2;
    wire c1047;
    assign in1047_1 = {pp48[29]};
    assign in1047_2 = {pp49[28]};
    Full_Adder FA_1047(s1047, c1047, in1047_1, in1047_2, pp47[30]);
    wire[0:0] s1048, in1048_1, in1048_2;
    wire c1048;
    assign in1048_1 = {pp51[26]};
    assign in1048_2 = {pp52[25]};
    Full_Adder FA_1048(s1048, c1048, in1048_1, in1048_2, pp50[27]);
    wire[0:0] s1049, in1049_1, in1049_2;
    wire c1049;
    assign in1049_1 = {pp54[23]};
    assign in1049_2 = {pp55[22]};
    Full_Adder FA_1049(s1049, c1049, in1049_1, in1049_2, pp53[24]);
    wire[0:0] s1050, in1050_1, in1050_2;
    wire c1050;
    assign in1050_1 = {pp57[20]};
    assign in1050_2 = {pp58[19]};
    Full_Adder FA_1050(s1050, c1050, in1050_1, in1050_2, pp56[21]);
    wire[0:0] s1051, in1051_1, in1051_2;
    wire c1051;
    assign in1051_1 = {pp60[17]};
    assign in1051_2 = {pp61[16]};
    Full_Adder FA_1051(s1051, c1051, in1051_1, in1051_2, pp59[18]);
    wire[0:0] s1052, in1052_1, in1052_2;
    wire c1052;
    assign in1052_1 = {pp63[14]};
    assign in1052_2 = {c418};
    Full_Adder FA_1052(s1052, c1052, in1052_1, in1052_2, pp62[15]);
    wire[0:0] s1053, in1053_1, in1053_2;
    wire c1053;
    assign in1053_1 = {c420};
    assign in1053_2 = {c421};
    Full_Adder FA_1053(s1053, c1053, in1053_1, in1053_2, c419);
    wire[0:0] s1054, in1054_1, in1054_2;
    wire c1054;
    assign in1054_1 = {c423};
    assign in1054_2 = {c424};
    Full_Adder FA_1054(s1054, c1054, in1054_1, in1054_2, c422);
    wire[0:0] s1055, in1055_1, in1055_2;
    wire c1055;
    assign in1055_1 = {c426};
    assign in1055_2 = {s427[0]};
    Full_Adder FA_1055(s1055, c1055, in1055_1, in1055_2, c425);
    wire[0:0] s1056, in1056_1, in1056_2;
    wire c1056;
    assign in1056_1 = {s429[0]};
    assign in1056_2 = {s430[0]};
    Full_Adder FA_1056(s1056, c1056, in1056_1, in1056_2, s428[0]);
    wire[0:0] s1057, in1057_1, in1057_2;
    wire c1057;
    assign in1057_1 = {s432[0]};
    assign in1057_2 = {s433[0]};
    Full_Adder FA_1057(s1057, c1057, in1057_1, in1057_2, s431[0]);
    wire[0:0] s1058, in1058_1, in1058_2;
    wire c1058;
    assign in1058_1 = {pp37[41]};
    assign in1058_2 = {pp38[40]};
    Full_Adder FA_1058(s1058, c1058, in1058_1, in1058_2, pp36[42]);
    wire[0:0] s1059, in1059_1, in1059_2;
    wire c1059;
    assign in1059_1 = {pp40[38]};
    assign in1059_2 = {pp41[37]};
    Full_Adder FA_1059(s1059, c1059, in1059_1, in1059_2, pp39[39]);
    wire[0:0] s1060, in1060_1, in1060_2;
    wire c1060;
    assign in1060_1 = {pp43[35]};
    assign in1060_2 = {pp44[34]};
    Full_Adder FA_1060(s1060, c1060, in1060_1, in1060_2, pp42[36]);
    wire[0:0] s1061, in1061_1, in1061_2;
    wire c1061;
    assign in1061_1 = {pp46[32]};
    assign in1061_2 = {pp47[31]};
    Full_Adder FA_1061(s1061, c1061, in1061_1, in1061_2, pp45[33]);
    wire[0:0] s1062, in1062_1, in1062_2;
    wire c1062;
    assign in1062_1 = {pp49[29]};
    assign in1062_2 = {pp50[28]};
    Full_Adder FA_1062(s1062, c1062, in1062_1, in1062_2, pp48[30]);
    wire[0:0] s1063, in1063_1, in1063_2;
    wire c1063;
    assign in1063_1 = {pp52[26]};
    assign in1063_2 = {pp53[25]};
    Full_Adder FA_1063(s1063, c1063, in1063_1, in1063_2, pp51[27]);
    wire[0:0] s1064, in1064_1, in1064_2;
    wire c1064;
    assign in1064_1 = {pp55[23]};
    assign in1064_2 = {pp56[22]};
    Full_Adder FA_1064(s1064, c1064, in1064_1, in1064_2, pp54[24]);
    wire[0:0] s1065, in1065_1, in1065_2;
    wire c1065;
    assign in1065_1 = {pp58[20]};
    assign in1065_2 = {pp59[19]};
    Full_Adder FA_1065(s1065, c1065, in1065_1, in1065_2, pp57[21]);
    wire[0:0] s1066, in1066_1, in1066_2;
    wire c1066;
    assign in1066_1 = {pp61[17]};
    assign in1066_2 = {pp62[16]};
    Full_Adder FA_1066(s1066, c1066, in1066_1, in1066_2, pp60[18]);
    wire[0:0] s1067, in1067_1, in1067_2;
    wire c1067;
    assign in1067_1 = {c427};
    assign in1067_2 = {c428};
    Full_Adder FA_1067(s1067, c1067, in1067_1, in1067_2, pp63[15]);
    wire[0:0] s1068, in1068_1, in1068_2;
    wire c1068;
    assign in1068_1 = {c430};
    assign in1068_2 = {c431};
    Full_Adder FA_1068(s1068, c1068, in1068_1, in1068_2, c429);
    wire[0:0] s1069, in1069_1, in1069_2;
    wire c1069;
    assign in1069_1 = {c433};
    assign in1069_2 = {c434};
    Full_Adder FA_1069(s1069, c1069, in1069_1, in1069_2, c432);
    wire[0:0] s1070, in1070_1, in1070_2;
    wire c1070;
    assign in1070_1 = {s436[0]};
    assign in1070_2 = {s437[0]};
    Full_Adder FA_1070(s1070, c1070, in1070_1, in1070_2, s435[0]);
    wire[0:0] s1071, in1071_1, in1071_2;
    wire c1071;
    assign in1071_1 = {s439[0]};
    assign in1071_2 = {s440[0]};
    Full_Adder FA_1071(s1071, c1071, in1071_1, in1071_2, s438[0]);
    wire[0:0] s1072, in1072_1, in1072_2;
    wire c1072;
    assign in1072_1 = {pp35[44]};
    assign in1072_2 = {pp36[43]};
    Full_Adder FA_1072(s1072, c1072, in1072_1, in1072_2, pp34[45]);
    wire[0:0] s1073, in1073_1, in1073_2;
    wire c1073;
    assign in1073_1 = {pp38[41]};
    assign in1073_2 = {pp39[40]};
    Full_Adder FA_1073(s1073, c1073, in1073_1, in1073_2, pp37[42]);
    wire[0:0] s1074, in1074_1, in1074_2;
    wire c1074;
    assign in1074_1 = {pp41[38]};
    assign in1074_2 = {pp42[37]};
    Full_Adder FA_1074(s1074, c1074, in1074_1, in1074_2, pp40[39]);
    wire[0:0] s1075, in1075_1, in1075_2;
    wire c1075;
    assign in1075_1 = {pp44[35]};
    assign in1075_2 = {pp45[34]};
    Full_Adder FA_1075(s1075, c1075, in1075_1, in1075_2, pp43[36]);
    wire[0:0] s1076, in1076_1, in1076_2;
    wire c1076;
    assign in1076_1 = {pp47[32]};
    assign in1076_2 = {pp48[31]};
    Full_Adder FA_1076(s1076, c1076, in1076_1, in1076_2, pp46[33]);
    wire[0:0] s1077, in1077_1, in1077_2;
    wire c1077;
    assign in1077_1 = {pp50[29]};
    assign in1077_2 = {pp51[28]};
    Full_Adder FA_1077(s1077, c1077, in1077_1, in1077_2, pp49[30]);
    wire[0:0] s1078, in1078_1, in1078_2;
    wire c1078;
    assign in1078_1 = {pp53[26]};
    assign in1078_2 = {pp54[25]};
    Full_Adder FA_1078(s1078, c1078, in1078_1, in1078_2, pp52[27]);
    wire[0:0] s1079, in1079_1, in1079_2;
    wire c1079;
    assign in1079_1 = {pp56[23]};
    assign in1079_2 = {pp57[22]};
    Full_Adder FA_1079(s1079, c1079, in1079_1, in1079_2, pp55[24]);
    wire[0:0] s1080, in1080_1, in1080_2;
    wire c1080;
    assign in1080_1 = {pp59[20]};
    assign in1080_2 = {pp60[19]};
    Full_Adder FA_1080(s1080, c1080, in1080_1, in1080_2, pp58[21]);
    wire[0:0] s1081, in1081_1, in1081_2;
    wire c1081;
    assign in1081_1 = {pp62[17]};
    assign in1081_2 = {pp63[16]};
    Full_Adder FA_1081(s1081, c1081, in1081_1, in1081_2, pp61[18]);
    wire[0:0] s1082, in1082_1, in1082_2;
    wire c1082;
    assign in1082_1 = {c436};
    assign in1082_2 = {c437};
    Full_Adder FA_1082(s1082, c1082, in1082_1, in1082_2, c435);
    wire[0:0] s1083, in1083_1, in1083_2;
    wire c1083;
    assign in1083_1 = {c439};
    assign in1083_2 = {c440};
    Full_Adder FA_1083(s1083, c1083, in1083_1, in1083_2, c438);
    wire[0:0] s1084, in1084_1, in1084_2;
    wire c1084;
    assign in1084_1 = {s442[0]};
    assign in1084_2 = {s443[0]};
    Full_Adder FA_1084(s1084, c1084, in1084_1, in1084_2, c441);
    wire[0:0] s1085, in1085_1, in1085_2;
    wire c1085;
    assign in1085_1 = {s445[0]};
    assign in1085_2 = {s446[0]};
    Full_Adder FA_1085(s1085, c1085, in1085_1, in1085_2, s444[0]);
    wire[0:0] s1086, in1086_1, in1086_2;
    wire c1086;
    assign in1086_1 = {pp33[47]};
    assign in1086_2 = {pp34[46]};
    Full_Adder FA_1086(s1086, c1086, in1086_1, in1086_2, pp32[48]);
    wire[0:0] s1087, in1087_1, in1087_2;
    wire c1087;
    assign in1087_1 = {pp36[44]};
    assign in1087_2 = {pp37[43]};
    Full_Adder FA_1087(s1087, c1087, in1087_1, in1087_2, pp35[45]);
    wire[0:0] s1088, in1088_1, in1088_2;
    wire c1088;
    assign in1088_1 = {pp39[41]};
    assign in1088_2 = {pp40[40]};
    Full_Adder FA_1088(s1088, c1088, in1088_1, in1088_2, pp38[42]);
    wire[0:0] s1089, in1089_1, in1089_2;
    wire c1089;
    assign in1089_1 = {pp42[38]};
    assign in1089_2 = {pp43[37]};
    Full_Adder FA_1089(s1089, c1089, in1089_1, in1089_2, pp41[39]);
    wire[0:0] s1090, in1090_1, in1090_2;
    wire c1090;
    assign in1090_1 = {pp45[35]};
    assign in1090_2 = {pp46[34]};
    Full_Adder FA_1090(s1090, c1090, in1090_1, in1090_2, pp44[36]);
    wire[0:0] s1091, in1091_1, in1091_2;
    wire c1091;
    assign in1091_1 = {pp48[32]};
    assign in1091_2 = {pp49[31]};
    Full_Adder FA_1091(s1091, c1091, in1091_1, in1091_2, pp47[33]);
    wire[0:0] s1092, in1092_1, in1092_2;
    wire c1092;
    assign in1092_1 = {pp51[29]};
    assign in1092_2 = {pp52[28]};
    Full_Adder FA_1092(s1092, c1092, in1092_1, in1092_2, pp50[30]);
    wire[0:0] s1093, in1093_1, in1093_2;
    wire c1093;
    assign in1093_1 = {pp54[26]};
    assign in1093_2 = {pp55[25]};
    Full_Adder FA_1093(s1093, c1093, in1093_1, in1093_2, pp53[27]);
    wire[0:0] s1094, in1094_1, in1094_2;
    wire c1094;
    assign in1094_1 = {pp57[23]};
    assign in1094_2 = {pp58[22]};
    Full_Adder FA_1094(s1094, c1094, in1094_1, in1094_2, pp56[24]);
    wire[0:0] s1095, in1095_1, in1095_2;
    wire c1095;
    assign in1095_1 = {pp60[20]};
    assign in1095_2 = {pp61[19]};
    Full_Adder FA_1095(s1095, c1095, in1095_1, in1095_2, pp59[21]);
    wire[0:0] s1096, in1096_1, in1096_2;
    wire c1096;
    assign in1096_1 = {pp63[17]};
    assign in1096_2 = {c442};
    Full_Adder FA_1096(s1096, c1096, in1096_1, in1096_2, pp62[18]);
    wire[0:0] s1097, in1097_1, in1097_2;
    wire c1097;
    assign in1097_1 = {c444};
    assign in1097_2 = {c445};
    Full_Adder FA_1097(s1097, c1097, in1097_1, in1097_2, c443);
    wire[0:0] s1098, in1098_1, in1098_2;
    wire c1098;
    assign in1098_1 = {c447};
    assign in1098_2 = {s448[0]};
    Full_Adder FA_1098(s1098, c1098, in1098_1, in1098_2, c446);
    wire[0:0] s1099, in1099_1, in1099_2;
    wire c1099;
    assign in1099_1 = {s450[0]};
    assign in1099_2 = {s451[0]};
    Full_Adder FA_1099(s1099, c1099, in1099_1, in1099_2, s449[0]);
    wire[0:0] s1100, in1100_1, in1100_2;
    wire c1100;
    assign in1100_1 = {pp31[50]};
    assign in1100_2 = {pp32[49]};
    Full_Adder FA_1100(s1100, c1100, in1100_1, in1100_2, pp30[51]);
    wire[0:0] s1101, in1101_1, in1101_2;
    wire c1101;
    assign in1101_1 = {pp34[47]};
    assign in1101_2 = {pp35[46]};
    Full_Adder FA_1101(s1101, c1101, in1101_1, in1101_2, pp33[48]);
    wire[0:0] s1102, in1102_1, in1102_2;
    wire c1102;
    assign in1102_1 = {pp37[44]};
    assign in1102_2 = {pp38[43]};
    Full_Adder FA_1102(s1102, c1102, in1102_1, in1102_2, pp36[45]);
    wire[0:0] s1103, in1103_1, in1103_2;
    wire c1103;
    assign in1103_1 = {pp40[41]};
    assign in1103_2 = {pp41[40]};
    Full_Adder FA_1103(s1103, c1103, in1103_1, in1103_2, pp39[42]);
    wire[0:0] s1104, in1104_1, in1104_2;
    wire c1104;
    assign in1104_1 = {pp43[38]};
    assign in1104_2 = {pp44[37]};
    Full_Adder FA_1104(s1104, c1104, in1104_1, in1104_2, pp42[39]);
    wire[0:0] s1105, in1105_1, in1105_2;
    wire c1105;
    assign in1105_1 = {pp46[35]};
    assign in1105_2 = {pp47[34]};
    Full_Adder FA_1105(s1105, c1105, in1105_1, in1105_2, pp45[36]);
    wire[0:0] s1106, in1106_1, in1106_2;
    wire c1106;
    assign in1106_1 = {pp49[32]};
    assign in1106_2 = {pp50[31]};
    Full_Adder FA_1106(s1106, c1106, in1106_1, in1106_2, pp48[33]);
    wire[0:0] s1107, in1107_1, in1107_2;
    wire c1107;
    assign in1107_1 = {pp52[29]};
    assign in1107_2 = {pp53[28]};
    Full_Adder FA_1107(s1107, c1107, in1107_1, in1107_2, pp51[30]);
    wire[0:0] s1108, in1108_1, in1108_2;
    wire c1108;
    assign in1108_1 = {pp55[26]};
    assign in1108_2 = {pp56[25]};
    Full_Adder FA_1108(s1108, c1108, in1108_1, in1108_2, pp54[27]);
    wire[0:0] s1109, in1109_1, in1109_2;
    wire c1109;
    assign in1109_1 = {pp58[23]};
    assign in1109_2 = {pp59[22]};
    Full_Adder FA_1109(s1109, c1109, in1109_1, in1109_2, pp57[24]);
    wire[0:0] s1110, in1110_1, in1110_2;
    wire c1110;
    assign in1110_1 = {pp61[20]};
    assign in1110_2 = {pp62[19]};
    Full_Adder FA_1110(s1110, c1110, in1110_1, in1110_2, pp60[21]);
    wire[0:0] s1111, in1111_1, in1111_2;
    wire c1111;
    assign in1111_1 = {c448};
    assign in1111_2 = {c449};
    Full_Adder FA_1111(s1111, c1111, in1111_1, in1111_2, pp63[18]);
    wire[0:0] s1112, in1112_1, in1112_2;
    wire c1112;
    assign in1112_1 = {c451};
    assign in1112_2 = {c452};
    Full_Adder FA_1112(s1112, c1112, in1112_1, in1112_2, c450);
    wire[0:0] s1113, in1113_1, in1113_2;
    wire c1113;
    assign in1113_1 = {s454[0]};
    assign in1113_2 = {s455[0]};
    Full_Adder FA_1113(s1113, c1113, in1113_1, in1113_2, s453[0]);
    wire[0:0] s1114, in1114_1, in1114_2;
    wire c1114;
    assign in1114_1 = {pp29[53]};
    assign in1114_2 = {pp30[52]};
    Full_Adder FA_1114(s1114, c1114, in1114_1, in1114_2, pp28[54]);
    wire[0:0] s1115, in1115_1, in1115_2;
    wire c1115;
    assign in1115_1 = {pp32[50]};
    assign in1115_2 = {pp33[49]};
    Full_Adder FA_1115(s1115, c1115, in1115_1, in1115_2, pp31[51]);
    wire[0:0] s1116, in1116_1, in1116_2;
    wire c1116;
    assign in1116_1 = {pp35[47]};
    assign in1116_2 = {pp36[46]};
    Full_Adder FA_1116(s1116, c1116, in1116_1, in1116_2, pp34[48]);
    wire[0:0] s1117, in1117_1, in1117_2;
    wire c1117;
    assign in1117_1 = {pp38[44]};
    assign in1117_2 = {pp39[43]};
    Full_Adder FA_1117(s1117, c1117, in1117_1, in1117_2, pp37[45]);
    wire[0:0] s1118, in1118_1, in1118_2;
    wire c1118;
    assign in1118_1 = {pp41[41]};
    assign in1118_2 = {pp42[40]};
    Full_Adder FA_1118(s1118, c1118, in1118_1, in1118_2, pp40[42]);
    wire[0:0] s1119, in1119_1, in1119_2;
    wire c1119;
    assign in1119_1 = {pp44[38]};
    assign in1119_2 = {pp45[37]};
    Full_Adder FA_1119(s1119, c1119, in1119_1, in1119_2, pp43[39]);
    wire[0:0] s1120, in1120_1, in1120_2;
    wire c1120;
    assign in1120_1 = {pp47[35]};
    assign in1120_2 = {pp48[34]};
    Full_Adder FA_1120(s1120, c1120, in1120_1, in1120_2, pp46[36]);
    wire[0:0] s1121, in1121_1, in1121_2;
    wire c1121;
    assign in1121_1 = {pp50[32]};
    assign in1121_2 = {pp51[31]};
    Full_Adder FA_1121(s1121, c1121, in1121_1, in1121_2, pp49[33]);
    wire[0:0] s1122, in1122_1, in1122_2;
    wire c1122;
    assign in1122_1 = {pp53[29]};
    assign in1122_2 = {pp54[28]};
    Full_Adder FA_1122(s1122, c1122, in1122_1, in1122_2, pp52[30]);
    wire[0:0] s1123, in1123_1, in1123_2;
    wire c1123;
    assign in1123_1 = {pp56[26]};
    assign in1123_2 = {pp57[25]};
    Full_Adder FA_1123(s1123, c1123, in1123_1, in1123_2, pp55[27]);
    wire[0:0] s1124, in1124_1, in1124_2;
    wire c1124;
    assign in1124_1 = {pp59[23]};
    assign in1124_2 = {pp60[22]};
    Full_Adder FA_1124(s1124, c1124, in1124_1, in1124_2, pp58[24]);
    wire[0:0] s1125, in1125_1, in1125_2;
    wire c1125;
    assign in1125_1 = {pp62[20]};
    assign in1125_2 = {pp63[19]};
    Full_Adder FA_1125(s1125, c1125, in1125_1, in1125_2, pp61[21]);
    wire[0:0] s1126, in1126_1, in1126_2;
    wire c1126;
    assign in1126_1 = {c454};
    assign in1126_2 = {c455};
    Full_Adder FA_1126(s1126, c1126, in1126_1, in1126_2, c453);
    wire[0:0] s1127, in1127_1, in1127_2;
    wire c1127;
    assign in1127_1 = {s457[0]};
    assign in1127_2 = {s458[0]};
    Full_Adder FA_1127(s1127, c1127, in1127_1, in1127_2, c456);
    wire[0:0] s1128, in1128_1, in1128_2;
    wire c1128;
    assign in1128_1 = {pp27[56]};
    assign in1128_2 = {pp28[55]};
    Full_Adder FA_1128(s1128, c1128, in1128_1, in1128_2, pp26[57]);
    wire[0:0] s1129, in1129_1, in1129_2;
    wire c1129;
    assign in1129_1 = {pp30[53]};
    assign in1129_2 = {pp31[52]};
    Full_Adder FA_1129(s1129, c1129, in1129_1, in1129_2, pp29[54]);
    wire[0:0] s1130, in1130_1, in1130_2;
    wire c1130;
    assign in1130_1 = {pp33[50]};
    assign in1130_2 = {pp34[49]};
    Full_Adder FA_1130(s1130, c1130, in1130_1, in1130_2, pp32[51]);
    wire[0:0] s1131, in1131_1, in1131_2;
    wire c1131;
    assign in1131_1 = {pp36[47]};
    assign in1131_2 = {pp37[46]};
    Full_Adder FA_1131(s1131, c1131, in1131_1, in1131_2, pp35[48]);
    wire[0:0] s1132, in1132_1, in1132_2;
    wire c1132;
    assign in1132_1 = {pp39[44]};
    assign in1132_2 = {pp40[43]};
    Full_Adder FA_1132(s1132, c1132, in1132_1, in1132_2, pp38[45]);
    wire[0:0] s1133, in1133_1, in1133_2;
    wire c1133;
    assign in1133_1 = {pp42[41]};
    assign in1133_2 = {pp43[40]};
    Full_Adder FA_1133(s1133, c1133, in1133_1, in1133_2, pp41[42]);
    wire[0:0] s1134, in1134_1, in1134_2;
    wire c1134;
    assign in1134_1 = {pp45[38]};
    assign in1134_2 = {pp46[37]};
    Full_Adder FA_1134(s1134, c1134, in1134_1, in1134_2, pp44[39]);
    wire[0:0] s1135, in1135_1, in1135_2;
    wire c1135;
    assign in1135_1 = {pp48[35]};
    assign in1135_2 = {pp49[34]};
    Full_Adder FA_1135(s1135, c1135, in1135_1, in1135_2, pp47[36]);
    wire[0:0] s1136, in1136_1, in1136_2;
    wire c1136;
    assign in1136_1 = {pp51[32]};
    assign in1136_2 = {pp52[31]};
    Full_Adder FA_1136(s1136, c1136, in1136_1, in1136_2, pp50[33]);
    wire[0:0] s1137, in1137_1, in1137_2;
    wire c1137;
    assign in1137_1 = {pp54[29]};
    assign in1137_2 = {pp55[28]};
    Full_Adder FA_1137(s1137, c1137, in1137_1, in1137_2, pp53[30]);
    wire[0:0] s1138, in1138_1, in1138_2;
    wire c1138;
    assign in1138_1 = {pp57[26]};
    assign in1138_2 = {pp58[25]};
    Full_Adder FA_1138(s1138, c1138, in1138_1, in1138_2, pp56[27]);
    wire[0:0] s1139, in1139_1, in1139_2;
    wire c1139;
    assign in1139_1 = {pp60[23]};
    assign in1139_2 = {pp61[22]};
    Full_Adder FA_1139(s1139, c1139, in1139_1, in1139_2, pp59[24]);
    wire[0:0] s1140, in1140_1, in1140_2;
    wire c1140;
    assign in1140_1 = {pp63[20]};
    assign in1140_2 = {c457};
    Full_Adder FA_1140(s1140, c1140, in1140_1, in1140_2, pp62[21]);
    wire[0:0] s1141, in1141_1, in1141_2;
    wire c1141;
    assign in1141_1 = {c459};
    assign in1141_2 = {s460[0]};
    Full_Adder FA_1141(s1141, c1141, in1141_1, in1141_2, c458);
    wire[0:0] s1142, in1142_1, in1142_2;
    wire c1142;
    assign in1142_1 = {pp25[59]};
    assign in1142_2 = {pp26[58]};
    Full_Adder FA_1142(s1142, c1142, in1142_1, in1142_2, pp24[60]);
    wire[0:0] s1143, in1143_1, in1143_2;
    wire c1143;
    assign in1143_1 = {pp28[56]};
    assign in1143_2 = {pp29[55]};
    Full_Adder FA_1143(s1143, c1143, in1143_1, in1143_2, pp27[57]);
    wire[0:0] s1144, in1144_1, in1144_2;
    wire c1144;
    assign in1144_1 = {pp31[53]};
    assign in1144_2 = {pp32[52]};
    Full_Adder FA_1144(s1144, c1144, in1144_1, in1144_2, pp30[54]);
    wire[0:0] s1145, in1145_1, in1145_2;
    wire c1145;
    assign in1145_1 = {pp34[50]};
    assign in1145_2 = {pp35[49]};
    Full_Adder FA_1145(s1145, c1145, in1145_1, in1145_2, pp33[51]);
    wire[0:0] s1146, in1146_1, in1146_2;
    wire c1146;
    assign in1146_1 = {pp37[47]};
    assign in1146_2 = {pp38[46]};
    Full_Adder FA_1146(s1146, c1146, in1146_1, in1146_2, pp36[48]);
    wire[0:0] s1147, in1147_1, in1147_2;
    wire c1147;
    assign in1147_1 = {pp40[44]};
    assign in1147_2 = {pp41[43]};
    Full_Adder FA_1147(s1147, c1147, in1147_1, in1147_2, pp39[45]);
    wire[0:0] s1148, in1148_1, in1148_2;
    wire c1148;
    assign in1148_1 = {pp43[41]};
    assign in1148_2 = {pp44[40]};
    Full_Adder FA_1148(s1148, c1148, in1148_1, in1148_2, pp42[42]);
    wire[0:0] s1149, in1149_1, in1149_2;
    wire c1149;
    assign in1149_1 = {pp46[38]};
    assign in1149_2 = {pp47[37]};
    Full_Adder FA_1149(s1149, c1149, in1149_1, in1149_2, pp45[39]);
    wire[0:0] s1150, in1150_1, in1150_2;
    wire c1150;
    assign in1150_1 = {pp49[35]};
    assign in1150_2 = {pp50[34]};
    Full_Adder FA_1150(s1150, c1150, in1150_1, in1150_2, pp48[36]);
    wire[0:0] s1151, in1151_1, in1151_2;
    wire c1151;
    assign in1151_1 = {pp52[32]};
    assign in1151_2 = {pp53[31]};
    Full_Adder FA_1151(s1151, c1151, in1151_1, in1151_2, pp51[33]);
    wire[0:0] s1152, in1152_1, in1152_2;
    wire c1152;
    assign in1152_1 = {pp55[29]};
    assign in1152_2 = {pp56[28]};
    Full_Adder FA_1152(s1152, c1152, in1152_1, in1152_2, pp54[30]);
    wire[0:0] s1153, in1153_1, in1153_2;
    wire c1153;
    assign in1153_1 = {pp58[26]};
    assign in1153_2 = {pp59[25]};
    Full_Adder FA_1153(s1153, c1153, in1153_1, in1153_2, pp57[27]);
    wire[0:0] s1154, in1154_1, in1154_2;
    wire c1154;
    assign in1154_1 = {pp61[23]};
    assign in1154_2 = {pp62[22]};
    Full_Adder FA_1154(s1154, c1154, in1154_1, in1154_2, pp60[24]);
    wire[0:0] s1155, in1155_1, in1155_2;
    wire c1155;
    assign in1155_1 = {c460};
    assign in1155_2 = {c461};
    Full_Adder FA_1155(s1155, c1155, in1155_1, in1155_2, pp63[21]);
    wire[0:0] s1156, in1156_1, in1156_2;
    wire c1156;
    assign in1156_1 = {pp23[62]};
    assign in1156_2 = {pp24[61]};
    Full_Adder FA_1156(s1156, c1156, in1156_1, in1156_2, pp22[63]);
    wire[0:0] s1157, in1157_1, in1157_2;
    wire c1157;
    assign in1157_1 = {pp26[59]};
    assign in1157_2 = {pp27[58]};
    Full_Adder FA_1157(s1157, c1157, in1157_1, in1157_2, pp25[60]);
    wire[0:0] s1158, in1158_1, in1158_2;
    wire c1158;
    assign in1158_1 = {pp29[56]};
    assign in1158_2 = {pp30[55]};
    Full_Adder FA_1158(s1158, c1158, in1158_1, in1158_2, pp28[57]);
    wire[0:0] s1159, in1159_1, in1159_2;
    wire c1159;
    assign in1159_1 = {pp32[53]};
    assign in1159_2 = {pp33[52]};
    Full_Adder FA_1159(s1159, c1159, in1159_1, in1159_2, pp31[54]);
    wire[0:0] s1160, in1160_1, in1160_2;
    wire c1160;
    assign in1160_1 = {pp35[50]};
    assign in1160_2 = {pp36[49]};
    Full_Adder FA_1160(s1160, c1160, in1160_1, in1160_2, pp34[51]);
    wire[0:0] s1161, in1161_1, in1161_2;
    wire c1161;
    assign in1161_1 = {pp38[47]};
    assign in1161_2 = {pp39[46]};
    Full_Adder FA_1161(s1161, c1161, in1161_1, in1161_2, pp37[48]);
    wire[0:0] s1162, in1162_1, in1162_2;
    wire c1162;
    assign in1162_1 = {pp41[44]};
    assign in1162_2 = {pp42[43]};
    Full_Adder FA_1162(s1162, c1162, in1162_1, in1162_2, pp40[45]);
    wire[0:0] s1163, in1163_1, in1163_2;
    wire c1163;
    assign in1163_1 = {pp44[41]};
    assign in1163_2 = {pp45[40]};
    Full_Adder FA_1163(s1163, c1163, in1163_1, in1163_2, pp43[42]);
    wire[0:0] s1164, in1164_1, in1164_2;
    wire c1164;
    assign in1164_1 = {pp47[38]};
    assign in1164_2 = {pp48[37]};
    Full_Adder FA_1164(s1164, c1164, in1164_1, in1164_2, pp46[39]);
    wire[0:0] s1165, in1165_1, in1165_2;
    wire c1165;
    assign in1165_1 = {pp50[35]};
    assign in1165_2 = {pp51[34]};
    Full_Adder FA_1165(s1165, c1165, in1165_1, in1165_2, pp49[36]);
    wire[0:0] s1166, in1166_1, in1166_2;
    wire c1166;
    assign in1166_1 = {pp53[32]};
    assign in1166_2 = {pp54[31]};
    Full_Adder FA_1166(s1166, c1166, in1166_1, in1166_2, pp52[33]);
    wire[0:0] s1167, in1167_1, in1167_2;
    wire c1167;
    assign in1167_1 = {pp56[29]};
    assign in1167_2 = {pp57[28]};
    Full_Adder FA_1167(s1167, c1167, in1167_1, in1167_2, pp55[30]);
    wire[0:0] s1168, in1168_1, in1168_2;
    wire c1168;
    assign in1168_1 = {pp59[26]};
    assign in1168_2 = {pp60[25]};
    Full_Adder FA_1168(s1168, c1168, in1168_1, in1168_2, pp58[27]);
    wire[0:0] s1169, in1169_1, in1169_2;
    wire c1169;
    assign in1169_1 = {pp62[23]};
    assign in1169_2 = {pp63[22]};
    Full_Adder FA_1169(s1169, c1169, in1169_1, in1169_2, pp61[24]);
    wire[0:0] s1170, in1170_1, in1170_2;
    wire c1170;
    assign in1170_1 = {pp24[62]};
    assign in1170_2 = {pp25[61]};
    Full_Adder FA_1170(s1170, c1170, in1170_1, in1170_2, pp23[63]);
    wire[0:0] s1171, in1171_1, in1171_2;
    wire c1171;
    assign in1171_1 = {pp27[59]};
    assign in1171_2 = {pp28[58]};
    Full_Adder FA_1171(s1171, c1171, in1171_1, in1171_2, pp26[60]);
    wire[0:0] s1172, in1172_1, in1172_2;
    wire c1172;
    assign in1172_1 = {pp30[56]};
    assign in1172_2 = {pp31[55]};
    Full_Adder FA_1172(s1172, c1172, in1172_1, in1172_2, pp29[57]);
    wire[0:0] s1173, in1173_1, in1173_2;
    wire c1173;
    assign in1173_1 = {pp33[53]};
    assign in1173_2 = {pp34[52]};
    Full_Adder FA_1173(s1173, c1173, in1173_1, in1173_2, pp32[54]);
    wire[0:0] s1174, in1174_1, in1174_2;
    wire c1174;
    assign in1174_1 = {pp36[50]};
    assign in1174_2 = {pp37[49]};
    Full_Adder FA_1174(s1174, c1174, in1174_1, in1174_2, pp35[51]);
    wire[0:0] s1175, in1175_1, in1175_2;
    wire c1175;
    assign in1175_1 = {pp39[47]};
    assign in1175_2 = {pp40[46]};
    Full_Adder FA_1175(s1175, c1175, in1175_1, in1175_2, pp38[48]);
    wire[0:0] s1176, in1176_1, in1176_2;
    wire c1176;
    assign in1176_1 = {pp42[44]};
    assign in1176_2 = {pp43[43]};
    Full_Adder FA_1176(s1176, c1176, in1176_1, in1176_2, pp41[45]);
    wire[0:0] s1177, in1177_1, in1177_2;
    wire c1177;
    assign in1177_1 = {pp45[41]};
    assign in1177_2 = {pp46[40]};
    Full_Adder FA_1177(s1177, c1177, in1177_1, in1177_2, pp44[42]);
    wire[0:0] s1178, in1178_1, in1178_2;
    wire c1178;
    assign in1178_1 = {pp48[38]};
    assign in1178_2 = {pp49[37]};
    Full_Adder FA_1178(s1178, c1178, in1178_1, in1178_2, pp47[39]);
    wire[0:0] s1179, in1179_1, in1179_2;
    wire c1179;
    assign in1179_1 = {pp51[35]};
    assign in1179_2 = {pp52[34]};
    Full_Adder FA_1179(s1179, c1179, in1179_1, in1179_2, pp50[36]);
    wire[0:0] s1180, in1180_1, in1180_2;
    wire c1180;
    assign in1180_1 = {pp54[32]};
    assign in1180_2 = {pp55[31]};
    Full_Adder FA_1180(s1180, c1180, in1180_1, in1180_2, pp53[33]);
    wire[0:0] s1181, in1181_1, in1181_2;
    wire c1181;
    assign in1181_1 = {pp57[29]};
    assign in1181_2 = {pp58[28]};
    Full_Adder FA_1181(s1181, c1181, in1181_1, in1181_2, pp56[30]);
    wire[0:0] s1182, in1182_1, in1182_2;
    wire c1182;
    assign in1182_1 = {pp60[26]};
    assign in1182_2 = {pp61[25]};
    Full_Adder FA_1182(s1182, c1182, in1182_1, in1182_2, pp59[27]);
    wire[0:0] s1183, in1183_1, in1183_2;
    wire c1183;
    assign in1183_1 = {pp25[62]};
    assign in1183_2 = {pp26[61]};
    Full_Adder FA_1183(s1183, c1183, in1183_1, in1183_2, pp24[63]);
    wire[0:0] s1184, in1184_1, in1184_2;
    wire c1184;
    assign in1184_1 = {pp28[59]};
    assign in1184_2 = {pp29[58]};
    Full_Adder FA_1184(s1184, c1184, in1184_1, in1184_2, pp27[60]);
    wire[0:0] s1185, in1185_1, in1185_2;
    wire c1185;
    assign in1185_1 = {pp31[56]};
    assign in1185_2 = {pp32[55]};
    Full_Adder FA_1185(s1185, c1185, in1185_1, in1185_2, pp30[57]);
    wire[0:0] s1186, in1186_1, in1186_2;
    wire c1186;
    assign in1186_1 = {pp34[53]};
    assign in1186_2 = {pp35[52]};
    Full_Adder FA_1186(s1186, c1186, in1186_1, in1186_2, pp33[54]);
    wire[0:0] s1187, in1187_1, in1187_2;
    wire c1187;
    assign in1187_1 = {pp37[50]};
    assign in1187_2 = {pp38[49]};
    Full_Adder FA_1187(s1187, c1187, in1187_1, in1187_2, pp36[51]);
    wire[0:0] s1188, in1188_1, in1188_2;
    wire c1188;
    assign in1188_1 = {pp40[47]};
    assign in1188_2 = {pp41[46]};
    Full_Adder FA_1188(s1188, c1188, in1188_1, in1188_2, pp39[48]);
    wire[0:0] s1189, in1189_1, in1189_2;
    wire c1189;
    assign in1189_1 = {pp43[44]};
    assign in1189_2 = {pp44[43]};
    Full_Adder FA_1189(s1189, c1189, in1189_1, in1189_2, pp42[45]);
    wire[0:0] s1190, in1190_1, in1190_2;
    wire c1190;
    assign in1190_1 = {pp46[41]};
    assign in1190_2 = {pp47[40]};
    Full_Adder FA_1190(s1190, c1190, in1190_1, in1190_2, pp45[42]);
    wire[0:0] s1191, in1191_1, in1191_2;
    wire c1191;
    assign in1191_1 = {pp49[38]};
    assign in1191_2 = {pp50[37]};
    Full_Adder FA_1191(s1191, c1191, in1191_1, in1191_2, pp48[39]);
    wire[0:0] s1192, in1192_1, in1192_2;
    wire c1192;
    assign in1192_1 = {pp52[35]};
    assign in1192_2 = {pp53[34]};
    Full_Adder FA_1192(s1192, c1192, in1192_1, in1192_2, pp51[36]);
    wire[0:0] s1193, in1193_1, in1193_2;
    wire c1193;
    assign in1193_1 = {pp55[32]};
    assign in1193_2 = {pp56[31]};
    Full_Adder FA_1193(s1193, c1193, in1193_1, in1193_2, pp54[33]);
    wire[0:0] s1194, in1194_1, in1194_2;
    wire c1194;
    assign in1194_1 = {pp58[29]};
    assign in1194_2 = {pp59[28]};
    Full_Adder FA_1194(s1194, c1194, in1194_1, in1194_2, pp57[30]);
    wire[0:0] s1195, in1195_1, in1195_2;
    wire c1195;
    assign in1195_1 = {pp26[62]};
    assign in1195_2 = {pp27[61]};
    Full_Adder FA_1195(s1195, c1195, in1195_1, in1195_2, pp25[63]);
    wire[0:0] s1196, in1196_1, in1196_2;
    wire c1196;
    assign in1196_1 = {pp29[59]};
    assign in1196_2 = {pp30[58]};
    Full_Adder FA_1196(s1196, c1196, in1196_1, in1196_2, pp28[60]);
    wire[0:0] s1197, in1197_1, in1197_2;
    wire c1197;
    assign in1197_1 = {pp32[56]};
    assign in1197_2 = {pp33[55]};
    Full_Adder FA_1197(s1197, c1197, in1197_1, in1197_2, pp31[57]);
    wire[0:0] s1198, in1198_1, in1198_2;
    wire c1198;
    assign in1198_1 = {pp35[53]};
    assign in1198_2 = {pp36[52]};
    Full_Adder FA_1198(s1198, c1198, in1198_1, in1198_2, pp34[54]);
    wire[0:0] s1199, in1199_1, in1199_2;
    wire c1199;
    assign in1199_1 = {pp38[50]};
    assign in1199_2 = {pp39[49]};
    Full_Adder FA_1199(s1199, c1199, in1199_1, in1199_2, pp37[51]);
    wire[0:0] s1200, in1200_1, in1200_2;
    wire c1200;
    assign in1200_1 = {pp41[47]};
    assign in1200_2 = {pp42[46]};
    Full_Adder FA_1200(s1200, c1200, in1200_1, in1200_2, pp40[48]);
    wire[0:0] s1201, in1201_1, in1201_2;
    wire c1201;
    assign in1201_1 = {pp44[44]};
    assign in1201_2 = {pp45[43]};
    Full_Adder FA_1201(s1201, c1201, in1201_1, in1201_2, pp43[45]);
    wire[0:0] s1202, in1202_1, in1202_2;
    wire c1202;
    assign in1202_1 = {pp47[41]};
    assign in1202_2 = {pp48[40]};
    Full_Adder FA_1202(s1202, c1202, in1202_1, in1202_2, pp46[42]);
    wire[0:0] s1203, in1203_1, in1203_2;
    wire c1203;
    assign in1203_1 = {pp50[38]};
    assign in1203_2 = {pp51[37]};
    Full_Adder FA_1203(s1203, c1203, in1203_1, in1203_2, pp49[39]);
    wire[0:0] s1204, in1204_1, in1204_2;
    wire c1204;
    assign in1204_1 = {pp53[35]};
    assign in1204_2 = {pp54[34]};
    Full_Adder FA_1204(s1204, c1204, in1204_1, in1204_2, pp52[36]);
    wire[0:0] s1205, in1205_1, in1205_2;
    wire c1205;
    assign in1205_1 = {pp56[32]};
    assign in1205_2 = {pp57[31]};
    Full_Adder FA_1205(s1205, c1205, in1205_1, in1205_2, pp55[33]);
    wire[0:0] s1206, in1206_1, in1206_2;
    wire c1206;
    assign in1206_1 = {pp27[62]};
    assign in1206_2 = {pp28[61]};
    Full_Adder FA_1206(s1206, c1206, in1206_1, in1206_2, pp26[63]);
    wire[0:0] s1207, in1207_1, in1207_2;
    wire c1207;
    assign in1207_1 = {pp30[59]};
    assign in1207_2 = {pp31[58]};
    Full_Adder FA_1207(s1207, c1207, in1207_1, in1207_2, pp29[60]);
    wire[0:0] s1208, in1208_1, in1208_2;
    wire c1208;
    assign in1208_1 = {pp33[56]};
    assign in1208_2 = {pp34[55]};
    Full_Adder FA_1208(s1208, c1208, in1208_1, in1208_2, pp32[57]);
    wire[0:0] s1209, in1209_1, in1209_2;
    wire c1209;
    assign in1209_1 = {pp36[53]};
    assign in1209_2 = {pp37[52]};
    Full_Adder FA_1209(s1209, c1209, in1209_1, in1209_2, pp35[54]);
    wire[0:0] s1210, in1210_1, in1210_2;
    wire c1210;
    assign in1210_1 = {pp39[50]};
    assign in1210_2 = {pp40[49]};
    Full_Adder FA_1210(s1210, c1210, in1210_1, in1210_2, pp38[51]);
    wire[0:0] s1211, in1211_1, in1211_2;
    wire c1211;
    assign in1211_1 = {pp42[47]};
    assign in1211_2 = {pp43[46]};
    Full_Adder FA_1211(s1211, c1211, in1211_1, in1211_2, pp41[48]);
    wire[0:0] s1212, in1212_1, in1212_2;
    wire c1212;
    assign in1212_1 = {pp45[44]};
    assign in1212_2 = {pp46[43]};
    Full_Adder FA_1212(s1212, c1212, in1212_1, in1212_2, pp44[45]);
    wire[0:0] s1213, in1213_1, in1213_2;
    wire c1213;
    assign in1213_1 = {pp48[41]};
    assign in1213_2 = {pp49[40]};
    Full_Adder FA_1213(s1213, c1213, in1213_1, in1213_2, pp47[42]);
    wire[0:0] s1214, in1214_1, in1214_2;
    wire c1214;
    assign in1214_1 = {pp51[38]};
    assign in1214_2 = {pp52[37]};
    Full_Adder FA_1214(s1214, c1214, in1214_1, in1214_2, pp50[39]);
    wire[0:0] s1215, in1215_1, in1215_2;
    wire c1215;
    assign in1215_1 = {pp54[35]};
    assign in1215_2 = {pp55[34]};
    Full_Adder FA_1215(s1215, c1215, in1215_1, in1215_2, pp53[36]);
    wire[0:0] s1216, in1216_1, in1216_2;
    wire c1216;
    assign in1216_1 = {pp28[62]};
    assign in1216_2 = {pp29[61]};
    Full_Adder FA_1216(s1216, c1216, in1216_1, in1216_2, pp27[63]);
    wire[0:0] s1217, in1217_1, in1217_2;
    wire c1217;
    assign in1217_1 = {pp31[59]};
    assign in1217_2 = {pp32[58]};
    Full_Adder FA_1217(s1217, c1217, in1217_1, in1217_2, pp30[60]);
    wire[0:0] s1218, in1218_1, in1218_2;
    wire c1218;
    assign in1218_1 = {pp34[56]};
    assign in1218_2 = {pp35[55]};
    Full_Adder FA_1218(s1218, c1218, in1218_1, in1218_2, pp33[57]);
    wire[0:0] s1219, in1219_1, in1219_2;
    wire c1219;
    assign in1219_1 = {pp37[53]};
    assign in1219_2 = {pp38[52]};
    Full_Adder FA_1219(s1219, c1219, in1219_1, in1219_2, pp36[54]);
    wire[0:0] s1220, in1220_1, in1220_2;
    wire c1220;
    assign in1220_1 = {pp40[50]};
    assign in1220_2 = {pp41[49]};
    Full_Adder FA_1220(s1220, c1220, in1220_1, in1220_2, pp39[51]);
    wire[0:0] s1221, in1221_1, in1221_2;
    wire c1221;
    assign in1221_1 = {pp43[47]};
    assign in1221_2 = {pp44[46]};
    Full_Adder FA_1221(s1221, c1221, in1221_1, in1221_2, pp42[48]);
    wire[0:0] s1222, in1222_1, in1222_2;
    wire c1222;
    assign in1222_1 = {pp46[44]};
    assign in1222_2 = {pp47[43]};
    Full_Adder FA_1222(s1222, c1222, in1222_1, in1222_2, pp45[45]);
    wire[0:0] s1223, in1223_1, in1223_2;
    wire c1223;
    assign in1223_1 = {pp49[41]};
    assign in1223_2 = {pp50[40]};
    Full_Adder FA_1223(s1223, c1223, in1223_1, in1223_2, pp48[42]);
    wire[0:0] s1224, in1224_1, in1224_2;
    wire c1224;
    assign in1224_1 = {pp52[38]};
    assign in1224_2 = {pp53[37]};
    Full_Adder FA_1224(s1224, c1224, in1224_1, in1224_2, pp51[39]);
    wire[0:0] s1225, in1225_1, in1225_2;
    wire c1225;
    assign in1225_1 = {pp29[62]};
    assign in1225_2 = {pp30[61]};
    Full_Adder FA_1225(s1225, c1225, in1225_1, in1225_2, pp28[63]);
    wire[0:0] s1226, in1226_1, in1226_2;
    wire c1226;
    assign in1226_1 = {pp32[59]};
    assign in1226_2 = {pp33[58]};
    Full_Adder FA_1226(s1226, c1226, in1226_1, in1226_2, pp31[60]);
    wire[0:0] s1227, in1227_1, in1227_2;
    wire c1227;
    assign in1227_1 = {pp35[56]};
    assign in1227_2 = {pp36[55]};
    Full_Adder FA_1227(s1227, c1227, in1227_1, in1227_2, pp34[57]);
    wire[0:0] s1228, in1228_1, in1228_2;
    wire c1228;
    assign in1228_1 = {pp38[53]};
    assign in1228_2 = {pp39[52]};
    Full_Adder FA_1228(s1228, c1228, in1228_1, in1228_2, pp37[54]);
    wire[0:0] s1229, in1229_1, in1229_2;
    wire c1229;
    assign in1229_1 = {pp41[50]};
    assign in1229_2 = {pp42[49]};
    Full_Adder FA_1229(s1229, c1229, in1229_1, in1229_2, pp40[51]);
    wire[0:0] s1230, in1230_1, in1230_2;
    wire c1230;
    assign in1230_1 = {pp44[47]};
    assign in1230_2 = {pp45[46]};
    Full_Adder FA_1230(s1230, c1230, in1230_1, in1230_2, pp43[48]);
    wire[0:0] s1231, in1231_1, in1231_2;
    wire c1231;
    assign in1231_1 = {pp47[44]};
    assign in1231_2 = {pp48[43]};
    Full_Adder FA_1231(s1231, c1231, in1231_1, in1231_2, pp46[45]);
    wire[0:0] s1232, in1232_1, in1232_2;
    wire c1232;
    assign in1232_1 = {pp50[41]};
    assign in1232_2 = {pp51[40]};
    Full_Adder FA_1232(s1232, c1232, in1232_1, in1232_2, pp49[42]);
    wire[0:0] s1233, in1233_1, in1233_2;
    wire c1233;
    assign in1233_1 = {pp30[62]};
    assign in1233_2 = {pp31[61]};
    Full_Adder FA_1233(s1233, c1233, in1233_1, in1233_2, pp29[63]);
    wire[0:0] s1234, in1234_1, in1234_2;
    wire c1234;
    assign in1234_1 = {pp33[59]};
    assign in1234_2 = {pp34[58]};
    Full_Adder FA_1234(s1234, c1234, in1234_1, in1234_2, pp32[60]);
    wire[0:0] s1235, in1235_1, in1235_2;
    wire c1235;
    assign in1235_1 = {pp36[56]};
    assign in1235_2 = {pp37[55]};
    Full_Adder FA_1235(s1235, c1235, in1235_1, in1235_2, pp35[57]);
    wire[0:0] s1236, in1236_1, in1236_2;
    wire c1236;
    assign in1236_1 = {pp39[53]};
    assign in1236_2 = {pp40[52]};
    Full_Adder FA_1236(s1236, c1236, in1236_1, in1236_2, pp38[54]);
    wire[0:0] s1237, in1237_1, in1237_2;
    wire c1237;
    assign in1237_1 = {pp42[50]};
    assign in1237_2 = {pp43[49]};
    Full_Adder FA_1237(s1237, c1237, in1237_1, in1237_2, pp41[51]);
    wire[0:0] s1238, in1238_1, in1238_2;
    wire c1238;
    assign in1238_1 = {pp45[47]};
    assign in1238_2 = {pp46[46]};
    Full_Adder FA_1238(s1238, c1238, in1238_1, in1238_2, pp44[48]);
    wire[0:0] s1239, in1239_1, in1239_2;
    wire c1239;
    assign in1239_1 = {pp48[44]};
    assign in1239_2 = {pp49[43]};
    Full_Adder FA_1239(s1239, c1239, in1239_1, in1239_2, pp47[45]);
    wire[0:0] s1240, in1240_1, in1240_2;
    wire c1240;
    assign in1240_1 = {pp31[62]};
    assign in1240_2 = {pp32[61]};
    Full_Adder FA_1240(s1240, c1240, in1240_1, in1240_2, pp30[63]);
    wire[0:0] s1241, in1241_1, in1241_2;
    wire c1241;
    assign in1241_1 = {pp34[59]};
    assign in1241_2 = {pp35[58]};
    Full_Adder FA_1241(s1241, c1241, in1241_1, in1241_2, pp33[60]);
    wire[0:0] s1242, in1242_1, in1242_2;
    wire c1242;
    assign in1242_1 = {pp37[56]};
    assign in1242_2 = {pp38[55]};
    Full_Adder FA_1242(s1242, c1242, in1242_1, in1242_2, pp36[57]);
    wire[0:0] s1243, in1243_1, in1243_2;
    wire c1243;
    assign in1243_1 = {pp40[53]};
    assign in1243_2 = {pp41[52]};
    Full_Adder FA_1243(s1243, c1243, in1243_1, in1243_2, pp39[54]);
    wire[0:0] s1244, in1244_1, in1244_2;
    wire c1244;
    assign in1244_1 = {pp43[50]};
    assign in1244_2 = {pp44[49]};
    Full_Adder FA_1244(s1244, c1244, in1244_1, in1244_2, pp42[51]);
    wire[0:0] s1245, in1245_1, in1245_2;
    wire c1245;
    assign in1245_1 = {pp46[47]};
    assign in1245_2 = {pp47[46]};
    Full_Adder FA_1245(s1245, c1245, in1245_1, in1245_2, pp45[48]);
    wire[0:0] s1246, in1246_1, in1246_2;
    wire c1246;
    assign in1246_1 = {pp32[62]};
    assign in1246_2 = {pp33[61]};
    Full_Adder FA_1246(s1246, c1246, in1246_1, in1246_2, pp31[63]);
    wire[0:0] s1247, in1247_1, in1247_2;
    wire c1247;
    assign in1247_1 = {pp35[59]};
    assign in1247_2 = {pp36[58]};
    Full_Adder FA_1247(s1247, c1247, in1247_1, in1247_2, pp34[60]);
    wire[0:0] s1248, in1248_1, in1248_2;
    wire c1248;
    assign in1248_1 = {pp38[56]};
    assign in1248_2 = {pp39[55]};
    Full_Adder FA_1248(s1248, c1248, in1248_1, in1248_2, pp37[57]);
    wire[0:0] s1249, in1249_1, in1249_2;
    wire c1249;
    assign in1249_1 = {pp41[53]};
    assign in1249_2 = {pp42[52]};
    Full_Adder FA_1249(s1249, c1249, in1249_1, in1249_2, pp40[54]);
    wire[0:0] s1250, in1250_1, in1250_2;
    wire c1250;
    assign in1250_1 = {pp44[50]};
    assign in1250_2 = {pp45[49]};
    Full_Adder FA_1250(s1250, c1250, in1250_1, in1250_2, pp43[51]);
    wire[0:0] s1251, in1251_1, in1251_2;
    wire c1251;
    assign in1251_1 = {pp33[62]};
    assign in1251_2 = {pp34[61]};
    Full_Adder FA_1251(s1251, c1251, in1251_1, in1251_2, pp32[63]);
    wire[0:0] s1252, in1252_1, in1252_2;
    wire c1252;
    assign in1252_1 = {pp36[59]};
    assign in1252_2 = {pp37[58]};
    Full_Adder FA_1252(s1252, c1252, in1252_1, in1252_2, pp35[60]);
    wire[0:0] s1253, in1253_1, in1253_2;
    wire c1253;
    assign in1253_1 = {pp39[56]};
    assign in1253_2 = {pp40[55]};
    Full_Adder FA_1253(s1253, c1253, in1253_1, in1253_2, pp38[57]);
    wire[0:0] s1254, in1254_1, in1254_2;
    wire c1254;
    assign in1254_1 = {pp42[53]};
    assign in1254_2 = {pp43[52]};
    Full_Adder FA_1254(s1254, c1254, in1254_1, in1254_2, pp41[54]);
    wire[0:0] s1255, in1255_1, in1255_2;
    wire c1255;
    assign in1255_1 = {pp34[62]};
    assign in1255_2 = {pp35[61]};
    Full_Adder FA_1255(s1255, c1255, in1255_1, in1255_2, pp33[63]);
    wire[0:0] s1256, in1256_1, in1256_2;
    wire c1256;
    assign in1256_1 = {pp37[59]};
    assign in1256_2 = {pp38[58]};
    Full_Adder FA_1256(s1256, c1256, in1256_1, in1256_2, pp36[60]);
    wire[0:0] s1257, in1257_1, in1257_2;
    wire c1257;
    assign in1257_1 = {pp40[56]};
    assign in1257_2 = {pp41[55]};
    Full_Adder FA_1257(s1257, c1257, in1257_1, in1257_2, pp39[57]);
    wire[0:0] s1258, in1258_1, in1258_2;
    wire c1258;
    assign in1258_1 = {pp35[62]};
    assign in1258_2 = {pp36[61]};
    Full_Adder FA_1258(s1258, c1258, in1258_1, in1258_2, pp34[63]);
    wire[0:0] s1259, in1259_1, in1259_2;
    wire c1259;
    assign in1259_1 = {pp38[59]};
    assign in1259_2 = {pp39[58]};
    Full_Adder FA_1259(s1259, c1259, in1259_1, in1259_2, pp37[60]);
    wire[0:0] s1260, in1260_1, in1260_2;
    wire c1260;
    assign in1260_1 = {pp36[62]};
    assign in1260_2 = {pp37[61]};
    Full_Adder FA_1260(s1260, c1260, in1260_1, in1260_2, pp35[63]);

    /*Stage 3*/
    wire[0:0] s1261, in1261_1, in1261_2;
    wire c1261;
    assign in1261_1 = {pp0[20]};
    assign in1261_2 = {pp1[19]};
    Half_Adder HA_1261(s1261, c1261, in1261_1, in1261_2);
    wire[0:0] s1262, in1262_1, in1262_2;
    wire c1262;
    assign in1262_1 = {pp1[20]};
    assign in1262_2 = {pp2[19]};
    Full_Adder FA_1262(s1262, c1262, in1262_1, in1262_2, pp0[21]);
    wire[0:0] s1263, in1263_1, in1263_2;
    wire c1263;
    assign in1263_1 = {pp3[18]};
    assign in1263_2 = {pp4[17]};
    Half_Adder HA_1263(s1263, c1263, in1263_1, in1263_2);
    wire[0:0] s1264, in1264_1, in1264_2;
    wire c1264;
    assign in1264_1 = {pp1[21]};
    assign in1264_2 = {pp2[20]};
    Full_Adder FA_1264(s1264, c1264, in1264_1, in1264_2, pp0[22]);
    wire[0:0] s1265, in1265_1, in1265_2;
    wire c1265;
    assign in1265_1 = {pp4[18]};
    assign in1265_2 = {pp5[17]};
    Full_Adder FA_1265(s1265, c1265, in1265_1, in1265_2, pp3[19]);
    wire[0:0] s1266, in1266_1, in1266_2;
    wire c1266;
    assign in1266_1 = {pp6[16]};
    assign in1266_2 = {pp7[15]};
    Half_Adder HA_1266(s1266, c1266, in1266_1, in1266_2);
    wire[0:0] s1267, in1267_1, in1267_2;
    wire c1267;
    assign in1267_1 = {pp1[22]};
    assign in1267_2 = {pp2[21]};
    Full_Adder FA_1267(s1267, c1267, in1267_1, in1267_2, pp0[23]);
    wire[0:0] s1268, in1268_1, in1268_2;
    wire c1268;
    assign in1268_1 = {pp4[19]};
    assign in1268_2 = {pp5[18]};
    Full_Adder FA_1268(s1268, c1268, in1268_1, in1268_2, pp3[20]);
    wire[0:0] s1269, in1269_1, in1269_2;
    wire c1269;
    assign in1269_1 = {pp7[16]};
    assign in1269_2 = {pp8[15]};
    Full_Adder FA_1269(s1269, c1269, in1269_1, in1269_2, pp6[17]);
    wire[0:0] s1270, in1270_1, in1270_2;
    wire c1270;
    assign in1270_1 = {pp9[14]};
    assign in1270_2 = {pp10[13]};
    Half_Adder HA_1270(s1270, c1270, in1270_1, in1270_2);
    wire[0:0] s1271, in1271_1, in1271_2;
    wire c1271;
    assign in1271_1 = {pp1[23]};
    assign in1271_2 = {pp2[22]};
    Full_Adder FA_1271(s1271, c1271, in1271_1, in1271_2, pp0[24]);
    wire[0:0] s1272, in1272_1, in1272_2;
    wire c1272;
    assign in1272_1 = {pp4[20]};
    assign in1272_2 = {pp5[19]};
    Full_Adder FA_1272(s1272, c1272, in1272_1, in1272_2, pp3[21]);
    wire[0:0] s1273, in1273_1, in1273_2;
    wire c1273;
    assign in1273_1 = {pp7[17]};
    assign in1273_2 = {pp8[16]};
    Full_Adder FA_1273(s1273, c1273, in1273_1, in1273_2, pp6[18]);
    wire[0:0] s1274, in1274_1, in1274_2;
    wire c1274;
    assign in1274_1 = {pp10[14]};
    assign in1274_2 = {pp11[13]};
    Full_Adder FA_1274(s1274, c1274, in1274_1, in1274_2, pp9[15]);
    wire[0:0] s1275, in1275_1, in1275_2;
    wire c1275;
    assign in1275_1 = {pp12[12]};
    assign in1275_2 = {pp13[11]};
    Half_Adder HA_1275(s1275, c1275, in1275_1, in1275_2);
    wire[0:0] s1276, in1276_1, in1276_2;
    wire c1276;
    assign in1276_1 = {pp1[24]};
    assign in1276_2 = {pp2[23]};
    Full_Adder FA_1276(s1276, c1276, in1276_1, in1276_2, pp0[25]);
    wire[0:0] s1277, in1277_1, in1277_2;
    wire c1277;
    assign in1277_1 = {pp4[21]};
    assign in1277_2 = {pp5[20]};
    Full_Adder FA_1277(s1277, c1277, in1277_1, in1277_2, pp3[22]);
    wire[0:0] s1278, in1278_1, in1278_2;
    wire c1278;
    assign in1278_1 = {pp7[18]};
    assign in1278_2 = {pp8[17]};
    Full_Adder FA_1278(s1278, c1278, in1278_1, in1278_2, pp6[19]);
    wire[0:0] s1279, in1279_1, in1279_2;
    wire c1279;
    assign in1279_1 = {pp10[15]};
    assign in1279_2 = {pp11[14]};
    Full_Adder FA_1279(s1279, c1279, in1279_1, in1279_2, pp9[16]);
    wire[0:0] s1280, in1280_1, in1280_2;
    wire c1280;
    assign in1280_1 = {pp13[12]};
    assign in1280_2 = {pp14[11]};
    Full_Adder FA_1280(s1280, c1280, in1280_1, in1280_2, pp12[13]);
    wire[0:0] s1281, in1281_1, in1281_2;
    wire c1281;
    assign in1281_1 = {pp15[10]};
    assign in1281_2 = {pp16[9]};
    Half_Adder HA_1281(s1281, c1281, in1281_1, in1281_2);
    wire[0:0] s1282, in1282_1, in1282_2;
    wire c1282;
    assign in1282_1 = {pp1[25]};
    assign in1282_2 = {pp2[24]};
    Full_Adder FA_1282(s1282, c1282, in1282_1, in1282_2, pp0[26]);
    wire[0:0] s1283, in1283_1, in1283_2;
    wire c1283;
    assign in1283_1 = {pp4[22]};
    assign in1283_2 = {pp5[21]};
    Full_Adder FA_1283(s1283, c1283, in1283_1, in1283_2, pp3[23]);
    wire[0:0] s1284, in1284_1, in1284_2;
    wire c1284;
    assign in1284_1 = {pp7[19]};
    assign in1284_2 = {pp8[18]};
    Full_Adder FA_1284(s1284, c1284, in1284_1, in1284_2, pp6[20]);
    wire[0:0] s1285, in1285_1, in1285_2;
    wire c1285;
    assign in1285_1 = {pp10[16]};
    assign in1285_2 = {pp11[15]};
    Full_Adder FA_1285(s1285, c1285, in1285_1, in1285_2, pp9[17]);
    wire[0:0] s1286, in1286_1, in1286_2;
    wire c1286;
    assign in1286_1 = {pp13[13]};
    assign in1286_2 = {pp14[12]};
    Full_Adder FA_1286(s1286, c1286, in1286_1, in1286_2, pp12[14]);
    wire[0:0] s1287, in1287_1, in1287_2;
    wire c1287;
    assign in1287_1 = {pp16[10]};
    assign in1287_2 = {pp17[9]};
    Full_Adder FA_1287(s1287, c1287, in1287_1, in1287_2, pp15[11]);
    wire[0:0] s1288, in1288_1, in1288_2;
    wire c1288;
    assign in1288_1 = {pp18[8]};
    assign in1288_2 = {pp19[7]};
    Half_Adder HA_1288(s1288, c1288, in1288_1, in1288_2);
    wire[0:0] s1289, in1289_1, in1289_2;
    wire c1289;
    assign in1289_1 = {pp1[26]};
    assign in1289_2 = {pp2[25]};
    Full_Adder FA_1289(s1289, c1289, in1289_1, in1289_2, pp0[27]);
    wire[0:0] s1290, in1290_1, in1290_2;
    wire c1290;
    assign in1290_1 = {pp4[23]};
    assign in1290_2 = {pp5[22]};
    Full_Adder FA_1290(s1290, c1290, in1290_1, in1290_2, pp3[24]);
    wire[0:0] s1291, in1291_1, in1291_2;
    wire c1291;
    assign in1291_1 = {pp7[20]};
    assign in1291_2 = {pp8[19]};
    Full_Adder FA_1291(s1291, c1291, in1291_1, in1291_2, pp6[21]);
    wire[0:0] s1292, in1292_1, in1292_2;
    wire c1292;
    assign in1292_1 = {pp10[17]};
    assign in1292_2 = {pp11[16]};
    Full_Adder FA_1292(s1292, c1292, in1292_1, in1292_2, pp9[18]);
    wire[0:0] s1293, in1293_1, in1293_2;
    wire c1293;
    assign in1293_1 = {pp13[14]};
    assign in1293_2 = {pp14[13]};
    Full_Adder FA_1293(s1293, c1293, in1293_1, in1293_2, pp12[15]);
    wire[0:0] s1294, in1294_1, in1294_2;
    wire c1294;
    assign in1294_1 = {pp16[11]};
    assign in1294_2 = {pp17[10]};
    Full_Adder FA_1294(s1294, c1294, in1294_1, in1294_2, pp15[12]);
    wire[0:0] s1295, in1295_1, in1295_2;
    wire c1295;
    assign in1295_1 = {pp19[8]};
    assign in1295_2 = {pp20[7]};
    Full_Adder FA_1295(s1295, c1295, in1295_1, in1295_2, pp18[9]);
    wire[0:0] s1296, in1296_1, in1296_2;
    wire c1296;
    assign in1296_1 = {pp21[6]};
    assign in1296_2 = {pp22[5]};
    Half_Adder HA_1296(s1296, c1296, in1296_1, in1296_2);
    wire[0:0] s1297, in1297_1, in1297_2;
    wire c1297;
    assign in1297_1 = {pp1[27]};
    assign in1297_2 = {pp2[26]};
    Full_Adder FA_1297(s1297, c1297, in1297_1, in1297_2, pp0[28]);
    wire[0:0] s1298, in1298_1, in1298_2;
    wire c1298;
    assign in1298_1 = {pp4[24]};
    assign in1298_2 = {pp5[23]};
    Full_Adder FA_1298(s1298, c1298, in1298_1, in1298_2, pp3[25]);
    wire[0:0] s1299, in1299_1, in1299_2;
    wire c1299;
    assign in1299_1 = {pp7[21]};
    assign in1299_2 = {pp8[20]};
    Full_Adder FA_1299(s1299, c1299, in1299_1, in1299_2, pp6[22]);
    wire[0:0] s1300, in1300_1, in1300_2;
    wire c1300;
    assign in1300_1 = {pp10[18]};
    assign in1300_2 = {pp11[17]};
    Full_Adder FA_1300(s1300, c1300, in1300_1, in1300_2, pp9[19]);
    wire[0:0] s1301, in1301_1, in1301_2;
    wire c1301;
    assign in1301_1 = {pp13[15]};
    assign in1301_2 = {pp14[14]};
    Full_Adder FA_1301(s1301, c1301, in1301_1, in1301_2, pp12[16]);
    wire[0:0] s1302, in1302_1, in1302_2;
    wire c1302;
    assign in1302_1 = {pp16[12]};
    assign in1302_2 = {pp17[11]};
    Full_Adder FA_1302(s1302, c1302, in1302_1, in1302_2, pp15[13]);
    wire[0:0] s1303, in1303_1, in1303_2;
    wire c1303;
    assign in1303_1 = {pp19[9]};
    assign in1303_2 = {pp20[8]};
    Full_Adder FA_1303(s1303, c1303, in1303_1, in1303_2, pp18[10]);
    wire[0:0] s1304, in1304_1, in1304_2;
    wire c1304;
    assign in1304_1 = {pp22[6]};
    assign in1304_2 = {pp23[5]};
    Full_Adder FA_1304(s1304, c1304, in1304_1, in1304_2, pp21[7]);
    wire[0:0] s1305, in1305_1, in1305_2;
    wire c1305;
    assign in1305_1 = {pp24[4]};
    assign in1305_2 = {pp25[3]};
    Half_Adder HA_1305(s1305, c1305, in1305_1, in1305_2);
    wire[0:0] s1306, in1306_1, in1306_2;
    wire c1306;
    assign in1306_1 = {pp3[26]};
    assign in1306_2 = {pp4[25]};
    Full_Adder FA_1306(s1306, c1306, in1306_1, in1306_2, pp2[27]);
    wire[0:0] s1307, in1307_1, in1307_2;
    wire c1307;
    assign in1307_1 = {pp6[23]};
    assign in1307_2 = {pp7[22]};
    Full_Adder FA_1307(s1307, c1307, in1307_1, in1307_2, pp5[24]);
    wire[0:0] s1308, in1308_1, in1308_2;
    wire c1308;
    assign in1308_1 = {pp9[20]};
    assign in1308_2 = {pp10[19]};
    Full_Adder FA_1308(s1308, c1308, in1308_1, in1308_2, pp8[21]);
    wire[0:0] s1309, in1309_1, in1309_2;
    wire c1309;
    assign in1309_1 = {pp12[17]};
    assign in1309_2 = {pp13[16]};
    Full_Adder FA_1309(s1309, c1309, in1309_1, in1309_2, pp11[18]);
    wire[0:0] s1310, in1310_1, in1310_2;
    wire c1310;
    assign in1310_1 = {pp15[14]};
    assign in1310_2 = {pp16[13]};
    Full_Adder FA_1310(s1310, c1310, in1310_1, in1310_2, pp14[15]);
    wire[0:0] s1311, in1311_1, in1311_2;
    wire c1311;
    assign in1311_1 = {pp18[11]};
    assign in1311_2 = {pp19[10]};
    Full_Adder FA_1311(s1311, c1311, in1311_1, in1311_2, pp17[12]);
    wire[0:0] s1312, in1312_1, in1312_2;
    wire c1312;
    assign in1312_1 = {pp21[8]};
    assign in1312_2 = {pp22[7]};
    Full_Adder FA_1312(s1312, c1312, in1312_1, in1312_2, pp20[9]);
    wire[0:0] s1313, in1313_1, in1313_2;
    wire c1313;
    assign in1313_1 = {pp24[5]};
    assign in1313_2 = {pp25[4]};
    Full_Adder FA_1313(s1313, c1313, in1313_1, in1313_2, pp23[6]);
    wire[0:0] s1314, in1314_1, in1314_2;
    wire c1314;
    assign in1314_1 = {pp27[2]};
    assign in1314_2 = {pp28[1]};
    Full_Adder FA_1314(s1314, c1314, in1314_1, in1314_2, pp26[3]);
    wire[0:0] s1315, in1315_1, in1315_2;
    wire c1315;
    assign in1315_1 = {pp6[24]};
    assign in1315_2 = {pp7[23]};
    Full_Adder FA_1315(s1315, c1315, in1315_1, in1315_2, pp5[25]);
    wire[0:0] s1316, in1316_1, in1316_2;
    wire c1316;
    assign in1316_1 = {pp9[21]};
    assign in1316_2 = {pp10[20]};
    Full_Adder FA_1316(s1316, c1316, in1316_1, in1316_2, pp8[22]);
    wire[0:0] s1317, in1317_1, in1317_2;
    wire c1317;
    assign in1317_1 = {pp12[18]};
    assign in1317_2 = {pp13[17]};
    Full_Adder FA_1317(s1317, c1317, in1317_1, in1317_2, pp11[19]);
    wire[0:0] s1318, in1318_1, in1318_2;
    wire c1318;
    assign in1318_1 = {pp15[15]};
    assign in1318_2 = {pp16[14]};
    Full_Adder FA_1318(s1318, c1318, in1318_1, in1318_2, pp14[16]);
    wire[0:0] s1319, in1319_1, in1319_2;
    wire c1319;
    assign in1319_1 = {pp18[12]};
    assign in1319_2 = {pp19[11]};
    Full_Adder FA_1319(s1319, c1319, in1319_1, in1319_2, pp17[13]);
    wire[0:0] s1320, in1320_1, in1320_2;
    wire c1320;
    assign in1320_1 = {pp21[9]};
    assign in1320_2 = {pp22[8]};
    Full_Adder FA_1320(s1320, c1320, in1320_1, in1320_2, pp20[10]);
    wire[0:0] s1321, in1321_1, in1321_2;
    wire c1321;
    assign in1321_1 = {pp24[6]};
    assign in1321_2 = {pp25[5]};
    Full_Adder FA_1321(s1321, c1321, in1321_1, in1321_2, pp23[7]);
    wire[0:0] s1322, in1322_1, in1322_2;
    wire c1322;
    assign in1322_1 = {pp27[3]};
    assign in1322_2 = {pp28[2]};
    Full_Adder FA_1322(s1322, c1322, in1322_1, in1322_2, pp26[4]);
    wire[0:0] s1323, in1323_1, in1323_2;
    wire c1323;
    assign in1323_1 = {pp30[0]};
    assign in1323_2 = {c463};
    Full_Adder FA_1323(s1323, c1323, in1323_1, in1323_2, pp29[1]);
    wire[0:0] s1324, in1324_1, in1324_2;
    wire c1324;
    assign in1324_1 = {pp9[22]};
    assign in1324_2 = {pp10[21]};
    Full_Adder FA_1324(s1324, c1324, in1324_1, in1324_2, pp8[23]);
    wire[0:0] s1325, in1325_1, in1325_2;
    wire c1325;
    assign in1325_1 = {pp12[19]};
    assign in1325_2 = {pp13[18]};
    Full_Adder FA_1325(s1325, c1325, in1325_1, in1325_2, pp11[20]);
    wire[0:0] s1326, in1326_1, in1326_2;
    wire c1326;
    assign in1326_1 = {pp15[16]};
    assign in1326_2 = {pp16[15]};
    Full_Adder FA_1326(s1326, c1326, in1326_1, in1326_2, pp14[17]);
    wire[0:0] s1327, in1327_1, in1327_2;
    wire c1327;
    assign in1327_1 = {pp18[13]};
    assign in1327_2 = {pp19[12]};
    Full_Adder FA_1327(s1327, c1327, in1327_1, in1327_2, pp17[14]);
    wire[0:0] s1328, in1328_1, in1328_2;
    wire c1328;
    assign in1328_1 = {pp21[10]};
    assign in1328_2 = {pp22[9]};
    Full_Adder FA_1328(s1328, c1328, in1328_1, in1328_2, pp20[11]);
    wire[0:0] s1329, in1329_1, in1329_2;
    wire c1329;
    assign in1329_1 = {pp24[7]};
    assign in1329_2 = {pp25[6]};
    Full_Adder FA_1329(s1329, c1329, in1329_1, in1329_2, pp23[8]);
    wire[0:0] s1330, in1330_1, in1330_2;
    wire c1330;
    assign in1330_1 = {pp27[4]};
    assign in1330_2 = {pp28[3]};
    Full_Adder FA_1330(s1330, c1330, in1330_1, in1330_2, pp26[5]);
    wire[0:0] s1331, in1331_1, in1331_2;
    wire c1331;
    assign in1331_1 = {pp30[1]};
    assign in1331_2 = {pp31[0]};
    Full_Adder FA_1331(s1331, c1331, in1331_1, in1331_2, pp29[2]);
    wire[0:0] s1332, in1332_1, in1332_2;
    wire c1332;
    assign in1332_1 = {c465};
    assign in1332_2 = {s466[0]};
    Full_Adder FA_1332(s1332, c1332, in1332_1, in1332_2, c464);
    wire[0:0] s1333, in1333_1, in1333_2;
    wire c1333;
    assign in1333_1 = {pp12[20]};
    assign in1333_2 = {pp13[19]};
    Full_Adder FA_1333(s1333, c1333, in1333_1, in1333_2, pp11[21]);
    wire[0:0] s1334, in1334_1, in1334_2;
    wire c1334;
    assign in1334_1 = {pp15[17]};
    assign in1334_2 = {pp16[16]};
    Full_Adder FA_1334(s1334, c1334, in1334_1, in1334_2, pp14[18]);
    wire[0:0] s1335, in1335_1, in1335_2;
    wire c1335;
    assign in1335_1 = {pp18[14]};
    assign in1335_2 = {pp19[13]};
    Full_Adder FA_1335(s1335, c1335, in1335_1, in1335_2, pp17[15]);
    wire[0:0] s1336, in1336_1, in1336_2;
    wire c1336;
    assign in1336_1 = {pp21[11]};
    assign in1336_2 = {pp22[10]};
    Full_Adder FA_1336(s1336, c1336, in1336_1, in1336_2, pp20[12]);
    wire[0:0] s1337, in1337_1, in1337_2;
    wire c1337;
    assign in1337_1 = {pp24[8]};
    assign in1337_2 = {pp25[7]};
    Full_Adder FA_1337(s1337, c1337, in1337_1, in1337_2, pp23[9]);
    wire[0:0] s1338, in1338_1, in1338_2;
    wire c1338;
    assign in1338_1 = {pp27[5]};
    assign in1338_2 = {pp28[4]};
    Full_Adder FA_1338(s1338, c1338, in1338_1, in1338_2, pp26[6]);
    wire[0:0] s1339, in1339_1, in1339_2;
    wire c1339;
    assign in1339_1 = {pp30[2]};
    assign in1339_2 = {pp31[1]};
    Full_Adder FA_1339(s1339, c1339, in1339_1, in1339_2, pp29[3]);
    wire[0:0] s1340, in1340_1, in1340_2;
    wire c1340;
    assign in1340_1 = {c466};
    assign in1340_2 = {c467};
    Full_Adder FA_1340(s1340, c1340, in1340_1, in1340_2, pp32[0]);
    wire[0:0] s1341, in1341_1, in1341_2;
    wire c1341;
    assign in1341_1 = {s469[0]};
    assign in1341_2 = {s470[0]};
    Full_Adder FA_1341(s1341, c1341, in1341_1, in1341_2, c468);
    wire[0:0] s1342, in1342_1, in1342_2;
    wire c1342;
    assign in1342_1 = {pp15[18]};
    assign in1342_2 = {pp16[17]};
    Full_Adder FA_1342(s1342, c1342, in1342_1, in1342_2, pp14[19]);
    wire[0:0] s1343, in1343_1, in1343_2;
    wire c1343;
    assign in1343_1 = {pp18[15]};
    assign in1343_2 = {pp19[14]};
    Full_Adder FA_1343(s1343, c1343, in1343_1, in1343_2, pp17[16]);
    wire[0:0] s1344, in1344_1, in1344_2;
    wire c1344;
    assign in1344_1 = {pp21[12]};
    assign in1344_2 = {pp22[11]};
    Full_Adder FA_1344(s1344, c1344, in1344_1, in1344_2, pp20[13]);
    wire[0:0] s1345, in1345_1, in1345_2;
    wire c1345;
    assign in1345_1 = {pp24[9]};
    assign in1345_2 = {pp25[8]};
    Full_Adder FA_1345(s1345, c1345, in1345_1, in1345_2, pp23[10]);
    wire[0:0] s1346, in1346_1, in1346_2;
    wire c1346;
    assign in1346_1 = {pp27[6]};
    assign in1346_2 = {pp28[5]};
    Full_Adder FA_1346(s1346, c1346, in1346_1, in1346_2, pp26[7]);
    wire[0:0] s1347, in1347_1, in1347_2;
    wire c1347;
    assign in1347_1 = {pp30[3]};
    assign in1347_2 = {pp31[2]};
    Full_Adder FA_1347(s1347, c1347, in1347_1, in1347_2, pp29[4]);
    wire[0:0] s1348, in1348_1, in1348_2;
    wire c1348;
    assign in1348_1 = {pp33[0]};
    assign in1348_2 = {c469};
    Full_Adder FA_1348(s1348, c1348, in1348_1, in1348_2, pp32[1]);
    wire[0:0] s1349, in1349_1, in1349_2;
    wire c1349;
    assign in1349_1 = {c471};
    assign in1349_2 = {c472};
    Full_Adder FA_1349(s1349, c1349, in1349_1, in1349_2, c470);
    wire[0:0] s1350, in1350_1, in1350_2;
    wire c1350;
    assign in1350_1 = {s474[0]};
    assign in1350_2 = {s475[0]};
    Full_Adder FA_1350(s1350, c1350, in1350_1, in1350_2, s473[0]);
    wire[0:0] s1351, in1351_1, in1351_2;
    wire c1351;
    assign in1351_1 = {pp18[16]};
    assign in1351_2 = {pp19[15]};
    Full_Adder FA_1351(s1351, c1351, in1351_1, in1351_2, pp17[17]);
    wire[0:0] s1352, in1352_1, in1352_2;
    wire c1352;
    assign in1352_1 = {pp21[13]};
    assign in1352_2 = {pp22[12]};
    Full_Adder FA_1352(s1352, c1352, in1352_1, in1352_2, pp20[14]);
    wire[0:0] s1353, in1353_1, in1353_2;
    wire c1353;
    assign in1353_1 = {pp24[10]};
    assign in1353_2 = {pp25[9]};
    Full_Adder FA_1353(s1353, c1353, in1353_1, in1353_2, pp23[11]);
    wire[0:0] s1354, in1354_1, in1354_2;
    wire c1354;
    assign in1354_1 = {pp27[7]};
    assign in1354_2 = {pp28[6]};
    Full_Adder FA_1354(s1354, c1354, in1354_1, in1354_2, pp26[8]);
    wire[0:0] s1355, in1355_1, in1355_2;
    wire c1355;
    assign in1355_1 = {pp30[4]};
    assign in1355_2 = {pp31[3]};
    Full_Adder FA_1355(s1355, c1355, in1355_1, in1355_2, pp29[5]);
    wire[0:0] s1356, in1356_1, in1356_2;
    wire c1356;
    assign in1356_1 = {pp33[1]};
    assign in1356_2 = {pp34[0]};
    Full_Adder FA_1356(s1356, c1356, in1356_1, in1356_2, pp32[2]);
    wire[0:0] s1357, in1357_1, in1357_2;
    wire c1357;
    assign in1357_1 = {c474};
    assign in1357_2 = {c475};
    Full_Adder FA_1357(s1357, c1357, in1357_1, in1357_2, c473);
    wire[0:0] s1358, in1358_1, in1358_2;
    wire c1358;
    assign in1358_1 = {c477};
    assign in1358_2 = {s478[0]};
    Full_Adder FA_1358(s1358, c1358, in1358_1, in1358_2, c476);
    wire[0:0] s1359, in1359_1, in1359_2;
    wire c1359;
    assign in1359_1 = {s480[0]};
    assign in1359_2 = {s481[0]};
    Full_Adder FA_1359(s1359, c1359, in1359_1, in1359_2, s479[0]);
    wire[0:0] s1360, in1360_1, in1360_2;
    wire c1360;
    assign in1360_1 = {pp21[14]};
    assign in1360_2 = {pp22[13]};
    Full_Adder FA_1360(s1360, c1360, in1360_1, in1360_2, pp20[15]);
    wire[0:0] s1361, in1361_1, in1361_2;
    wire c1361;
    assign in1361_1 = {pp24[11]};
    assign in1361_2 = {pp25[10]};
    Full_Adder FA_1361(s1361, c1361, in1361_1, in1361_2, pp23[12]);
    wire[0:0] s1362, in1362_1, in1362_2;
    wire c1362;
    assign in1362_1 = {pp27[8]};
    assign in1362_2 = {pp28[7]};
    Full_Adder FA_1362(s1362, c1362, in1362_1, in1362_2, pp26[9]);
    wire[0:0] s1363, in1363_1, in1363_2;
    wire c1363;
    assign in1363_1 = {pp30[5]};
    assign in1363_2 = {pp31[4]};
    Full_Adder FA_1363(s1363, c1363, in1363_1, in1363_2, pp29[6]);
    wire[0:0] s1364, in1364_1, in1364_2;
    wire c1364;
    assign in1364_1 = {pp33[2]};
    assign in1364_2 = {pp34[1]};
    Full_Adder FA_1364(s1364, c1364, in1364_1, in1364_2, pp32[3]);
    wire[0:0] s1365, in1365_1, in1365_2;
    wire c1365;
    assign in1365_1 = {c478};
    assign in1365_2 = {c479};
    Full_Adder FA_1365(s1365, c1365, in1365_1, in1365_2, pp35[0]);
    wire[0:0] s1366, in1366_1, in1366_2;
    wire c1366;
    assign in1366_1 = {c481};
    assign in1366_2 = {c482};
    Full_Adder FA_1366(s1366, c1366, in1366_1, in1366_2, c480);
    wire[0:0] s1367, in1367_1, in1367_2;
    wire c1367;
    assign in1367_1 = {s484[0]};
    assign in1367_2 = {s485[0]};
    Full_Adder FA_1367(s1367, c1367, in1367_1, in1367_2, c483);
    wire[0:0] s1368, in1368_1, in1368_2;
    wire c1368;
    assign in1368_1 = {s487[0]};
    assign in1368_2 = {s488[0]};
    Full_Adder FA_1368(s1368, c1368, in1368_1, in1368_2, s486[0]);
    wire[0:0] s1369, in1369_1, in1369_2;
    wire c1369;
    assign in1369_1 = {pp24[12]};
    assign in1369_2 = {pp25[11]};
    Full_Adder FA_1369(s1369, c1369, in1369_1, in1369_2, pp23[13]);
    wire[0:0] s1370, in1370_1, in1370_2;
    wire c1370;
    assign in1370_1 = {pp27[9]};
    assign in1370_2 = {pp28[8]};
    Full_Adder FA_1370(s1370, c1370, in1370_1, in1370_2, pp26[10]);
    wire[0:0] s1371, in1371_1, in1371_2;
    wire c1371;
    assign in1371_1 = {pp30[6]};
    assign in1371_2 = {pp31[5]};
    Full_Adder FA_1371(s1371, c1371, in1371_1, in1371_2, pp29[7]);
    wire[0:0] s1372, in1372_1, in1372_2;
    wire c1372;
    assign in1372_1 = {pp33[3]};
    assign in1372_2 = {pp34[2]};
    Full_Adder FA_1372(s1372, c1372, in1372_1, in1372_2, pp32[4]);
    wire[0:0] s1373, in1373_1, in1373_2;
    wire c1373;
    assign in1373_1 = {pp36[0]};
    assign in1373_2 = {c484};
    Full_Adder FA_1373(s1373, c1373, in1373_1, in1373_2, pp35[1]);
    wire[0:0] s1374, in1374_1, in1374_2;
    wire c1374;
    assign in1374_1 = {c486};
    assign in1374_2 = {c487};
    Full_Adder FA_1374(s1374, c1374, in1374_1, in1374_2, c485);
    wire[0:0] s1375, in1375_1, in1375_2;
    wire c1375;
    assign in1375_1 = {c489};
    assign in1375_2 = {c490};
    Full_Adder FA_1375(s1375, c1375, in1375_1, in1375_2, c488);
    wire[0:0] s1376, in1376_1, in1376_2;
    wire c1376;
    assign in1376_1 = {s492[0]};
    assign in1376_2 = {s493[0]};
    Full_Adder FA_1376(s1376, c1376, in1376_1, in1376_2, s491[0]);
    wire[0:0] s1377, in1377_1, in1377_2;
    wire c1377;
    assign in1377_1 = {s495[0]};
    assign in1377_2 = {s496[0]};
    Full_Adder FA_1377(s1377, c1377, in1377_1, in1377_2, s494[0]);
    wire[0:0] s1378, in1378_1, in1378_2;
    wire c1378;
    assign in1378_1 = {pp27[10]};
    assign in1378_2 = {pp28[9]};
    Full_Adder FA_1378(s1378, c1378, in1378_1, in1378_2, pp26[11]);
    wire[0:0] s1379, in1379_1, in1379_2;
    wire c1379;
    assign in1379_1 = {pp30[7]};
    assign in1379_2 = {pp31[6]};
    Full_Adder FA_1379(s1379, c1379, in1379_1, in1379_2, pp29[8]);
    wire[0:0] s1380, in1380_1, in1380_2;
    wire c1380;
    assign in1380_1 = {pp33[4]};
    assign in1380_2 = {pp34[3]};
    Full_Adder FA_1380(s1380, c1380, in1380_1, in1380_2, pp32[5]);
    wire[0:0] s1381, in1381_1, in1381_2;
    wire c1381;
    assign in1381_1 = {pp36[1]};
    assign in1381_2 = {pp37[0]};
    Full_Adder FA_1381(s1381, c1381, in1381_1, in1381_2, pp35[2]);
    wire[0:0] s1382, in1382_1, in1382_2;
    wire c1382;
    assign in1382_1 = {c492};
    assign in1382_2 = {c493};
    Full_Adder FA_1382(s1382, c1382, in1382_1, in1382_2, c491);
    wire[0:0] s1383, in1383_1, in1383_2;
    wire c1383;
    assign in1383_1 = {c495};
    assign in1383_2 = {c496};
    Full_Adder FA_1383(s1383, c1383, in1383_1, in1383_2, c494);
    wire[0:0] s1384, in1384_1, in1384_2;
    wire c1384;
    assign in1384_1 = {c498};
    assign in1384_2 = {s499[0]};
    Full_Adder FA_1384(s1384, c1384, in1384_1, in1384_2, c497);
    wire[0:0] s1385, in1385_1, in1385_2;
    wire c1385;
    assign in1385_1 = {s501[0]};
    assign in1385_2 = {s502[0]};
    Full_Adder FA_1385(s1385, c1385, in1385_1, in1385_2, s500[0]);
    wire[0:0] s1386, in1386_1, in1386_2;
    wire c1386;
    assign in1386_1 = {s504[0]};
    assign in1386_2 = {s505[0]};
    Full_Adder FA_1386(s1386, c1386, in1386_1, in1386_2, s503[0]);
    wire[0:0] s1387, in1387_1, in1387_2;
    wire c1387;
    assign in1387_1 = {pp30[8]};
    assign in1387_2 = {pp31[7]};
    Full_Adder FA_1387(s1387, c1387, in1387_1, in1387_2, pp29[9]);
    wire[0:0] s1388, in1388_1, in1388_2;
    wire c1388;
    assign in1388_1 = {pp33[5]};
    assign in1388_2 = {pp34[4]};
    Full_Adder FA_1388(s1388, c1388, in1388_1, in1388_2, pp32[6]);
    wire[0:0] s1389, in1389_1, in1389_2;
    wire c1389;
    assign in1389_1 = {pp36[2]};
    assign in1389_2 = {pp37[1]};
    Full_Adder FA_1389(s1389, c1389, in1389_1, in1389_2, pp35[3]);
    wire[0:0] s1390, in1390_1, in1390_2;
    wire c1390;
    assign in1390_1 = {c499};
    assign in1390_2 = {c500};
    Full_Adder FA_1390(s1390, c1390, in1390_1, in1390_2, pp38[0]);
    wire[0:0] s1391, in1391_1, in1391_2;
    wire c1391;
    assign in1391_1 = {c502};
    assign in1391_2 = {c503};
    Full_Adder FA_1391(s1391, c1391, in1391_1, in1391_2, c501);
    wire[0:0] s1392, in1392_1, in1392_2;
    wire c1392;
    assign in1392_1 = {c505};
    assign in1392_2 = {c506};
    Full_Adder FA_1392(s1392, c1392, in1392_1, in1392_2, c504);
    wire[0:0] s1393, in1393_1, in1393_2;
    wire c1393;
    assign in1393_1 = {s508[0]};
    assign in1393_2 = {s509[0]};
    Full_Adder FA_1393(s1393, c1393, in1393_1, in1393_2, c507);
    wire[0:0] s1394, in1394_1, in1394_2;
    wire c1394;
    assign in1394_1 = {s511[0]};
    assign in1394_2 = {s512[0]};
    Full_Adder FA_1394(s1394, c1394, in1394_1, in1394_2, s510[0]);
    wire[0:0] s1395, in1395_1, in1395_2;
    wire c1395;
    assign in1395_1 = {s514[0]};
    assign in1395_2 = {s515[0]};
    Full_Adder FA_1395(s1395, c1395, in1395_1, in1395_2, s513[0]);
    wire[0:0] s1396, in1396_1, in1396_2;
    wire c1396;
    assign in1396_1 = {pp33[6]};
    assign in1396_2 = {pp34[5]};
    Full_Adder FA_1396(s1396, c1396, in1396_1, in1396_2, pp32[7]);
    wire[0:0] s1397, in1397_1, in1397_2;
    wire c1397;
    assign in1397_1 = {pp36[3]};
    assign in1397_2 = {pp37[2]};
    Full_Adder FA_1397(s1397, c1397, in1397_1, in1397_2, pp35[4]);
    wire[0:0] s1398, in1398_1, in1398_2;
    wire c1398;
    assign in1398_1 = {pp39[0]};
    assign in1398_2 = {c508};
    Full_Adder FA_1398(s1398, c1398, in1398_1, in1398_2, pp38[1]);
    wire[0:0] s1399, in1399_1, in1399_2;
    wire c1399;
    assign in1399_1 = {c510};
    assign in1399_2 = {c511};
    Full_Adder FA_1399(s1399, c1399, in1399_1, in1399_2, c509);
    wire[0:0] s1400, in1400_1, in1400_2;
    wire c1400;
    assign in1400_1 = {c513};
    assign in1400_2 = {c514};
    Full_Adder FA_1400(s1400, c1400, in1400_1, in1400_2, c512);
    wire[0:0] s1401, in1401_1, in1401_2;
    wire c1401;
    assign in1401_1 = {c516};
    assign in1401_2 = {c517};
    Full_Adder FA_1401(s1401, c1401, in1401_1, in1401_2, c515);
    wire[0:0] s1402, in1402_1, in1402_2;
    wire c1402;
    assign in1402_1 = {s519[0]};
    assign in1402_2 = {s520[0]};
    Full_Adder FA_1402(s1402, c1402, in1402_1, in1402_2, s518[0]);
    wire[0:0] s1403, in1403_1, in1403_2;
    wire c1403;
    assign in1403_1 = {s522[0]};
    assign in1403_2 = {s523[0]};
    Full_Adder FA_1403(s1403, c1403, in1403_1, in1403_2, s521[0]);
    wire[0:0] s1404, in1404_1, in1404_2;
    wire c1404;
    assign in1404_1 = {s525[0]};
    assign in1404_2 = {s526[0]};
    Full_Adder FA_1404(s1404, c1404, in1404_1, in1404_2, s524[0]);
    wire[0:0] s1405, in1405_1, in1405_2;
    wire c1405;
    assign in1405_1 = {pp36[4]};
    assign in1405_2 = {pp37[3]};
    Full_Adder FA_1405(s1405, c1405, in1405_1, in1405_2, pp35[5]);
    wire[0:0] s1406, in1406_1, in1406_2;
    wire c1406;
    assign in1406_1 = {pp39[1]};
    assign in1406_2 = {pp40[0]};
    Full_Adder FA_1406(s1406, c1406, in1406_1, in1406_2, pp38[2]);
    wire[0:0] s1407, in1407_1, in1407_2;
    wire c1407;
    assign in1407_1 = {c519};
    assign in1407_2 = {c520};
    Full_Adder FA_1407(s1407, c1407, in1407_1, in1407_2, c518);
    wire[0:0] s1408, in1408_1, in1408_2;
    wire c1408;
    assign in1408_1 = {c522};
    assign in1408_2 = {c523};
    Full_Adder FA_1408(s1408, c1408, in1408_1, in1408_2, c521);
    wire[0:0] s1409, in1409_1, in1409_2;
    wire c1409;
    assign in1409_1 = {c525};
    assign in1409_2 = {c526};
    Full_Adder FA_1409(s1409, c1409, in1409_1, in1409_2, c524);
    wire[0:0] s1410, in1410_1, in1410_2;
    wire c1410;
    assign in1410_1 = {c528};
    assign in1410_2 = {s529[0]};
    Full_Adder FA_1410(s1410, c1410, in1410_1, in1410_2, c527);
    wire[0:0] s1411, in1411_1, in1411_2;
    wire c1411;
    assign in1411_1 = {s531[0]};
    assign in1411_2 = {s532[0]};
    Full_Adder FA_1411(s1411, c1411, in1411_1, in1411_2, s530[0]);
    wire[0:0] s1412, in1412_1, in1412_2;
    wire c1412;
    assign in1412_1 = {s534[0]};
    assign in1412_2 = {s535[0]};
    Full_Adder FA_1412(s1412, c1412, in1412_1, in1412_2, s533[0]);
    wire[0:0] s1413, in1413_1, in1413_2;
    wire c1413;
    assign in1413_1 = {s537[0]};
    assign in1413_2 = {s538[0]};
    Full_Adder FA_1413(s1413, c1413, in1413_1, in1413_2, s536[0]);
    wire[0:0] s1414, in1414_1, in1414_2;
    wire c1414;
    assign in1414_1 = {pp39[2]};
    assign in1414_2 = {pp40[1]};
    Full_Adder FA_1414(s1414, c1414, in1414_1, in1414_2, pp38[3]);
    wire[0:0] s1415, in1415_1, in1415_2;
    wire c1415;
    assign in1415_1 = {c529};
    assign in1415_2 = {c530};
    Full_Adder FA_1415(s1415, c1415, in1415_1, in1415_2, pp41[0]);
    wire[0:0] s1416, in1416_1, in1416_2;
    wire c1416;
    assign in1416_1 = {c532};
    assign in1416_2 = {c533};
    Full_Adder FA_1416(s1416, c1416, in1416_1, in1416_2, c531);
    wire[0:0] s1417, in1417_1, in1417_2;
    wire c1417;
    assign in1417_1 = {c535};
    assign in1417_2 = {c536};
    Full_Adder FA_1417(s1417, c1417, in1417_1, in1417_2, c534);
    wire[0:0] s1418, in1418_1, in1418_2;
    wire c1418;
    assign in1418_1 = {c538};
    assign in1418_2 = {c539};
    Full_Adder FA_1418(s1418, c1418, in1418_1, in1418_2, c537);
    wire[0:0] s1419, in1419_1, in1419_2;
    wire c1419;
    assign in1419_1 = {s541[0]};
    assign in1419_2 = {s542[0]};
    Full_Adder FA_1419(s1419, c1419, in1419_1, in1419_2, c540);
    wire[0:0] s1420, in1420_1, in1420_2;
    wire c1420;
    assign in1420_1 = {s544[0]};
    assign in1420_2 = {s545[0]};
    Full_Adder FA_1420(s1420, c1420, in1420_1, in1420_2, s543[0]);
    wire[0:0] s1421, in1421_1, in1421_2;
    wire c1421;
    assign in1421_1 = {s547[0]};
    assign in1421_2 = {s548[0]};
    Full_Adder FA_1421(s1421, c1421, in1421_1, in1421_2, s546[0]);
    wire[0:0] s1422, in1422_1, in1422_2;
    wire c1422;
    assign in1422_1 = {s550[0]};
    assign in1422_2 = {s551[0]};
    Full_Adder FA_1422(s1422, c1422, in1422_1, in1422_2, s549[0]);
    wire[0:0] s1423, in1423_1, in1423_2;
    wire c1423;
    assign in1423_1 = {pp42[0]};
    assign in1423_2 = {c541};
    Full_Adder FA_1423(s1423, c1423, in1423_1, in1423_2, pp41[1]);
    wire[0:0] s1424, in1424_1, in1424_2;
    wire c1424;
    assign in1424_1 = {c543};
    assign in1424_2 = {c544};
    Full_Adder FA_1424(s1424, c1424, in1424_1, in1424_2, c542);
    wire[0:0] s1425, in1425_1, in1425_2;
    wire c1425;
    assign in1425_1 = {c546};
    assign in1425_2 = {c547};
    Full_Adder FA_1425(s1425, c1425, in1425_1, in1425_2, c545);
    wire[0:0] s1426, in1426_1, in1426_2;
    wire c1426;
    assign in1426_1 = {c549};
    assign in1426_2 = {c550};
    Full_Adder FA_1426(s1426, c1426, in1426_1, in1426_2, c548);
    wire[0:0] s1427, in1427_1, in1427_2;
    wire c1427;
    assign in1427_1 = {c552};
    assign in1427_2 = {c553};
    Full_Adder FA_1427(s1427, c1427, in1427_1, in1427_2, c551);
    wire[0:0] s1428, in1428_1, in1428_2;
    wire c1428;
    assign in1428_1 = {s555[0]};
    assign in1428_2 = {s556[0]};
    Full_Adder FA_1428(s1428, c1428, in1428_1, in1428_2, s554[0]);
    wire[0:0] s1429, in1429_1, in1429_2;
    wire c1429;
    assign in1429_1 = {s558[0]};
    assign in1429_2 = {s559[0]};
    Full_Adder FA_1429(s1429, c1429, in1429_1, in1429_2, s557[0]);
    wire[0:0] s1430, in1430_1, in1430_2;
    wire c1430;
    assign in1430_1 = {s561[0]};
    assign in1430_2 = {s562[0]};
    Full_Adder FA_1430(s1430, c1430, in1430_1, in1430_2, s560[0]);
    wire[0:0] s1431, in1431_1, in1431_2;
    wire c1431;
    assign in1431_1 = {s564[0]};
    assign in1431_2 = {s565[0]};
    Full_Adder FA_1431(s1431, c1431, in1431_1, in1431_2, s563[0]);
    wire[0:0] s1432, in1432_1, in1432_2;
    wire c1432;
    assign in1432_1 = {c554};
    assign in1432_2 = {c555};
    Full_Adder FA_1432(s1432, c1432, in1432_1, in1432_2, s1[0]);
    wire[0:0] s1433, in1433_1, in1433_2;
    wire c1433;
    assign in1433_1 = {c557};
    assign in1433_2 = {c558};
    Full_Adder FA_1433(s1433, c1433, in1433_1, in1433_2, c556);
    wire[0:0] s1434, in1434_1, in1434_2;
    wire c1434;
    assign in1434_1 = {c560};
    assign in1434_2 = {c561};
    Full_Adder FA_1434(s1434, c1434, in1434_1, in1434_2, c559);
    wire[0:0] s1435, in1435_1, in1435_2;
    wire c1435;
    assign in1435_1 = {c563};
    assign in1435_2 = {c564};
    Full_Adder FA_1435(s1435, c1435, in1435_1, in1435_2, c562);
    wire[0:0] s1436, in1436_1, in1436_2;
    wire c1436;
    assign in1436_1 = {c566};
    assign in1436_2 = {c567};
    Full_Adder FA_1436(s1436, c1436, in1436_1, in1436_2, c565);
    wire[0:0] s1437, in1437_1, in1437_2;
    wire c1437;
    assign in1437_1 = {s569[0]};
    assign in1437_2 = {s570[0]};
    Full_Adder FA_1437(s1437, c1437, in1437_1, in1437_2, s568[0]);
    wire[0:0] s1438, in1438_1, in1438_2;
    wire c1438;
    assign in1438_1 = {s572[0]};
    assign in1438_2 = {s573[0]};
    Full_Adder FA_1438(s1438, c1438, in1438_1, in1438_2, s571[0]);
    wire[0:0] s1439, in1439_1, in1439_2;
    wire c1439;
    assign in1439_1 = {s575[0]};
    assign in1439_2 = {s576[0]};
    Full_Adder FA_1439(s1439, c1439, in1439_1, in1439_2, s574[0]);
    wire[0:0] s1440, in1440_1, in1440_2;
    wire c1440;
    assign in1440_1 = {s578[0]};
    assign in1440_2 = {s579[0]};
    Full_Adder FA_1440(s1440, c1440, in1440_1, in1440_2, s577[0]);
    wire[0:0] s1441, in1441_1, in1441_2;
    wire c1441;
    assign in1441_1 = {c568};
    assign in1441_2 = {c569};
    Full_Adder FA_1441(s1441, c1441, in1441_1, in1441_2, s3[0]);
    wire[0:0] s1442, in1442_1, in1442_2;
    wire c1442;
    assign in1442_1 = {c571};
    assign in1442_2 = {c572};
    Full_Adder FA_1442(s1442, c1442, in1442_1, in1442_2, c570);
    wire[0:0] s1443, in1443_1, in1443_2;
    wire c1443;
    assign in1443_1 = {c574};
    assign in1443_2 = {c575};
    Full_Adder FA_1443(s1443, c1443, in1443_1, in1443_2, c573);
    wire[0:0] s1444, in1444_1, in1444_2;
    wire c1444;
    assign in1444_1 = {c577};
    assign in1444_2 = {c578};
    Full_Adder FA_1444(s1444, c1444, in1444_1, in1444_2, c576);
    wire[0:0] s1445, in1445_1, in1445_2;
    wire c1445;
    assign in1445_1 = {c580};
    assign in1445_2 = {c581};
    Full_Adder FA_1445(s1445, c1445, in1445_1, in1445_2, c579);
    wire[0:0] s1446, in1446_1, in1446_2;
    wire c1446;
    assign in1446_1 = {s583[0]};
    assign in1446_2 = {s584[0]};
    Full_Adder FA_1446(s1446, c1446, in1446_1, in1446_2, s582[0]);
    wire[0:0] s1447, in1447_1, in1447_2;
    wire c1447;
    assign in1447_1 = {s586[0]};
    assign in1447_2 = {s587[0]};
    Full_Adder FA_1447(s1447, c1447, in1447_1, in1447_2, s585[0]);
    wire[0:0] s1448, in1448_1, in1448_2;
    wire c1448;
    assign in1448_1 = {s589[0]};
    assign in1448_2 = {s590[0]};
    Full_Adder FA_1448(s1448, c1448, in1448_1, in1448_2, s588[0]);
    wire[0:0] s1449, in1449_1, in1449_2;
    wire c1449;
    assign in1449_1 = {s592[0]};
    assign in1449_2 = {s593[0]};
    Full_Adder FA_1449(s1449, c1449, in1449_1, in1449_2, s591[0]);
    wire[0:0] s1450, in1450_1, in1450_2;
    wire c1450;
    assign in1450_1 = {c582};
    assign in1450_2 = {c583};
    Full_Adder FA_1450(s1450, c1450, in1450_1, in1450_2, s6[0]);
    wire[0:0] s1451, in1451_1, in1451_2;
    wire c1451;
    assign in1451_1 = {c585};
    assign in1451_2 = {c586};
    Full_Adder FA_1451(s1451, c1451, in1451_1, in1451_2, c584);
    wire[0:0] s1452, in1452_1, in1452_2;
    wire c1452;
    assign in1452_1 = {c588};
    assign in1452_2 = {c589};
    Full_Adder FA_1452(s1452, c1452, in1452_1, in1452_2, c587);
    wire[0:0] s1453, in1453_1, in1453_2;
    wire c1453;
    assign in1453_1 = {c591};
    assign in1453_2 = {c592};
    Full_Adder FA_1453(s1453, c1453, in1453_1, in1453_2, c590);
    wire[0:0] s1454, in1454_1, in1454_2;
    wire c1454;
    assign in1454_1 = {c594};
    assign in1454_2 = {c595};
    Full_Adder FA_1454(s1454, c1454, in1454_1, in1454_2, c593);
    wire[0:0] s1455, in1455_1, in1455_2;
    wire c1455;
    assign in1455_1 = {s597[0]};
    assign in1455_2 = {s598[0]};
    Full_Adder FA_1455(s1455, c1455, in1455_1, in1455_2, s596[0]);
    wire[0:0] s1456, in1456_1, in1456_2;
    wire c1456;
    assign in1456_1 = {s600[0]};
    assign in1456_2 = {s601[0]};
    Full_Adder FA_1456(s1456, c1456, in1456_1, in1456_2, s599[0]);
    wire[0:0] s1457, in1457_1, in1457_2;
    wire c1457;
    assign in1457_1 = {s603[0]};
    assign in1457_2 = {s604[0]};
    Full_Adder FA_1457(s1457, c1457, in1457_1, in1457_2, s602[0]);
    wire[0:0] s1458, in1458_1, in1458_2;
    wire c1458;
    assign in1458_1 = {s606[0]};
    assign in1458_2 = {s607[0]};
    Full_Adder FA_1458(s1458, c1458, in1458_1, in1458_2, s605[0]);
    wire[0:0] s1459, in1459_1, in1459_2;
    wire c1459;
    assign in1459_1 = {c596};
    assign in1459_2 = {c597};
    Full_Adder FA_1459(s1459, c1459, in1459_1, in1459_2, s10[0]);
    wire[0:0] s1460, in1460_1, in1460_2;
    wire c1460;
    assign in1460_1 = {c599};
    assign in1460_2 = {c600};
    Full_Adder FA_1460(s1460, c1460, in1460_1, in1460_2, c598);
    wire[0:0] s1461, in1461_1, in1461_2;
    wire c1461;
    assign in1461_1 = {c602};
    assign in1461_2 = {c603};
    Full_Adder FA_1461(s1461, c1461, in1461_1, in1461_2, c601);
    wire[0:0] s1462, in1462_1, in1462_2;
    wire c1462;
    assign in1462_1 = {c605};
    assign in1462_2 = {c606};
    Full_Adder FA_1462(s1462, c1462, in1462_1, in1462_2, c604);
    wire[0:0] s1463, in1463_1, in1463_2;
    wire c1463;
    assign in1463_1 = {c608};
    assign in1463_2 = {c609};
    Full_Adder FA_1463(s1463, c1463, in1463_1, in1463_2, c607);
    wire[0:0] s1464, in1464_1, in1464_2;
    wire c1464;
    assign in1464_1 = {s611[0]};
    assign in1464_2 = {s612[0]};
    Full_Adder FA_1464(s1464, c1464, in1464_1, in1464_2, s610[0]);
    wire[0:0] s1465, in1465_1, in1465_2;
    wire c1465;
    assign in1465_1 = {s614[0]};
    assign in1465_2 = {s615[0]};
    Full_Adder FA_1465(s1465, c1465, in1465_1, in1465_2, s613[0]);
    wire[0:0] s1466, in1466_1, in1466_2;
    wire c1466;
    assign in1466_1 = {s617[0]};
    assign in1466_2 = {s618[0]};
    Full_Adder FA_1466(s1466, c1466, in1466_1, in1466_2, s616[0]);
    wire[0:0] s1467, in1467_1, in1467_2;
    wire c1467;
    assign in1467_1 = {s620[0]};
    assign in1467_2 = {s621[0]};
    Full_Adder FA_1467(s1467, c1467, in1467_1, in1467_2, s619[0]);
    wire[0:0] s1468, in1468_1, in1468_2;
    wire c1468;
    assign in1468_1 = {c610};
    assign in1468_2 = {c611};
    Full_Adder FA_1468(s1468, c1468, in1468_1, in1468_2, s15[0]);
    wire[0:0] s1469, in1469_1, in1469_2;
    wire c1469;
    assign in1469_1 = {c613};
    assign in1469_2 = {c614};
    Full_Adder FA_1469(s1469, c1469, in1469_1, in1469_2, c612);
    wire[0:0] s1470, in1470_1, in1470_2;
    wire c1470;
    assign in1470_1 = {c616};
    assign in1470_2 = {c617};
    Full_Adder FA_1470(s1470, c1470, in1470_1, in1470_2, c615);
    wire[0:0] s1471, in1471_1, in1471_2;
    wire c1471;
    assign in1471_1 = {c619};
    assign in1471_2 = {c620};
    Full_Adder FA_1471(s1471, c1471, in1471_1, in1471_2, c618);
    wire[0:0] s1472, in1472_1, in1472_2;
    wire c1472;
    assign in1472_1 = {c622};
    assign in1472_2 = {c623};
    Full_Adder FA_1472(s1472, c1472, in1472_1, in1472_2, c621);
    wire[0:0] s1473, in1473_1, in1473_2;
    wire c1473;
    assign in1473_1 = {s625[0]};
    assign in1473_2 = {s626[0]};
    Full_Adder FA_1473(s1473, c1473, in1473_1, in1473_2, s624[0]);
    wire[0:0] s1474, in1474_1, in1474_2;
    wire c1474;
    assign in1474_1 = {s628[0]};
    assign in1474_2 = {s629[0]};
    Full_Adder FA_1474(s1474, c1474, in1474_1, in1474_2, s627[0]);
    wire[0:0] s1475, in1475_1, in1475_2;
    wire c1475;
    assign in1475_1 = {s631[0]};
    assign in1475_2 = {s632[0]};
    Full_Adder FA_1475(s1475, c1475, in1475_1, in1475_2, s630[0]);
    wire[0:0] s1476, in1476_1, in1476_2;
    wire c1476;
    assign in1476_1 = {s634[0]};
    assign in1476_2 = {s635[0]};
    Full_Adder FA_1476(s1476, c1476, in1476_1, in1476_2, s633[0]);
    wire[0:0] s1477, in1477_1, in1477_2;
    wire c1477;
    assign in1477_1 = {c624};
    assign in1477_2 = {c625};
    Full_Adder FA_1477(s1477, c1477, in1477_1, in1477_2, s21[0]);
    wire[0:0] s1478, in1478_1, in1478_2;
    wire c1478;
    assign in1478_1 = {c627};
    assign in1478_2 = {c628};
    Full_Adder FA_1478(s1478, c1478, in1478_1, in1478_2, c626);
    wire[0:0] s1479, in1479_1, in1479_2;
    wire c1479;
    assign in1479_1 = {c630};
    assign in1479_2 = {c631};
    Full_Adder FA_1479(s1479, c1479, in1479_1, in1479_2, c629);
    wire[0:0] s1480, in1480_1, in1480_2;
    wire c1480;
    assign in1480_1 = {c633};
    assign in1480_2 = {c634};
    Full_Adder FA_1480(s1480, c1480, in1480_1, in1480_2, c632);
    wire[0:0] s1481, in1481_1, in1481_2;
    wire c1481;
    assign in1481_1 = {c636};
    assign in1481_2 = {c637};
    Full_Adder FA_1481(s1481, c1481, in1481_1, in1481_2, c635);
    wire[0:0] s1482, in1482_1, in1482_2;
    wire c1482;
    assign in1482_1 = {s639[0]};
    assign in1482_2 = {s640[0]};
    Full_Adder FA_1482(s1482, c1482, in1482_1, in1482_2, s638[0]);
    wire[0:0] s1483, in1483_1, in1483_2;
    wire c1483;
    assign in1483_1 = {s642[0]};
    assign in1483_2 = {s643[0]};
    Full_Adder FA_1483(s1483, c1483, in1483_1, in1483_2, s641[0]);
    wire[0:0] s1484, in1484_1, in1484_2;
    wire c1484;
    assign in1484_1 = {s645[0]};
    assign in1484_2 = {s646[0]};
    Full_Adder FA_1484(s1484, c1484, in1484_1, in1484_2, s644[0]);
    wire[0:0] s1485, in1485_1, in1485_2;
    wire c1485;
    assign in1485_1 = {s648[0]};
    assign in1485_2 = {s649[0]};
    Full_Adder FA_1485(s1485, c1485, in1485_1, in1485_2, s647[0]);
    wire[0:0] s1486, in1486_1, in1486_2;
    wire c1486;
    assign in1486_1 = {c638};
    assign in1486_2 = {c639};
    Full_Adder FA_1486(s1486, c1486, in1486_1, in1486_2, s28[0]);
    wire[0:0] s1487, in1487_1, in1487_2;
    wire c1487;
    assign in1487_1 = {c641};
    assign in1487_2 = {c642};
    Full_Adder FA_1487(s1487, c1487, in1487_1, in1487_2, c640);
    wire[0:0] s1488, in1488_1, in1488_2;
    wire c1488;
    assign in1488_1 = {c644};
    assign in1488_2 = {c645};
    Full_Adder FA_1488(s1488, c1488, in1488_1, in1488_2, c643);
    wire[0:0] s1489, in1489_1, in1489_2;
    wire c1489;
    assign in1489_1 = {c647};
    assign in1489_2 = {c648};
    Full_Adder FA_1489(s1489, c1489, in1489_1, in1489_2, c646);
    wire[0:0] s1490, in1490_1, in1490_2;
    wire c1490;
    assign in1490_1 = {c650};
    assign in1490_2 = {c651};
    Full_Adder FA_1490(s1490, c1490, in1490_1, in1490_2, c649);
    wire[0:0] s1491, in1491_1, in1491_2;
    wire c1491;
    assign in1491_1 = {s653[0]};
    assign in1491_2 = {s654[0]};
    Full_Adder FA_1491(s1491, c1491, in1491_1, in1491_2, s652[0]);
    wire[0:0] s1492, in1492_1, in1492_2;
    wire c1492;
    assign in1492_1 = {s656[0]};
    assign in1492_2 = {s657[0]};
    Full_Adder FA_1492(s1492, c1492, in1492_1, in1492_2, s655[0]);
    wire[0:0] s1493, in1493_1, in1493_2;
    wire c1493;
    assign in1493_1 = {s659[0]};
    assign in1493_2 = {s660[0]};
    Full_Adder FA_1493(s1493, c1493, in1493_1, in1493_2, s658[0]);
    wire[0:0] s1494, in1494_1, in1494_2;
    wire c1494;
    assign in1494_1 = {s662[0]};
    assign in1494_2 = {s663[0]};
    Full_Adder FA_1494(s1494, c1494, in1494_1, in1494_2, s661[0]);
    wire[0:0] s1495, in1495_1, in1495_2;
    wire c1495;
    assign in1495_1 = {c652};
    assign in1495_2 = {c653};
    Full_Adder FA_1495(s1495, c1495, in1495_1, in1495_2, s36[0]);
    wire[0:0] s1496, in1496_1, in1496_2;
    wire c1496;
    assign in1496_1 = {c655};
    assign in1496_2 = {c656};
    Full_Adder FA_1496(s1496, c1496, in1496_1, in1496_2, c654);
    wire[0:0] s1497, in1497_1, in1497_2;
    wire c1497;
    assign in1497_1 = {c658};
    assign in1497_2 = {c659};
    Full_Adder FA_1497(s1497, c1497, in1497_1, in1497_2, c657);
    wire[0:0] s1498, in1498_1, in1498_2;
    wire c1498;
    assign in1498_1 = {c661};
    assign in1498_2 = {c662};
    Full_Adder FA_1498(s1498, c1498, in1498_1, in1498_2, c660);
    wire[0:0] s1499, in1499_1, in1499_2;
    wire c1499;
    assign in1499_1 = {c664};
    assign in1499_2 = {c665};
    Full_Adder FA_1499(s1499, c1499, in1499_1, in1499_2, c663);
    wire[0:0] s1500, in1500_1, in1500_2;
    wire c1500;
    assign in1500_1 = {s667[0]};
    assign in1500_2 = {s668[0]};
    Full_Adder FA_1500(s1500, c1500, in1500_1, in1500_2, s666[0]);
    wire[0:0] s1501, in1501_1, in1501_2;
    wire c1501;
    assign in1501_1 = {s670[0]};
    assign in1501_2 = {s671[0]};
    Full_Adder FA_1501(s1501, c1501, in1501_1, in1501_2, s669[0]);
    wire[0:0] s1502, in1502_1, in1502_2;
    wire c1502;
    assign in1502_1 = {s673[0]};
    assign in1502_2 = {s674[0]};
    Full_Adder FA_1502(s1502, c1502, in1502_1, in1502_2, s672[0]);
    wire[0:0] s1503, in1503_1, in1503_2;
    wire c1503;
    assign in1503_1 = {s676[0]};
    assign in1503_2 = {s677[0]};
    Full_Adder FA_1503(s1503, c1503, in1503_1, in1503_2, s675[0]);
    wire[0:0] s1504, in1504_1, in1504_2;
    wire c1504;
    assign in1504_1 = {c666};
    assign in1504_2 = {c667};
    Full_Adder FA_1504(s1504, c1504, in1504_1, in1504_2, s45[0]);
    wire[0:0] s1505, in1505_1, in1505_2;
    wire c1505;
    assign in1505_1 = {c669};
    assign in1505_2 = {c670};
    Full_Adder FA_1505(s1505, c1505, in1505_1, in1505_2, c668);
    wire[0:0] s1506, in1506_1, in1506_2;
    wire c1506;
    assign in1506_1 = {c672};
    assign in1506_2 = {c673};
    Full_Adder FA_1506(s1506, c1506, in1506_1, in1506_2, c671);
    wire[0:0] s1507, in1507_1, in1507_2;
    wire c1507;
    assign in1507_1 = {c675};
    assign in1507_2 = {c676};
    Full_Adder FA_1507(s1507, c1507, in1507_1, in1507_2, c674);
    wire[0:0] s1508, in1508_1, in1508_2;
    wire c1508;
    assign in1508_1 = {c678};
    assign in1508_2 = {c679};
    Full_Adder FA_1508(s1508, c1508, in1508_1, in1508_2, c677);
    wire[0:0] s1509, in1509_1, in1509_2;
    wire c1509;
    assign in1509_1 = {s681[0]};
    assign in1509_2 = {s682[0]};
    Full_Adder FA_1509(s1509, c1509, in1509_1, in1509_2, s680[0]);
    wire[0:0] s1510, in1510_1, in1510_2;
    wire c1510;
    assign in1510_1 = {s684[0]};
    assign in1510_2 = {s685[0]};
    Full_Adder FA_1510(s1510, c1510, in1510_1, in1510_2, s683[0]);
    wire[0:0] s1511, in1511_1, in1511_2;
    wire c1511;
    assign in1511_1 = {s687[0]};
    assign in1511_2 = {s688[0]};
    Full_Adder FA_1511(s1511, c1511, in1511_1, in1511_2, s686[0]);
    wire[0:0] s1512, in1512_1, in1512_2;
    wire c1512;
    assign in1512_1 = {s690[0]};
    assign in1512_2 = {s691[0]};
    Full_Adder FA_1512(s1512, c1512, in1512_1, in1512_2, s689[0]);
    wire[0:0] s1513, in1513_1, in1513_2;
    wire c1513;
    assign in1513_1 = {c680};
    assign in1513_2 = {c681};
    Full_Adder FA_1513(s1513, c1513, in1513_1, in1513_2, s55[0]);
    wire[0:0] s1514, in1514_1, in1514_2;
    wire c1514;
    assign in1514_1 = {c683};
    assign in1514_2 = {c684};
    Full_Adder FA_1514(s1514, c1514, in1514_1, in1514_2, c682);
    wire[0:0] s1515, in1515_1, in1515_2;
    wire c1515;
    assign in1515_1 = {c686};
    assign in1515_2 = {c687};
    Full_Adder FA_1515(s1515, c1515, in1515_1, in1515_2, c685);
    wire[0:0] s1516, in1516_1, in1516_2;
    wire c1516;
    assign in1516_1 = {c689};
    assign in1516_2 = {c690};
    Full_Adder FA_1516(s1516, c1516, in1516_1, in1516_2, c688);
    wire[0:0] s1517, in1517_1, in1517_2;
    wire c1517;
    assign in1517_1 = {c692};
    assign in1517_2 = {c693};
    Full_Adder FA_1517(s1517, c1517, in1517_1, in1517_2, c691);
    wire[0:0] s1518, in1518_1, in1518_2;
    wire c1518;
    assign in1518_1 = {s695[0]};
    assign in1518_2 = {s696[0]};
    Full_Adder FA_1518(s1518, c1518, in1518_1, in1518_2, s694[0]);
    wire[0:0] s1519, in1519_1, in1519_2;
    wire c1519;
    assign in1519_1 = {s698[0]};
    assign in1519_2 = {s699[0]};
    Full_Adder FA_1519(s1519, c1519, in1519_1, in1519_2, s697[0]);
    wire[0:0] s1520, in1520_1, in1520_2;
    wire c1520;
    assign in1520_1 = {s701[0]};
    assign in1520_2 = {s702[0]};
    Full_Adder FA_1520(s1520, c1520, in1520_1, in1520_2, s700[0]);
    wire[0:0] s1521, in1521_1, in1521_2;
    wire c1521;
    assign in1521_1 = {s704[0]};
    assign in1521_2 = {s705[0]};
    Full_Adder FA_1521(s1521, c1521, in1521_1, in1521_2, s703[0]);
    wire[0:0] s1522, in1522_1, in1522_2;
    wire c1522;
    assign in1522_1 = {c694};
    assign in1522_2 = {c695};
    Full_Adder FA_1522(s1522, c1522, in1522_1, in1522_2, s66[0]);
    wire[0:0] s1523, in1523_1, in1523_2;
    wire c1523;
    assign in1523_1 = {c697};
    assign in1523_2 = {c698};
    Full_Adder FA_1523(s1523, c1523, in1523_1, in1523_2, c696);
    wire[0:0] s1524, in1524_1, in1524_2;
    wire c1524;
    assign in1524_1 = {c700};
    assign in1524_2 = {c701};
    Full_Adder FA_1524(s1524, c1524, in1524_1, in1524_2, c699);
    wire[0:0] s1525, in1525_1, in1525_2;
    wire c1525;
    assign in1525_1 = {c703};
    assign in1525_2 = {c704};
    Full_Adder FA_1525(s1525, c1525, in1525_1, in1525_2, c702);
    wire[0:0] s1526, in1526_1, in1526_2;
    wire c1526;
    assign in1526_1 = {c706};
    assign in1526_2 = {c707};
    Full_Adder FA_1526(s1526, c1526, in1526_1, in1526_2, c705);
    wire[0:0] s1527, in1527_1, in1527_2;
    wire c1527;
    assign in1527_1 = {s709[0]};
    assign in1527_2 = {s710[0]};
    Full_Adder FA_1527(s1527, c1527, in1527_1, in1527_2, s708[0]);
    wire[0:0] s1528, in1528_1, in1528_2;
    wire c1528;
    assign in1528_1 = {s712[0]};
    assign in1528_2 = {s713[0]};
    Full_Adder FA_1528(s1528, c1528, in1528_1, in1528_2, s711[0]);
    wire[0:0] s1529, in1529_1, in1529_2;
    wire c1529;
    assign in1529_1 = {s715[0]};
    assign in1529_2 = {s716[0]};
    Full_Adder FA_1529(s1529, c1529, in1529_1, in1529_2, s714[0]);
    wire[0:0] s1530, in1530_1, in1530_2;
    wire c1530;
    assign in1530_1 = {s718[0]};
    assign in1530_2 = {s719[0]};
    Full_Adder FA_1530(s1530, c1530, in1530_1, in1530_2, s717[0]);
    wire[0:0] s1531, in1531_1, in1531_2;
    wire c1531;
    assign in1531_1 = {c708};
    assign in1531_2 = {c709};
    Full_Adder FA_1531(s1531, c1531, in1531_1, in1531_2, s78[0]);
    wire[0:0] s1532, in1532_1, in1532_2;
    wire c1532;
    assign in1532_1 = {c711};
    assign in1532_2 = {c712};
    Full_Adder FA_1532(s1532, c1532, in1532_1, in1532_2, c710);
    wire[0:0] s1533, in1533_1, in1533_2;
    wire c1533;
    assign in1533_1 = {c714};
    assign in1533_2 = {c715};
    Full_Adder FA_1533(s1533, c1533, in1533_1, in1533_2, c713);
    wire[0:0] s1534, in1534_1, in1534_2;
    wire c1534;
    assign in1534_1 = {c717};
    assign in1534_2 = {c718};
    Full_Adder FA_1534(s1534, c1534, in1534_1, in1534_2, c716);
    wire[0:0] s1535, in1535_1, in1535_2;
    wire c1535;
    assign in1535_1 = {c720};
    assign in1535_2 = {c721};
    Full_Adder FA_1535(s1535, c1535, in1535_1, in1535_2, c719);
    wire[0:0] s1536, in1536_1, in1536_2;
    wire c1536;
    assign in1536_1 = {s723[0]};
    assign in1536_2 = {s724[0]};
    Full_Adder FA_1536(s1536, c1536, in1536_1, in1536_2, s722[0]);
    wire[0:0] s1537, in1537_1, in1537_2;
    wire c1537;
    assign in1537_1 = {s726[0]};
    assign in1537_2 = {s727[0]};
    Full_Adder FA_1537(s1537, c1537, in1537_1, in1537_2, s725[0]);
    wire[0:0] s1538, in1538_1, in1538_2;
    wire c1538;
    assign in1538_1 = {s729[0]};
    assign in1538_2 = {s730[0]};
    Full_Adder FA_1538(s1538, c1538, in1538_1, in1538_2, s728[0]);
    wire[0:0] s1539, in1539_1, in1539_2;
    wire c1539;
    assign in1539_1 = {s732[0]};
    assign in1539_2 = {s733[0]};
    Full_Adder FA_1539(s1539, c1539, in1539_1, in1539_2, s731[0]);
    wire[0:0] s1540, in1540_1, in1540_2;
    wire c1540;
    assign in1540_1 = {c722};
    assign in1540_2 = {c723};
    Full_Adder FA_1540(s1540, c1540, in1540_1, in1540_2, s91[0]);
    wire[0:0] s1541, in1541_1, in1541_2;
    wire c1541;
    assign in1541_1 = {c725};
    assign in1541_2 = {c726};
    Full_Adder FA_1541(s1541, c1541, in1541_1, in1541_2, c724);
    wire[0:0] s1542, in1542_1, in1542_2;
    wire c1542;
    assign in1542_1 = {c728};
    assign in1542_2 = {c729};
    Full_Adder FA_1542(s1542, c1542, in1542_1, in1542_2, c727);
    wire[0:0] s1543, in1543_1, in1543_2;
    wire c1543;
    assign in1543_1 = {c731};
    assign in1543_2 = {c732};
    Full_Adder FA_1543(s1543, c1543, in1543_1, in1543_2, c730);
    wire[0:0] s1544, in1544_1, in1544_2;
    wire c1544;
    assign in1544_1 = {c734};
    assign in1544_2 = {c735};
    Full_Adder FA_1544(s1544, c1544, in1544_1, in1544_2, c733);
    wire[0:0] s1545, in1545_1, in1545_2;
    wire c1545;
    assign in1545_1 = {s737[0]};
    assign in1545_2 = {s738[0]};
    Full_Adder FA_1545(s1545, c1545, in1545_1, in1545_2, s736[0]);
    wire[0:0] s1546, in1546_1, in1546_2;
    wire c1546;
    assign in1546_1 = {s740[0]};
    assign in1546_2 = {s741[0]};
    Full_Adder FA_1546(s1546, c1546, in1546_1, in1546_2, s739[0]);
    wire[0:0] s1547, in1547_1, in1547_2;
    wire c1547;
    assign in1547_1 = {s743[0]};
    assign in1547_2 = {s744[0]};
    Full_Adder FA_1547(s1547, c1547, in1547_1, in1547_2, s742[0]);
    wire[0:0] s1548, in1548_1, in1548_2;
    wire c1548;
    assign in1548_1 = {s746[0]};
    assign in1548_2 = {s747[0]};
    Full_Adder FA_1548(s1548, c1548, in1548_1, in1548_2, s745[0]);
    wire[0:0] s1549, in1549_1, in1549_2;
    wire c1549;
    assign in1549_1 = {c736};
    assign in1549_2 = {c737};
    Full_Adder FA_1549(s1549, c1549, in1549_1, in1549_2, s105[0]);
    wire[0:0] s1550, in1550_1, in1550_2;
    wire c1550;
    assign in1550_1 = {c739};
    assign in1550_2 = {c740};
    Full_Adder FA_1550(s1550, c1550, in1550_1, in1550_2, c738);
    wire[0:0] s1551, in1551_1, in1551_2;
    wire c1551;
    assign in1551_1 = {c742};
    assign in1551_2 = {c743};
    Full_Adder FA_1551(s1551, c1551, in1551_1, in1551_2, c741);
    wire[0:0] s1552, in1552_1, in1552_2;
    wire c1552;
    assign in1552_1 = {c745};
    assign in1552_2 = {c746};
    Full_Adder FA_1552(s1552, c1552, in1552_1, in1552_2, c744);
    wire[0:0] s1553, in1553_1, in1553_2;
    wire c1553;
    assign in1553_1 = {c748};
    assign in1553_2 = {c749};
    Full_Adder FA_1553(s1553, c1553, in1553_1, in1553_2, c747);
    wire[0:0] s1554, in1554_1, in1554_2;
    wire c1554;
    assign in1554_1 = {s751[0]};
    assign in1554_2 = {s752[0]};
    Full_Adder FA_1554(s1554, c1554, in1554_1, in1554_2, s750[0]);
    wire[0:0] s1555, in1555_1, in1555_2;
    wire c1555;
    assign in1555_1 = {s754[0]};
    assign in1555_2 = {s755[0]};
    Full_Adder FA_1555(s1555, c1555, in1555_1, in1555_2, s753[0]);
    wire[0:0] s1556, in1556_1, in1556_2;
    wire c1556;
    assign in1556_1 = {s757[0]};
    assign in1556_2 = {s758[0]};
    Full_Adder FA_1556(s1556, c1556, in1556_1, in1556_2, s756[0]);
    wire[0:0] s1557, in1557_1, in1557_2;
    wire c1557;
    assign in1557_1 = {s760[0]};
    assign in1557_2 = {s761[0]};
    Full_Adder FA_1557(s1557, c1557, in1557_1, in1557_2, s759[0]);
    wire[0:0] s1558, in1558_1, in1558_2;
    wire c1558;
    assign in1558_1 = {c750};
    assign in1558_2 = {c751};
    Full_Adder FA_1558(s1558, c1558, in1558_1, in1558_2, s120[0]);
    wire[0:0] s1559, in1559_1, in1559_2;
    wire c1559;
    assign in1559_1 = {c753};
    assign in1559_2 = {c754};
    Full_Adder FA_1559(s1559, c1559, in1559_1, in1559_2, c752);
    wire[0:0] s1560, in1560_1, in1560_2;
    wire c1560;
    assign in1560_1 = {c756};
    assign in1560_2 = {c757};
    Full_Adder FA_1560(s1560, c1560, in1560_1, in1560_2, c755);
    wire[0:0] s1561, in1561_1, in1561_2;
    wire c1561;
    assign in1561_1 = {c759};
    assign in1561_2 = {c760};
    Full_Adder FA_1561(s1561, c1561, in1561_1, in1561_2, c758);
    wire[0:0] s1562, in1562_1, in1562_2;
    wire c1562;
    assign in1562_1 = {c762};
    assign in1562_2 = {c763};
    Full_Adder FA_1562(s1562, c1562, in1562_1, in1562_2, c761);
    wire[0:0] s1563, in1563_1, in1563_2;
    wire c1563;
    assign in1563_1 = {s765[0]};
    assign in1563_2 = {s766[0]};
    Full_Adder FA_1563(s1563, c1563, in1563_1, in1563_2, s764[0]);
    wire[0:0] s1564, in1564_1, in1564_2;
    wire c1564;
    assign in1564_1 = {s768[0]};
    assign in1564_2 = {s769[0]};
    Full_Adder FA_1564(s1564, c1564, in1564_1, in1564_2, s767[0]);
    wire[0:0] s1565, in1565_1, in1565_2;
    wire c1565;
    assign in1565_1 = {s771[0]};
    assign in1565_2 = {s772[0]};
    Full_Adder FA_1565(s1565, c1565, in1565_1, in1565_2, s770[0]);
    wire[0:0] s1566, in1566_1, in1566_2;
    wire c1566;
    assign in1566_1 = {s774[0]};
    assign in1566_2 = {s775[0]};
    Full_Adder FA_1566(s1566, c1566, in1566_1, in1566_2, s773[0]);
    wire[0:0] s1567, in1567_1, in1567_2;
    wire c1567;
    assign in1567_1 = {c764};
    assign in1567_2 = {c765};
    Full_Adder FA_1567(s1567, c1567, in1567_1, in1567_2, s136[0]);
    wire[0:0] s1568, in1568_1, in1568_2;
    wire c1568;
    assign in1568_1 = {c767};
    assign in1568_2 = {c768};
    Full_Adder FA_1568(s1568, c1568, in1568_1, in1568_2, c766);
    wire[0:0] s1569, in1569_1, in1569_2;
    wire c1569;
    assign in1569_1 = {c770};
    assign in1569_2 = {c771};
    Full_Adder FA_1569(s1569, c1569, in1569_1, in1569_2, c769);
    wire[0:0] s1570, in1570_1, in1570_2;
    wire c1570;
    assign in1570_1 = {c773};
    assign in1570_2 = {c774};
    Full_Adder FA_1570(s1570, c1570, in1570_1, in1570_2, c772);
    wire[0:0] s1571, in1571_1, in1571_2;
    wire c1571;
    assign in1571_1 = {c776};
    assign in1571_2 = {c777};
    Full_Adder FA_1571(s1571, c1571, in1571_1, in1571_2, c775);
    wire[0:0] s1572, in1572_1, in1572_2;
    wire c1572;
    assign in1572_1 = {s779[0]};
    assign in1572_2 = {s780[0]};
    Full_Adder FA_1572(s1572, c1572, in1572_1, in1572_2, s778[0]);
    wire[0:0] s1573, in1573_1, in1573_2;
    wire c1573;
    assign in1573_1 = {s782[0]};
    assign in1573_2 = {s783[0]};
    Full_Adder FA_1573(s1573, c1573, in1573_1, in1573_2, s781[0]);
    wire[0:0] s1574, in1574_1, in1574_2;
    wire c1574;
    assign in1574_1 = {s785[0]};
    assign in1574_2 = {s786[0]};
    Full_Adder FA_1574(s1574, c1574, in1574_1, in1574_2, s784[0]);
    wire[0:0] s1575, in1575_1, in1575_2;
    wire c1575;
    assign in1575_1 = {s788[0]};
    assign in1575_2 = {s789[0]};
    Full_Adder FA_1575(s1575, c1575, in1575_1, in1575_2, s787[0]);
    wire[0:0] s1576, in1576_1, in1576_2;
    wire c1576;
    assign in1576_1 = {c778};
    assign in1576_2 = {c779};
    Full_Adder FA_1576(s1576, c1576, in1576_1, in1576_2, s153[0]);
    wire[0:0] s1577, in1577_1, in1577_2;
    wire c1577;
    assign in1577_1 = {c781};
    assign in1577_2 = {c782};
    Full_Adder FA_1577(s1577, c1577, in1577_1, in1577_2, c780);
    wire[0:0] s1578, in1578_1, in1578_2;
    wire c1578;
    assign in1578_1 = {c784};
    assign in1578_2 = {c785};
    Full_Adder FA_1578(s1578, c1578, in1578_1, in1578_2, c783);
    wire[0:0] s1579, in1579_1, in1579_2;
    wire c1579;
    assign in1579_1 = {c787};
    assign in1579_2 = {c788};
    Full_Adder FA_1579(s1579, c1579, in1579_1, in1579_2, c786);
    wire[0:0] s1580, in1580_1, in1580_2;
    wire c1580;
    assign in1580_1 = {c790};
    assign in1580_2 = {c791};
    Full_Adder FA_1580(s1580, c1580, in1580_1, in1580_2, c789);
    wire[0:0] s1581, in1581_1, in1581_2;
    wire c1581;
    assign in1581_1 = {s793[0]};
    assign in1581_2 = {s794[0]};
    Full_Adder FA_1581(s1581, c1581, in1581_1, in1581_2, s792[0]);
    wire[0:0] s1582, in1582_1, in1582_2;
    wire c1582;
    assign in1582_1 = {s796[0]};
    assign in1582_2 = {s797[0]};
    Full_Adder FA_1582(s1582, c1582, in1582_1, in1582_2, s795[0]);
    wire[0:0] s1583, in1583_1, in1583_2;
    wire c1583;
    assign in1583_1 = {s799[0]};
    assign in1583_2 = {s800[0]};
    Full_Adder FA_1583(s1583, c1583, in1583_1, in1583_2, s798[0]);
    wire[0:0] s1584, in1584_1, in1584_2;
    wire c1584;
    assign in1584_1 = {s802[0]};
    assign in1584_2 = {s803[0]};
    Full_Adder FA_1584(s1584, c1584, in1584_1, in1584_2, s801[0]);
    wire[0:0] s1585, in1585_1, in1585_2;
    wire c1585;
    assign in1585_1 = {c792};
    assign in1585_2 = {c793};
    Full_Adder FA_1585(s1585, c1585, in1585_1, in1585_2, s171[0]);
    wire[0:0] s1586, in1586_1, in1586_2;
    wire c1586;
    assign in1586_1 = {c795};
    assign in1586_2 = {c796};
    Full_Adder FA_1586(s1586, c1586, in1586_1, in1586_2, c794);
    wire[0:0] s1587, in1587_1, in1587_2;
    wire c1587;
    assign in1587_1 = {c798};
    assign in1587_2 = {c799};
    Full_Adder FA_1587(s1587, c1587, in1587_1, in1587_2, c797);
    wire[0:0] s1588, in1588_1, in1588_2;
    wire c1588;
    assign in1588_1 = {c801};
    assign in1588_2 = {c802};
    Full_Adder FA_1588(s1588, c1588, in1588_1, in1588_2, c800);
    wire[0:0] s1589, in1589_1, in1589_2;
    wire c1589;
    assign in1589_1 = {c804};
    assign in1589_2 = {c805};
    Full_Adder FA_1589(s1589, c1589, in1589_1, in1589_2, c803);
    wire[0:0] s1590, in1590_1, in1590_2;
    wire c1590;
    assign in1590_1 = {s807[0]};
    assign in1590_2 = {s808[0]};
    Full_Adder FA_1590(s1590, c1590, in1590_1, in1590_2, s806[0]);
    wire[0:0] s1591, in1591_1, in1591_2;
    wire c1591;
    assign in1591_1 = {s810[0]};
    assign in1591_2 = {s811[0]};
    Full_Adder FA_1591(s1591, c1591, in1591_1, in1591_2, s809[0]);
    wire[0:0] s1592, in1592_1, in1592_2;
    wire c1592;
    assign in1592_1 = {s813[0]};
    assign in1592_2 = {s814[0]};
    Full_Adder FA_1592(s1592, c1592, in1592_1, in1592_2, s812[0]);
    wire[0:0] s1593, in1593_1, in1593_2;
    wire c1593;
    assign in1593_1 = {s816[0]};
    assign in1593_2 = {s817[0]};
    Full_Adder FA_1593(s1593, c1593, in1593_1, in1593_2, s815[0]);
    wire[0:0] s1594, in1594_1, in1594_2;
    wire c1594;
    assign in1594_1 = {c806};
    assign in1594_2 = {c807};
    Full_Adder FA_1594(s1594, c1594, in1594_1, in1594_2, s190[0]);
    wire[0:0] s1595, in1595_1, in1595_2;
    wire c1595;
    assign in1595_1 = {c809};
    assign in1595_2 = {c810};
    Full_Adder FA_1595(s1595, c1595, in1595_1, in1595_2, c808);
    wire[0:0] s1596, in1596_1, in1596_2;
    wire c1596;
    assign in1596_1 = {c812};
    assign in1596_2 = {c813};
    Full_Adder FA_1596(s1596, c1596, in1596_1, in1596_2, c811);
    wire[0:0] s1597, in1597_1, in1597_2;
    wire c1597;
    assign in1597_1 = {c815};
    assign in1597_2 = {c816};
    Full_Adder FA_1597(s1597, c1597, in1597_1, in1597_2, c814);
    wire[0:0] s1598, in1598_1, in1598_2;
    wire c1598;
    assign in1598_1 = {c818};
    assign in1598_2 = {c819};
    Full_Adder FA_1598(s1598, c1598, in1598_1, in1598_2, c817);
    wire[0:0] s1599, in1599_1, in1599_2;
    wire c1599;
    assign in1599_1 = {s821[0]};
    assign in1599_2 = {s822[0]};
    Full_Adder FA_1599(s1599, c1599, in1599_1, in1599_2, s820[0]);
    wire[0:0] s1600, in1600_1, in1600_2;
    wire c1600;
    assign in1600_1 = {s824[0]};
    assign in1600_2 = {s825[0]};
    Full_Adder FA_1600(s1600, c1600, in1600_1, in1600_2, s823[0]);
    wire[0:0] s1601, in1601_1, in1601_2;
    wire c1601;
    assign in1601_1 = {s827[0]};
    assign in1601_2 = {s828[0]};
    Full_Adder FA_1601(s1601, c1601, in1601_1, in1601_2, s826[0]);
    wire[0:0] s1602, in1602_1, in1602_2;
    wire c1602;
    assign in1602_1 = {s830[0]};
    assign in1602_2 = {s831[0]};
    Full_Adder FA_1602(s1602, c1602, in1602_1, in1602_2, s829[0]);
    wire[0:0] s1603, in1603_1, in1603_2;
    wire c1603;
    assign in1603_1 = {c820};
    assign in1603_2 = {c821};
    Full_Adder FA_1603(s1603, c1603, in1603_1, in1603_2, s210[0]);
    wire[0:0] s1604, in1604_1, in1604_2;
    wire c1604;
    assign in1604_1 = {c823};
    assign in1604_2 = {c824};
    Full_Adder FA_1604(s1604, c1604, in1604_1, in1604_2, c822);
    wire[0:0] s1605, in1605_1, in1605_2;
    wire c1605;
    assign in1605_1 = {c826};
    assign in1605_2 = {c827};
    Full_Adder FA_1605(s1605, c1605, in1605_1, in1605_2, c825);
    wire[0:0] s1606, in1606_1, in1606_2;
    wire c1606;
    assign in1606_1 = {c829};
    assign in1606_2 = {c830};
    Full_Adder FA_1606(s1606, c1606, in1606_1, in1606_2, c828);
    wire[0:0] s1607, in1607_1, in1607_2;
    wire c1607;
    assign in1607_1 = {c832};
    assign in1607_2 = {c833};
    Full_Adder FA_1607(s1607, c1607, in1607_1, in1607_2, c831);
    wire[0:0] s1608, in1608_1, in1608_2;
    wire c1608;
    assign in1608_1 = {s835[0]};
    assign in1608_2 = {s836[0]};
    Full_Adder FA_1608(s1608, c1608, in1608_1, in1608_2, s834[0]);
    wire[0:0] s1609, in1609_1, in1609_2;
    wire c1609;
    assign in1609_1 = {s838[0]};
    assign in1609_2 = {s839[0]};
    Full_Adder FA_1609(s1609, c1609, in1609_1, in1609_2, s837[0]);
    wire[0:0] s1610, in1610_1, in1610_2;
    wire c1610;
    assign in1610_1 = {s841[0]};
    assign in1610_2 = {s842[0]};
    Full_Adder FA_1610(s1610, c1610, in1610_1, in1610_2, s840[0]);
    wire[0:0] s1611, in1611_1, in1611_2;
    wire c1611;
    assign in1611_1 = {s844[0]};
    assign in1611_2 = {s845[0]};
    Full_Adder FA_1611(s1611, c1611, in1611_1, in1611_2, s843[0]);
    wire[0:0] s1612, in1612_1, in1612_2;
    wire c1612;
    assign in1612_1 = {c834};
    assign in1612_2 = {c835};
    Full_Adder FA_1612(s1612, c1612, in1612_1, in1612_2, s231[0]);
    wire[0:0] s1613, in1613_1, in1613_2;
    wire c1613;
    assign in1613_1 = {c837};
    assign in1613_2 = {c838};
    Full_Adder FA_1613(s1613, c1613, in1613_1, in1613_2, c836);
    wire[0:0] s1614, in1614_1, in1614_2;
    wire c1614;
    assign in1614_1 = {c840};
    assign in1614_2 = {c841};
    Full_Adder FA_1614(s1614, c1614, in1614_1, in1614_2, c839);
    wire[0:0] s1615, in1615_1, in1615_2;
    wire c1615;
    assign in1615_1 = {c843};
    assign in1615_2 = {c844};
    Full_Adder FA_1615(s1615, c1615, in1615_1, in1615_2, c842);
    wire[0:0] s1616, in1616_1, in1616_2;
    wire c1616;
    assign in1616_1 = {c846};
    assign in1616_2 = {c847};
    Full_Adder FA_1616(s1616, c1616, in1616_1, in1616_2, c845);
    wire[0:0] s1617, in1617_1, in1617_2;
    wire c1617;
    assign in1617_1 = {s849[0]};
    assign in1617_2 = {s850[0]};
    Full_Adder FA_1617(s1617, c1617, in1617_1, in1617_2, s848[0]);
    wire[0:0] s1618, in1618_1, in1618_2;
    wire c1618;
    assign in1618_1 = {s852[0]};
    assign in1618_2 = {s853[0]};
    Full_Adder FA_1618(s1618, c1618, in1618_1, in1618_2, s851[0]);
    wire[0:0] s1619, in1619_1, in1619_2;
    wire c1619;
    assign in1619_1 = {s855[0]};
    assign in1619_2 = {s856[0]};
    Full_Adder FA_1619(s1619, c1619, in1619_1, in1619_2, s854[0]);
    wire[0:0] s1620, in1620_1, in1620_2;
    wire c1620;
    assign in1620_1 = {s858[0]};
    assign in1620_2 = {s859[0]};
    Full_Adder FA_1620(s1620, c1620, in1620_1, in1620_2, s857[0]);
    wire[0:0] s1621, in1621_1, in1621_2;
    wire c1621;
    assign in1621_1 = {c848};
    assign in1621_2 = {c849};
    Full_Adder FA_1621(s1621, c1621, in1621_1, in1621_2, s252[0]);
    wire[0:0] s1622, in1622_1, in1622_2;
    wire c1622;
    assign in1622_1 = {c851};
    assign in1622_2 = {c852};
    Full_Adder FA_1622(s1622, c1622, in1622_1, in1622_2, c850);
    wire[0:0] s1623, in1623_1, in1623_2;
    wire c1623;
    assign in1623_1 = {c854};
    assign in1623_2 = {c855};
    Full_Adder FA_1623(s1623, c1623, in1623_1, in1623_2, c853);
    wire[0:0] s1624, in1624_1, in1624_2;
    wire c1624;
    assign in1624_1 = {c857};
    assign in1624_2 = {c858};
    Full_Adder FA_1624(s1624, c1624, in1624_1, in1624_2, c856);
    wire[0:0] s1625, in1625_1, in1625_2;
    wire c1625;
    assign in1625_1 = {c860};
    assign in1625_2 = {c861};
    Full_Adder FA_1625(s1625, c1625, in1625_1, in1625_2, c859);
    wire[0:0] s1626, in1626_1, in1626_2;
    wire c1626;
    assign in1626_1 = {s863[0]};
    assign in1626_2 = {s864[0]};
    Full_Adder FA_1626(s1626, c1626, in1626_1, in1626_2, s862[0]);
    wire[0:0] s1627, in1627_1, in1627_2;
    wire c1627;
    assign in1627_1 = {s866[0]};
    assign in1627_2 = {s867[0]};
    Full_Adder FA_1627(s1627, c1627, in1627_1, in1627_2, s865[0]);
    wire[0:0] s1628, in1628_1, in1628_2;
    wire c1628;
    assign in1628_1 = {s869[0]};
    assign in1628_2 = {s870[0]};
    Full_Adder FA_1628(s1628, c1628, in1628_1, in1628_2, s868[0]);
    wire[0:0] s1629, in1629_1, in1629_2;
    wire c1629;
    assign in1629_1 = {s872[0]};
    assign in1629_2 = {s873[0]};
    Full_Adder FA_1629(s1629, c1629, in1629_1, in1629_2, s871[0]);
    wire[0:0] s1630, in1630_1, in1630_2;
    wire c1630;
    assign in1630_1 = {c862};
    assign in1630_2 = {c863};
    Full_Adder FA_1630(s1630, c1630, in1630_1, in1630_2, s272[0]);
    wire[0:0] s1631, in1631_1, in1631_2;
    wire c1631;
    assign in1631_1 = {c865};
    assign in1631_2 = {c866};
    Full_Adder FA_1631(s1631, c1631, in1631_1, in1631_2, c864);
    wire[0:0] s1632, in1632_1, in1632_2;
    wire c1632;
    assign in1632_1 = {c868};
    assign in1632_2 = {c869};
    Full_Adder FA_1632(s1632, c1632, in1632_1, in1632_2, c867);
    wire[0:0] s1633, in1633_1, in1633_2;
    wire c1633;
    assign in1633_1 = {c871};
    assign in1633_2 = {c872};
    Full_Adder FA_1633(s1633, c1633, in1633_1, in1633_2, c870);
    wire[0:0] s1634, in1634_1, in1634_2;
    wire c1634;
    assign in1634_1 = {c874};
    assign in1634_2 = {c875};
    Full_Adder FA_1634(s1634, c1634, in1634_1, in1634_2, c873);
    wire[0:0] s1635, in1635_1, in1635_2;
    wire c1635;
    assign in1635_1 = {s877[0]};
    assign in1635_2 = {s878[0]};
    Full_Adder FA_1635(s1635, c1635, in1635_1, in1635_2, s876[0]);
    wire[0:0] s1636, in1636_1, in1636_2;
    wire c1636;
    assign in1636_1 = {s880[0]};
    assign in1636_2 = {s881[0]};
    Full_Adder FA_1636(s1636, c1636, in1636_1, in1636_2, s879[0]);
    wire[0:0] s1637, in1637_1, in1637_2;
    wire c1637;
    assign in1637_1 = {s883[0]};
    assign in1637_2 = {s884[0]};
    Full_Adder FA_1637(s1637, c1637, in1637_1, in1637_2, s882[0]);
    wire[0:0] s1638, in1638_1, in1638_2;
    wire c1638;
    assign in1638_1 = {s886[0]};
    assign in1638_2 = {s887[0]};
    Full_Adder FA_1638(s1638, c1638, in1638_1, in1638_2, s885[0]);
    wire[0:0] s1639, in1639_1, in1639_2;
    wire c1639;
    assign in1639_1 = {c876};
    assign in1639_2 = {c877};
    Full_Adder FA_1639(s1639, c1639, in1639_1, in1639_2, s291[0]);
    wire[0:0] s1640, in1640_1, in1640_2;
    wire c1640;
    assign in1640_1 = {c879};
    assign in1640_2 = {c880};
    Full_Adder FA_1640(s1640, c1640, in1640_1, in1640_2, c878);
    wire[0:0] s1641, in1641_1, in1641_2;
    wire c1641;
    assign in1641_1 = {c882};
    assign in1641_2 = {c883};
    Full_Adder FA_1641(s1641, c1641, in1641_1, in1641_2, c881);
    wire[0:0] s1642, in1642_1, in1642_2;
    wire c1642;
    assign in1642_1 = {c885};
    assign in1642_2 = {c886};
    Full_Adder FA_1642(s1642, c1642, in1642_1, in1642_2, c884);
    wire[0:0] s1643, in1643_1, in1643_2;
    wire c1643;
    assign in1643_1 = {c888};
    assign in1643_2 = {c889};
    Full_Adder FA_1643(s1643, c1643, in1643_1, in1643_2, c887);
    wire[0:0] s1644, in1644_1, in1644_2;
    wire c1644;
    assign in1644_1 = {s891[0]};
    assign in1644_2 = {s892[0]};
    Full_Adder FA_1644(s1644, c1644, in1644_1, in1644_2, s890[0]);
    wire[0:0] s1645, in1645_1, in1645_2;
    wire c1645;
    assign in1645_1 = {s894[0]};
    assign in1645_2 = {s895[0]};
    Full_Adder FA_1645(s1645, c1645, in1645_1, in1645_2, s893[0]);
    wire[0:0] s1646, in1646_1, in1646_2;
    wire c1646;
    assign in1646_1 = {s897[0]};
    assign in1646_2 = {s898[0]};
    Full_Adder FA_1646(s1646, c1646, in1646_1, in1646_2, s896[0]);
    wire[0:0] s1647, in1647_1, in1647_2;
    wire c1647;
    assign in1647_1 = {s900[0]};
    assign in1647_2 = {s901[0]};
    Full_Adder FA_1647(s1647, c1647, in1647_1, in1647_2, s899[0]);
    wire[0:0] s1648, in1648_1, in1648_2;
    wire c1648;
    assign in1648_1 = {c890};
    assign in1648_2 = {c891};
    Full_Adder FA_1648(s1648, c1648, in1648_1, in1648_2, s309[0]);
    wire[0:0] s1649, in1649_1, in1649_2;
    wire c1649;
    assign in1649_1 = {c893};
    assign in1649_2 = {c894};
    Full_Adder FA_1649(s1649, c1649, in1649_1, in1649_2, c892);
    wire[0:0] s1650, in1650_1, in1650_2;
    wire c1650;
    assign in1650_1 = {c896};
    assign in1650_2 = {c897};
    Full_Adder FA_1650(s1650, c1650, in1650_1, in1650_2, c895);
    wire[0:0] s1651, in1651_1, in1651_2;
    wire c1651;
    assign in1651_1 = {c899};
    assign in1651_2 = {c900};
    Full_Adder FA_1651(s1651, c1651, in1651_1, in1651_2, c898);
    wire[0:0] s1652, in1652_1, in1652_2;
    wire c1652;
    assign in1652_1 = {c902};
    assign in1652_2 = {c903};
    Full_Adder FA_1652(s1652, c1652, in1652_1, in1652_2, c901);
    wire[0:0] s1653, in1653_1, in1653_2;
    wire c1653;
    assign in1653_1 = {s905[0]};
    assign in1653_2 = {s906[0]};
    Full_Adder FA_1653(s1653, c1653, in1653_1, in1653_2, s904[0]);
    wire[0:0] s1654, in1654_1, in1654_2;
    wire c1654;
    assign in1654_1 = {s908[0]};
    assign in1654_2 = {s909[0]};
    Full_Adder FA_1654(s1654, c1654, in1654_1, in1654_2, s907[0]);
    wire[0:0] s1655, in1655_1, in1655_2;
    wire c1655;
    assign in1655_1 = {s911[0]};
    assign in1655_2 = {s912[0]};
    Full_Adder FA_1655(s1655, c1655, in1655_1, in1655_2, s910[0]);
    wire[0:0] s1656, in1656_1, in1656_2;
    wire c1656;
    assign in1656_1 = {s914[0]};
    assign in1656_2 = {s915[0]};
    Full_Adder FA_1656(s1656, c1656, in1656_1, in1656_2, s913[0]);
    wire[0:0] s1657, in1657_1, in1657_2;
    wire c1657;
    assign in1657_1 = {c904};
    assign in1657_2 = {c905};
    Full_Adder FA_1657(s1657, c1657, in1657_1, in1657_2, s326[0]);
    wire[0:0] s1658, in1658_1, in1658_2;
    wire c1658;
    assign in1658_1 = {c907};
    assign in1658_2 = {c908};
    Full_Adder FA_1658(s1658, c1658, in1658_1, in1658_2, c906);
    wire[0:0] s1659, in1659_1, in1659_2;
    wire c1659;
    assign in1659_1 = {c910};
    assign in1659_2 = {c911};
    Full_Adder FA_1659(s1659, c1659, in1659_1, in1659_2, c909);
    wire[0:0] s1660, in1660_1, in1660_2;
    wire c1660;
    assign in1660_1 = {c913};
    assign in1660_2 = {c914};
    Full_Adder FA_1660(s1660, c1660, in1660_1, in1660_2, c912);
    wire[0:0] s1661, in1661_1, in1661_2;
    wire c1661;
    assign in1661_1 = {c916};
    assign in1661_2 = {c917};
    Full_Adder FA_1661(s1661, c1661, in1661_1, in1661_2, c915);
    wire[0:0] s1662, in1662_1, in1662_2;
    wire c1662;
    assign in1662_1 = {s919[0]};
    assign in1662_2 = {s920[0]};
    Full_Adder FA_1662(s1662, c1662, in1662_1, in1662_2, s918[0]);
    wire[0:0] s1663, in1663_1, in1663_2;
    wire c1663;
    assign in1663_1 = {s922[0]};
    assign in1663_2 = {s923[0]};
    Full_Adder FA_1663(s1663, c1663, in1663_1, in1663_2, s921[0]);
    wire[0:0] s1664, in1664_1, in1664_2;
    wire c1664;
    assign in1664_1 = {s925[0]};
    assign in1664_2 = {s926[0]};
    Full_Adder FA_1664(s1664, c1664, in1664_1, in1664_2, s924[0]);
    wire[0:0] s1665, in1665_1, in1665_2;
    wire c1665;
    assign in1665_1 = {s928[0]};
    assign in1665_2 = {s929[0]};
    Full_Adder FA_1665(s1665, c1665, in1665_1, in1665_2, s927[0]);
    wire[0:0] s1666, in1666_1, in1666_2;
    wire c1666;
    assign in1666_1 = {c918};
    assign in1666_2 = {c919};
    Full_Adder FA_1666(s1666, c1666, in1666_1, in1666_2, s342[0]);
    wire[0:0] s1667, in1667_1, in1667_2;
    wire c1667;
    assign in1667_1 = {c921};
    assign in1667_2 = {c922};
    Full_Adder FA_1667(s1667, c1667, in1667_1, in1667_2, c920);
    wire[0:0] s1668, in1668_1, in1668_2;
    wire c1668;
    assign in1668_1 = {c924};
    assign in1668_2 = {c925};
    Full_Adder FA_1668(s1668, c1668, in1668_1, in1668_2, c923);
    wire[0:0] s1669, in1669_1, in1669_2;
    wire c1669;
    assign in1669_1 = {c927};
    assign in1669_2 = {c928};
    Full_Adder FA_1669(s1669, c1669, in1669_1, in1669_2, c926);
    wire[0:0] s1670, in1670_1, in1670_2;
    wire c1670;
    assign in1670_1 = {c930};
    assign in1670_2 = {c931};
    Full_Adder FA_1670(s1670, c1670, in1670_1, in1670_2, c929);
    wire[0:0] s1671, in1671_1, in1671_2;
    wire c1671;
    assign in1671_1 = {s933[0]};
    assign in1671_2 = {s934[0]};
    Full_Adder FA_1671(s1671, c1671, in1671_1, in1671_2, s932[0]);
    wire[0:0] s1672, in1672_1, in1672_2;
    wire c1672;
    assign in1672_1 = {s936[0]};
    assign in1672_2 = {s937[0]};
    Full_Adder FA_1672(s1672, c1672, in1672_1, in1672_2, s935[0]);
    wire[0:0] s1673, in1673_1, in1673_2;
    wire c1673;
    assign in1673_1 = {s939[0]};
    assign in1673_2 = {s940[0]};
    Full_Adder FA_1673(s1673, c1673, in1673_1, in1673_2, s938[0]);
    wire[0:0] s1674, in1674_1, in1674_2;
    wire c1674;
    assign in1674_1 = {s942[0]};
    assign in1674_2 = {s943[0]};
    Full_Adder FA_1674(s1674, c1674, in1674_1, in1674_2, s941[0]);
    wire[0:0] s1675, in1675_1, in1675_2;
    wire c1675;
    assign in1675_1 = {c932};
    assign in1675_2 = {c933};
    Full_Adder FA_1675(s1675, c1675, in1675_1, in1675_2, s357[0]);
    wire[0:0] s1676, in1676_1, in1676_2;
    wire c1676;
    assign in1676_1 = {c935};
    assign in1676_2 = {c936};
    Full_Adder FA_1676(s1676, c1676, in1676_1, in1676_2, c934);
    wire[0:0] s1677, in1677_1, in1677_2;
    wire c1677;
    assign in1677_1 = {c938};
    assign in1677_2 = {c939};
    Full_Adder FA_1677(s1677, c1677, in1677_1, in1677_2, c937);
    wire[0:0] s1678, in1678_1, in1678_2;
    wire c1678;
    assign in1678_1 = {c941};
    assign in1678_2 = {c942};
    Full_Adder FA_1678(s1678, c1678, in1678_1, in1678_2, c940);
    wire[0:0] s1679, in1679_1, in1679_2;
    wire c1679;
    assign in1679_1 = {c944};
    assign in1679_2 = {c945};
    Full_Adder FA_1679(s1679, c1679, in1679_1, in1679_2, c943);
    wire[0:0] s1680, in1680_1, in1680_2;
    wire c1680;
    assign in1680_1 = {s947[0]};
    assign in1680_2 = {s948[0]};
    Full_Adder FA_1680(s1680, c1680, in1680_1, in1680_2, s946[0]);
    wire[0:0] s1681, in1681_1, in1681_2;
    wire c1681;
    assign in1681_1 = {s950[0]};
    assign in1681_2 = {s951[0]};
    Full_Adder FA_1681(s1681, c1681, in1681_1, in1681_2, s949[0]);
    wire[0:0] s1682, in1682_1, in1682_2;
    wire c1682;
    assign in1682_1 = {s953[0]};
    assign in1682_2 = {s954[0]};
    Full_Adder FA_1682(s1682, c1682, in1682_1, in1682_2, s952[0]);
    wire[0:0] s1683, in1683_1, in1683_2;
    wire c1683;
    assign in1683_1 = {s956[0]};
    assign in1683_2 = {s957[0]};
    Full_Adder FA_1683(s1683, c1683, in1683_1, in1683_2, s955[0]);
    wire[0:0] s1684, in1684_1, in1684_2;
    wire c1684;
    assign in1684_1 = {c946};
    assign in1684_2 = {c947};
    Full_Adder FA_1684(s1684, c1684, in1684_1, in1684_2, s371[0]);
    wire[0:0] s1685, in1685_1, in1685_2;
    wire c1685;
    assign in1685_1 = {c949};
    assign in1685_2 = {c950};
    Full_Adder FA_1685(s1685, c1685, in1685_1, in1685_2, c948);
    wire[0:0] s1686, in1686_1, in1686_2;
    wire c1686;
    assign in1686_1 = {c952};
    assign in1686_2 = {c953};
    Full_Adder FA_1686(s1686, c1686, in1686_1, in1686_2, c951);
    wire[0:0] s1687, in1687_1, in1687_2;
    wire c1687;
    assign in1687_1 = {c955};
    assign in1687_2 = {c956};
    Full_Adder FA_1687(s1687, c1687, in1687_1, in1687_2, c954);
    wire[0:0] s1688, in1688_1, in1688_2;
    wire c1688;
    assign in1688_1 = {c958};
    assign in1688_2 = {c959};
    Full_Adder FA_1688(s1688, c1688, in1688_1, in1688_2, c957);
    wire[0:0] s1689, in1689_1, in1689_2;
    wire c1689;
    assign in1689_1 = {s961[0]};
    assign in1689_2 = {s962[0]};
    Full_Adder FA_1689(s1689, c1689, in1689_1, in1689_2, s960[0]);
    wire[0:0] s1690, in1690_1, in1690_2;
    wire c1690;
    assign in1690_1 = {s964[0]};
    assign in1690_2 = {s965[0]};
    Full_Adder FA_1690(s1690, c1690, in1690_1, in1690_2, s963[0]);
    wire[0:0] s1691, in1691_1, in1691_2;
    wire c1691;
    assign in1691_1 = {s967[0]};
    assign in1691_2 = {s968[0]};
    Full_Adder FA_1691(s1691, c1691, in1691_1, in1691_2, s966[0]);
    wire[0:0] s1692, in1692_1, in1692_2;
    wire c1692;
    assign in1692_1 = {s970[0]};
    assign in1692_2 = {s971[0]};
    Full_Adder FA_1692(s1692, c1692, in1692_1, in1692_2, s969[0]);
    wire[0:0] s1693, in1693_1, in1693_2;
    wire c1693;
    assign in1693_1 = {c960};
    assign in1693_2 = {c961};
    Full_Adder FA_1693(s1693, c1693, in1693_1, in1693_2, s384[0]);
    wire[0:0] s1694, in1694_1, in1694_2;
    wire c1694;
    assign in1694_1 = {c963};
    assign in1694_2 = {c964};
    Full_Adder FA_1694(s1694, c1694, in1694_1, in1694_2, c962);
    wire[0:0] s1695, in1695_1, in1695_2;
    wire c1695;
    assign in1695_1 = {c966};
    assign in1695_2 = {c967};
    Full_Adder FA_1695(s1695, c1695, in1695_1, in1695_2, c965);
    wire[0:0] s1696, in1696_1, in1696_2;
    wire c1696;
    assign in1696_1 = {c969};
    assign in1696_2 = {c970};
    Full_Adder FA_1696(s1696, c1696, in1696_1, in1696_2, c968);
    wire[0:0] s1697, in1697_1, in1697_2;
    wire c1697;
    assign in1697_1 = {c972};
    assign in1697_2 = {c973};
    Full_Adder FA_1697(s1697, c1697, in1697_1, in1697_2, c971);
    wire[0:0] s1698, in1698_1, in1698_2;
    wire c1698;
    assign in1698_1 = {s975[0]};
    assign in1698_2 = {s976[0]};
    Full_Adder FA_1698(s1698, c1698, in1698_1, in1698_2, s974[0]);
    wire[0:0] s1699, in1699_1, in1699_2;
    wire c1699;
    assign in1699_1 = {s978[0]};
    assign in1699_2 = {s979[0]};
    Full_Adder FA_1699(s1699, c1699, in1699_1, in1699_2, s977[0]);
    wire[0:0] s1700, in1700_1, in1700_2;
    wire c1700;
    assign in1700_1 = {s981[0]};
    assign in1700_2 = {s982[0]};
    Full_Adder FA_1700(s1700, c1700, in1700_1, in1700_2, s980[0]);
    wire[0:0] s1701, in1701_1, in1701_2;
    wire c1701;
    assign in1701_1 = {s984[0]};
    assign in1701_2 = {s985[0]};
    Full_Adder FA_1701(s1701, c1701, in1701_1, in1701_2, s983[0]);
    wire[0:0] s1702, in1702_1, in1702_2;
    wire c1702;
    assign in1702_1 = {c974};
    assign in1702_2 = {c975};
    Full_Adder FA_1702(s1702, c1702, in1702_1, in1702_2, s396[0]);
    wire[0:0] s1703, in1703_1, in1703_2;
    wire c1703;
    assign in1703_1 = {c977};
    assign in1703_2 = {c978};
    Full_Adder FA_1703(s1703, c1703, in1703_1, in1703_2, c976);
    wire[0:0] s1704, in1704_1, in1704_2;
    wire c1704;
    assign in1704_1 = {c980};
    assign in1704_2 = {c981};
    Full_Adder FA_1704(s1704, c1704, in1704_1, in1704_2, c979);
    wire[0:0] s1705, in1705_1, in1705_2;
    wire c1705;
    assign in1705_1 = {c983};
    assign in1705_2 = {c984};
    Full_Adder FA_1705(s1705, c1705, in1705_1, in1705_2, c982);
    wire[0:0] s1706, in1706_1, in1706_2;
    wire c1706;
    assign in1706_1 = {c986};
    assign in1706_2 = {c987};
    Full_Adder FA_1706(s1706, c1706, in1706_1, in1706_2, c985);
    wire[0:0] s1707, in1707_1, in1707_2;
    wire c1707;
    assign in1707_1 = {s989[0]};
    assign in1707_2 = {s990[0]};
    Full_Adder FA_1707(s1707, c1707, in1707_1, in1707_2, s988[0]);
    wire[0:0] s1708, in1708_1, in1708_2;
    wire c1708;
    assign in1708_1 = {s992[0]};
    assign in1708_2 = {s993[0]};
    Full_Adder FA_1708(s1708, c1708, in1708_1, in1708_2, s991[0]);
    wire[0:0] s1709, in1709_1, in1709_2;
    wire c1709;
    assign in1709_1 = {s995[0]};
    assign in1709_2 = {s996[0]};
    Full_Adder FA_1709(s1709, c1709, in1709_1, in1709_2, s994[0]);
    wire[0:0] s1710, in1710_1, in1710_2;
    wire c1710;
    assign in1710_1 = {s998[0]};
    assign in1710_2 = {s999[0]};
    Full_Adder FA_1710(s1710, c1710, in1710_1, in1710_2, s997[0]);
    wire[0:0] s1711, in1711_1, in1711_2;
    wire c1711;
    assign in1711_1 = {c988};
    assign in1711_2 = {c989};
    Full_Adder FA_1711(s1711, c1711, in1711_1, in1711_2, s407[0]);
    wire[0:0] s1712, in1712_1, in1712_2;
    wire c1712;
    assign in1712_1 = {c991};
    assign in1712_2 = {c992};
    Full_Adder FA_1712(s1712, c1712, in1712_1, in1712_2, c990);
    wire[0:0] s1713, in1713_1, in1713_2;
    wire c1713;
    assign in1713_1 = {c994};
    assign in1713_2 = {c995};
    Full_Adder FA_1713(s1713, c1713, in1713_1, in1713_2, c993);
    wire[0:0] s1714, in1714_1, in1714_2;
    wire c1714;
    assign in1714_1 = {c997};
    assign in1714_2 = {c998};
    Full_Adder FA_1714(s1714, c1714, in1714_1, in1714_2, c996);
    wire[0:0] s1715, in1715_1, in1715_2;
    wire c1715;
    assign in1715_1 = {c1000};
    assign in1715_2 = {c1001};
    Full_Adder FA_1715(s1715, c1715, in1715_1, in1715_2, c999);
    wire[0:0] s1716, in1716_1, in1716_2;
    wire c1716;
    assign in1716_1 = {s1003[0]};
    assign in1716_2 = {s1004[0]};
    Full_Adder FA_1716(s1716, c1716, in1716_1, in1716_2, s1002[0]);
    wire[0:0] s1717, in1717_1, in1717_2;
    wire c1717;
    assign in1717_1 = {s1006[0]};
    assign in1717_2 = {s1007[0]};
    Full_Adder FA_1717(s1717, c1717, in1717_1, in1717_2, s1005[0]);
    wire[0:0] s1718, in1718_1, in1718_2;
    wire c1718;
    assign in1718_1 = {s1009[0]};
    assign in1718_2 = {s1010[0]};
    Full_Adder FA_1718(s1718, c1718, in1718_1, in1718_2, s1008[0]);
    wire[0:0] s1719, in1719_1, in1719_2;
    wire c1719;
    assign in1719_1 = {s1012[0]};
    assign in1719_2 = {s1013[0]};
    Full_Adder FA_1719(s1719, c1719, in1719_1, in1719_2, s1011[0]);
    wire[0:0] s1720, in1720_1, in1720_2;
    wire c1720;
    assign in1720_1 = {c1002};
    assign in1720_2 = {c1003};
    Full_Adder FA_1720(s1720, c1720, in1720_1, in1720_2, s417[0]);
    wire[0:0] s1721, in1721_1, in1721_2;
    wire c1721;
    assign in1721_1 = {c1005};
    assign in1721_2 = {c1006};
    Full_Adder FA_1721(s1721, c1721, in1721_1, in1721_2, c1004);
    wire[0:0] s1722, in1722_1, in1722_2;
    wire c1722;
    assign in1722_1 = {c1008};
    assign in1722_2 = {c1009};
    Full_Adder FA_1722(s1722, c1722, in1722_1, in1722_2, c1007);
    wire[0:0] s1723, in1723_1, in1723_2;
    wire c1723;
    assign in1723_1 = {c1011};
    assign in1723_2 = {c1012};
    Full_Adder FA_1723(s1723, c1723, in1723_1, in1723_2, c1010);
    wire[0:0] s1724, in1724_1, in1724_2;
    wire c1724;
    assign in1724_1 = {c1014};
    assign in1724_2 = {c1015};
    Full_Adder FA_1724(s1724, c1724, in1724_1, in1724_2, c1013);
    wire[0:0] s1725, in1725_1, in1725_2;
    wire c1725;
    assign in1725_1 = {s1017[0]};
    assign in1725_2 = {s1018[0]};
    Full_Adder FA_1725(s1725, c1725, in1725_1, in1725_2, s1016[0]);
    wire[0:0] s1726, in1726_1, in1726_2;
    wire c1726;
    assign in1726_1 = {s1020[0]};
    assign in1726_2 = {s1021[0]};
    Full_Adder FA_1726(s1726, c1726, in1726_1, in1726_2, s1019[0]);
    wire[0:0] s1727, in1727_1, in1727_2;
    wire c1727;
    assign in1727_1 = {s1023[0]};
    assign in1727_2 = {s1024[0]};
    Full_Adder FA_1727(s1727, c1727, in1727_1, in1727_2, s1022[0]);
    wire[0:0] s1728, in1728_1, in1728_2;
    wire c1728;
    assign in1728_1 = {s1026[0]};
    assign in1728_2 = {s1027[0]};
    Full_Adder FA_1728(s1728, c1728, in1728_1, in1728_2, s1025[0]);
    wire[0:0] s1729, in1729_1, in1729_2;
    wire c1729;
    assign in1729_1 = {c1016};
    assign in1729_2 = {c1017};
    Full_Adder FA_1729(s1729, c1729, in1729_1, in1729_2, s426[0]);
    wire[0:0] s1730, in1730_1, in1730_2;
    wire c1730;
    assign in1730_1 = {c1019};
    assign in1730_2 = {c1020};
    Full_Adder FA_1730(s1730, c1730, in1730_1, in1730_2, c1018);
    wire[0:0] s1731, in1731_1, in1731_2;
    wire c1731;
    assign in1731_1 = {c1022};
    assign in1731_2 = {c1023};
    Full_Adder FA_1731(s1731, c1731, in1731_1, in1731_2, c1021);
    wire[0:0] s1732, in1732_1, in1732_2;
    wire c1732;
    assign in1732_1 = {c1025};
    assign in1732_2 = {c1026};
    Full_Adder FA_1732(s1732, c1732, in1732_1, in1732_2, c1024);
    wire[0:0] s1733, in1733_1, in1733_2;
    wire c1733;
    assign in1733_1 = {c1028};
    assign in1733_2 = {c1029};
    Full_Adder FA_1733(s1733, c1733, in1733_1, in1733_2, c1027);
    wire[0:0] s1734, in1734_1, in1734_2;
    wire c1734;
    assign in1734_1 = {s1031[0]};
    assign in1734_2 = {s1032[0]};
    Full_Adder FA_1734(s1734, c1734, in1734_1, in1734_2, s1030[0]);
    wire[0:0] s1735, in1735_1, in1735_2;
    wire c1735;
    assign in1735_1 = {s1034[0]};
    assign in1735_2 = {s1035[0]};
    Full_Adder FA_1735(s1735, c1735, in1735_1, in1735_2, s1033[0]);
    wire[0:0] s1736, in1736_1, in1736_2;
    wire c1736;
    assign in1736_1 = {s1037[0]};
    assign in1736_2 = {s1038[0]};
    Full_Adder FA_1736(s1736, c1736, in1736_1, in1736_2, s1036[0]);
    wire[0:0] s1737, in1737_1, in1737_2;
    wire c1737;
    assign in1737_1 = {s1040[0]};
    assign in1737_2 = {s1041[0]};
    Full_Adder FA_1737(s1737, c1737, in1737_1, in1737_2, s1039[0]);
    wire[0:0] s1738, in1738_1, in1738_2;
    wire c1738;
    assign in1738_1 = {c1030};
    assign in1738_2 = {c1031};
    Full_Adder FA_1738(s1738, c1738, in1738_1, in1738_2, s434[0]);
    wire[0:0] s1739, in1739_1, in1739_2;
    wire c1739;
    assign in1739_1 = {c1033};
    assign in1739_2 = {c1034};
    Full_Adder FA_1739(s1739, c1739, in1739_1, in1739_2, c1032);
    wire[0:0] s1740, in1740_1, in1740_2;
    wire c1740;
    assign in1740_1 = {c1036};
    assign in1740_2 = {c1037};
    Full_Adder FA_1740(s1740, c1740, in1740_1, in1740_2, c1035);
    wire[0:0] s1741, in1741_1, in1741_2;
    wire c1741;
    assign in1741_1 = {c1039};
    assign in1741_2 = {c1040};
    Full_Adder FA_1741(s1741, c1741, in1741_1, in1741_2, c1038);
    wire[0:0] s1742, in1742_1, in1742_2;
    wire c1742;
    assign in1742_1 = {c1042};
    assign in1742_2 = {c1043};
    Full_Adder FA_1742(s1742, c1742, in1742_1, in1742_2, c1041);
    wire[0:0] s1743, in1743_1, in1743_2;
    wire c1743;
    assign in1743_1 = {s1045[0]};
    assign in1743_2 = {s1046[0]};
    Full_Adder FA_1743(s1743, c1743, in1743_1, in1743_2, s1044[0]);
    wire[0:0] s1744, in1744_1, in1744_2;
    wire c1744;
    assign in1744_1 = {s1048[0]};
    assign in1744_2 = {s1049[0]};
    Full_Adder FA_1744(s1744, c1744, in1744_1, in1744_2, s1047[0]);
    wire[0:0] s1745, in1745_1, in1745_2;
    wire c1745;
    assign in1745_1 = {s1051[0]};
    assign in1745_2 = {s1052[0]};
    Full_Adder FA_1745(s1745, c1745, in1745_1, in1745_2, s1050[0]);
    wire[0:0] s1746, in1746_1, in1746_2;
    wire c1746;
    assign in1746_1 = {s1054[0]};
    assign in1746_2 = {s1055[0]};
    Full_Adder FA_1746(s1746, c1746, in1746_1, in1746_2, s1053[0]);
    wire[0:0] s1747, in1747_1, in1747_2;
    wire c1747;
    assign in1747_1 = {c1044};
    assign in1747_2 = {c1045};
    Full_Adder FA_1747(s1747, c1747, in1747_1, in1747_2, s441[0]);
    wire[0:0] s1748, in1748_1, in1748_2;
    wire c1748;
    assign in1748_1 = {c1047};
    assign in1748_2 = {c1048};
    Full_Adder FA_1748(s1748, c1748, in1748_1, in1748_2, c1046);
    wire[0:0] s1749, in1749_1, in1749_2;
    wire c1749;
    assign in1749_1 = {c1050};
    assign in1749_2 = {c1051};
    Full_Adder FA_1749(s1749, c1749, in1749_1, in1749_2, c1049);
    wire[0:0] s1750, in1750_1, in1750_2;
    wire c1750;
    assign in1750_1 = {c1053};
    assign in1750_2 = {c1054};
    Full_Adder FA_1750(s1750, c1750, in1750_1, in1750_2, c1052);
    wire[0:0] s1751, in1751_1, in1751_2;
    wire c1751;
    assign in1751_1 = {c1056};
    assign in1751_2 = {c1057};
    Full_Adder FA_1751(s1751, c1751, in1751_1, in1751_2, c1055);
    wire[0:0] s1752, in1752_1, in1752_2;
    wire c1752;
    assign in1752_1 = {s1059[0]};
    assign in1752_2 = {s1060[0]};
    Full_Adder FA_1752(s1752, c1752, in1752_1, in1752_2, s1058[0]);
    wire[0:0] s1753, in1753_1, in1753_2;
    wire c1753;
    assign in1753_1 = {s1062[0]};
    assign in1753_2 = {s1063[0]};
    Full_Adder FA_1753(s1753, c1753, in1753_1, in1753_2, s1061[0]);
    wire[0:0] s1754, in1754_1, in1754_2;
    wire c1754;
    assign in1754_1 = {s1065[0]};
    assign in1754_2 = {s1066[0]};
    Full_Adder FA_1754(s1754, c1754, in1754_1, in1754_2, s1064[0]);
    wire[0:0] s1755, in1755_1, in1755_2;
    wire c1755;
    assign in1755_1 = {s1068[0]};
    assign in1755_2 = {s1069[0]};
    Full_Adder FA_1755(s1755, c1755, in1755_1, in1755_2, s1067[0]);
    wire[0:0] s1756, in1756_1, in1756_2;
    wire c1756;
    assign in1756_1 = {c1058};
    assign in1756_2 = {c1059};
    Full_Adder FA_1756(s1756, c1756, in1756_1, in1756_2, s447[0]);
    wire[0:0] s1757, in1757_1, in1757_2;
    wire c1757;
    assign in1757_1 = {c1061};
    assign in1757_2 = {c1062};
    Full_Adder FA_1757(s1757, c1757, in1757_1, in1757_2, c1060);
    wire[0:0] s1758, in1758_1, in1758_2;
    wire c1758;
    assign in1758_1 = {c1064};
    assign in1758_2 = {c1065};
    Full_Adder FA_1758(s1758, c1758, in1758_1, in1758_2, c1063);
    wire[0:0] s1759, in1759_1, in1759_2;
    wire c1759;
    assign in1759_1 = {c1067};
    assign in1759_2 = {c1068};
    Full_Adder FA_1759(s1759, c1759, in1759_1, in1759_2, c1066);
    wire[0:0] s1760, in1760_1, in1760_2;
    wire c1760;
    assign in1760_1 = {c1070};
    assign in1760_2 = {c1071};
    Full_Adder FA_1760(s1760, c1760, in1760_1, in1760_2, c1069);
    wire[0:0] s1761, in1761_1, in1761_2;
    wire c1761;
    assign in1761_1 = {s1073[0]};
    assign in1761_2 = {s1074[0]};
    Full_Adder FA_1761(s1761, c1761, in1761_1, in1761_2, s1072[0]);
    wire[0:0] s1762, in1762_1, in1762_2;
    wire c1762;
    assign in1762_1 = {s1076[0]};
    assign in1762_2 = {s1077[0]};
    Full_Adder FA_1762(s1762, c1762, in1762_1, in1762_2, s1075[0]);
    wire[0:0] s1763, in1763_1, in1763_2;
    wire c1763;
    assign in1763_1 = {s1079[0]};
    assign in1763_2 = {s1080[0]};
    Full_Adder FA_1763(s1763, c1763, in1763_1, in1763_2, s1078[0]);
    wire[0:0] s1764, in1764_1, in1764_2;
    wire c1764;
    assign in1764_1 = {s1082[0]};
    assign in1764_2 = {s1083[0]};
    Full_Adder FA_1764(s1764, c1764, in1764_1, in1764_2, s1081[0]);
    wire[0:0] s1765, in1765_1, in1765_2;
    wire c1765;
    assign in1765_1 = {c1072};
    assign in1765_2 = {c1073};
    Full_Adder FA_1765(s1765, c1765, in1765_1, in1765_2, s452[0]);
    wire[0:0] s1766, in1766_1, in1766_2;
    wire c1766;
    assign in1766_1 = {c1075};
    assign in1766_2 = {c1076};
    Full_Adder FA_1766(s1766, c1766, in1766_1, in1766_2, c1074);
    wire[0:0] s1767, in1767_1, in1767_2;
    wire c1767;
    assign in1767_1 = {c1078};
    assign in1767_2 = {c1079};
    Full_Adder FA_1767(s1767, c1767, in1767_1, in1767_2, c1077);
    wire[0:0] s1768, in1768_1, in1768_2;
    wire c1768;
    assign in1768_1 = {c1081};
    assign in1768_2 = {c1082};
    Full_Adder FA_1768(s1768, c1768, in1768_1, in1768_2, c1080);
    wire[0:0] s1769, in1769_1, in1769_2;
    wire c1769;
    assign in1769_1 = {c1084};
    assign in1769_2 = {c1085};
    Full_Adder FA_1769(s1769, c1769, in1769_1, in1769_2, c1083);
    wire[0:0] s1770, in1770_1, in1770_2;
    wire c1770;
    assign in1770_1 = {s1087[0]};
    assign in1770_2 = {s1088[0]};
    Full_Adder FA_1770(s1770, c1770, in1770_1, in1770_2, s1086[0]);
    wire[0:0] s1771, in1771_1, in1771_2;
    wire c1771;
    assign in1771_1 = {s1090[0]};
    assign in1771_2 = {s1091[0]};
    Full_Adder FA_1771(s1771, c1771, in1771_1, in1771_2, s1089[0]);
    wire[0:0] s1772, in1772_1, in1772_2;
    wire c1772;
    assign in1772_1 = {s1093[0]};
    assign in1772_2 = {s1094[0]};
    Full_Adder FA_1772(s1772, c1772, in1772_1, in1772_2, s1092[0]);
    wire[0:0] s1773, in1773_1, in1773_2;
    wire c1773;
    assign in1773_1 = {s1096[0]};
    assign in1773_2 = {s1097[0]};
    Full_Adder FA_1773(s1773, c1773, in1773_1, in1773_2, s1095[0]);
    wire[0:0] s1774, in1774_1, in1774_2;
    wire c1774;
    assign in1774_1 = {c1086};
    assign in1774_2 = {c1087};
    Full_Adder FA_1774(s1774, c1774, in1774_1, in1774_2, s456[0]);
    wire[0:0] s1775, in1775_1, in1775_2;
    wire c1775;
    assign in1775_1 = {c1089};
    assign in1775_2 = {c1090};
    Full_Adder FA_1775(s1775, c1775, in1775_1, in1775_2, c1088);
    wire[0:0] s1776, in1776_1, in1776_2;
    wire c1776;
    assign in1776_1 = {c1092};
    assign in1776_2 = {c1093};
    Full_Adder FA_1776(s1776, c1776, in1776_1, in1776_2, c1091);
    wire[0:0] s1777, in1777_1, in1777_2;
    wire c1777;
    assign in1777_1 = {c1095};
    assign in1777_2 = {c1096};
    Full_Adder FA_1777(s1777, c1777, in1777_1, in1777_2, c1094);
    wire[0:0] s1778, in1778_1, in1778_2;
    wire c1778;
    assign in1778_1 = {c1098};
    assign in1778_2 = {c1099};
    Full_Adder FA_1778(s1778, c1778, in1778_1, in1778_2, c1097);
    wire[0:0] s1779, in1779_1, in1779_2;
    wire c1779;
    assign in1779_1 = {s1101[0]};
    assign in1779_2 = {s1102[0]};
    Full_Adder FA_1779(s1779, c1779, in1779_1, in1779_2, s1100[0]);
    wire[0:0] s1780, in1780_1, in1780_2;
    wire c1780;
    assign in1780_1 = {s1104[0]};
    assign in1780_2 = {s1105[0]};
    Full_Adder FA_1780(s1780, c1780, in1780_1, in1780_2, s1103[0]);
    wire[0:0] s1781, in1781_1, in1781_2;
    wire c1781;
    assign in1781_1 = {s1107[0]};
    assign in1781_2 = {s1108[0]};
    Full_Adder FA_1781(s1781, c1781, in1781_1, in1781_2, s1106[0]);
    wire[0:0] s1782, in1782_1, in1782_2;
    wire c1782;
    assign in1782_1 = {s1110[0]};
    assign in1782_2 = {s1111[0]};
    Full_Adder FA_1782(s1782, c1782, in1782_1, in1782_2, s1109[0]);
    wire[0:0] s1783, in1783_1, in1783_2;
    wire c1783;
    assign in1783_1 = {c1100};
    assign in1783_2 = {c1101};
    Full_Adder FA_1783(s1783, c1783, in1783_1, in1783_2, s459[0]);
    wire[0:0] s1784, in1784_1, in1784_2;
    wire c1784;
    assign in1784_1 = {c1103};
    assign in1784_2 = {c1104};
    Full_Adder FA_1784(s1784, c1784, in1784_1, in1784_2, c1102);
    wire[0:0] s1785, in1785_1, in1785_2;
    wire c1785;
    assign in1785_1 = {c1106};
    assign in1785_2 = {c1107};
    Full_Adder FA_1785(s1785, c1785, in1785_1, in1785_2, c1105);
    wire[0:0] s1786, in1786_1, in1786_2;
    wire c1786;
    assign in1786_1 = {c1109};
    assign in1786_2 = {c1110};
    Full_Adder FA_1786(s1786, c1786, in1786_1, in1786_2, c1108);
    wire[0:0] s1787, in1787_1, in1787_2;
    wire c1787;
    assign in1787_1 = {c1112};
    assign in1787_2 = {c1113};
    Full_Adder FA_1787(s1787, c1787, in1787_1, in1787_2, c1111);
    wire[0:0] s1788, in1788_1, in1788_2;
    wire c1788;
    assign in1788_1 = {s1115[0]};
    assign in1788_2 = {s1116[0]};
    Full_Adder FA_1788(s1788, c1788, in1788_1, in1788_2, s1114[0]);
    wire[0:0] s1789, in1789_1, in1789_2;
    wire c1789;
    assign in1789_1 = {s1118[0]};
    assign in1789_2 = {s1119[0]};
    Full_Adder FA_1789(s1789, c1789, in1789_1, in1789_2, s1117[0]);
    wire[0:0] s1790, in1790_1, in1790_2;
    wire c1790;
    assign in1790_1 = {s1121[0]};
    assign in1790_2 = {s1122[0]};
    Full_Adder FA_1790(s1790, c1790, in1790_1, in1790_2, s1120[0]);
    wire[0:0] s1791, in1791_1, in1791_2;
    wire c1791;
    assign in1791_1 = {s1124[0]};
    assign in1791_2 = {s1125[0]};
    Full_Adder FA_1791(s1791, c1791, in1791_1, in1791_2, s1123[0]);
    wire[0:0] s1792, in1792_1, in1792_2;
    wire c1792;
    assign in1792_1 = {c1114};
    assign in1792_2 = {c1115};
    Full_Adder FA_1792(s1792, c1792, in1792_1, in1792_2, s461[0]);
    wire[0:0] s1793, in1793_1, in1793_2;
    wire c1793;
    assign in1793_1 = {c1117};
    assign in1793_2 = {c1118};
    Full_Adder FA_1793(s1793, c1793, in1793_1, in1793_2, c1116);
    wire[0:0] s1794, in1794_1, in1794_2;
    wire c1794;
    assign in1794_1 = {c1120};
    assign in1794_2 = {c1121};
    Full_Adder FA_1794(s1794, c1794, in1794_1, in1794_2, c1119);
    wire[0:0] s1795, in1795_1, in1795_2;
    wire c1795;
    assign in1795_1 = {c1123};
    assign in1795_2 = {c1124};
    Full_Adder FA_1795(s1795, c1795, in1795_1, in1795_2, c1122);
    wire[0:0] s1796, in1796_1, in1796_2;
    wire c1796;
    assign in1796_1 = {c1126};
    assign in1796_2 = {c1127};
    Full_Adder FA_1796(s1796, c1796, in1796_1, in1796_2, c1125);
    wire[0:0] s1797, in1797_1, in1797_2;
    wire c1797;
    assign in1797_1 = {s1129[0]};
    assign in1797_2 = {s1130[0]};
    Full_Adder FA_1797(s1797, c1797, in1797_1, in1797_2, s1128[0]);
    wire[0:0] s1798, in1798_1, in1798_2;
    wire c1798;
    assign in1798_1 = {s1132[0]};
    assign in1798_2 = {s1133[0]};
    Full_Adder FA_1798(s1798, c1798, in1798_1, in1798_2, s1131[0]);
    wire[0:0] s1799, in1799_1, in1799_2;
    wire c1799;
    assign in1799_1 = {s1135[0]};
    assign in1799_2 = {s1136[0]};
    Full_Adder FA_1799(s1799, c1799, in1799_1, in1799_2, s1134[0]);
    wire[0:0] s1800, in1800_1, in1800_2;
    wire c1800;
    assign in1800_1 = {s1138[0]};
    assign in1800_2 = {s1139[0]};
    Full_Adder FA_1800(s1800, c1800, in1800_1, in1800_2, s1137[0]);
    wire[0:0] s1801, in1801_1, in1801_2;
    wire c1801;
    assign in1801_1 = {c1128};
    assign in1801_2 = {c1129};
    Full_Adder FA_1801(s1801, c1801, in1801_1, in1801_2, s462[0]);
    wire[0:0] s1802, in1802_1, in1802_2;
    wire c1802;
    assign in1802_1 = {c1131};
    assign in1802_2 = {c1132};
    Full_Adder FA_1802(s1802, c1802, in1802_1, in1802_2, c1130);
    wire[0:0] s1803, in1803_1, in1803_2;
    wire c1803;
    assign in1803_1 = {c1134};
    assign in1803_2 = {c1135};
    Full_Adder FA_1803(s1803, c1803, in1803_1, in1803_2, c1133);
    wire[0:0] s1804, in1804_1, in1804_2;
    wire c1804;
    assign in1804_1 = {c1137};
    assign in1804_2 = {c1138};
    Full_Adder FA_1804(s1804, c1804, in1804_1, in1804_2, c1136);
    wire[0:0] s1805, in1805_1, in1805_2;
    wire c1805;
    assign in1805_1 = {c1140};
    assign in1805_2 = {c1141};
    Full_Adder FA_1805(s1805, c1805, in1805_1, in1805_2, c1139);
    wire[0:0] s1806, in1806_1, in1806_2;
    wire c1806;
    assign in1806_1 = {s1143[0]};
    assign in1806_2 = {s1144[0]};
    Full_Adder FA_1806(s1806, c1806, in1806_1, in1806_2, s1142[0]);
    wire[0:0] s1807, in1807_1, in1807_2;
    wire c1807;
    assign in1807_1 = {s1146[0]};
    assign in1807_2 = {s1147[0]};
    Full_Adder FA_1807(s1807, c1807, in1807_1, in1807_2, s1145[0]);
    wire[0:0] s1808, in1808_1, in1808_2;
    wire c1808;
    assign in1808_1 = {s1149[0]};
    assign in1808_2 = {s1150[0]};
    Full_Adder FA_1808(s1808, c1808, in1808_1, in1808_2, s1148[0]);
    wire[0:0] s1809, in1809_1, in1809_2;
    wire c1809;
    assign in1809_1 = {s1152[0]};
    assign in1809_2 = {s1153[0]};
    Full_Adder FA_1809(s1809, c1809, in1809_1, in1809_2, s1151[0]);
    wire[0:0] s1810, in1810_1, in1810_2;
    wire c1810;
    assign in1810_1 = {c1142};
    assign in1810_2 = {c1143};
    Full_Adder FA_1810(s1810, c1810, in1810_1, in1810_2, c462);
    wire[0:0] s1811, in1811_1, in1811_2;
    wire c1811;
    assign in1811_1 = {c1145};
    assign in1811_2 = {c1146};
    Full_Adder FA_1811(s1811, c1811, in1811_1, in1811_2, c1144);
    wire[0:0] s1812, in1812_1, in1812_2;
    wire c1812;
    assign in1812_1 = {c1148};
    assign in1812_2 = {c1149};
    Full_Adder FA_1812(s1812, c1812, in1812_1, in1812_2, c1147);
    wire[0:0] s1813, in1813_1, in1813_2;
    wire c1813;
    assign in1813_1 = {c1151};
    assign in1813_2 = {c1152};
    Full_Adder FA_1813(s1813, c1813, in1813_1, in1813_2, c1150);
    wire[0:0] s1814, in1814_1, in1814_2;
    wire c1814;
    assign in1814_1 = {c1154};
    assign in1814_2 = {c1155};
    Full_Adder FA_1814(s1814, c1814, in1814_1, in1814_2, c1153);
    wire[0:0] s1815, in1815_1, in1815_2;
    wire c1815;
    assign in1815_1 = {s1157[0]};
    assign in1815_2 = {s1158[0]};
    Full_Adder FA_1815(s1815, c1815, in1815_1, in1815_2, s1156[0]);
    wire[0:0] s1816, in1816_1, in1816_2;
    wire c1816;
    assign in1816_1 = {s1160[0]};
    assign in1816_2 = {s1161[0]};
    Full_Adder FA_1816(s1816, c1816, in1816_1, in1816_2, s1159[0]);
    wire[0:0] s1817, in1817_1, in1817_2;
    wire c1817;
    assign in1817_1 = {s1163[0]};
    assign in1817_2 = {s1164[0]};
    Full_Adder FA_1817(s1817, c1817, in1817_1, in1817_2, s1162[0]);
    wire[0:0] s1818, in1818_1, in1818_2;
    wire c1818;
    assign in1818_1 = {s1166[0]};
    assign in1818_2 = {s1167[0]};
    Full_Adder FA_1818(s1818, c1818, in1818_1, in1818_2, s1165[0]);
    wire[0:0] s1819, in1819_1, in1819_2;
    wire c1819;
    assign in1819_1 = {pp63[23]};
    assign in1819_2 = {c1156};
    Full_Adder FA_1819(s1819, c1819, in1819_1, in1819_2, pp62[24]);
    wire[0:0] s1820, in1820_1, in1820_2;
    wire c1820;
    assign in1820_1 = {c1158};
    assign in1820_2 = {c1159};
    Full_Adder FA_1820(s1820, c1820, in1820_1, in1820_2, c1157);
    wire[0:0] s1821, in1821_1, in1821_2;
    wire c1821;
    assign in1821_1 = {c1161};
    assign in1821_2 = {c1162};
    Full_Adder FA_1821(s1821, c1821, in1821_1, in1821_2, c1160);
    wire[0:0] s1822, in1822_1, in1822_2;
    wire c1822;
    assign in1822_1 = {c1164};
    assign in1822_2 = {c1165};
    Full_Adder FA_1822(s1822, c1822, in1822_1, in1822_2, c1163);
    wire[0:0] s1823, in1823_1, in1823_2;
    wire c1823;
    assign in1823_1 = {c1167};
    assign in1823_2 = {c1168};
    Full_Adder FA_1823(s1823, c1823, in1823_1, in1823_2, c1166);
    wire[0:0] s1824, in1824_1, in1824_2;
    wire c1824;
    assign in1824_1 = {s1170[0]};
    assign in1824_2 = {s1171[0]};
    Full_Adder FA_1824(s1824, c1824, in1824_1, in1824_2, c1169);
    wire[0:0] s1825, in1825_1, in1825_2;
    wire c1825;
    assign in1825_1 = {s1173[0]};
    assign in1825_2 = {s1174[0]};
    Full_Adder FA_1825(s1825, c1825, in1825_1, in1825_2, s1172[0]);
    wire[0:0] s1826, in1826_1, in1826_2;
    wire c1826;
    assign in1826_1 = {s1176[0]};
    assign in1826_2 = {s1177[0]};
    Full_Adder FA_1826(s1826, c1826, in1826_1, in1826_2, s1175[0]);
    wire[0:0] s1827, in1827_1, in1827_2;
    wire c1827;
    assign in1827_1 = {s1179[0]};
    assign in1827_2 = {s1180[0]};
    Full_Adder FA_1827(s1827, c1827, in1827_1, in1827_2, s1178[0]);
    wire[0:0] s1828, in1828_1, in1828_2;
    wire c1828;
    assign in1828_1 = {pp61[26]};
    assign in1828_2 = {pp62[25]};
    Full_Adder FA_1828(s1828, c1828, in1828_1, in1828_2, pp60[27]);
    wire[0:0] s1829, in1829_1, in1829_2;
    wire c1829;
    assign in1829_1 = {c1170};
    assign in1829_2 = {c1171};
    Full_Adder FA_1829(s1829, c1829, in1829_1, in1829_2, pp63[24]);
    wire[0:0] s1830, in1830_1, in1830_2;
    wire c1830;
    assign in1830_1 = {c1173};
    assign in1830_2 = {c1174};
    Full_Adder FA_1830(s1830, c1830, in1830_1, in1830_2, c1172);
    wire[0:0] s1831, in1831_1, in1831_2;
    wire c1831;
    assign in1831_1 = {c1176};
    assign in1831_2 = {c1177};
    Full_Adder FA_1831(s1831, c1831, in1831_1, in1831_2, c1175);
    wire[0:0] s1832, in1832_1, in1832_2;
    wire c1832;
    assign in1832_1 = {c1179};
    assign in1832_2 = {c1180};
    Full_Adder FA_1832(s1832, c1832, in1832_1, in1832_2, c1178);
    wire[0:0] s1833, in1833_1, in1833_2;
    wire c1833;
    assign in1833_1 = {c1182};
    assign in1833_2 = {s1183[0]};
    Full_Adder FA_1833(s1833, c1833, in1833_1, in1833_2, c1181);
    wire[0:0] s1834, in1834_1, in1834_2;
    wire c1834;
    assign in1834_1 = {s1185[0]};
    assign in1834_2 = {s1186[0]};
    Full_Adder FA_1834(s1834, c1834, in1834_1, in1834_2, s1184[0]);
    wire[0:0] s1835, in1835_1, in1835_2;
    wire c1835;
    assign in1835_1 = {s1188[0]};
    assign in1835_2 = {s1189[0]};
    Full_Adder FA_1835(s1835, c1835, in1835_1, in1835_2, s1187[0]);
    wire[0:0] s1836, in1836_1, in1836_2;
    wire c1836;
    assign in1836_1 = {s1191[0]};
    assign in1836_2 = {s1192[0]};
    Full_Adder FA_1836(s1836, c1836, in1836_1, in1836_2, s1190[0]);
    wire[0:0] s1837, in1837_1, in1837_2;
    wire c1837;
    assign in1837_1 = {pp59[29]};
    assign in1837_2 = {pp60[28]};
    Full_Adder FA_1837(s1837, c1837, in1837_1, in1837_2, pp58[30]);
    wire[0:0] s1838, in1838_1, in1838_2;
    wire c1838;
    assign in1838_1 = {pp62[26]};
    assign in1838_2 = {pp63[25]};
    Full_Adder FA_1838(s1838, c1838, in1838_1, in1838_2, pp61[27]);
    wire[0:0] s1839, in1839_1, in1839_2;
    wire c1839;
    assign in1839_1 = {c1184};
    assign in1839_2 = {c1185};
    Full_Adder FA_1839(s1839, c1839, in1839_1, in1839_2, c1183);
    wire[0:0] s1840, in1840_1, in1840_2;
    wire c1840;
    assign in1840_1 = {c1187};
    assign in1840_2 = {c1188};
    Full_Adder FA_1840(s1840, c1840, in1840_1, in1840_2, c1186);
    wire[0:0] s1841, in1841_1, in1841_2;
    wire c1841;
    assign in1841_1 = {c1190};
    assign in1841_2 = {c1191};
    Full_Adder FA_1841(s1841, c1841, in1841_1, in1841_2, c1189);
    wire[0:0] s1842, in1842_1, in1842_2;
    wire c1842;
    assign in1842_1 = {c1193};
    assign in1842_2 = {c1194};
    Full_Adder FA_1842(s1842, c1842, in1842_1, in1842_2, c1192);
    wire[0:0] s1843, in1843_1, in1843_2;
    wire c1843;
    assign in1843_1 = {s1196[0]};
    assign in1843_2 = {s1197[0]};
    Full_Adder FA_1843(s1843, c1843, in1843_1, in1843_2, s1195[0]);
    wire[0:0] s1844, in1844_1, in1844_2;
    wire c1844;
    assign in1844_1 = {s1199[0]};
    assign in1844_2 = {s1200[0]};
    Full_Adder FA_1844(s1844, c1844, in1844_1, in1844_2, s1198[0]);
    wire[0:0] s1845, in1845_1, in1845_2;
    wire c1845;
    assign in1845_1 = {s1202[0]};
    assign in1845_2 = {s1203[0]};
    Full_Adder FA_1845(s1845, c1845, in1845_1, in1845_2, s1201[0]);
    wire[0:0] s1846, in1846_1, in1846_2;
    wire c1846;
    assign in1846_1 = {pp57[32]};
    assign in1846_2 = {pp58[31]};
    Full_Adder FA_1846(s1846, c1846, in1846_1, in1846_2, pp56[33]);
    wire[0:0] s1847, in1847_1, in1847_2;
    wire c1847;
    assign in1847_1 = {pp60[29]};
    assign in1847_2 = {pp61[28]};
    Full_Adder FA_1847(s1847, c1847, in1847_1, in1847_2, pp59[30]);
    wire[0:0] s1848, in1848_1, in1848_2;
    wire c1848;
    assign in1848_1 = {pp63[26]};
    assign in1848_2 = {c1195};
    Full_Adder FA_1848(s1848, c1848, in1848_1, in1848_2, pp62[27]);
    wire[0:0] s1849, in1849_1, in1849_2;
    wire c1849;
    assign in1849_1 = {c1197};
    assign in1849_2 = {c1198};
    Full_Adder FA_1849(s1849, c1849, in1849_1, in1849_2, c1196);
    wire[0:0] s1850, in1850_1, in1850_2;
    wire c1850;
    assign in1850_1 = {c1200};
    assign in1850_2 = {c1201};
    Full_Adder FA_1850(s1850, c1850, in1850_1, in1850_2, c1199);
    wire[0:0] s1851, in1851_1, in1851_2;
    wire c1851;
    assign in1851_1 = {c1203};
    assign in1851_2 = {c1204};
    Full_Adder FA_1851(s1851, c1851, in1851_1, in1851_2, c1202);
    wire[0:0] s1852, in1852_1, in1852_2;
    wire c1852;
    assign in1852_1 = {s1206[0]};
    assign in1852_2 = {s1207[0]};
    Full_Adder FA_1852(s1852, c1852, in1852_1, in1852_2, c1205);
    wire[0:0] s1853, in1853_1, in1853_2;
    wire c1853;
    assign in1853_1 = {s1209[0]};
    assign in1853_2 = {s1210[0]};
    Full_Adder FA_1853(s1853, c1853, in1853_1, in1853_2, s1208[0]);
    wire[0:0] s1854, in1854_1, in1854_2;
    wire c1854;
    assign in1854_1 = {s1212[0]};
    assign in1854_2 = {s1213[0]};
    Full_Adder FA_1854(s1854, c1854, in1854_1, in1854_2, s1211[0]);
    wire[0:0] s1855, in1855_1, in1855_2;
    wire c1855;
    assign in1855_1 = {pp55[35]};
    assign in1855_2 = {pp56[34]};
    Full_Adder FA_1855(s1855, c1855, in1855_1, in1855_2, pp54[36]);
    wire[0:0] s1856, in1856_1, in1856_2;
    wire c1856;
    assign in1856_1 = {pp58[32]};
    assign in1856_2 = {pp59[31]};
    Full_Adder FA_1856(s1856, c1856, in1856_1, in1856_2, pp57[33]);
    wire[0:0] s1857, in1857_1, in1857_2;
    wire c1857;
    assign in1857_1 = {pp61[29]};
    assign in1857_2 = {pp62[28]};
    Full_Adder FA_1857(s1857, c1857, in1857_1, in1857_2, pp60[30]);
    wire[0:0] s1858, in1858_1, in1858_2;
    wire c1858;
    assign in1858_1 = {c1206};
    assign in1858_2 = {c1207};
    Full_Adder FA_1858(s1858, c1858, in1858_1, in1858_2, pp63[27]);
    wire[0:0] s1859, in1859_1, in1859_2;
    wire c1859;
    assign in1859_1 = {c1209};
    assign in1859_2 = {c1210};
    Full_Adder FA_1859(s1859, c1859, in1859_1, in1859_2, c1208);
    wire[0:0] s1860, in1860_1, in1860_2;
    wire c1860;
    assign in1860_1 = {c1212};
    assign in1860_2 = {c1213};
    Full_Adder FA_1860(s1860, c1860, in1860_1, in1860_2, c1211);
    wire[0:0] s1861, in1861_1, in1861_2;
    wire c1861;
    assign in1861_1 = {c1215};
    assign in1861_2 = {s1216[0]};
    Full_Adder FA_1861(s1861, c1861, in1861_1, in1861_2, c1214);
    wire[0:0] s1862, in1862_1, in1862_2;
    wire c1862;
    assign in1862_1 = {s1218[0]};
    assign in1862_2 = {s1219[0]};
    Full_Adder FA_1862(s1862, c1862, in1862_1, in1862_2, s1217[0]);
    wire[0:0] s1863, in1863_1, in1863_2;
    wire c1863;
    assign in1863_1 = {s1221[0]};
    assign in1863_2 = {s1222[0]};
    Full_Adder FA_1863(s1863, c1863, in1863_1, in1863_2, s1220[0]);
    wire[0:0] s1864, in1864_1, in1864_2;
    wire c1864;
    assign in1864_1 = {pp53[38]};
    assign in1864_2 = {pp54[37]};
    Full_Adder FA_1864(s1864, c1864, in1864_1, in1864_2, pp52[39]);
    wire[0:0] s1865, in1865_1, in1865_2;
    wire c1865;
    assign in1865_1 = {pp56[35]};
    assign in1865_2 = {pp57[34]};
    Full_Adder FA_1865(s1865, c1865, in1865_1, in1865_2, pp55[36]);
    wire[0:0] s1866, in1866_1, in1866_2;
    wire c1866;
    assign in1866_1 = {pp59[32]};
    assign in1866_2 = {pp60[31]};
    Full_Adder FA_1866(s1866, c1866, in1866_1, in1866_2, pp58[33]);
    wire[0:0] s1867, in1867_1, in1867_2;
    wire c1867;
    assign in1867_1 = {pp62[29]};
    assign in1867_2 = {pp63[28]};
    Full_Adder FA_1867(s1867, c1867, in1867_1, in1867_2, pp61[30]);
    wire[0:0] s1868, in1868_1, in1868_2;
    wire c1868;
    assign in1868_1 = {c1217};
    assign in1868_2 = {c1218};
    Full_Adder FA_1868(s1868, c1868, in1868_1, in1868_2, c1216);
    wire[0:0] s1869, in1869_1, in1869_2;
    wire c1869;
    assign in1869_1 = {c1220};
    assign in1869_2 = {c1221};
    Full_Adder FA_1869(s1869, c1869, in1869_1, in1869_2, c1219);
    wire[0:0] s1870, in1870_1, in1870_2;
    wire c1870;
    assign in1870_1 = {c1223};
    assign in1870_2 = {c1224};
    Full_Adder FA_1870(s1870, c1870, in1870_1, in1870_2, c1222);
    wire[0:0] s1871, in1871_1, in1871_2;
    wire c1871;
    assign in1871_1 = {s1226[0]};
    assign in1871_2 = {s1227[0]};
    Full_Adder FA_1871(s1871, c1871, in1871_1, in1871_2, s1225[0]);
    wire[0:0] s1872, in1872_1, in1872_2;
    wire c1872;
    assign in1872_1 = {s1229[0]};
    assign in1872_2 = {s1230[0]};
    Full_Adder FA_1872(s1872, c1872, in1872_1, in1872_2, s1228[0]);
    wire[0:0] s1873, in1873_1, in1873_2;
    wire c1873;
    assign in1873_1 = {pp51[41]};
    assign in1873_2 = {pp52[40]};
    Full_Adder FA_1873(s1873, c1873, in1873_1, in1873_2, pp50[42]);
    wire[0:0] s1874, in1874_1, in1874_2;
    wire c1874;
    assign in1874_1 = {pp54[38]};
    assign in1874_2 = {pp55[37]};
    Full_Adder FA_1874(s1874, c1874, in1874_1, in1874_2, pp53[39]);
    wire[0:0] s1875, in1875_1, in1875_2;
    wire c1875;
    assign in1875_1 = {pp57[35]};
    assign in1875_2 = {pp58[34]};
    Full_Adder FA_1875(s1875, c1875, in1875_1, in1875_2, pp56[36]);
    wire[0:0] s1876, in1876_1, in1876_2;
    wire c1876;
    assign in1876_1 = {pp60[32]};
    assign in1876_2 = {pp61[31]};
    Full_Adder FA_1876(s1876, c1876, in1876_1, in1876_2, pp59[33]);
    wire[0:0] s1877, in1877_1, in1877_2;
    wire c1877;
    assign in1877_1 = {pp63[29]};
    assign in1877_2 = {c1225};
    Full_Adder FA_1877(s1877, c1877, in1877_1, in1877_2, pp62[30]);
    wire[0:0] s1878, in1878_1, in1878_2;
    wire c1878;
    assign in1878_1 = {c1227};
    assign in1878_2 = {c1228};
    Full_Adder FA_1878(s1878, c1878, in1878_1, in1878_2, c1226);
    wire[0:0] s1879, in1879_1, in1879_2;
    wire c1879;
    assign in1879_1 = {c1230};
    assign in1879_2 = {c1231};
    Full_Adder FA_1879(s1879, c1879, in1879_1, in1879_2, c1229);
    wire[0:0] s1880, in1880_1, in1880_2;
    wire c1880;
    assign in1880_1 = {s1233[0]};
    assign in1880_2 = {s1234[0]};
    Full_Adder FA_1880(s1880, c1880, in1880_1, in1880_2, c1232);
    wire[0:0] s1881, in1881_1, in1881_2;
    wire c1881;
    assign in1881_1 = {s1236[0]};
    assign in1881_2 = {s1237[0]};
    Full_Adder FA_1881(s1881, c1881, in1881_1, in1881_2, s1235[0]);
    wire[0:0] s1882, in1882_1, in1882_2;
    wire c1882;
    assign in1882_1 = {pp49[44]};
    assign in1882_2 = {pp50[43]};
    Full_Adder FA_1882(s1882, c1882, in1882_1, in1882_2, pp48[45]);
    wire[0:0] s1883, in1883_1, in1883_2;
    wire c1883;
    assign in1883_1 = {pp52[41]};
    assign in1883_2 = {pp53[40]};
    Full_Adder FA_1883(s1883, c1883, in1883_1, in1883_2, pp51[42]);
    wire[0:0] s1884, in1884_1, in1884_2;
    wire c1884;
    assign in1884_1 = {pp55[38]};
    assign in1884_2 = {pp56[37]};
    Full_Adder FA_1884(s1884, c1884, in1884_1, in1884_2, pp54[39]);
    wire[0:0] s1885, in1885_1, in1885_2;
    wire c1885;
    assign in1885_1 = {pp58[35]};
    assign in1885_2 = {pp59[34]};
    Full_Adder FA_1885(s1885, c1885, in1885_1, in1885_2, pp57[36]);
    wire[0:0] s1886, in1886_1, in1886_2;
    wire c1886;
    assign in1886_1 = {pp61[32]};
    assign in1886_2 = {pp62[31]};
    Full_Adder FA_1886(s1886, c1886, in1886_1, in1886_2, pp60[33]);
    wire[0:0] s1887, in1887_1, in1887_2;
    wire c1887;
    assign in1887_1 = {c1233};
    assign in1887_2 = {c1234};
    Full_Adder FA_1887(s1887, c1887, in1887_1, in1887_2, pp63[30]);
    wire[0:0] s1888, in1888_1, in1888_2;
    wire c1888;
    assign in1888_1 = {c1236};
    assign in1888_2 = {c1237};
    Full_Adder FA_1888(s1888, c1888, in1888_1, in1888_2, c1235);
    wire[0:0] s1889, in1889_1, in1889_2;
    wire c1889;
    assign in1889_1 = {c1239};
    assign in1889_2 = {s1240[0]};
    Full_Adder FA_1889(s1889, c1889, in1889_1, in1889_2, c1238);
    wire[0:0] s1890, in1890_1, in1890_2;
    wire c1890;
    assign in1890_1 = {s1242[0]};
    assign in1890_2 = {s1243[0]};
    Full_Adder FA_1890(s1890, c1890, in1890_1, in1890_2, s1241[0]);
    wire[0:0] s1891, in1891_1, in1891_2;
    wire c1891;
    assign in1891_1 = {pp47[47]};
    assign in1891_2 = {pp48[46]};
    Full_Adder FA_1891(s1891, c1891, in1891_1, in1891_2, pp46[48]);
    wire[0:0] s1892, in1892_1, in1892_2;
    wire c1892;
    assign in1892_1 = {pp50[44]};
    assign in1892_2 = {pp51[43]};
    Full_Adder FA_1892(s1892, c1892, in1892_1, in1892_2, pp49[45]);
    wire[0:0] s1893, in1893_1, in1893_2;
    wire c1893;
    assign in1893_1 = {pp53[41]};
    assign in1893_2 = {pp54[40]};
    Full_Adder FA_1893(s1893, c1893, in1893_1, in1893_2, pp52[42]);
    wire[0:0] s1894, in1894_1, in1894_2;
    wire c1894;
    assign in1894_1 = {pp56[38]};
    assign in1894_2 = {pp57[37]};
    Full_Adder FA_1894(s1894, c1894, in1894_1, in1894_2, pp55[39]);
    wire[0:0] s1895, in1895_1, in1895_2;
    wire c1895;
    assign in1895_1 = {pp59[35]};
    assign in1895_2 = {pp60[34]};
    Full_Adder FA_1895(s1895, c1895, in1895_1, in1895_2, pp58[36]);
    wire[0:0] s1896, in1896_1, in1896_2;
    wire c1896;
    assign in1896_1 = {pp62[32]};
    assign in1896_2 = {pp63[31]};
    Full_Adder FA_1896(s1896, c1896, in1896_1, in1896_2, pp61[33]);
    wire[0:0] s1897, in1897_1, in1897_2;
    wire c1897;
    assign in1897_1 = {c1241};
    assign in1897_2 = {c1242};
    Full_Adder FA_1897(s1897, c1897, in1897_1, in1897_2, c1240);
    wire[0:0] s1898, in1898_1, in1898_2;
    wire c1898;
    assign in1898_1 = {c1244};
    assign in1898_2 = {c1245};
    Full_Adder FA_1898(s1898, c1898, in1898_1, in1898_2, c1243);
    wire[0:0] s1899, in1899_1, in1899_2;
    wire c1899;
    assign in1899_1 = {s1247[0]};
    assign in1899_2 = {s1248[0]};
    Full_Adder FA_1899(s1899, c1899, in1899_1, in1899_2, s1246[0]);
    wire[0:0] s1900, in1900_1, in1900_2;
    wire c1900;
    assign in1900_1 = {pp45[50]};
    assign in1900_2 = {pp46[49]};
    Full_Adder FA_1900(s1900, c1900, in1900_1, in1900_2, pp44[51]);
    wire[0:0] s1901, in1901_1, in1901_2;
    wire c1901;
    assign in1901_1 = {pp48[47]};
    assign in1901_2 = {pp49[46]};
    Full_Adder FA_1901(s1901, c1901, in1901_1, in1901_2, pp47[48]);
    wire[0:0] s1902, in1902_1, in1902_2;
    wire c1902;
    assign in1902_1 = {pp51[44]};
    assign in1902_2 = {pp52[43]};
    Full_Adder FA_1902(s1902, c1902, in1902_1, in1902_2, pp50[45]);
    wire[0:0] s1903, in1903_1, in1903_2;
    wire c1903;
    assign in1903_1 = {pp54[41]};
    assign in1903_2 = {pp55[40]};
    Full_Adder FA_1903(s1903, c1903, in1903_1, in1903_2, pp53[42]);
    wire[0:0] s1904, in1904_1, in1904_2;
    wire c1904;
    assign in1904_1 = {pp57[38]};
    assign in1904_2 = {pp58[37]};
    Full_Adder FA_1904(s1904, c1904, in1904_1, in1904_2, pp56[39]);
    wire[0:0] s1905, in1905_1, in1905_2;
    wire c1905;
    assign in1905_1 = {pp60[35]};
    assign in1905_2 = {pp61[34]};
    Full_Adder FA_1905(s1905, c1905, in1905_1, in1905_2, pp59[36]);
    wire[0:0] s1906, in1906_1, in1906_2;
    wire c1906;
    assign in1906_1 = {pp63[32]};
    assign in1906_2 = {c1246};
    Full_Adder FA_1906(s1906, c1906, in1906_1, in1906_2, pp62[33]);
    wire[0:0] s1907, in1907_1, in1907_2;
    wire c1907;
    assign in1907_1 = {c1248};
    assign in1907_2 = {c1249};
    Full_Adder FA_1907(s1907, c1907, in1907_1, in1907_2, c1247);
    wire[0:0] s1908, in1908_1, in1908_2;
    wire c1908;
    assign in1908_1 = {s1251[0]};
    assign in1908_2 = {s1252[0]};
    Full_Adder FA_1908(s1908, c1908, in1908_1, in1908_2, c1250);
    wire[0:0] s1909, in1909_1, in1909_2;
    wire c1909;
    assign in1909_1 = {pp43[53]};
    assign in1909_2 = {pp44[52]};
    Full_Adder FA_1909(s1909, c1909, in1909_1, in1909_2, pp42[54]);
    wire[0:0] s1910, in1910_1, in1910_2;
    wire c1910;
    assign in1910_1 = {pp46[50]};
    assign in1910_2 = {pp47[49]};
    Full_Adder FA_1910(s1910, c1910, in1910_1, in1910_2, pp45[51]);
    wire[0:0] s1911, in1911_1, in1911_2;
    wire c1911;
    assign in1911_1 = {pp49[47]};
    assign in1911_2 = {pp50[46]};
    Full_Adder FA_1911(s1911, c1911, in1911_1, in1911_2, pp48[48]);
    wire[0:0] s1912, in1912_1, in1912_2;
    wire c1912;
    assign in1912_1 = {pp52[44]};
    assign in1912_2 = {pp53[43]};
    Full_Adder FA_1912(s1912, c1912, in1912_1, in1912_2, pp51[45]);
    wire[0:0] s1913, in1913_1, in1913_2;
    wire c1913;
    assign in1913_1 = {pp55[41]};
    assign in1913_2 = {pp56[40]};
    Full_Adder FA_1913(s1913, c1913, in1913_1, in1913_2, pp54[42]);
    wire[0:0] s1914, in1914_1, in1914_2;
    wire c1914;
    assign in1914_1 = {pp58[38]};
    assign in1914_2 = {pp59[37]};
    Full_Adder FA_1914(s1914, c1914, in1914_1, in1914_2, pp57[39]);
    wire[0:0] s1915, in1915_1, in1915_2;
    wire c1915;
    assign in1915_1 = {pp61[35]};
    assign in1915_2 = {pp62[34]};
    Full_Adder FA_1915(s1915, c1915, in1915_1, in1915_2, pp60[36]);
    wire[0:0] s1916, in1916_1, in1916_2;
    wire c1916;
    assign in1916_1 = {c1251};
    assign in1916_2 = {c1252};
    Full_Adder FA_1916(s1916, c1916, in1916_1, in1916_2, pp63[33]);
    wire[0:0] s1917, in1917_1, in1917_2;
    wire c1917;
    assign in1917_1 = {c1254};
    assign in1917_2 = {s1255[0]};
    Full_Adder FA_1917(s1917, c1917, in1917_1, in1917_2, c1253);
    wire[0:0] s1918, in1918_1, in1918_2;
    wire c1918;
    assign in1918_1 = {pp41[56]};
    assign in1918_2 = {pp42[55]};
    Full_Adder FA_1918(s1918, c1918, in1918_1, in1918_2, pp40[57]);
    wire[0:0] s1919, in1919_1, in1919_2;
    wire c1919;
    assign in1919_1 = {pp44[53]};
    assign in1919_2 = {pp45[52]};
    Full_Adder FA_1919(s1919, c1919, in1919_1, in1919_2, pp43[54]);
    wire[0:0] s1920, in1920_1, in1920_2;
    wire c1920;
    assign in1920_1 = {pp47[50]};
    assign in1920_2 = {pp48[49]};
    Full_Adder FA_1920(s1920, c1920, in1920_1, in1920_2, pp46[51]);
    wire[0:0] s1921, in1921_1, in1921_2;
    wire c1921;
    assign in1921_1 = {pp50[47]};
    assign in1921_2 = {pp51[46]};
    Full_Adder FA_1921(s1921, c1921, in1921_1, in1921_2, pp49[48]);
    wire[0:0] s1922, in1922_1, in1922_2;
    wire c1922;
    assign in1922_1 = {pp53[44]};
    assign in1922_2 = {pp54[43]};
    Full_Adder FA_1922(s1922, c1922, in1922_1, in1922_2, pp52[45]);
    wire[0:0] s1923, in1923_1, in1923_2;
    wire c1923;
    assign in1923_1 = {pp56[41]};
    assign in1923_2 = {pp57[40]};
    Full_Adder FA_1923(s1923, c1923, in1923_1, in1923_2, pp55[42]);
    wire[0:0] s1924, in1924_1, in1924_2;
    wire c1924;
    assign in1924_1 = {pp59[38]};
    assign in1924_2 = {pp60[37]};
    Full_Adder FA_1924(s1924, c1924, in1924_1, in1924_2, pp58[39]);
    wire[0:0] s1925, in1925_1, in1925_2;
    wire c1925;
    assign in1925_1 = {pp62[35]};
    assign in1925_2 = {pp63[34]};
    Full_Adder FA_1925(s1925, c1925, in1925_1, in1925_2, pp61[36]);
    wire[0:0] s1926, in1926_1, in1926_2;
    wire c1926;
    assign in1926_1 = {c1256};
    assign in1926_2 = {c1257};
    Full_Adder FA_1926(s1926, c1926, in1926_1, in1926_2, c1255);
    wire[0:0] s1927, in1927_1, in1927_2;
    wire c1927;
    assign in1927_1 = {pp39[59]};
    assign in1927_2 = {pp40[58]};
    Full_Adder FA_1927(s1927, c1927, in1927_1, in1927_2, pp38[60]);
    wire[0:0] s1928, in1928_1, in1928_2;
    wire c1928;
    assign in1928_1 = {pp42[56]};
    assign in1928_2 = {pp43[55]};
    Full_Adder FA_1928(s1928, c1928, in1928_1, in1928_2, pp41[57]);
    wire[0:0] s1929, in1929_1, in1929_2;
    wire c1929;
    assign in1929_1 = {pp45[53]};
    assign in1929_2 = {pp46[52]};
    Full_Adder FA_1929(s1929, c1929, in1929_1, in1929_2, pp44[54]);
    wire[0:0] s1930, in1930_1, in1930_2;
    wire c1930;
    assign in1930_1 = {pp48[50]};
    assign in1930_2 = {pp49[49]};
    Full_Adder FA_1930(s1930, c1930, in1930_1, in1930_2, pp47[51]);
    wire[0:0] s1931, in1931_1, in1931_2;
    wire c1931;
    assign in1931_1 = {pp51[47]};
    assign in1931_2 = {pp52[46]};
    Full_Adder FA_1931(s1931, c1931, in1931_1, in1931_2, pp50[48]);
    wire[0:0] s1932, in1932_1, in1932_2;
    wire c1932;
    assign in1932_1 = {pp54[44]};
    assign in1932_2 = {pp55[43]};
    Full_Adder FA_1932(s1932, c1932, in1932_1, in1932_2, pp53[45]);
    wire[0:0] s1933, in1933_1, in1933_2;
    wire c1933;
    assign in1933_1 = {pp57[41]};
    assign in1933_2 = {pp58[40]};
    Full_Adder FA_1933(s1933, c1933, in1933_1, in1933_2, pp56[42]);
    wire[0:0] s1934, in1934_1, in1934_2;
    wire c1934;
    assign in1934_1 = {pp60[38]};
    assign in1934_2 = {pp61[37]};
    Full_Adder FA_1934(s1934, c1934, in1934_1, in1934_2, pp59[39]);
    wire[0:0] s1935, in1935_1, in1935_2;
    wire c1935;
    assign in1935_1 = {pp63[35]};
    assign in1935_2 = {c1258};
    Full_Adder FA_1935(s1935, c1935, in1935_1, in1935_2, pp62[36]);
    wire[0:0] s1936, in1936_1, in1936_2;
    wire c1936;
    assign in1936_1 = {pp37[62]};
    assign in1936_2 = {pp38[61]};
    Full_Adder FA_1936(s1936, c1936, in1936_1, in1936_2, pp36[63]);
    wire[0:0] s1937, in1937_1, in1937_2;
    wire c1937;
    assign in1937_1 = {pp40[59]};
    assign in1937_2 = {pp41[58]};
    Full_Adder FA_1937(s1937, c1937, in1937_1, in1937_2, pp39[60]);
    wire[0:0] s1938, in1938_1, in1938_2;
    wire c1938;
    assign in1938_1 = {pp43[56]};
    assign in1938_2 = {pp44[55]};
    Full_Adder FA_1938(s1938, c1938, in1938_1, in1938_2, pp42[57]);
    wire[0:0] s1939, in1939_1, in1939_2;
    wire c1939;
    assign in1939_1 = {pp46[53]};
    assign in1939_2 = {pp47[52]};
    Full_Adder FA_1939(s1939, c1939, in1939_1, in1939_2, pp45[54]);
    wire[0:0] s1940, in1940_1, in1940_2;
    wire c1940;
    assign in1940_1 = {pp49[50]};
    assign in1940_2 = {pp50[49]};
    Full_Adder FA_1940(s1940, c1940, in1940_1, in1940_2, pp48[51]);
    wire[0:0] s1941, in1941_1, in1941_2;
    wire c1941;
    assign in1941_1 = {pp52[47]};
    assign in1941_2 = {pp53[46]};
    Full_Adder FA_1941(s1941, c1941, in1941_1, in1941_2, pp51[48]);
    wire[0:0] s1942, in1942_1, in1942_2;
    wire c1942;
    assign in1942_1 = {pp55[44]};
    assign in1942_2 = {pp56[43]};
    Full_Adder FA_1942(s1942, c1942, in1942_1, in1942_2, pp54[45]);
    wire[0:0] s1943, in1943_1, in1943_2;
    wire c1943;
    assign in1943_1 = {pp58[41]};
    assign in1943_2 = {pp59[40]};
    Full_Adder FA_1943(s1943, c1943, in1943_1, in1943_2, pp57[42]);
    wire[0:0] s1944, in1944_1, in1944_2;
    wire c1944;
    assign in1944_1 = {pp61[38]};
    assign in1944_2 = {pp62[37]};
    Full_Adder FA_1944(s1944, c1944, in1944_1, in1944_2, pp60[39]);
    wire[0:0] s1945, in1945_1, in1945_2;
    wire c1945;
    assign in1945_1 = {pp38[62]};
    assign in1945_2 = {pp39[61]};
    Full_Adder FA_1945(s1945, c1945, in1945_1, in1945_2, pp37[63]);
    wire[0:0] s1946, in1946_1, in1946_2;
    wire c1946;
    assign in1946_1 = {pp41[59]};
    assign in1946_2 = {pp42[58]};
    Full_Adder FA_1946(s1946, c1946, in1946_1, in1946_2, pp40[60]);
    wire[0:0] s1947, in1947_1, in1947_2;
    wire c1947;
    assign in1947_1 = {pp44[56]};
    assign in1947_2 = {pp45[55]};
    Full_Adder FA_1947(s1947, c1947, in1947_1, in1947_2, pp43[57]);
    wire[0:0] s1948, in1948_1, in1948_2;
    wire c1948;
    assign in1948_1 = {pp47[53]};
    assign in1948_2 = {pp48[52]};
    Full_Adder FA_1948(s1948, c1948, in1948_1, in1948_2, pp46[54]);
    wire[0:0] s1949, in1949_1, in1949_2;
    wire c1949;
    assign in1949_1 = {pp50[50]};
    assign in1949_2 = {pp51[49]};
    Full_Adder FA_1949(s1949, c1949, in1949_1, in1949_2, pp49[51]);
    wire[0:0] s1950, in1950_1, in1950_2;
    wire c1950;
    assign in1950_1 = {pp53[47]};
    assign in1950_2 = {pp54[46]};
    Full_Adder FA_1950(s1950, c1950, in1950_1, in1950_2, pp52[48]);
    wire[0:0] s1951, in1951_1, in1951_2;
    wire c1951;
    assign in1951_1 = {pp56[44]};
    assign in1951_2 = {pp57[43]};
    Full_Adder FA_1951(s1951, c1951, in1951_1, in1951_2, pp55[45]);
    wire[0:0] s1952, in1952_1, in1952_2;
    wire c1952;
    assign in1952_1 = {pp59[41]};
    assign in1952_2 = {pp60[40]};
    Full_Adder FA_1952(s1952, c1952, in1952_1, in1952_2, pp58[42]);
    wire[0:0] s1953, in1953_1, in1953_2;
    wire c1953;
    assign in1953_1 = {pp39[62]};
    assign in1953_2 = {pp40[61]};
    Full_Adder FA_1953(s1953, c1953, in1953_1, in1953_2, pp38[63]);
    wire[0:0] s1954, in1954_1, in1954_2;
    wire c1954;
    assign in1954_1 = {pp42[59]};
    assign in1954_2 = {pp43[58]};
    Full_Adder FA_1954(s1954, c1954, in1954_1, in1954_2, pp41[60]);
    wire[0:0] s1955, in1955_1, in1955_2;
    wire c1955;
    assign in1955_1 = {pp45[56]};
    assign in1955_2 = {pp46[55]};
    Full_Adder FA_1955(s1955, c1955, in1955_1, in1955_2, pp44[57]);
    wire[0:0] s1956, in1956_1, in1956_2;
    wire c1956;
    assign in1956_1 = {pp48[53]};
    assign in1956_2 = {pp49[52]};
    Full_Adder FA_1956(s1956, c1956, in1956_1, in1956_2, pp47[54]);
    wire[0:0] s1957, in1957_1, in1957_2;
    wire c1957;
    assign in1957_1 = {pp51[50]};
    assign in1957_2 = {pp52[49]};
    Full_Adder FA_1957(s1957, c1957, in1957_1, in1957_2, pp50[51]);
    wire[0:0] s1958, in1958_1, in1958_2;
    wire c1958;
    assign in1958_1 = {pp54[47]};
    assign in1958_2 = {pp55[46]};
    Full_Adder FA_1958(s1958, c1958, in1958_1, in1958_2, pp53[48]);
    wire[0:0] s1959, in1959_1, in1959_2;
    wire c1959;
    assign in1959_1 = {pp57[44]};
    assign in1959_2 = {pp58[43]};
    Full_Adder FA_1959(s1959, c1959, in1959_1, in1959_2, pp56[45]);
    wire[0:0] s1960, in1960_1, in1960_2;
    wire c1960;
    assign in1960_1 = {pp40[62]};
    assign in1960_2 = {pp41[61]};
    Full_Adder FA_1960(s1960, c1960, in1960_1, in1960_2, pp39[63]);
    wire[0:0] s1961, in1961_1, in1961_2;
    wire c1961;
    assign in1961_1 = {pp43[59]};
    assign in1961_2 = {pp44[58]};
    Full_Adder FA_1961(s1961, c1961, in1961_1, in1961_2, pp42[60]);
    wire[0:0] s1962, in1962_1, in1962_2;
    wire c1962;
    assign in1962_1 = {pp46[56]};
    assign in1962_2 = {pp47[55]};
    Full_Adder FA_1962(s1962, c1962, in1962_1, in1962_2, pp45[57]);
    wire[0:0] s1963, in1963_1, in1963_2;
    wire c1963;
    assign in1963_1 = {pp49[53]};
    assign in1963_2 = {pp50[52]};
    Full_Adder FA_1963(s1963, c1963, in1963_1, in1963_2, pp48[54]);
    wire[0:0] s1964, in1964_1, in1964_2;
    wire c1964;
    assign in1964_1 = {pp52[50]};
    assign in1964_2 = {pp53[49]};
    Full_Adder FA_1964(s1964, c1964, in1964_1, in1964_2, pp51[51]);
    wire[0:0] s1965, in1965_1, in1965_2;
    wire c1965;
    assign in1965_1 = {pp55[47]};
    assign in1965_2 = {pp56[46]};
    Full_Adder FA_1965(s1965, c1965, in1965_1, in1965_2, pp54[48]);
    wire[0:0] s1966, in1966_1, in1966_2;
    wire c1966;
    assign in1966_1 = {pp41[62]};
    assign in1966_2 = {pp42[61]};
    Full_Adder FA_1966(s1966, c1966, in1966_1, in1966_2, pp40[63]);
    wire[0:0] s1967, in1967_1, in1967_2;
    wire c1967;
    assign in1967_1 = {pp44[59]};
    assign in1967_2 = {pp45[58]};
    Full_Adder FA_1967(s1967, c1967, in1967_1, in1967_2, pp43[60]);
    wire[0:0] s1968, in1968_1, in1968_2;
    wire c1968;
    assign in1968_1 = {pp47[56]};
    assign in1968_2 = {pp48[55]};
    Full_Adder FA_1968(s1968, c1968, in1968_1, in1968_2, pp46[57]);
    wire[0:0] s1969, in1969_1, in1969_2;
    wire c1969;
    assign in1969_1 = {pp50[53]};
    assign in1969_2 = {pp51[52]};
    Full_Adder FA_1969(s1969, c1969, in1969_1, in1969_2, pp49[54]);
    wire[0:0] s1970, in1970_1, in1970_2;
    wire c1970;
    assign in1970_1 = {pp53[50]};
    assign in1970_2 = {pp54[49]};
    Full_Adder FA_1970(s1970, c1970, in1970_1, in1970_2, pp52[51]);
    wire[0:0] s1971, in1971_1, in1971_2;
    wire c1971;
    assign in1971_1 = {pp42[62]};
    assign in1971_2 = {pp43[61]};
    Full_Adder FA_1971(s1971, c1971, in1971_1, in1971_2, pp41[63]);
    wire[0:0] s1972, in1972_1, in1972_2;
    wire c1972;
    assign in1972_1 = {pp45[59]};
    assign in1972_2 = {pp46[58]};
    Full_Adder FA_1972(s1972, c1972, in1972_1, in1972_2, pp44[60]);
    wire[0:0] s1973, in1973_1, in1973_2;
    wire c1973;
    assign in1973_1 = {pp48[56]};
    assign in1973_2 = {pp49[55]};
    Full_Adder FA_1973(s1973, c1973, in1973_1, in1973_2, pp47[57]);
    wire[0:0] s1974, in1974_1, in1974_2;
    wire c1974;
    assign in1974_1 = {pp51[53]};
    assign in1974_2 = {pp52[52]};
    Full_Adder FA_1974(s1974, c1974, in1974_1, in1974_2, pp50[54]);
    wire[0:0] s1975, in1975_1, in1975_2;
    wire c1975;
    assign in1975_1 = {pp43[62]};
    assign in1975_2 = {pp44[61]};
    Full_Adder FA_1975(s1975, c1975, in1975_1, in1975_2, pp42[63]);
    wire[0:0] s1976, in1976_1, in1976_2;
    wire c1976;
    assign in1976_1 = {pp46[59]};
    assign in1976_2 = {pp47[58]};
    Full_Adder FA_1976(s1976, c1976, in1976_1, in1976_2, pp45[60]);
    wire[0:0] s1977, in1977_1, in1977_2;
    wire c1977;
    assign in1977_1 = {pp49[56]};
    assign in1977_2 = {pp50[55]};
    Full_Adder FA_1977(s1977, c1977, in1977_1, in1977_2, pp48[57]);
    wire[0:0] s1978, in1978_1, in1978_2;
    wire c1978;
    assign in1978_1 = {pp44[62]};
    assign in1978_2 = {pp45[61]};
    Full_Adder FA_1978(s1978, c1978, in1978_1, in1978_2, pp43[63]);
    wire[0:0] s1979, in1979_1, in1979_2;
    wire c1979;
    assign in1979_1 = {pp47[59]};
    assign in1979_2 = {pp48[58]};
    Full_Adder FA_1979(s1979, c1979, in1979_1, in1979_2, pp46[60]);
    wire[0:0] s1980, in1980_1, in1980_2;
    wire c1980;
    assign in1980_1 = {pp45[62]};
    assign in1980_2 = {pp46[61]};
    Full_Adder FA_1980(s1980, c1980, in1980_1, in1980_2, pp44[63]);

    /*Stage 4*/
    wire[0:0] s1981, in1981_1, in1981_2;
    wire c1981;
    assign in1981_1 = {pp0[14]};
    assign in1981_2 = {pp1[13]};
    Half_Adder HA_1981(s1981, c1981, in1981_1, in1981_2);
    wire[0:0] s1982, in1982_1, in1982_2;
    wire c1982;
    assign in1982_1 = {pp1[14]};
    assign in1982_2 = {pp2[13]};
    Full_Adder FA_1982(s1982, c1982, in1982_1, in1982_2, pp0[15]);
    wire[0:0] s1983, in1983_1, in1983_2;
    wire c1983;
    assign in1983_1 = {pp3[12]};
    assign in1983_2 = {pp4[11]};
    Half_Adder HA_1983(s1983, c1983, in1983_1, in1983_2);
    wire[0:0] s1984, in1984_1, in1984_2;
    wire c1984;
    assign in1984_1 = {pp1[15]};
    assign in1984_2 = {pp2[14]};
    Full_Adder FA_1984(s1984, c1984, in1984_1, in1984_2, pp0[16]);
    wire[0:0] s1985, in1985_1, in1985_2;
    wire c1985;
    assign in1985_1 = {pp4[12]};
    assign in1985_2 = {pp5[11]};
    Full_Adder FA_1985(s1985, c1985, in1985_1, in1985_2, pp3[13]);
    wire[0:0] s1986, in1986_1, in1986_2;
    wire c1986;
    assign in1986_1 = {pp6[10]};
    assign in1986_2 = {pp7[9]};
    Half_Adder HA_1986(s1986, c1986, in1986_1, in1986_2);
    wire[0:0] s1987, in1987_1, in1987_2;
    wire c1987;
    assign in1987_1 = {pp1[16]};
    assign in1987_2 = {pp2[15]};
    Full_Adder FA_1987(s1987, c1987, in1987_1, in1987_2, pp0[17]);
    wire[0:0] s1988, in1988_1, in1988_2;
    wire c1988;
    assign in1988_1 = {pp4[13]};
    assign in1988_2 = {pp5[12]};
    Full_Adder FA_1988(s1988, c1988, in1988_1, in1988_2, pp3[14]);
    wire[0:0] s1989, in1989_1, in1989_2;
    wire c1989;
    assign in1989_1 = {pp7[10]};
    assign in1989_2 = {pp8[9]};
    Full_Adder FA_1989(s1989, c1989, in1989_1, in1989_2, pp6[11]);
    wire[0:0] s1990, in1990_1, in1990_2;
    wire c1990;
    assign in1990_1 = {pp9[8]};
    assign in1990_2 = {pp10[7]};
    Half_Adder HA_1990(s1990, c1990, in1990_1, in1990_2);
    wire[0:0] s1991, in1991_1, in1991_2;
    wire c1991;
    assign in1991_1 = {pp1[17]};
    assign in1991_2 = {pp2[16]};
    Full_Adder FA_1991(s1991, c1991, in1991_1, in1991_2, pp0[18]);
    wire[0:0] s1992, in1992_1, in1992_2;
    wire c1992;
    assign in1992_1 = {pp4[14]};
    assign in1992_2 = {pp5[13]};
    Full_Adder FA_1992(s1992, c1992, in1992_1, in1992_2, pp3[15]);
    wire[0:0] s1993, in1993_1, in1993_2;
    wire c1993;
    assign in1993_1 = {pp7[11]};
    assign in1993_2 = {pp8[10]};
    Full_Adder FA_1993(s1993, c1993, in1993_1, in1993_2, pp6[12]);
    wire[0:0] s1994, in1994_1, in1994_2;
    wire c1994;
    assign in1994_1 = {pp10[8]};
    assign in1994_2 = {pp11[7]};
    Full_Adder FA_1994(s1994, c1994, in1994_1, in1994_2, pp9[9]);
    wire[0:0] s1995, in1995_1, in1995_2;
    wire c1995;
    assign in1995_1 = {pp12[6]};
    assign in1995_2 = {pp13[5]};
    Half_Adder HA_1995(s1995, c1995, in1995_1, in1995_2);
    wire[0:0] s1996, in1996_1, in1996_2;
    wire c1996;
    assign in1996_1 = {pp1[18]};
    assign in1996_2 = {pp2[17]};
    Full_Adder FA_1996(s1996, c1996, in1996_1, in1996_2, pp0[19]);
    wire[0:0] s1997, in1997_1, in1997_2;
    wire c1997;
    assign in1997_1 = {pp4[15]};
    assign in1997_2 = {pp5[14]};
    Full_Adder FA_1997(s1997, c1997, in1997_1, in1997_2, pp3[16]);
    wire[0:0] s1998, in1998_1, in1998_2;
    wire c1998;
    assign in1998_1 = {pp7[12]};
    assign in1998_2 = {pp8[11]};
    Full_Adder FA_1998(s1998, c1998, in1998_1, in1998_2, pp6[13]);
    wire[0:0] s1999, in1999_1, in1999_2;
    wire c1999;
    assign in1999_1 = {pp10[9]};
    assign in1999_2 = {pp11[8]};
    Full_Adder FA_1999(s1999, c1999, in1999_1, in1999_2, pp9[10]);
    wire[0:0] s2000, in2000_1, in2000_2;
    wire c2000;
    assign in2000_1 = {pp13[6]};
    assign in2000_2 = {pp14[5]};
    Full_Adder FA_2000(s2000, c2000, in2000_1, in2000_2, pp12[7]);
    wire[0:0] s2001, in2001_1, in2001_2;
    wire c2001;
    assign in2001_1 = {pp15[4]};
    assign in2001_2 = {pp16[3]};
    Half_Adder HA_2001(s2001, c2001, in2001_1, in2001_2);
    wire[0:0] s2002, in2002_1, in2002_2;
    wire c2002;
    assign in2002_1 = {pp3[17]};
    assign in2002_2 = {pp4[16]};
    Full_Adder FA_2002(s2002, c2002, in2002_1, in2002_2, pp2[18]);
    wire[0:0] s2003, in2003_1, in2003_2;
    wire c2003;
    assign in2003_1 = {pp6[14]};
    assign in2003_2 = {pp7[13]};
    Full_Adder FA_2003(s2003, c2003, in2003_1, in2003_2, pp5[15]);
    wire[0:0] s2004, in2004_1, in2004_2;
    wire c2004;
    assign in2004_1 = {pp9[11]};
    assign in2004_2 = {pp10[10]};
    Full_Adder FA_2004(s2004, c2004, in2004_1, in2004_2, pp8[12]);
    wire[0:0] s2005, in2005_1, in2005_2;
    wire c2005;
    assign in2005_1 = {pp12[8]};
    assign in2005_2 = {pp13[7]};
    Full_Adder FA_2005(s2005, c2005, in2005_1, in2005_2, pp11[9]);
    wire[0:0] s2006, in2006_1, in2006_2;
    wire c2006;
    assign in2006_1 = {pp15[5]};
    assign in2006_2 = {pp16[4]};
    Full_Adder FA_2006(s2006, c2006, in2006_1, in2006_2, pp14[6]);
    wire[0:0] s2007, in2007_1, in2007_2;
    wire c2007;
    assign in2007_1 = {pp18[2]};
    assign in2007_2 = {pp19[1]};
    Full_Adder FA_2007(s2007, c2007, in2007_1, in2007_2, pp17[3]);
    wire[0:0] s2008, in2008_1, in2008_2;
    wire c2008;
    assign in2008_1 = {pp6[15]};
    assign in2008_2 = {pp7[14]};
    Full_Adder FA_2008(s2008, c2008, in2008_1, in2008_2, pp5[16]);
    wire[0:0] s2009, in2009_1, in2009_2;
    wire c2009;
    assign in2009_1 = {pp9[12]};
    assign in2009_2 = {pp10[11]};
    Full_Adder FA_2009(s2009, c2009, in2009_1, in2009_2, pp8[13]);
    wire[0:0] s2010, in2010_1, in2010_2;
    wire c2010;
    assign in2010_1 = {pp12[9]};
    assign in2010_2 = {pp13[8]};
    Full_Adder FA_2010(s2010, c2010, in2010_1, in2010_2, pp11[10]);
    wire[0:0] s2011, in2011_1, in2011_2;
    wire c2011;
    assign in2011_1 = {pp15[6]};
    assign in2011_2 = {pp16[5]};
    Full_Adder FA_2011(s2011, c2011, in2011_1, in2011_2, pp14[7]);
    wire[0:0] s2012, in2012_1, in2012_2;
    wire c2012;
    assign in2012_1 = {pp18[3]};
    assign in2012_2 = {pp19[2]};
    Full_Adder FA_2012(s2012, c2012, in2012_1, in2012_2, pp17[4]);
    wire[0:0] s2013, in2013_1, in2013_2;
    wire c2013;
    assign in2013_1 = {pp21[0]};
    assign in2013_2 = {c1261};
    Full_Adder FA_2013(s2013, c2013, in2013_1, in2013_2, pp20[1]);
    wire[0:0] s2014, in2014_1, in2014_2;
    wire c2014;
    assign in2014_1 = {pp9[13]};
    assign in2014_2 = {pp10[12]};
    Full_Adder FA_2014(s2014, c2014, in2014_1, in2014_2, pp8[14]);
    wire[0:0] s2015, in2015_1, in2015_2;
    wire c2015;
    assign in2015_1 = {pp12[10]};
    assign in2015_2 = {pp13[9]};
    Full_Adder FA_2015(s2015, c2015, in2015_1, in2015_2, pp11[11]);
    wire[0:0] s2016, in2016_1, in2016_2;
    wire c2016;
    assign in2016_1 = {pp15[7]};
    assign in2016_2 = {pp16[6]};
    Full_Adder FA_2016(s2016, c2016, in2016_1, in2016_2, pp14[8]);
    wire[0:0] s2017, in2017_1, in2017_2;
    wire c2017;
    assign in2017_1 = {pp18[4]};
    assign in2017_2 = {pp19[3]};
    Full_Adder FA_2017(s2017, c2017, in2017_1, in2017_2, pp17[5]);
    wire[0:0] s2018, in2018_1, in2018_2;
    wire c2018;
    assign in2018_1 = {pp21[1]};
    assign in2018_2 = {pp22[0]};
    Full_Adder FA_2018(s2018, c2018, in2018_1, in2018_2, pp20[2]);
    wire[0:0] s2019, in2019_1, in2019_2;
    wire c2019;
    assign in2019_1 = {c1263};
    assign in2019_2 = {s1264[0]};
    Full_Adder FA_2019(s2019, c2019, in2019_1, in2019_2, c1262);
    wire[0:0] s2020, in2020_1, in2020_2;
    wire c2020;
    assign in2020_1 = {pp12[11]};
    assign in2020_2 = {pp13[10]};
    Full_Adder FA_2020(s2020, c2020, in2020_1, in2020_2, pp11[12]);
    wire[0:0] s2021, in2021_1, in2021_2;
    wire c2021;
    assign in2021_1 = {pp15[8]};
    assign in2021_2 = {pp16[7]};
    Full_Adder FA_2021(s2021, c2021, in2021_1, in2021_2, pp14[9]);
    wire[0:0] s2022, in2022_1, in2022_2;
    wire c2022;
    assign in2022_1 = {pp18[5]};
    assign in2022_2 = {pp19[4]};
    Full_Adder FA_2022(s2022, c2022, in2022_1, in2022_2, pp17[6]);
    wire[0:0] s2023, in2023_1, in2023_2;
    wire c2023;
    assign in2023_1 = {pp21[2]};
    assign in2023_2 = {pp22[1]};
    Full_Adder FA_2023(s2023, c2023, in2023_1, in2023_2, pp20[3]);
    wire[0:0] s2024, in2024_1, in2024_2;
    wire c2024;
    assign in2024_1 = {c1264};
    assign in2024_2 = {c1265};
    Full_Adder FA_2024(s2024, c2024, in2024_1, in2024_2, pp23[0]);
    wire[0:0] s2025, in2025_1, in2025_2;
    wire c2025;
    assign in2025_1 = {s1267[0]};
    assign in2025_2 = {s1268[0]};
    Full_Adder FA_2025(s2025, c2025, in2025_1, in2025_2, c1266);
    wire[0:0] s2026, in2026_1, in2026_2;
    wire c2026;
    assign in2026_1 = {pp15[9]};
    assign in2026_2 = {pp16[8]};
    Full_Adder FA_2026(s2026, c2026, in2026_1, in2026_2, pp14[10]);
    wire[0:0] s2027, in2027_1, in2027_2;
    wire c2027;
    assign in2027_1 = {pp18[6]};
    assign in2027_2 = {pp19[5]};
    Full_Adder FA_2027(s2027, c2027, in2027_1, in2027_2, pp17[7]);
    wire[0:0] s2028, in2028_1, in2028_2;
    wire c2028;
    assign in2028_1 = {pp21[3]};
    assign in2028_2 = {pp22[2]};
    Full_Adder FA_2028(s2028, c2028, in2028_1, in2028_2, pp20[4]);
    wire[0:0] s2029, in2029_1, in2029_2;
    wire c2029;
    assign in2029_1 = {pp24[0]};
    assign in2029_2 = {c1267};
    Full_Adder FA_2029(s2029, c2029, in2029_1, in2029_2, pp23[1]);
    wire[0:0] s2030, in2030_1, in2030_2;
    wire c2030;
    assign in2030_1 = {c1269};
    assign in2030_2 = {c1270};
    Full_Adder FA_2030(s2030, c2030, in2030_1, in2030_2, c1268);
    wire[0:0] s2031, in2031_1, in2031_2;
    wire c2031;
    assign in2031_1 = {s1272[0]};
    assign in2031_2 = {s1273[0]};
    Full_Adder FA_2031(s2031, c2031, in2031_1, in2031_2, s1271[0]);
    wire[0:0] s2032, in2032_1, in2032_2;
    wire c2032;
    assign in2032_1 = {pp18[7]};
    assign in2032_2 = {pp19[6]};
    Full_Adder FA_2032(s2032, c2032, in2032_1, in2032_2, pp17[8]);
    wire[0:0] s2033, in2033_1, in2033_2;
    wire c2033;
    assign in2033_1 = {pp21[4]};
    assign in2033_2 = {pp22[3]};
    Full_Adder FA_2033(s2033, c2033, in2033_1, in2033_2, pp20[5]);
    wire[0:0] s2034, in2034_1, in2034_2;
    wire c2034;
    assign in2034_1 = {pp24[1]};
    assign in2034_2 = {pp25[0]};
    Full_Adder FA_2034(s2034, c2034, in2034_1, in2034_2, pp23[2]);
    wire[0:0] s2035, in2035_1, in2035_2;
    wire c2035;
    assign in2035_1 = {c1272};
    assign in2035_2 = {c1273};
    Full_Adder FA_2035(s2035, c2035, in2035_1, in2035_2, c1271);
    wire[0:0] s2036, in2036_1, in2036_2;
    wire c2036;
    assign in2036_1 = {c1275};
    assign in2036_2 = {s1276[0]};
    Full_Adder FA_2036(s2036, c2036, in2036_1, in2036_2, c1274);
    wire[0:0] s2037, in2037_1, in2037_2;
    wire c2037;
    assign in2037_1 = {s1278[0]};
    assign in2037_2 = {s1279[0]};
    Full_Adder FA_2037(s2037, c2037, in2037_1, in2037_2, s1277[0]);
    wire[0:0] s2038, in2038_1, in2038_2;
    wire c2038;
    assign in2038_1 = {pp21[5]};
    assign in2038_2 = {pp22[4]};
    Full_Adder FA_2038(s2038, c2038, in2038_1, in2038_2, pp20[6]);
    wire[0:0] s2039, in2039_1, in2039_2;
    wire c2039;
    assign in2039_1 = {pp24[2]};
    assign in2039_2 = {pp25[1]};
    Full_Adder FA_2039(s2039, c2039, in2039_1, in2039_2, pp23[3]);
    wire[0:0] s2040, in2040_1, in2040_2;
    wire c2040;
    assign in2040_1 = {c1276};
    assign in2040_2 = {c1277};
    Full_Adder FA_2040(s2040, c2040, in2040_1, in2040_2, pp26[0]);
    wire[0:0] s2041, in2041_1, in2041_2;
    wire c2041;
    assign in2041_1 = {c1279};
    assign in2041_2 = {c1280};
    Full_Adder FA_2041(s2041, c2041, in2041_1, in2041_2, c1278);
    wire[0:0] s2042, in2042_1, in2042_2;
    wire c2042;
    assign in2042_1 = {s1282[0]};
    assign in2042_2 = {s1283[0]};
    Full_Adder FA_2042(s2042, c2042, in2042_1, in2042_2, c1281);
    wire[0:0] s2043, in2043_1, in2043_2;
    wire c2043;
    assign in2043_1 = {s1285[0]};
    assign in2043_2 = {s1286[0]};
    Full_Adder FA_2043(s2043, c2043, in2043_1, in2043_2, s1284[0]);
    wire[0:0] s2044, in2044_1, in2044_2;
    wire c2044;
    assign in2044_1 = {pp24[3]};
    assign in2044_2 = {pp25[2]};
    Full_Adder FA_2044(s2044, c2044, in2044_1, in2044_2, pp23[4]);
    wire[0:0] s2045, in2045_1, in2045_2;
    wire c2045;
    assign in2045_1 = {pp27[0]};
    assign in2045_2 = {c1282};
    Full_Adder FA_2045(s2045, c2045, in2045_1, in2045_2, pp26[1]);
    wire[0:0] s2046, in2046_1, in2046_2;
    wire c2046;
    assign in2046_1 = {c1284};
    assign in2046_2 = {c1285};
    Full_Adder FA_2046(s2046, c2046, in2046_1, in2046_2, c1283);
    wire[0:0] s2047, in2047_1, in2047_2;
    wire c2047;
    assign in2047_1 = {c1287};
    assign in2047_2 = {c1288};
    Full_Adder FA_2047(s2047, c2047, in2047_1, in2047_2, c1286);
    wire[0:0] s2048, in2048_1, in2048_2;
    wire c2048;
    assign in2048_1 = {s1290[0]};
    assign in2048_2 = {s1291[0]};
    Full_Adder FA_2048(s2048, c2048, in2048_1, in2048_2, s1289[0]);
    wire[0:0] s2049, in2049_1, in2049_2;
    wire c2049;
    assign in2049_1 = {s1293[0]};
    assign in2049_2 = {s1294[0]};
    Full_Adder FA_2049(s2049, c2049, in2049_1, in2049_2, s1292[0]);
    wire[0:0] s2050, in2050_1, in2050_2;
    wire c2050;
    assign in2050_1 = {pp27[1]};
    assign in2050_2 = {pp28[0]};
    Full_Adder FA_2050(s2050, c2050, in2050_1, in2050_2, pp26[2]);
    wire[0:0] s2051, in2051_1, in2051_2;
    wire c2051;
    assign in2051_1 = {c1290};
    assign in2051_2 = {c1291};
    Full_Adder FA_2051(s2051, c2051, in2051_1, in2051_2, c1289);
    wire[0:0] s2052, in2052_1, in2052_2;
    wire c2052;
    assign in2052_1 = {c1293};
    assign in2052_2 = {c1294};
    Full_Adder FA_2052(s2052, c2052, in2052_1, in2052_2, c1292);
    wire[0:0] s2053, in2053_1, in2053_2;
    wire c2053;
    assign in2053_1 = {c1296};
    assign in2053_2 = {s1297[0]};
    Full_Adder FA_2053(s2053, c2053, in2053_1, in2053_2, c1295);
    wire[0:0] s2054, in2054_1, in2054_2;
    wire c2054;
    assign in2054_1 = {s1299[0]};
    assign in2054_2 = {s1300[0]};
    Full_Adder FA_2054(s2054, c2054, in2054_1, in2054_2, s1298[0]);
    wire[0:0] s2055, in2055_1, in2055_2;
    wire c2055;
    assign in2055_1 = {s1302[0]};
    assign in2055_2 = {s1303[0]};
    Full_Adder FA_2055(s2055, c2055, in2055_1, in2055_2, s1301[0]);
    wire[0:0] s2056, in2056_1, in2056_2;
    wire c2056;
    assign in2056_1 = {s463[0]};
    assign in2056_2 = {c1297};
    Full_Adder FA_2056(s2056, c2056, in2056_1, in2056_2, pp29[0]);
    wire[0:0] s2057, in2057_1, in2057_2;
    wire c2057;
    assign in2057_1 = {c1299};
    assign in2057_2 = {c1300};
    Full_Adder FA_2057(s2057, c2057, in2057_1, in2057_2, c1298);
    wire[0:0] s2058, in2058_1, in2058_2;
    wire c2058;
    assign in2058_1 = {c1302};
    assign in2058_2 = {c1303};
    Full_Adder FA_2058(s2058, c2058, in2058_1, in2058_2, c1301);
    wire[0:0] s2059, in2059_1, in2059_2;
    wire c2059;
    assign in2059_1 = {c1305};
    assign in2059_2 = {s1306[0]};
    Full_Adder FA_2059(s2059, c2059, in2059_1, in2059_2, c1304);
    wire[0:0] s2060, in2060_1, in2060_2;
    wire c2060;
    assign in2060_1 = {s1308[0]};
    assign in2060_2 = {s1309[0]};
    Full_Adder FA_2060(s2060, c2060, in2060_1, in2060_2, s1307[0]);
    wire[0:0] s2061, in2061_1, in2061_2;
    wire c2061;
    assign in2061_1 = {s1311[0]};
    assign in2061_2 = {s1312[0]};
    Full_Adder FA_2061(s2061, c2061, in2061_1, in2061_2, s1310[0]);
    wire[0:0] s2062, in2062_1, in2062_2;
    wire c2062;
    assign in2062_1 = {s465[0]};
    assign in2062_2 = {c1306};
    Full_Adder FA_2062(s2062, c2062, in2062_1, in2062_2, s464[0]);
    wire[0:0] s2063, in2063_1, in2063_2;
    wire c2063;
    assign in2063_1 = {c1308};
    assign in2063_2 = {c1309};
    Full_Adder FA_2063(s2063, c2063, in2063_1, in2063_2, c1307);
    wire[0:0] s2064, in2064_1, in2064_2;
    wire c2064;
    assign in2064_1 = {c1311};
    assign in2064_2 = {c1312};
    Full_Adder FA_2064(s2064, c2064, in2064_1, in2064_2, c1310);
    wire[0:0] s2065, in2065_1, in2065_2;
    wire c2065;
    assign in2065_1 = {c1314};
    assign in2065_2 = {s1315[0]};
    Full_Adder FA_2065(s2065, c2065, in2065_1, in2065_2, c1313);
    wire[0:0] s2066, in2066_1, in2066_2;
    wire c2066;
    assign in2066_1 = {s1317[0]};
    assign in2066_2 = {s1318[0]};
    Full_Adder FA_2066(s2066, c2066, in2066_1, in2066_2, s1316[0]);
    wire[0:0] s2067, in2067_1, in2067_2;
    wire c2067;
    assign in2067_1 = {s1320[0]};
    assign in2067_2 = {s1321[0]};
    Full_Adder FA_2067(s2067, c2067, in2067_1, in2067_2, s1319[0]);
    wire[0:0] s2068, in2068_1, in2068_2;
    wire c2068;
    assign in2068_1 = {s468[0]};
    assign in2068_2 = {c1315};
    Full_Adder FA_2068(s2068, c2068, in2068_1, in2068_2, s467[0]);
    wire[0:0] s2069, in2069_1, in2069_2;
    wire c2069;
    assign in2069_1 = {c1317};
    assign in2069_2 = {c1318};
    Full_Adder FA_2069(s2069, c2069, in2069_1, in2069_2, c1316);
    wire[0:0] s2070, in2070_1, in2070_2;
    wire c2070;
    assign in2070_1 = {c1320};
    assign in2070_2 = {c1321};
    Full_Adder FA_2070(s2070, c2070, in2070_1, in2070_2, c1319);
    wire[0:0] s2071, in2071_1, in2071_2;
    wire c2071;
    assign in2071_1 = {c1323};
    assign in2071_2 = {s1324[0]};
    Full_Adder FA_2071(s2071, c2071, in2071_1, in2071_2, c1322);
    wire[0:0] s2072, in2072_1, in2072_2;
    wire c2072;
    assign in2072_1 = {s1326[0]};
    assign in2072_2 = {s1327[0]};
    Full_Adder FA_2072(s2072, c2072, in2072_1, in2072_2, s1325[0]);
    wire[0:0] s2073, in2073_1, in2073_2;
    wire c2073;
    assign in2073_1 = {s1329[0]};
    assign in2073_2 = {s1330[0]};
    Full_Adder FA_2073(s2073, c2073, in2073_1, in2073_2, s1328[0]);
    wire[0:0] s2074, in2074_1, in2074_2;
    wire c2074;
    assign in2074_1 = {s472[0]};
    assign in2074_2 = {c1324};
    Full_Adder FA_2074(s2074, c2074, in2074_1, in2074_2, s471[0]);
    wire[0:0] s2075, in2075_1, in2075_2;
    wire c2075;
    assign in2075_1 = {c1326};
    assign in2075_2 = {c1327};
    Full_Adder FA_2075(s2075, c2075, in2075_1, in2075_2, c1325);
    wire[0:0] s2076, in2076_1, in2076_2;
    wire c2076;
    assign in2076_1 = {c1329};
    assign in2076_2 = {c1330};
    Full_Adder FA_2076(s2076, c2076, in2076_1, in2076_2, c1328);
    wire[0:0] s2077, in2077_1, in2077_2;
    wire c2077;
    assign in2077_1 = {c1332};
    assign in2077_2 = {s1333[0]};
    Full_Adder FA_2077(s2077, c2077, in2077_1, in2077_2, c1331);
    wire[0:0] s2078, in2078_1, in2078_2;
    wire c2078;
    assign in2078_1 = {s1335[0]};
    assign in2078_2 = {s1336[0]};
    Full_Adder FA_2078(s2078, c2078, in2078_1, in2078_2, s1334[0]);
    wire[0:0] s2079, in2079_1, in2079_2;
    wire c2079;
    assign in2079_1 = {s1338[0]};
    assign in2079_2 = {s1339[0]};
    Full_Adder FA_2079(s2079, c2079, in2079_1, in2079_2, s1337[0]);
    wire[0:0] s2080, in2080_1, in2080_2;
    wire c2080;
    assign in2080_1 = {s477[0]};
    assign in2080_2 = {c1333};
    Full_Adder FA_2080(s2080, c2080, in2080_1, in2080_2, s476[0]);
    wire[0:0] s2081, in2081_1, in2081_2;
    wire c2081;
    assign in2081_1 = {c1335};
    assign in2081_2 = {c1336};
    Full_Adder FA_2081(s2081, c2081, in2081_1, in2081_2, c1334);
    wire[0:0] s2082, in2082_1, in2082_2;
    wire c2082;
    assign in2082_1 = {c1338};
    assign in2082_2 = {c1339};
    Full_Adder FA_2082(s2082, c2082, in2082_1, in2082_2, c1337);
    wire[0:0] s2083, in2083_1, in2083_2;
    wire c2083;
    assign in2083_1 = {c1341};
    assign in2083_2 = {s1342[0]};
    Full_Adder FA_2083(s2083, c2083, in2083_1, in2083_2, c1340);
    wire[0:0] s2084, in2084_1, in2084_2;
    wire c2084;
    assign in2084_1 = {s1344[0]};
    assign in2084_2 = {s1345[0]};
    Full_Adder FA_2084(s2084, c2084, in2084_1, in2084_2, s1343[0]);
    wire[0:0] s2085, in2085_1, in2085_2;
    wire c2085;
    assign in2085_1 = {s1347[0]};
    assign in2085_2 = {s1348[0]};
    Full_Adder FA_2085(s2085, c2085, in2085_1, in2085_2, s1346[0]);
    wire[0:0] s2086, in2086_1, in2086_2;
    wire c2086;
    assign in2086_1 = {s483[0]};
    assign in2086_2 = {c1342};
    Full_Adder FA_2086(s2086, c2086, in2086_1, in2086_2, s482[0]);
    wire[0:0] s2087, in2087_1, in2087_2;
    wire c2087;
    assign in2087_1 = {c1344};
    assign in2087_2 = {c1345};
    Full_Adder FA_2087(s2087, c2087, in2087_1, in2087_2, c1343);
    wire[0:0] s2088, in2088_1, in2088_2;
    wire c2088;
    assign in2088_1 = {c1347};
    assign in2088_2 = {c1348};
    Full_Adder FA_2088(s2088, c2088, in2088_1, in2088_2, c1346);
    wire[0:0] s2089, in2089_1, in2089_2;
    wire c2089;
    assign in2089_1 = {c1350};
    assign in2089_2 = {s1351[0]};
    Full_Adder FA_2089(s2089, c2089, in2089_1, in2089_2, c1349);
    wire[0:0] s2090, in2090_1, in2090_2;
    wire c2090;
    assign in2090_1 = {s1353[0]};
    assign in2090_2 = {s1354[0]};
    Full_Adder FA_2090(s2090, c2090, in2090_1, in2090_2, s1352[0]);
    wire[0:0] s2091, in2091_1, in2091_2;
    wire c2091;
    assign in2091_1 = {s1356[0]};
    assign in2091_2 = {s1357[0]};
    Full_Adder FA_2091(s2091, c2091, in2091_1, in2091_2, s1355[0]);
    wire[0:0] s2092, in2092_1, in2092_2;
    wire c2092;
    assign in2092_1 = {s490[0]};
    assign in2092_2 = {c1351};
    Full_Adder FA_2092(s2092, c2092, in2092_1, in2092_2, s489[0]);
    wire[0:0] s2093, in2093_1, in2093_2;
    wire c2093;
    assign in2093_1 = {c1353};
    assign in2093_2 = {c1354};
    Full_Adder FA_2093(s2093, c2093, in2093_1, in2093_2, c1352);
    wire[0:0] s2094, in2094_1, in2094_2;
    wire c2094;
    assign in2094_1 = {c1356};
    assign in2094_2 = {c1357};
    Full_Adder FA_2094(s2094, c2094, in2094_1, in2094_2, c1355);
    wire[0:0] s2095, in2095_1, in2095_2;
    wire c2095;
    assign in2095_1 = {c1359};
    assign in2095_2 = {s1360[0]};
    Full_Adder FA_2095(s2095, c2095, in2095_1, in2095_2, c1358);
    wire[0:0] s2096, in2096_1, in2096_2;
    wire c2096;
    assign in2096_1 = {s1362[0]};
    assign in2096_2 = {s1363[0]};
    Full_Adder FA_2096(s2096, c2096, in2096_1, in2096_2, s1361[0]);
    wire[0:0] s2097, in2097_1, in2097_2;
    wire c2097;
    assign in2097_1 = {s1365[0]};
    assign in2097_2 = {s1366[0]};
    Full_Adder FA_2097(s2097, c2097, in2097_1, in2097_2, s1364[0]);
    wire[0:0] s2098, in2098_1, in2098_2;
    wire c2098;
    assign in2098_1 = {s498[0]};
    assign in2098_2 = {c1360};
    Full_Adder FA_2098(s2098, c2098, in2098_1, in2098_2, s497[0]);
    wire[0:0] s2099, in2099_1, in2099_2;
    wire c2099;
    assign in2099_1 = {c1362};
    assign in2099_2 = {c1363};
    Full_Adder FA_2099(s2099, c2099, in2099_1, in2099_2, c1361);
    wire[0:0] s2100, in2100_1, in2100_2;
    wire c2100;
    assign in2100_1 = {c1365};
    assign in2100_2 = {c1366};
    Full_Adder FA_2100(s2100, c2100, in2100_1, in2100_2, c1364);
    wire[0:0] s2101, in2101_1, in2101_2;
    wire c2101;
    assign in2101_1 = {c1368};
    assign in2101_2 = {s1369[0]};
    Full_Adder FA_2101(s2101, c2101, in2101_1, in2101_2, c1367);
    wire[0:0] s2102, in2102_1, in2102_2;
    wire c2102;
    assign in2102_1 = {s1371[0]};
    assign in2102_2 = {s1372[0]};
    Full_Adder FA_2102(s2102, c2102, in2102_1, in2102_2, s1370[0]);
    wire[0:0] s2103, in2103_1, in2103_2;
    wire c2103;
    assign in2103_1 = {s1374[0]};
    assign in2103_2 = {s1375[0]};
    Full_Adder FA_2103(s2103, c2103, in2103_1, in2103_2, s1373[0]);
    wire[0:0] s2104, in2104_1, in2104_2;
    wire c2104;
    assign in2104_1 = {s507[0]};
    assign in2104_2 = {c1369};
    Full_Adder FA_2104(s2104, c2104, in2104_1, in2104_2, s506[0]);
    wire[0:0] s2105, in2105_1, in2105_2;
    wire c2105;
    assign in2105_1 = {c1371};
    assign in2105_2 = {c1372};
    Full_Adder FA_2105(s2105, c2105, in2105_1, in2105_2, c1370);
    wire[0:0] s2106, in2106_1, in2106_2;
    wire c2106;
    assign in2106_1 = {c1374};
    assign in2106_2 = {c1375};
    Full_Adder FA_2106(s2106, c2106, in2106_1, in2106_2, c1373);
    wire[0:0] s2107, in2107_1, in2107_2;
    wire c2107;
    assign in2107_1 = {c1377};
    assign in2107_2 = {s1378[0]};
    Full_Adder FA_2107(s2107, c2107, in2107_1, in2107_2, c1376);
    wire[0:0] s2108, in2108_1, in2108_2;
    wire c2108;
    assign in2108_1 = {s1380[0]};
    assign in2108_2 = {s1381[0]};
    Full_Adder FA_2108(s2108, c2108, in2108_1, in2108_2, s1379[0]);
    wire[0:0] s2109, in2109_1, in2109_2;
    wire c2109;
    assign in2109_1 = {s1383[0]};
    assign in2109_2 = {s1384[0]};
    Full_Adder FA_2109(s2109, c2109, in2109_1, in2109_2, s1382[0]);
    wire[0:0] s2110, in2110_1, in2110_2;
    wire c2110;
    assign in2110_1 = {s517[0]};
    assign in2110_2 = {c1378};
    Full_Adder FA_2110(s2110, c2110, in2110_1, in2110_2, s516[0]);
    wire[0:0] s2111, in2111_1, in2111_2;
    wire c2111;
    assign in2111_1 = {c1380};
    assign in2111_2 = {c1381};
    Full_Adder FA_2111(s2111, c2111, in2111_1, in2111_2, c1379);
    wire[0:0] s2112, in2112_1, in2112_2;
    wire c2112;
    assign in2112_1 = {c1383};
    assign in2112_2 = {c1384};
    Full_Adder FA_2112(s2112, c2112, in2112_1, in2112_2, c1382);
    wire[0:0] s2113, in2113_1, in2113_2;
    wire c2113;
    assign in2113_1 = {c1386};
    assign in2113_2 = {s1387[0]};
    Full_Adder FA_2113(s2113, c2113, in2113_1, in2113_2, c1385);
    wire[0:0] s2114, in2114_1, in2114_2;
    wire c2114;
    assign in2114_1 = {s1389[0]};
    assign in2114_2 = {s1390[0]};
    Full_Adder FA_2114(s2114, c2114, in2114_1, in2114_2, s1388[0]);
    wire[0:0] s2115, in2115_1, in2115_2;
    wire c2115;
    assign in2115_1 = {s1392[0]};
    assign in2115_2 = {s1393[0]};
    Full_Adder FA_2115(s2115, c2115, in2115_1, in2115_2, s1391[0]);
    wire[0:0] s2116, in2116_1, in2116_2;
    wire c2116;
    assign in2116_1 = {s528[0]};
    assign in2116_2 = {c1387};
    Full_Adder FA_2116(s2116, c2116, in2116_1, in2116_2, s527[0]);
    wire[0:0] s2117, in2117_1, in2117_2;
    wire c2117;
    assign in2117_1 = {c1389};
    assign in2117_2 = {c1390};
    Full_Adder FA_2117(s2117, c2117, in2117_1, in2117_2, c1388);
    wire[0:0] s2118, in2118_1, in2118_2;
    wire c2118;
    assign in2118_1 = {c1392};
    assign in2118_2 = {c1393};
    Full_Adder FA_2118(s2118, c2118, in2118_1, in2118_2, c1391);
    wire[0:0] s2119, in2119_1, in2119_2;
    wire c2119;
    assign in2119_1 = {c1395};
    assign in2119_2 = {s1396[0]};
    Full_Adder FA_2119(s2119, c2119, in2119_1, in2119_2, c1394);
    wire[0:0] s2120, in2120_1, in2120_2;
    wire c2120;
    assign in2120_1 = {s1398[0]};
    assign in2120_2 = {s1399[0]};
    Full_Adder FA_2120(s2120, c2120, in2120_1, in2120_2, s1397[0]);
    wire[0:0] s2121, in2121_1, in2121_2;
    wire c2121;
    assign in2121_1 = {s1401[0]};
    assign in2121_2 = {s1402[0]};
    Full_Adder FA_2121(s2121, c2121, in2121_1, in2121_2, s1400[0]);
    wire[0:0] s2122, in2122_1, in2122_2;
    wire c2122;
    assign in2122_1 = {s540[0]};
    assign in2122_2 = {c1396};
    Full_Adder FA_2122(s2122, c2122, in2122_1, in2122_2, s539[0]);
    wire[0:0] s2123, in2123_1, in2123_2;
    wire c2123;
    assign in2123_1 = {c1398};
    assign in2123_2 = {c1399};
    Full_Adder FA_2123(s2123, c2123, in2123_1, in2123_2, c1397);
    wire[0:0] s2124, in2124_1, in2124_2;
    wire c2124;
    assign in2124_1 = {c1401};
    assign in2124_2 = {c1402};
    Full_Adder FA_2124(s2124, c2124, in2124_1, in2124_2, c1400);
    wire[0:0] s2125, in2125_1, in2125_2;
    wire c2125;
    assign in2125_1 = {c1404};
    assign in2125_2 = {s1405[0]};
    Full_Adder FA_2125(s2125, c2125, in2125_1, in2125_2, c1403);
    wire[0:0] s2126, in2126_1, in2126_2;
    wire c2126;
    assign in2126_1 = {s1407[0]};
    assign in2126_2 = {s1408[0]};
    Full_Adder FA_2126(s2126, c2126, in2126_1, in2126_2, s1406[0]);
    wire[0:0] s2127, in2127_1, in2127_2;
    wire c2127;
    assign in2127_1 = {s1410[0]};
    assign in2127_2 = {s1411[0]};
    Full_Adder FA_2127(s2127, c2127, in2127_1, in2127_2, s1409[0]);
    wire[0:0] s2128, in2128_1, in2128_2;
    wire c2128;
    assign in2128_1 = {s553[0]};
    assign in2128_2 = {c1405};
    Full_Adder FA_2128(s2128, c2128, in2128_1, in2128_2, s552[0]);
    wire[0:0] s2129, in2129_1, in2129_2;
    wire c2129;
    assign in2129_1 = {c1407};
    assign in2129_2 = {c1408};
    Full_Adder FA_2129(s2129, c2129, in2129_1, in2129_2, c1406);
    wire[0:0] s2130, in2130_1, in2130_2;
    wire c2130;
    assign in2130_1 = {c1410};
    assign in2130_2 = {c1411};
    Full_Adder FA_2130(s2130, c2130, in2130_1, in2130_2, c1409);
    wire[0:0] s2131, in2131_1, in2131_2;
    wire c2131;
    assign in2131_1 = {c1413};
    assign in2131_2 = {s1414[0]};
    Full_Adder FA_2131(s2131, c2131, in2131_1, in2131_2, c1412);
    wire[0:0] s2132, in2132_1, in2132_2;
    wire c2132;
    assign in2132_1 = {s1416[0]};
    assign in2132_2 = {s1417[0]};
    Full_Adder FA_2132(s2132, c2132, in2132_1, in2132_2, s1415[0]);
    wire[0:0] s2133, in2133_1, in2133_2;
    wire c2133;
    assign in2133_1 = {s1419[0]};
    assign in2133_2 = {s1420[0]};
    Full_Adder FA_2133(s2133, c2133, in2133_1, in2133_2, s1418[0]);
    wire[0:0] s2134, in2134_1, in2134_2;
    wire c2134;
    assign in2134_1 = {s567[0]};
    assign in2134_2 = {c1414};
    Full_Adder FA_2134(s2134, c2134, in2134_1, in2134_2, s566[0]);
    wire[0:0] s2135, in2135_1, in2135_2;
    wire c2135;
    assign in2135_1 = {c1416};
    assign in2135_2 = {c1417};
    Full_Adder FA_2135(s2135, c2135, in2135_1, in2135_2, c1415);
    wire[0:0] s2136, in2136_1, in2136_2;
    wire c2136;
    assign in2136_1 = {c1419};
    assign in2136_2 = {c1420};
    Full_Adder FA_2136(s2136, c2136, in2136_1, in2136_2, c1418);
    wire[0:0] s2137, in2137_1, in2137_2;
    wire c2137;
    assign in2137_1 = {c1422};
    assign in2137_2 = {s1423[0]};
    Full_Adder FA_2137(s2137, c2137, in2137_1, in2137_2, c1421);
    wire[0:0] s2138, in2138_1, in2138_2;
    wire c2138;
    assign in2138_1 = {s1425[0]};
    assign in2138_2 = {s1426[0]};
    Full_Adder FA_2138(s2138, c2138, in2138_1, in2138_2, s1424[0]);
    wire[0:0] s2139, in2139_1, in2139_2;
    wire c2139;
    assign in2139_1 = {s1428[0]};
    assign in2139_2 = {s1429[0]};
    Full_Adder FA_2139(s2139, c2139, in2139_1, in2139_2, s1427[0]);
    wire[0:0] s2140, in2140_1, in2140_2;
    wire c2140;
    assign in2140_1 = {s581[0]};
    assign in2140_2 = {c1423};
    Full_Adder FA_2140(s2140, c2140, in2140_1, in2140_2, s580[0]);
    wire[0:0] s2141, in2141_1, in2141_2;
    wire c2141;
    assign in2141_1 = {c1425};
    assign in2141_2 = {c1426};
    Full_Adder FA_2141(s2141, c2141, in2141_1, in2141_2, c1424);
    wire[0:0] s2142, in2142_1, in2142_2;
    wire c2142;
    assign in2142_1 = {c1428};
    assign in2142_2 = {c1429};
    Full_Adder FA_2142(s2142, c2142, in2142_1, in2142_2, c1427);
    wire[0:0] s2143, in2143_1, in2143_2;
    wire c2143;
    assign in2143_1 = {c1431};
    assign in2143_2 = {s1432[0]};
    Full_Adder FA_2143(s2143, c2143, in2143_1, in2143_2, c1430);
    wire[0:0] s2144, in2144_1, in2144_2;
    wire c2144;
    assign in2144_1 = {s1434[0]};
    assign in2144_2 = {s1435[0]};
    Full_Adder FA_2144(s2144, c2144, in2144_1, in2144_2, s1433[0]);
    wire[0:0] s2145, in2145_1, in2145_2;
    wire c2145;
    assign in2145_1 = {s1437[0]};
    assign in2145_2 = {s1438[0]};
    Full_Adder FA_2145(s2145, c2145, in2145_1, in2145_2, s1436[0]);
    wire[0:0] s2146, in2146_1, in2146_2;
    wire c2146;
    assign in2146_1 = {s595[0]};
    assign in2146_2 = {c1432};
    Full_Adder FA_2146(s2146, c2146, in2146_1, in2146_2, s594[0]);
    wire[0:0] s2147, in2147_1, in2147_2;
    wire c2147;
    assign in2147_1 = {c1434};
    assign in2147_2 = {c1435};
    Full_Adder FA_2147(s2147, c2147, in2147_1, in2147_2, c1433);
    wire[0:0] s2148, in2148_1, in2148_2;
    wire c2148;
    assign in2148_1 = {c1437};
    assign in2148_2 = {c1438};
    Full_Adder FA_2148(s2148, c2148, in2148_1, in2148_2, c1436);
    wire[0:0] s2149, in2149_1, in2149_2;
    wire c2149;
    assign in2149_1 = {c1440};
    assign in2149_2 = {s1441[0]};
    Full_Adder FA_2149(s2149, c2149, in2149_1, in2149_2, c1439);
    wire[0:0] s2150, in2150_1, in2150_2;
    wire c2150;
    assign in2150_1 = {s1443[0]};
    assign in2150_2 = {s1444[0]};
    Full_Adder FA_2150(s2150, c2150, in2150_1, in2150_2, s1442[0]);
    wire[0:0] s2151, in2151_1, in2151_2;
    wire c2151;
    assign in2151_1 = {s1446[0]};
    assign in2151_2 = {s1447[0]};
    Full_Adder FA_2151(s2151, c2151, in2151_1, in2151_2, s1445[0]);
    wire[0:0] s2152, in2152_1, in2152_2;
    wire c2152;
    assign in2152_1 = {s609[0]};
    assign in2152_2 = {c1441};
    Full_Adder FA_2152(s2152, c2152, in2152_1, in2152_2, s608[0]);
    wire[0:0] s2153, in2153_1, in2153_2;
    wire c2153;
    assign in2153_1 = {c1443};
    assign in2153_2 = {c1444};
    Full_Adder FA_2153(s2153, c2153, in2153_1, in2153_2, c1442);
    wire[0:0] s2154, in2154_1, in2154_2;
    wire c2154;
    assign in2154_1 = {c1446};
    assign in2154_2 = {c1447};
    Full_Adder FA_2154(s2154, c2154, in2154_1, in2154_2, c1445);
    wire[0:0] s2155, in2155_1, in2155_2;
    wire c2155;
    assign in2155_1 = {c1449};
    assign in2155_2 = {s1450[0]};
    Full_Adder FA_2155(s2155, c2155, in2155_1, in2155_2, c1448);
    wire[0:0] s2156, in2156_1, in2156_2;
    wire c2156;
    assign in2156_1 = {s1452[0]};
    assign in2156_2 = {s1453[0]};
    Full_Adder FA_2156(s2156, c2156, in2156_1, in2156_2, s1451[0]);
    wire[0:0] s2157, in2157_1, in2157_2;
    wire c2157;
    assign in2157_1 = {s1455[0]};
    assign in2157_2 = {s1456[0]};
    Full_Adder FA_2157(s2157, c2157, in2157_1, in2157_2, s1454[0]);
    wire[0:0] s2158, in2158_1, in2158_2;
    wire c2158;
    assign in2158_1 = {s623[0]};
    assign in2158_2 = {c1450};
    Full_Adder FA_2158(s2158, c2158, in2158_1, in2158_2, s622[0]);
    wire[0:0] s2159, in2159_1, in2159_2;
    wire c2159;
    assign in2159_1 = {c1452};
    assign in2159_2 = {c1453};
    Full_Adder FA_2159(s2159, c2159, in2159_1, in2159_2, c1451);
    wire[0:0] s2160, in2160_1, in2160_2;
    wire c2160;
    assign in2160_1 = {c1455};
    assign in2160_2 = {c1456};
    Full_Adder FA_2160(s2160, c2160, in2160_1, in2160_2, c1454);
    wire[0:0] s2161, in2161_1, in2161_2;
    wire c2161;
    assign in2161_1 = {c1458};
    assign in2161_2 = {s1459[0]};
    Full_Adder FA_2161(s2161, c2161, in2161_1, in2161_2, c1457);
    wire[0:0] s2162, in2162_1, in2162_2;
    wire c2162;
    assign in2162_1 = {s1461[0]};
    assign in2162_2 = {s1462[0]};
    Full_Adder FA_2162(s2162, c2162, in2162_1, in2162_2, s1460[0]);
    wire[0:0] s2163, in2163_1, in2163_2;
    wire c2163;
    assign in2163_1 = {s1464[0]};
    assign in2163_2 = {s1465[0]};
    Full_Adder FA_2163(s2163, c2163, in2163_1, in2163_2, s1463[0]);
    wire[0:0] s2164, in2164_1, in2164_2;
    wire c2164;
    assign in2164_1 = {s637[0]};
    assign in2164_2 = {c1459};
    Full_Adder FA_2164(s2164, c2164, in2164_1, in2164_2, s636[0]);
    wire[0:0] s2165, in2165_1, in2165_2;
    wire c2165;
    assign in2165_1 = {c1461};
    assign in2165_2 = {c1462};
    Full_Adder FA_2165(s2165, c2165, in2165_1, in2165_2, c1460);
    wire[0:0] s2166, in2166_1, in2166_2;
    wire c2166;
    assign in2166_1 = {c1464};
    assign in2166_2 = {c1465};
    Full_Adder FA_2166(s2166, c2166, in2166_1, in2166_2, c1463);
    wire[0:0] s2167, in2167_1, in2167_2;
    wire c2167;
    assign in2167_1 = {c1467};
    assign in2167_2 = {s1468[0]};
    Full_Adder FA_2167(s2167, c2167, in2167_1, in2167_2, c1466);
    wire[0:0] s2168, in2168_1, in2168_2;
    wire c2168;
    assign in2168_1 = {s1470[0]};
    assign in2168_2 = {s1471[0]};
    Full_Adder FA_2168(s2168, c2168, in2168_1, in2168_2, s1469[0]);
    wire[0:0] s2169, in2169_1, in2169_2;
    wire c2169;
    assign in2169_1 = {s1473[0]};
    assign in2169_2 = {s1474[0]};
    Full_Adder FA_2169(s2169, c2169, in2169_1, in2169_2, s1472[0]);
    wire[0:0] s2170, in2170_1, in2170_2;
    wire c2170;
    assign in2170_1 = {s651[0]};
    assign in2170_2 = {c1468};
    Full_Adder FA_2170(s2170, c2170, in2170_1, in2170_2, s650[0]);
    wire[0:0] s2171, in2171_1, in2171_2;
    wire c2171;
    assign in2171_1 = {c1470};
    assign in2171_2 = {c1471};
    Full_Adder FA_2171(s2171, c2171, in2171_1, in2171_2, c1469);
    wire[0:0] s2172, in2172_1, in2172_2;
    wire c2172;
    assign in2172_1 = {c1473};
    assign in2172_2 = {c1474};
    Full_Adder FA_2172(s2172, c2172, in2172_1, in2172_2, c1472);
    wire[0:0] s2173, in2173_1, in2173_2;
    wire c2173;
    assign in2173_1 = {c1476};
    assign in2173_2 = {s1477[0]};
    Full_Adder FA_2173(s2173, c2173, in2173_1, in2173_2, c1475);
    wire[0:0] s2174, in2174_1, in2174_2;
    wire c2174;
    assign in2174_1 = {s1479[0]};
    assign in2174_2 = {s1480[0]};
    Full_Adder FA_2174(s2174, c2174, in2174_1, in2174_2, s1478[0]);
    wire[0:0] s2175, in2175_1, in2175_2;
    wire c2175;
    assign in2175_1 = {s1482[0]};
    assign in2175_2 = {s1483[0]};
    Full_Adder FA_2175(s2175, c2175, in2175_1, in2175_2, s1481[0]);
    wire[0:0] s2176, in2176_1, in2176_2;
    wire c2176;
    assign in2176_1 = {s665[0]};
    assign in2176_2 = {c1477};
    Full_Adder FA_2176(s2176, c2176, in2176_1, in2176_2, s664[0]);
    wire[0:0] s2177, in2177_1, in2177_2;
    wire c2177;
    assign in2177_1 = {c1479};
    assign in2177_2 = {c1480};
    Full_Adder FA_2177(s2177, c2177, in2177_1, in2177_2, c1478);
    wire[0:0] s2178, in2178_1, in2178_2;
    wire c2178;
    assign in2178_1 = {c1482};
    assign in2178_2 = {c1483};
    Full_Adder FA_2178(s2178, c2178, in2178_1, in2178_2, c1481);
    wire[0:0] s2179, in2179_1, in2179_2;
    wire c2179;
    assign in2179_1 = {c1485};
    assign in2179_2 = {s1486[0]};
    Full_Adder FA_2179(s2179, c2179, in2179_1, in2179_2, c1484);
    wire[0:0] s2180, in2180_1, in2180_2;
    wire c2180;
    assign in2180_1 = {s1488[0]};
    assign in2180_2 = {s1489[0]};
    Full_Adder FA_2180(s2180, c2180, in2180_1, in2180_2, s1487[0]);
    wire[0:0] s2181, in2181_1, in2181_2;
    wire c2181;
    assign in2181_1 = {s1491[0]};
    assign in2181_2 = {s1492[0]};
    Full_Adder FA_2181(s2181, c2181, in2181_1, in2181_2, s1490[0]);
    wire[0:0] s2182, in2182_1, in2182_2;
    wire c2182;
    assign in2182_1 = {s679[0]};
    assign in2182_2 = {c1486};
    Full_Adder FA_2182(s2182, c2182, in2182_1, in2182_2, s678[0]);
    wire[0:0] s2183, in2183_1, in2183_2;
    wire c2183;
    assign in2183_1 = {c1488};
    assign in2183_2 = {c1489};
    Full_Adder FA_2183(s2183, c2183, in2183_1, in2183_2, c1487);
    wire[0:0] s2184, in2184_1, in2184_2;
    wire c2184;
    assign in2184_1 = {c1491};
    assign in2184_2 = {c1492};
    Full_Adder FA_2184(s2184, c2184, in2184_1, in2184_2, c1490);
    wire[0:0] s2185, in2185_1, in2185_2;
    wire c2185;
    assign in2185_1 = {c1494};
    assign in2185_2 = {s1495[0]};
    Full_Adder FA_2185(s2185, c2185, in2185_1, in2185_2, c1493);
    wire[0:0] s2186, in2186_1, in2186_2;
    wire c2186;
    assign in2186_1 = {s1497[0]};
    assign in2186_2 = {s1498[0]};
    Full_Adder FA_2186(s2186, c2186, in2186_1, in2186_2, s1496[0]);
    wire[0:0] s2187, in2187_1, in2187_2;
    wire c2187;
    assign in2187_1 = {s1500[0]};
    assign in2187_2 = {s1501[0]};
    Full_Adder FA_2187(s2187, c2187, in2187_1, in2187_2, s1499[0]);
    wire[0:0] s2188, in2188_1, in2188_2;
    wire c2188;
    assign in2188_1 = {s693[0]};
    assign in2188_2 = {c1495};
    Full_Adder FA_2188(s2188, c2188, in2188_1, in2188_2, s692[0]);
    wire[0:0] s2189, in2189_1, in2189_2;
    wire c2189;
    assign in2189_1 = {c1497};
    assign in2189_2 = {c1498};
    Full_Adder FA_2189(s2189, c2189, in2189_1, in2189_2, c1496);
    wire[0:0] s2190, in2190_1, in2190_2;
    wire c2190;
    assign in2190_1 = {c1500};
    assign in2190_2 = {c1501};
    Full_Adder FA_2190(s2190, c2190, in2190_1, in2190_2, c1499);
    wire[0:0] s2191, in2191_1, in2191_2;
    wire c2191;
    assign in2191_1 = {c1503};
    assign in2191_2 = {s1504[0]};
    Full_Adder FA_2191(s2191, c2191, in2191_1, in2191_2, c1502);
    wire[0:0] s2192, in2192_1, in2192_2;
    wire c2192;
    assign in2192_1 = {s1506[0]};
    assign in2192_2 = {s1507[0]};
    Full_Adder FA_2192(s2192, c2192, in2192_1, in2192_2, s1505[0]);
    wire[0:0] s2193, in2193_1, in2193_2;
    wire c2193;
    assign in2193_1 = {s1509[0]};
    assign in2193_2 = {s1510[0]};
    Full_Adder FA_2193(s2193, c2193, in2193_1, in2193_2, s1508[0]);
    wire[0:0] s2194, in2194_1, in2194_2;
    wire c2194;
    assign in2194_1 = {s707[0]};
    assign in2194_2 = {c1504};
    Full_Adder FA_2194(s2194, c2194, in2194_1, in2194_2, s706[0]);
    wire[0:0] s2195, in2195_1, in2195_2;
    wire c2195;
    assign in2195_1 = {c1506};
    assign in2195_2 = {c1507};
    Full_Adder FA_2195(s2195, c2195, in2195_1, in2195_2, c1505);
    wire[0:0] s2196, in2196_1, in2196_2;
    wire c2196;
    assign in2196_1 = {c1509};
    assign in2196_2 = {c1510};
    Full_Adder FA_2196(s2196, c2196, in2196_1, in2196_2, c1508);
    wire[0:0] s2197, in2197_1, in2197_2;
    wire c2197;
    assign in2197_1 = {c1512};
    assign in2197_2 = {s1513[0]};
    Full_Adder FA_2197(s2197, c2197, in2197_1, in2197_2, c1511);
    wire[0:0] s2198, in2198_1, in2198_2;
    wire c2198;
    assign in2198_1 = {s1515[0]};
    assign in2198_2 = {s1516[0]};
    Full_Adder FA_2198(s2198, c2198, in2198_1, in2198_2, s1514[0]);
    wire[0:0] s2199, in2199_1, in2199_2;
    wire c2199;
    assign in2199_1 = {s1518[0]};
    assign in2199_2 = {s1519[0]};
    Full_Adder FA_2199(s2199, c2199, in2199_1, in2199_2, s1517[0]);
    wire[0:0] s2200, in2200_1, in2200_2;
    wire c2200;
    assign in2200_1 = {s721[0]};
    assign in2200_2 = {c1513};
    Full_Adder FA_2200(s2200, c2200, in2200_1, in2200_2, s720[0]);
    wire[0:0] s2201, in2201_1, in2201_2;
    wire c2201;
    assign in2201_1 = {c1515};
    assign in2201_2 = {c1516};
    Full_Adder FA_2201(s2201, c2201, in2201_1, in2201_2, c1514);
    wire[0:0] s2202, in2202_1, in2202_2;
    wire c2202;
    assign in2202_1 = {c1518};
    assign in2202_2 = {c1519};
    Full_Adder FA_2202(s2202, c2202, in2202_1, in2202_2, c1517);
    wire[0:0] s2203, in2203_1, in2203_2;
    wire c2203;
    assign in2203_1 = {c1521};
    assign in2203_2 = {s1522[0]};
    Full_Adder FA_2203(s2203, c2203, in2203_1, in2203_2, c1520);
    wire[0:0] s2204, in2204_1, in2204_2;
    wire c2204;
    assign in2204_1 = {s1524[0]};
    assign in2204_2 = {s1525[0]};
    Full_Adder FA_2204(s2204, c2204, in2204_1, in2204_2, s1523[0]);
    wire[0:0] s2205, in2205_1, in2205_2;
    wire c2205;
    assign in2205_1 = {s1527[0]};
    assign in2205_2 = {s1528[0]};
    Full_Adder FA_2205(s2205, c2205, in2205_1, in2205_2, s1526[0]);
    wire[0:0] s2206, in2206_1, in2206_2;
    wire c2206;
    assign in2206_1 = {s735[0]};
    assign in2206_2 = {c1522};
    Full_Adder FA_2206(s2206, c2206, in2206_1, in2206_2, s734[0]);
    wire[0:0] s2207, in2207_1, in2207_2;
    wire c2207;
    assign in2207_1 = {c1524};
    assign in2207_2 = {c1525};
    Full_Adder FA_2207(s2207, c2207, in2207_1, in2207_2, c1523);
    wire[0:0] s2208, in2208_1, in2208_2;
    wire c2208;
    assign in2208_1 = {c1527};
    assign in2208_2 = {c1528};
    Full_Adder FA_2208(s2208, c2208, in2208_1, in2208_2, c1526);
    wire[0:0] s2209, in2209_1, in2209_2;
    wire c2209;
    assign in2209_1 = {c1530};
    assign in2209_2 = {s1531[0]};
    Full_Adder FA_2209(s2209, c2209, in2209_1, in2209_2, c1529);
    wire[0:0] s2210, in2210_1, in2210_2;
    wire c2210;
    assign in2210_1 = {s1533[0]};
    assign in2210_2 = {s1534[0]};
    Full_Adder FA_2210(s2210, c2210, in2210_1, in2210_2, s1532[0]);
    wire[0:0] s2211, in2211_1, in2211_2;
    wire c2211;
    assign in2211_1 = {s1536[0]};
    assign in2211_2 = {s1537[0]};
    Full_Adder FA_2211(s2211, c2211, in2211_1, in2211_2, s1535[0]);
    wire[0:0] s2212, in2212_1, in2212_2;
    wire c2212;
    assign in2212_1 = {s749[0]};
    assign in2212_2 = {c1531};
    Full_Adder FA_2212(s2212, c2212, in2212_1, in2212_2, s748[0]);
    wire[0:0] s2213, in2213_1, in2213_2;
    wire c2213;
    assign in2213_1 = {c1533};
    assign in2213_2 = {c1534};
    Full_Adder FA_2213(s2213, c2213, in2213_1, in2213_2, c1532);
    wire[0:0] s2214, in2214_1, in2214_2;
    wire c2214;
    assign in2214_1 = {c1536};
    assign in2214_2 = {c1537};
    Full_Adder FA_2214(s2214, c2214, in2214_1, in2214_2, c1535);
    wire[0:0] s2215, in2215_1, in2215_2;
    wire c2215;
    assign in2215_1 = {c1539};
    assign in2215_2 = {s1540[0]};
    Full_Adder FA_2215(s2215, c2215, in2215_1, in2215_2, c1538);
    wire[0:0] s2216, in2216_1, in2216_2;
    wire c2216;
    assign in2216_1 = {s1542[0]};
    assign in2216_2 = {s1543[0]};
    Full_Adder FA_2216(s2216, c2216, in2216_1, in2216_2, s1541[0]);
    wire[0:0] s2217, in2217_1, in2217_2;
    wire c2217;
    assign in2217_1 = {s1545[0]};
    assign in2217_2 = {s1546[0]};
    Full_Adder FA_2217(s2217, c2217, in2217_1, in2217_2, s1544[0]);
    wire[0:0] s2218, in2218_1, in2218_2;
    wire c2218;
    assign in2218_1 = {s763[0]};
    assign in2218_2 = {c1540};
    Full_Adder FA_2218(s2218, c2218, in2218_1, in2218_2, s762[0]);
    wire[0:0] s2219, in2219_1, in2219_2;
    wire c2219;
    assign in2219_1 = {c1542};
    assign in2219_2 = {c1543};
    Full_Adder FA_2219(s2219, c2219, in2219_1, in2219_2, c1541);
    wire[0:0] s2220, in2220_1, in2220_2;
    wire c2220;
    assign in2220_1 = {c1545};
    assign in2220_2 = {c1546};
    Full_Adder FA_2220(s2220, c2220, in2220_1, in2220_2, c1544);
    wire[0:0] s2221, in2221_1, in2221_2;
    wire c2221;
    assign in2221_1 = {c1548};
    assign in2221_2 = {s1549[0]};
    Full_Adder FA_2221(s2221, c2221, in2221_1, in2221_2, c1547);
    wire[0:0] s2222, in2222_1, in2222_2;
    wire c2222;
    assign in2222_1 = {s1551[0]};
    assign in2222_2 = {s1552[0]};
    Full_Adder FA_2222(s2222, c2222, in2222_1, in2222_2, s1550[0]);
    wire[0:0] s2223, in2223_1, in2223_2;
    wire c2223;
    assign in2223_1 = {s1554[0]};
    assign in2223_2 = {s1555[0]};
    Full_Adder FA_2223(s2223, c2223, in2223_1, in2223_2, s1553[0]);
    wire[0:0] s2224, in2224_1, in2224_2;
    wire c2224;
    assign in2224_1 = {s777[0]};
    assign in2224_2 = {c1549};
    Full_Adder FA_2224(s2224, c2224, in2224_1, in2224_2, s776[0]);
    wire[0:0] s2225, in2225_1, in2225_2;
    wire c2225;
    assign in2225_1 = {c1551};
    assign in2225_2 = {c1552};
    Full_Adder FA_2225(s2225, c2225, in2225_1, in2225_2, c1550);
    wire[0:0] s2226, in2226_1, in2226_2;
    wire c2226;
    assign in2226_1 = {c1554};
    assign in2226_2 = {c1555};
    Full_Adder FA_2226(s2226, c2226, in2226_1, in2226_2, c1553);
    wire[0:0] s2227, in2227_1, in2227_2;
    wire c2227;
    assign in2227_1 = {c1557};
    assign in2227_2 = {s1558[0]};
    Full_Adder FA_2227(s2227, c2227, in2227_1, in2227_2, c1556);
    wire[0:0] s2228, in2228_1, in2228_2;
    wire c2228;
    assign in2228_1 = {s1560[0]};
    assign in2228_2 = {s1561[0]};
    Full_Adder FA_2228(s2228, c2228, in2228_1, in2228_2, s1559[0]);
    wire[0:0] s2229, in2229_1, in2229_2;
    wire c2229;
    assign in2229_1 = {s1563[0]};
    assign in2229_2 = {s1564[0]};
    Full_Adder FA_2229(s2229, c2229, in2229_1, in2229_2, s1562[0]);
    wire[0:0] s2230, in2230_1, in2230_2;
    wire c2230;
    assign in2230_1 = {s791[0]};
    assign in2230_2 = {c1558};
    Full_Adder FA_2230(s2230, c2230, in2230_1, in2230_2, s790[0]);
    wire[0:0] s2231, in2231_1, in2231_2;
    wire c2231;
    assign in2231_1 = {c1560};
    assign in2231_2 = {c1561};
    Full_Adder FA_2231(s2231, c2231, in2231_1, in2231_2, c1559);
    wire[0:0] s2232, in2232_1, in2232_2;
    wire c2232;
    assign in2232_1 = {c1563};
    assign in2232_2 = {c1564};
    Full_Adder FA_2232(s2232, c2232, in2232_1, in2232_2, c1562);
    wire[0:0] s2233, in2233_1, in2233_2;
    wire c2233;
    assign in2233_1 = {c1566};
    assign in2233_2 = {s1567[0]};
    Full_Adder FA_2233(s2233, c2233, in2233_1, in2233_2, c1565);
    wire[0:0] s2234, in2234_1, in2234_2;
    wire c2234;
    assign in2234_1 = {s1569[0]};
    assign in2234_2 = {s1570[0]};
    Full_Adder FA_2234(s2234, c2234, in2234_1, in2234_2, s1568[0]);
    wire[0:0] s2235, in2235_1, in2235_2;
    wire c2235;
    assign in2235_1 = {s1572[0]};
    assign in2235_2 = {s1573[0]};
    Full_Adder FA_2235(s2235, c2235, in2235_1, in2235_2, s1571[0]);
    wire[0:0] s2236, in2236_1, in2236_2;
    wire c2236;
    assign in2236_1 = {s805[0]};
    assign in2236_2 = {c1567};
    Full_Adder FA_2236(s2236, c2236, in2236_1, in2236_2, s804[0]);
    wire[0:0] s2237, in2237_1, in2237_2;
    wire c2237;
    assign in2237_1 = {c1569};
    assign in2237_2 = {c1570};
    Full_Adder FA_2237(s2237, c2237, in2237_1, in2237_2, c1568);
    wire[0:0] s2238, in2238_1, in2238_2;
    wire c2238;
    assign in2238_1 = {c1572};
    assign in2238_2 = {c1573};
    Full_Adder FA_2238(s2238, c2238, in2238_1, in2238_2, c1571);
    wire[0:0] s2239, in2239_1, in2239_2;
    wire c2239;
    assign in2239_1 = {c1575};
    assign in2239_2 = {s1576[0]};
    Full_Adder FA_2239(s2239, c2239, in2239_1, in2239_2, c1574);
    wire[0:0] s2240, in2240_1, in2240_2;
    wire c2240;
    assign in2240_1 = {s1578[0]};
    assign in2240_2 = {s1579[0]};
    Full_Adder FA_2240(s2240, c2240, in2240_1, in2240_2, s1577[0]);
    wire[0:0] s2241, in2241_1, in2241_2;
    wire c2241;
    assign in2241_1 = {s1581[0]};
    assign in2241_2 = {s1582[0]};
    Full_Adder FA_2241(s2241, c2241, in2241_1, in2241_2, s1580[0]);
    wire[0:0] s2242, in2242_1, in2242_2;
    wire c2242;
    assign in2242_1 = {s819[0]};
    assign in2242_2 = {c1576};
    Full_Adder FA_2242(s2242, c2242, in2242_1, in2242_2, s818[0]);
    wire[0:0] s2243, in2243_1, in2243_2;
    wire c2243;
    assign in2243_1 = {c1578};
    assign in2243_2 = {c1579};
    Full_Adder FA_2243(s2243, c2243, in2243_1, in2243_2, c1577);
    wire[0:0] s2244, in2244_1, in2244_2;
    wire c2244;
    assign in2244_1 = {c1581};
    assign in2244_2 = {c1582};
    Full_Adder FA_2244(s2244, c2244, in2244_1, in2244_2, c1580);
    wire[0:0] s2245, in2245_1, in2245_2;
    wire c2245;
    assign in2245_1 = {c1584};
    assign in2245_2 = {s1585[0]};
    Full_Adder FA_2245(s2245, c2245, in2245_1, in2245_2, c1583);
    wire[0:0] s2246, in2246_1, in2246_2;
    wire c2246;
    assign in2246_1 = {s1587[0]};
    assign in2246_2 = {s1588[0]};
    Full_Adder FA_2246(s2246, c2246, in2246_1, in2246_2, s1586[0]);
    wire[0:0] s2247, in2247_1, in2247_2;
    wire c2247;
    assign in2247_1 = {s1590[0]};
    assign in2247_2 = {s1591[0]};
    Full_Adder FA_2247(s2247, c2247, in2247_1, in2247_2, s1589[0]);
    wire[0:0] s2248, in2248_1, in2248_2;
    wire c2248;
    assign in2248_1 = {s833[0]};
    assign in2248_2 = {c1585};
    Full_Adder FA_2248(s2248, c2248, in2248_1, in2248_2, s832[0]);
    wire[0:0] s2249, in2249_1, in2249_2;
    wire c2249;
    assign in2249_1 = {c1587};
    assign in2249_2 = {c1588};
    Full_Adder FA_2249(s2249, c2249, in2249_1, in2249_2, c1586);
    wire[0:0] s2250, in2250_1, in2250_2;
    wire c2250;
    assign in2250_1 = {c1590};
    assign in2250_2 = {c1591};
    Full_Adder FA_2250(s2250, c2250, in2250_1, in2250_2, c1589);
    wire[0:0] s2251, in2251_1, in2251_2;
    wire c2251;
    assign in2251_1 = {c1593};
    assign in2251_2 = {s1594[0]};
    Full_Adder FA_2251(s2251, c2251, in2251_1, in2251_2, c1592);
    wire[0:0] s2252, in2252_1, in2252_2;
    wire c2252;
    assign in2252_1 = {s1596[0]};
    assign in2252_2 = {s1597[0]};
    Full_Adder FA_2252(s2252, c2252, in2252_1, in2252_2, s1595[0]);
    wire[0:0] s2253, in2253_1, in2253_2;
    wire c2253;
    assign in2253_1 = {s1599[0]};
    assign in2253_2 = {s1600[0]};
    Full_Adder FA_2253(s2253, c2253, in2253_1, in2253_2, s1598[0]);
    wire[0:0] s2254, in2254_1, in2254_2;
    wire c2254;
    assign in2254_1 = {s847[0]};
    assign in2254_2 = {c1594};
    Full_Adder FA_2254(s2254, c2254, in2254_1, in2254_2, s846[0]);
    wire[0:0] s2255, in2255_1, in2255_2;
    wire c2255;
    assign in2255_1 = {c1596};
    assign in2255_2 = {c1597};
    Full_Adder FA_2255(s2255, c2255, in2255_1, in2255_2, c1595);
    wire[0:0] s2256, in2256_1, in2256_2;
    wire c2256;
    assign in2256_1 = {c1599};
    assign in2256_2 = {c1600};
    Full_Adder FA_2256(s2256, c2256, in2256_1, in2256_2, c1598);
    wire[0:0] s2257, in2257_1, in2257_2;
    wire c2257;
    assign in2257_1 = {c1602};
    assign in2257_2 = {s1603[0]};
    Full_Adder FA_2257(s2257, c2257, in2257_1, in2257_2, c1601);
    wire[0:0] s2258, in2258_1, in2258_2;
    wire c2258;
    assign in2258_1 = {s1605[0]};
    assign in2258_2 = {s1606[0]};
    Full_Adder FA_2258(s2258, c2258, in2258_1, in2258_2, s1604[0]);
    wire[0:0] s2259, in2259_1, in2259_2;
    wire c2259;
    assign in2259_1 = {s1608[0]};
    assign in2259_2 = {s1609[0]};
    Full_Adder FA_2259(s2259, c2259, in2259_1, in2259_2, s1607[0]);
    wire[0:0] s2260, in2260_1, in2260_2;
    wire c2260;
    assign in2260_1 = {s861[0]};
    assign in2260_2 = {c1603};
    Full_Adder FA_2260(s2260, c2260, in2260_1, in2260_2, s860[0]);
    wire[0:0] s2261, in2261_1, in2261_2;
    wire c2261;
    assign in2261_1 = {c1605};
    assign in2261_2 = {c1606};
    Full_Adder FA_2261(s2261, c2261, in2261_1, in2261_2, c1604);
    wire[0:0] s2262, in2262_1, in2262_2;
    wire c2262;
    assign in2262_1 = {c1608};
    assign in2262_2 = {c1609};
    Full_Adder FA_2262(s2262, c2262, in2262_1, in2262_2, c1607);
    wire[0:0] s2263, in2263_1, in2263_2;
    wire c2263;
    assign in2263_1 = {c1611};
    assign in2263_2 = {s1612[0]};
    Full_Adder FA_2263(s2263, c2263, in2263_1, in2263_2, c1610);
    wire[0:0] s2264, in2264_1, in2264_2;
    wire c2264;
    assign in2264_1 = {s1614[0]};
    assign in2264_2 = {s1615[0]};
    Full_Adder FA_2264(s2264, c2264, in2264_1, in2264_2, s1613[0]);
    wire[0:0] s2265, in2265_1, in2265_2;
    wire c2265;
    assign in2265_1 = {s1617[0]};
    assign in2265_2 = {s1618[0]};
    Full_Adder FA_2265(s2265, c2265, in2265_1, in2265_2, s1616[0]);
    wire[0:0] s2266, in2266_1, in2266_2;
    wire c2266;
    assign in2266_1 = {s875[0]};
    assign in2266_2 = {c1612};
    Full_Adder FA_2266(s2266, c2266, in2266_1, in2266_2, s874[0]);
    wire[0:0] s2267, in2267_1, in2267_2;
    wire c2267;
    assign in2267_1 = {c1614};
    assign in2267_2 = {c1615};
    Full_Adder FA_2267(s2267, c2267, in2267_1, in2267_2, c1613);
    wire[0:0] s2268, in2268_1, in2268_2;
    wire c2268;
    assign in2268_1 = {c1617};
    assign in2268_2 = {c1618};
    Full_Adder FA_2268(s2268, c2268, in2268_1, in2268_2, c1616);
    wire[0:0] s2269, in2269_1, in2269_2;
    wire c2269;
    assign in2269_1 = {c1620};
    assign in2269_2 = {s1621[0]};
    Full_Adder FA_2269(s2269, c2269, in2269_1, in2269_2, c1619);
    wire[0:0] s2270, in2270_1, in2270_2;
    wire c2270;
    assign in2270_1 = {s1623[0]};
    assign in2270_2 = {s1624[0]};
    Full_Adder FA_2270(s2270, c2270, in2270_1, in2270_2, s1622[0]);
    wire[0:0] s2271, in2271_1, in2271_2;
    wire c2271;
    assign in2271_1 = {s1626[0]};
    assign in2271_2 = {s1627[0]};
    Full_Adder FA_2271(s2271, c2271, in2271_1, in2271_2, s1625[0]);
    wire[0:0] s2272, in2272_1, in2272_2;
    wire c2272;
    assign in2272_1 = {s889[0]};
    assign in2272_2 = {c1621};
    Full_Adder FA_2272(s2272, c2272, in2272_1, in2272_2, s888[0]);
    wire[0:0] s2273, in2273_1, in2273_2;
    wire c2273;
    assign in2273_1 = {c1623};
    assign in2273_2 = {c1624};
    Full_Adder FA_2273(s2273, c2273, in2273_1, in2273_2, c1622);
    wire[0:0] s2274, in2274_1, in2274_2;
    wire c2274;
    assign in2274_1 = {c1626};
    assign in2274_2 = {c1627};
    Full_Adder FA_2274(s2274, c2274, in2274_1, in2274_2, c1625);
    wire[0:0] s2275, in2275_1, in2275_2;
    wire c2275;
    assign in2275_1 = {c1629};
    assign in2275_2 = {s1630[0]};
    Full_Adder FA_2275(s2275, c2275, in2275_1, in2275_2, c1628);
    wire[0:0] s2276, in2276_1, in2276_2;
    wire c2276;
    assign in2276_1 = {s1632[0]};
    assign in2276_2 = {s1633[0]};
    Full_Adder FA_2276(s2276, c2276, in2276_1, in2276_2, s1631[0]);
    wire[0:0] s2277, in2277_1, in2277_2;
    wire c2277;
    assign in2277_1 = {s1635[0]};
    assign in2277_2 = {s1636[0]};
    Full_Adder FA_2277(s2277, c2277, in2277_1, in2277_2, s1634[0]);
    wire[0:0] s2278, in2278_1, in2278_2;
    wire c2278;
    assign in2278_1 = {s903[0]};
    assign in2278_2 = {c1630};
    Full_Adder FA_2278(s2278, c2278, in2278_1, in2278_2, s902[0]);
    wire[0:0] s2279, in2279_1, in2279_2;
    wire c2279;
    assign in2279_1 = {c1632};
    assign in2279_2 = {c1633};
    Full_Adder FA_2279(s2279, c2279, in2279_1, in2279_2, c1631);
    wire[0:0] s2280, in2280_1, in2280_2;
    wire c2280;
    assign in2280_1 = {c1635};
    assign in2280_2 = {c1636};
    Full_Adder FA_2280(s2280, c2280, in2280_1, in2280_2, c1634);
    wire[0:0] s2281, in2281_1, in2281_2;
    wire c2281;
    assign in2281_1 = {c1638};
    assign in2281_2 = {s1639[0]};
    Full_Adder FA_2281(s2281, c2281, in2281_1, in2281_2, c1637);
    wire[0:0] s2282, in2282_1, in2282_2;
    wire c2282;
    assign in2282_1 = {s1641[0]};
    assign in2282_2 = {s1642[0]};
    Full_Adder FA_2282(s2282, c2282, in2282_1, in2282_2, s1640[0]);
    wire[0:0] s2283, in2283_1, in2283_2;
    wire c2283;
    assign in2283_1 = {s1644[0]};
    assign in2283_2 = {s1645[0]};
    Full_Adder FA_2283(s2283, c2283, in2283_1, in2283_2, s1643[0]);
    wire[0:0] s2284, in2284_1, in2284_2;
    wire c2284;
    assign in2284_1 = {s917[0]};
    assign in2284_2 = {c1639};
    Full_Adder FA_2284(s2284, c2284, in2284_1, in2284_2, s916[0]);
    wire[0:0] s2285, in2285_1, in2285_2;
    wire c2285;
    assign in2285_1 = {c1641};
    assign in2285_2 = {c1642};
    Full_Adder FA_2285(s2285, c2285, in2285_1, in2285_2, c1640);
    wire[0:0] s2286, in2286_1, in2286_2;
    wire c2286;
    assign in2286_1 = {c1644};
    assign in2286_2 = {c1645};
    Full_Adder FA_2286(s2286, c2286, in2286_1, in2286_2, c1643);
    wire[0:0] s2287, in2287_1, in2287_2;
    wire c2287;
    assign in2287_1 = {c1647};
    assign in2287_2 = {s1648[0]};
    Full_Adder FA_2287(s2287, c2287, in2287_1, in2287_2, c1646);
    wire[0:0] s2288, in2288_1, in2288_2;
    wire c2288;
    assign in2288_1 = {s1650[0]};
    assign in2288_2 = {s1651[0]};
    Full_Adder FA_2288(s2288, c2288, in2288_1, in2288_2, s1649[0]);
    wire[0:0] s2289, in2289_1, in2289_2;
    wire c2289;
    assign in2289_1 = {s1653[0]};
    assign in2289_2 = {s1654[0]};
    Full_Adder FA_2289(s2289, c2289, in2289_1, in2289_2, s1652[0]);
    wire[0:0] s2290, in2290_1, in2290_2;
    wire c2290;
    assign in2290_1 = {s931[0]};
    assign in2290_2 = {c1648};
    Full_Adder FA_2290(s2290, c2290, in2290_1, in2290_2, s930[0]);
    wire[0:0] s2291, in2291_1, in2291_2;
    wire c2291;
    assign in2291_1 = {c1650};
    assign in2291_2 = {c1651};
    Full_Adder FA_2291(s2291, c2291, in2291_1, in2291_2, c1649);
    wire[0:0] s2292, in2292_1, in2292_2;
    wire c2292;
    assign in2292_1 = {c1653};
    assign in2292_2 = {c1654};
    Full_Adder FA_2292(s2292, c2292, in2292_1, in2292_2, c1652);
    wire[0:0] s2293, in2293_1, in2293_2;
    wire c2293;
    assign in2293_1 = {c1656};
    assign in2293_2 = {s1657[0]};
    Full_Adder FA_2293(s2293, c2293, in2293_1, in2293_2, c1655);
    wire[0:0] s2294, in2294_1, in2294_2;
    wire c2294;
    assign in2294_1 = {s1659[0]};
    assign in2294_2 = {s1660[0]};
    Full_Adder FA_2294(s2294, c2294, in2294_1, in2294_2, s1658[0]);
    wire[0:0] s2295, in2295_1, in2295_2;
    wire c2295;
    assign in2295_1 = {s1662[0]};
    assign in2295_2 = {s1663[0]};
    Full_Adder FA_2295(s2295, c2295, in2295_1, in2295_2, s1661[0]);
    wire[0:0] s2296, in2296_1, in2296_2;
    wire c2296;
    assign in2296_1 = {s945[0]};
    assign in2296_2 = {c1657};
    Full_Adder FA_2296(s2296, c2296, in2296_1, in2296_2, s944[0]);
    wire[0:0] s2297, in2297_1, in2297_2;
    wire c2297;
    assign in2297_1 = {c1659};
    assign in2297_2 = {c1660};
    Full_Adder FA_2297(s2297, c2297, in2297_1, in2297_2, c1658);
    wire[0:0] s2298, in2298_1, in2298_2;
    wire c2298;
    assign in2298_1 = {c1662};
    assign in2298_2 = {c1663};
    Full_Adder FA_2298(s2298, c2298, in2298_1, in2298_2, c1661);
    wire[0:0] s2299, in2299_1, in2299_2;
    wire c2299;
    assign in2299_1 = {c1665};
    assign in2299_2 = {s1666[0]};
    Full_Adder FA_2299(s2299, c2299, in2299_1, in2299_2, c1664);
    wire[0:0] s2300, in2300_1, in2300_2;
    wire c2300;
    assign in2300_1 = {s1668[0]};
    assign in2300_2 = {s1669[0]};
    Full_Adder FA_2300(s2300, c2300, in2300_1, in2300_2, s1667[0]);
    wire[0:0] s2301, in2301_1, in2301_2;
    wire c2301;
    assign in2301_1 = {s1671[0]};
    assign in2301_2 = {s1672[0]};
    Full_Adder FA_2301(s2301, c2301, in2301_1, in2301_2, s1670[0]);
    wire[0:0] s2302, in2302_1, in2302_2;
    wire c2302;
    assign in2302_1 = {s959[0]};
    assign in2302_2 = {c1666};
    Full_Adder FA_2302(s2302, c2302, in2302_1, in2302_2, s958[0]);
    wire[0:0] s2303, in2303_1, in2303_2;
    wire c2303;
    assign in2303_1 = {c1668};
    assign in2303_2 = {c1669};
    Full_Adder FA_2303(s2303, c2303, in2303_1, in2303_2, c1667);
    wire[0:0] s2304, in2304_1, in2304_2;
    wire c2304;
    assign in2304_1 = {c1671};
    assign in2304_2 = {c1672};
    Full_Adder FA_2304(s2304, c2304, in2304_1, in2304_2, c1670);
    wire[0:0] s2305, in2305_1, in2305_2;
    wire c2305;
    assign in2305_1 = {c1674};
    assign in2305_2 = {s1675[0]};
    Full_Adder FA_2305(s2305, c2305, in2305_1, in2305_2, c1673);
    wire[0:0] s2306, in2306_1, in2306_2;
    wire c2306;
    assign in2306_1 = {s1677[0]};
    assign in2306_2 = {s1678[0]};
    Full_Adder FA_2306(s2306, c2306, in2306_1, in2306_2, s1676[0]);
    wire[0:0] s2307, in2307_1, in2307_2;
    wire c2307;
    assign in2307_1 = {s1680[0]};
    assign in2307_2 = {s1681[0]};
    Full_Adder FA_2307(s2307, c2307, in2307_1, in2307_2, s1679[0]);
    wire[0:0] s2308, in2308_1, in2308_2;
    wire c2308;
    assign in2308_1 = {s973[0]};
    assign in2308_2 = {c1675};
    Full_Adder FA_2308(s2308, c2308, in2308_1, in2308_2, s972[0]);
    wire[0:0] s2309, in2309_1, in2309_2;
    wire c2309;
    assign in2309_1 = {c1677};
    assign in2309_2 = {c1678};
    Full_Adder FA_2309(s2309, c2309, in2309_1, in2309_2, c1676);
    wire[0:0] s2310, in2310_1, in2310_2;
    wire c2310;
    assign in2310_1 = {c1680};
    assign in2310_2 = {c1681};
    Full_Adder FA_2310(s2310, c2310, in2310_1, in2310_2, c1679);
    wire[0:0] s2311, in2311_1, in2311_2;
    wire c2311;
    assign in2311_1 = {c1683};
    assign in2311_2 = {s1684[0]};
    Full_Adder FA_2311(s2311, c2311, in2311_1, in2311_2, c1682);
    wire[0:0] s2312, in2312_1, in2312_2;
    wire c2312;
    assign in2312_1 = {s1686[0]};
    assign in2312_2 = {s1687[0]};
    Full_Adder FA_2312(s2312, c2312, in2312_1, in2312_2, s1685[0]);
    wire[0:0] s2313, in2313_1, in2313_2;
    wire c2313;
    assign in2313_1 = {s1689[0]};
    assign in2313_2 = {s1690[0]};
    Full_Adder FA_2313(s2313, c2313, in2313_1, in2313_2, s1688[0]);
    wire[0:0] s2314, in2314_1, in2314_2;
    wire c2314;
    assign in2314_1 = {s987[0]};
    assign in2314_2 = {c1684};
    Full_Adder FA_2314(s2314, c2314, in2314_1, in2314_2, s986[0]);
    wire[0:0] s2315, in2315_1, in2315_2;
    wire c2315;
    assign in2315_1 = {c1686};
    assign in2315_2 = {c1687};
    Full_Adder FA_2315(s2315, c2315, in2315_1, in2315_2, c1685);
    wire[0:0] s2316, in2316_1, in2316_2;
    wire c2316;
    assign in2316_1 = {c1689};
    assign in2316_2 = {c1690};
    Full_Adder FA_2316(s2316, c2316, in2316_1, in2316_2, c1688);
    wire[0:0] s2317, in2317_1, in2317_2;
    wire c2317;
    assign in2317_1 = {c1692};
    assign in2317_2 = {s1693[0]};
    Full_Adder FA_2317(s2317, c2317, in2317_1, in2317_2, c1691);
    wire[0:0] s2318, in2318_1, in2318_2;
    wire c2318;
    assign in2318_1 = {s1695[0]};
    assign in2318_2 = {s1696[0]};
    Full_Adder FA_2318(s2318, c2318, in2318_1, in2318_2, s1694[0]);
    wire[0:0] s2319, in2319_1, in2319_2;
    wire c2319;
    assign in2319_1 = {s1698[0]};
    assign in2319_2 = {s1699[0]};
    Full_Adder FA_2319(s2319, c2319, in2319_1, in2319_2, s1697[0]);
    wire[0:0] s2320, in2320_1, in2320_2;
    wire c2320;
    assign in2320_1 = {s1001[0]};
    assign in2320_2 = {c1693};
    Full_Adder FA_2320(s2320, c2320, in2320_1, in2320_2, s1000[0]);
    wire[0:0] s2321, in2321_1, in2321_2;
    wire c2321;
    assign in2321_1 = {c1695};
    assign in2321_2 = {c1696};
    Full_Adder FA_2321(s2321, c2321, in2321_1, in2321_2, c1694);
    wire[0:0] s2322, in2322_1, in2322_2;
    wire c2322;
    assign in2322_1 = {c1698};
    assign in2322_2 = {c1699};
    Full_Adder FA_2322(s2322, c2322, in2322_1, in2322_2, c1697);
    wire[0:0] s2323, in2323_1, in2323_2;
    wire c2323;
    assign in2323_1 = {c1701};
    assign in2323_2 = {s1702[0]};
    Full_Adder FA_2323(s2323, c2323, in2323_1, in2323_2, c1700);
    wire[0:0] s2324, in2324_1, in2324_2;
    wire c2324;
    assign in2324_1 = {s1704[0]};
    assign in2324_2 = {s1705[0]};
    Full_Adder FA_2324(s2324, c2324, in2324_1, in2324_2, s1703[0]);
    wire[0:0] s2325, in2325_1, in2325_2;
    wire c2325;
    assign in2325_1 = {s1707[0]};
    assign in2325_2 = {s1708[0]};
    Full_Adder FA_2325(s2325, c2325, in2325_1, in2325_2, s1706[0]);
    wire[0:0] s2326, in2326_1, in2326_2;
    wire c2326;
    assign in2326_1 = {s1015[0]};
    assign in2326_2 = {c1702};
    Full_Adder FA_2326(s2326, c2326, in2326_1, in2326_2, s1014[0]);
    wire[0:0] s2327, in2327_1, in2327_2;
    wire c2327;
    assign in2327_1 = {c1704};
    assign in2327_2 = {c1705};
    Full_Adder FA_2327(s2327, c2327, in2327_1, in2327_2, c1703);
    wire[0:0] s2328, in2328_1, in2328_2;
    wire c2328;
    assign in2328_1 = {c1707};
    assign in2328_2 = {c1708};
    Full_Adder FA_2328(s2328, c2328, in2328_1, in2328_2, c1706);
    wire[0:0] s2329, in2329_1, in2329_2;
    wire c2329;
    assign in2329_1 = {c1710};
    assign in2329_2 = {s1711[0]};
    Full_Adder FA_2329(s2329, c2329, in2329_1, in2329_2, c1709);
    wire[0:0] s2330, in2330_1, in2330_2;
    wire c2330;
    assign in2330_1 = {s1713[0]};
    assign in2330_2 = {s1714[0]};
    Full_Adder FA_2330(s2330, c2330, in2330_1, in2330_2, s1712[0]);
    wire[0:0] s2331, in2331_1, in2331_2;
    wire c2331;
    assign in2331_1 = {s1716[0]};
    assign in2331_2 = {s1717[0]};
    Full_Adder FA_2331(s2331, c2331, in2331_1, in2331_2, s1715[0]);
    wire[0:0] s2332, in2332_1, in2332_2;
    wire c2332;
    assign in2332_1 = {s1029[0]};
    assign in2332_2 = {c1711};
    Full_Adder FA_2332(s2332, c2332, in2332_1, in2332_2, s1028[0]);
    wire[0:0] s2333, in2333_1, in2333_2;
    wire c2333;
    assign in2333_1 = {c1713};
    assign in2333_2 = {c1714};
    Full_Adder FA_2333(s2333, c2333, in2333_1, in2333_2, c1712);
    wire[0:0] s2334, in2334_1, in2334_2;
    wire c2334;
    assign in2334_1 = {c1716};
    assign in2334_2 = {c1717};
    Full_Adder FA_2334(s2334, c2334, in2334_1, in2334_2, c1715);
    wire[0:0] s2335, in2335_1, in2335_2;
    wire c2335;
    assign in2335_1 = {c1719};
    assign in2335_2 = {s1720[0]};
    Full_Adder FA_2335(s2335, c2335, in2335_1, in2335_2, c1718);
    wire[0:0] s2336, in2336_1, in2336_2;
    wire c2336;
    assign in2336_1 = {s1722[0]};
    assign in2336_2 = {s1723[0]};
    Full_Adder FA_2336(s2336, c2336, in2336_1, in2336_2, s1721[0]);
    wire[0:0] s2337, in2337_1, in2337_2;
    wire c2337;
    assign in2337_1 = {s1725[0]};
    assign in2337_2 = {s1726[0]};
    Full_Adder FA_2337(s2337, c2337, in2337_1, in2337_2, s1724[0]);
    wire[0:0] s2338, in2338_1, in2338_2;
    wire c2338;
    assign in2338_1 = {s1043[0]};
    assign in2338_2 = {c1720};
    Full_Adder FA_2338(s2338, c2338, in2338_1, in2338_2, s1042[0]);
    wire[0:0] s2339, in2339_1, in2339_2;
    wire c2339;
    assign in2339_1 = {c1722};
    assign in2339_2 = {c1723};
    Full_Adder FA_2339(s2339, c2339, in2339_1, in2339_2, c1721);
    wire[0:0] s2340, in2340_1, in2340_2;
    wire c2340;
    assign in2340_1 = {c1725};
    assign in2340_2 = {c1726};
    Full_Adder FA_2340(s2340, c2340, in2340_1, in2340_2, c1724);
    wire[0:0] s2341, in2341_1, in2341_2;
    wire c2341;
    assign in2341_1 = {c1728};
    assign in2341_2 = {s1729[0]};
    Full_Adder FA_2341(s2341, c2341, in2341_1, in2341_2, c1727);
    wire[0:0] s2342, in2342_1, in2342_2;
    wire c2342;
    assign in2342_1 = {s1731[0]};
    assign in2342_2 = {s1732[0]};
    Full_Adder FA_2342(s2342, c2342, in2342_1, in2342_2, s1730[0]);
    wire[0:0] s2343, in2343_1, in2343_2;
    wire c2343;
    assign in2343_1 = {s1734[0]};
    assign in2343_2 = {s1735[0]};
    Full_Adder FA_2343(s2343, c2343, in2343_1, in2343_2, s1733[0]);
    wire[0:0] s2344, in2344_1, in2344_2;
    wire c2344;
    assign in2344_1 = {s1057[0]};
    assign in2344_2 = {c1729};
    Full_Adder FA_2344(s2344, c2344, in2344_1, in2344_2, s1056[0]);
    wire[0:0] s2345, in2345_1, in2345_2;
    wire c2345;
    assign in2345_1 = {c1731};
    assign in2345_2 = {c1732};
    Full_Adder FA_2345(s2345, c2345, in2345_1, in2345_2, c1730);
    wire[0:0] s2346, in2346_1, in2346_2;
    wire c2346;
    assign in2346_1 = {c1734};
    assign in2346_2 = {c1735};
    Full_Adder FA_2346(s2346, c2346, in2346_1, in2346_2, c1733);
    wire[0:0] s2347, in2347_1, in2347_2;
    wire c2347;
    assign in2347_1 = {c1737};
    assign in2347_2 = {s1738[0]};
    Full_Adder FA_2347(s2347, c2347, in2347_1, in2347_2, c1736);
    wire[0:0] s2348, in2348_1, in2348_2;
    wire c2348;
    assign in2348_1 = {s1740[0]};
    assign in2348_2 = {s1741[0]};
    Full_Adder FA_2348(s2348, c2348, in2348_1, in2348_2, s1739[0]);
    wire[0:0] s2349, in2349_1, in2349_2;
    wire c2349;
    assign in2349_1 = {s1743[0]};
    assign in2349_2 = {s1744[0]};
    Full_Adder FA_2349(s2349, c2349, in2349_1, in2349_2, s1742[0]);
    wire[0:0] s2350, in2350_1, in2350_2;
    wire c2350;
    assign in2350_1 = {s1071[0]};
    assign in2350_2 = {c1738};
    Full_Adder FA_2350(s2350, c2350, in2350_1, in2350_2, s1070[0]);
    wire[0:0] s2351, in2351_1, in2351_2;
    wire c2351;
    assign in2351_1 = {c1740};
    assign in2351_2 = {c1741};
    Full_Adder FA_2351(s2351, c2351, in2351_1, in2351_2, c1739);
    wire[0:0] s2352, in2352_1, in2352_2;
    wire c2352;
    assign in2352_1 = {c1743};
    assign in2352_2 = {c1744};
    Full_Adder FA_2352(s2352, c2352, in2352_1, in2352_2, c1742);
    wire[0:0] s2353, in2353_1, in2353_2;
    wire c2353;
    assign in2353_1 = {c1746};
    assign in2353_2 = {s1747[0]};
    Full_Adder FA_2353(s2353, c2353, in2353_1, in2353_2, c1745);
    wire[0:0] s2354, in2354_1, in2354_2;
    wire c2354;
    assign in2354_1 = {s1749[0]};
    assign in2354_2 = {s1750[0]};
    Full_Adder FA_2354(s2354, c2354, in2354_1, in2354_2, s1748[0]);
    wire[0:0] s2355, in2355_1, in2355_2;
    wire c2355;
    assign in2355_1 = {s1752[0]};
    assign in2355_2 = {s1753[0]};
    Full_Adder FA_2355(s2355, c2355, in2355_1, in2355_2, s1751[0]);
    wire[0:0] s2356, in2356_1, in2356_2;
    wire c2356;
    assign in2356_1 = {s1085[0]};
    assign in2356_2 = {c1747};
    Full_Adder FA_2356(s2356, c2356, in2356_1, in2356_2, s1084[0]);
    wire[0:0] s2357, in2357_1, in2357_2;
    wire c2357;
    assign in2357_1 = {c1749};
    assign in2357_2 = {c1750};
    Full_Adder FA_2357(s2357, c2357, in2357_1, in2357_2, c1748);
    wire[0:0] s2358, in2358_1, in2358_2;
    wire c2358;
    assign in2358_1 = {c1752};
    assign in2358_2 = {c1753};
    Full_Adder FA_2358(s2358, c2358, in2358_1, in2358_2, c1751);
    wire[0:0] s2359, in2359_1, in2359_2;
    wire c2359;
    assign in2359_1 = {c1755};
    assign in2359_2 = {s1756[0]};
    Full_Adder FA_2359(s2359, c2359, in2359_1, in2359_2, c1754);
    wire[0:0] s2360, in2360_1, in2360_2;
    wire c2360;
    assign in2360_1 = {s1758[0]};
    assign in2360_2 = {s1759[0]};
    Full_Adder FA_2360(s2360, c2360, in2360_1, in2360_2, s1757[0]);
    wire[0:0] s2361, in2361_1, in2361_2;
    wire c2361;
    assign in2361_1 = {s1761[0]};
    assign in2361_2 = {s1762[0]};
    Full_Adder FA_2361(s2361, c2361, in2361_1, in2361_2, s1760[0]);
    wire[0:0] s2362, in2362_1, in2362_2;
    wire c2362;
    assign in2362_1 = {s1099[0]};
    assign in2362_2 = {c1756};
    Full_Adder FA_2362(s2362, c2362, in2362_1, in2362_2, s1098[0]);
    wire[0:0] s2363, in2363_1, in2363_2;
    wire c2363;
    assign in2363_1 = {c1758};
    assign in2363_2 = {c1759};
    Full_Adder FA_2363(s2363, c2363, in2363_1, in2363_2, c1757);
    wire[0:0] s2364, in2364_1, in2364_2;
    wire c2364;
    assign in2364_1 = {c1761};
    assign in2364_2 = {c1762};
    Full_Adder FA_2364(s2364, c2364, in2364_1, in2364_2, c1760);
    wire[0:0] s2365, in2365_1, in2365_2;
    wire c2365;
    assign in2365_1 = {c1764};
    assign in2365_2 = {s1765[0]};
    Full_Adder FA_2365(s2365, c2365, in2365_1, in2365_2, c1763);
    wire[0:0] s2366, in2366_1, in2366_2;
    wire c2366;
    assign in2366_1 = {s1767[0]};
    assign in2366_2 = {s1768[0]};
    Full_Adder FA_2366(s2366, c2366, in2366_1, in2366_2, s1766[0]);
    wire[0:0] s2367, in2367_1, in2367_2;
    wire c2367;
    assign in2367_1 = {s1770[0]};
    assign in2367_2 = {s1771[0]};
    Full_Adder FA_2367(s2367, c2367, in2367_1, in2367_2, s1769[0]);
    wire[0:0] s2368, in2368_1, in2368_2;
    wire c2368;
    assign in2368_1 = {s1113[0]};
    assign in2368_2 = {c1765};
    Full_Adder FA_2368(s2368, c2368, in2368_1, in2368_2, s1112[0]);
    wire[0:0] s2369, in2369_1, in2369_2;
    wire c2369;
    assign in2369_1 = {c1767};
    assign in2369_2 = {c1768};
    Full_Adder FA_2369(s2369, c2369, in2369_1, in2369_2, c1766);
    wire[0:0] s2370, in2370_1, in2370_2;
    wire c2370;
    assign in2370_1 = {c1770};
    assign in2370_2 = {c1771};
    Full_Adder FA_2370(s2370, c2370, in2370_1, in2370_2, c1769);
    wire[0:0] s2371, in2371_1, in2371_2;
    wire c2371;
    assign in2371_1 = {c1773};
    assign in2371_2 = {s1774[0]};
    Full_Adder FA_2371(s2371, c2371, in2371_1, in2371_2, c1772);
    wire[0:0] s2372, in2372_1, in2372_2;
    wire c2372;
    assign in2372_1 = {s1776[0]};
    assign in2372_2 = {s1777[0]};
    Full_Adder FA_2372(s2372, c2372, in2372_1, in2372_2, s1775[0]);
    wire[0:0] s2373, in2373_1, in2373_2;
    wire c2373;
    assign in2373_1 = {s1779[0]};
    assign in2373_2 = {s1780[0]};
    Full_Adder FA_2373(s2373, c2373, in2373_1, in2373_2, s1778[0]);
    wire[0:0] s2374, in2374_1, in2374_2;
    wire c2374;
    assign in2374_1 = {s1127[0]};
    assign in2374_2 = {c1774};
    Full_Adder FA_2374(s2374, c2374, in2374_1, in2374_2, s1126[0]);
    wire[0:0] s2375, in2375_1, in2375_2;
    wire c2375;
    assign in2375_1 = {c1776};
    assign in2375_2 = {c1777};
    Full_Adder FA_2375(s2375, c2375, in2375_1, in2375_2, c1775);
    wire[0:0] s2376, in2376_1, in2376_2;
    wire c2376;
    assign in2376_1 = {c1779};
    assign in2376_2 = {c1780};
    Full_Adder FA_2376(s2376, c2376, in2376_1, in2376_2, c1778);
    wire[0:0] s2377, in2377_1, in2377_2;
    wire c2377;
    assign in2377_1 = {c1782};
    assign in2377_2 = {s1783[0]};
    Full_Adder FA_2377(s2377, c2377, in2377_1, in2377_2, c1781);
    wire[0:0] s2378, in2378_1, in2378_2;
    wire c2378;
    assign in2378_1 = {s1785[0]};
    assign in2378_2 = {s1786[0]};
    Full_Adder FA_2378(s2378, c2378, in2378_1, in2378_2, s1784[0]);
    wire[0:0] s2379, in2379_1, in2379_2;
    wire c2379;
    assign in2379_1 = {s1788[0]};
    assign in2379_2 = {s1789[0]};
    Full_Adder FA_2379(s2379, c2379, in2379_1, in2379_2, s1787[0]);
    wire[0:0] s2380, in2380_1, in2380_2;
    wire c2380;
    assign in2380_1 = {s1141[0]};
    assign in2380_2 = {c1783};
    Full_Adder FA_2380(s2380, c2380, in2380_1, in2380_2, s1140[0]);
    wire[0:0] s2381, in2381_1, in2381_2;
    wire c2381;
    assign in2381_1 = {c1785};
    assign in2381_2 = {c1786};
    Full_Adder FA_2381(s2381, c2381, in2381_1, in2381_2, c1784);
    wire[0:0] s2382, in2382_1, in2382_2;
    wire c2382;
    assign in2382_1 = {c1788};
    assign in2382_2 = {c1789};
    Full_Adder FA_2382(s2382, c2382, in2382_1, in2382_2, c1787);
    wire[0:0] s2383, in2383_1, in2383_2;
    wire c2383;
    assign in2383_1 = {c1791};
    assign in2383_2 = {s1792[0]};
    Full_Adder FA_2383(s2383, c2383, in2383_1, in2383_2, c1790);
    wire[0:0] s2384, in2384_1, in2384_2;
    wire c2384;
    assign in2384_1 = {s1794[0]};
    assign in2384_2 = {s1795[0]};
    Full_Adder FA_2384(s2384, c2384, in2384_1, in2384_2, s1793[0]);
    wire[0:0] s2385, in2385_1, in2385_2;
    wire c2385;
    assign in2385_1 = {s1797[0]};
    assign in2385_2 = {s1798[0]};
    Full_Adder FA_2385(s2385, c2385, in2385_1, in2385_2, s1796[0]);
    wire[0:0] s2386, in2386_1, in2386_2;
    wire c2386;
    assign in2386_1 = {s1155[0]};
    assign in2386_2 = {c1792};
    Full_Adder FA_2386(s2386, c2386, in2386_1, in2386_2, s1154[0]);
    wire[0:0] s2387, in2387_1, in2387_2;
    wire c2387;
    assign in2387_1 = {c1794};
    assign in2387_2 = {c1795};
    Full_Adder FA_2387(s2387, c2387, in2387_1, in2387_2, c1793);
    wire[0:0] s2388, in2388_1, in2388_2;
    wire c2388;
    assign in2388_1 = {c1797};
    assign in2388_2 = {c1798};
    Full_Adder FA_2388(s2388, c2388, in2388_1, in2388_2, c1796);
    wire[0:0] s2389, in2389_1, in2389_2;
    wire c2389;
    assign in2389_1 = {c1800};
    assign in2389_2 = {s1801[0]};
    Full_Adder FA_2389(s2389, c2389, in2389_1, in2389_2, c1799);
    wire[0:0] s2390, in2390_1, in2390_2;
    wire c2390;
    assign in2390_1 = {s1803[0]};
    assign in2390_2 = {s1804[0]};
    Full_Adder FA_2390(s2390, c2390, in2390_1, in2390_2, s1802[0]);
    wire[0:0] s2391, in2391_1, in2391_2;
    wire c2391;
    assign in2391_1 = {s1806[0]};
    assign in2391_2 = {s1807[0]};
    Full_Adder FA_2391(s2391, c2391, in2391_1, in2391_2, s1805[0]);
    wire[0:0] s2392, in2392_1, in2392_2;
    wire c2392;
    assign in2392_1 = {s1169[0]};
    assign in2392_2 = {c1801};
    Full_Adder FA_2392(s2392, c2392, in2392_1, in2392_2, s1168[0]);
    wire[0:0] s2393, in2393_1, in2393_2;
    wire c2393;
    assign in2393_1 = {c1803};
    assign in2393_2 = {c1804};
    Full_Adder FA_2393(s2393, c2393, in2393_1, in2393_2, c1802);
    wire[0:0] s2394, in2394_1, in2394_2;
    wire c2394;
    assign in2394_1 = {c1806};
    assign in2394_2 = {c1807};
    Full_Adder FA_2394(s2394, c2394, in2394_1, in2394_2, c1805);
    wire[0:0] s2395, in2395_1, in2395_2;
    wire c2395;
    assign in2395_1 = {c1809};
    assign in2395_2 = {s1810[0]};
    Full_Adder FA_2395(s2395, c2395, in2395_1, in2395_2, c1808);
    wire[0:0] s2396, in2396_1, in2396_2;
    wire c2396;
    assign in2396_1 = {s1812[0]};
    assign in2396_2 = {s1813[0]};
    Full_Adder FA_2396(s2396, c2396, in2396_1, in2396_2, s1811[0]);
    wire[0:0] s2397, in2397_1, in2397_2;
    wire c2397;
    assign in2397_1 = {s1815[0]};
    assign in2397_2 = {s1816[0]};
    Full_Adder FA_2397(s2397, c2397, in2397_1, in2397_2, s1814[0]);
    wire[0:0] s2398, in2398_1, in2398_2;
    wire c2398;
    assign in2398_1 = {s1182[0]};
    assign in2398_2 = {c1810};
    Full_Adder FA_2398(s2398, c2398, in2398_1, in2398_2, s1181[0]);
    wire[0:0] s2399, in2399_1, in2399_2;
    wire c2399;
    assign in2399_1 = {c1812};
    assign in2399_2 = {c1813};
    Full_Adder FA_2399(s2399, c2399, in2399_1, in2399_2, c1811);
    wire[0:0] s2400, in2400_1, in2400_2;
    wire c2400;
    assign in2400_1 = {c1815};
    assign in2400_2 = {c1816};
    Full_Adder FA_2400(s2400, c2400, in2400_1, in2400_2, c1814);
    wire[0:0] s2401, in2401_1, in2401_2;
    wire c2401;
    assign in2401_1 = {c1818};
    assign in2401_2 = {s1819[0]};
    Full_Adder FA_2401(s2401, c2401, in2401_1, in2401_2, c1817);
    wire[0:0] s2402, in2402_1, in2402_2;
    wire c2402;
    assign in2402_1 = {s1821[0]};
    assign in2402_2 = {s1822[0]};
    Full_Adder FA_2402(s2402, c2402, in2402_1, in2402_2, s1820[0]);
    wire[0:0] s2403, in2403_1, in2403_2;
    wire c2403;
    assign in2403_1 = {s1824[0]};
    assign in2403_2 = {s1825[0]};
    Full_Adder FA_2403(s2403, c2403, in2403_1, in2403_2, s1823[0]);
    wire[0:0] s2404, in2404_1, in2404_2;
    wire c2404;
    assign in2404_1 = {s1194[0]};
    assign in2404_2 = {c1819};
    Full_Adder FA_2404(s2404, c2404, in2404_1, in2404_2, s1193[0]);
    wire[0:0] s2405, in2405_1, in2405_2;
    wire c2405;
    assign in2405_1 = {c1821};
    assign in2405_2 = {c1822};
    Full_Adder FA_2405(s2405, c2405, in2405_1, in2405_2, c1820);
    wire[0:0] s2406, in2406_1, in2406_2;
    wire c2406;
    assign in2406_1 = {c1824};
    assign in2406_2 = {c1825};
    Full_Adder FA_2406(s2406, c2406, in2406_1, in2406_2, c1823);
    wire[0:0] s2407, in2407_1, in2407_2;
    wire c2407;
    assign in2407_1 = {c1827};
    assign in2407_2 = {s1828[0]};
    Full_Adder FA_2407(s2407, c2407, in2407_1, in2407_2, c1826);
    wire[0:0] s2408, in2408_1, in2408_2;
    wire c2408;
    assign in2408_1 = {s1830[0]};
    assign in2408_2 = {s1831[0]};
    Full_Adder FA_2408(s2408, c2408, in2408_1, in2408_2, s1829[0]);
    wire[0:0] s2409, in2409_1, in2409_2;
    wire c2409;
    assign in2409_1 = {s1833[0]};
    assign in2409_2 = {s1834[0]};
    Full_Adder FA_2409(s2409, c2409, in2409_1, in2409_2, s1832[0]);
    wire[0:0] s2410, in2410_1, in2410_2;
    wire c2410;
    assign in2410_1 = {s1205[0]};
    assign in2410_2 = {c1828};
    Full_Adder FA_2410(s2410, c2410, in2410_1, in2410_2, s1204[0]);
    wire[0:0] s2411, in2411_1, in2411_2;
    wire c2411;
    assign in2411_1 = {c1830};
    assign in2411_2 = {c1831};
    Full_Adder FA_2411(s2411, c2411, in2411_1, in2411_2, c1829);
    wire[0:0] s2412, in2412_1, in2412_2;
    wire c2412;
    assign in2412_1 = {c1833};
    assign in2412_2 = {c1834};
    Full_Adder FA_2412(s2412, c2412, in2412_1, in2412_2, c1832);
    wire[0:0] s2413, in2413_1, in2413_2;
    wire c2413;
    assign in2413_1 = {c1836};
    assign in2413_2 = {s1837[0]};
    Full_Adder FA_2413(s2413, c2413, in2413_1, in2413_2, c1835);
    wire[0:0] s2414, in2414_1, in2414_2;
    wire c2414;
    assign in2414_1 = {s1839[0]};
    assign in2414_2 = {s1840[0]};
    Full_Adder FA_2414(s2414, c2414, in2414_1, in2414_2, s1838[0]);
    wire[0:0] s2415, in2415_1, in2415_2;
    wire c2415;
    assign in2415_1 = {s1842[0]};
    assign in2415_2 = {s1843[0]};
    Full_Adder FA_2415(s2415, c2415, in2415_1, in2415_2, s1841[0]);
    wire[0:0] s2416, in2416_1, in2416_2;
    wire c2416;
    assign in2416_1 = {s1215[0]};
    assign in2416_2 = {c1837};
    Full_Adder FA_2416(s2416, c2416, in2416_1, in2416_2, s1214[0]);
    wire[0:0] s2417, in2417_1, in2417_2;
    wire c2417;
    assign in2417_1 = {c1839};
    assign in2417_2 = {c1840};
    Full_Adder FA_2417(s2417, c2417, in2417_1, in2417_2, c1838);
    wire[0:0] s2418, in2418_1, in2418_2;
    wire c2418;
    assign in2418_1 = {c1842};
    assign in2418_2 = {c1843};
    Full_Adder FA_2418(s2418, c2418, in2418_1, in2418_2, c1841);
    wire[0:0] s2419, in2419_1, in2419_2;
    wire c2419;
    assign in2419_1 = {c1845};
    assign in2419_2 = {s1846[0]};
    Full_Adder FA_2419(s2419, c2419, in2419_1, in2419_2, c1844);
    wire[0:0] s2420, in2420_1, in2420_2;
    wire c2420;
    assign in2420_1 = {s1848[0]};
    assign in2420_2 = {s1849[0]};
    Full_Adder FA_2420(s2420, c2420, in2420_1, in2420_2, s1847[0]);
    wire[0:0] s2421, in2421_1, in2421_2;
    wire c2421;
    assign in2421_1 = {s1851[0]};
    assign in2421_2 = {s1852[0]};
    Full_Adder FA_2421(s2421, c2421, in2421_1, in2421_2, s1850[0]);
    wire[0:0] s2422, in2422_1, in2422_2;
    wire c2422;
    assign in2422_1 = {s1224[0]};
    assign in2422_2 = {c1846};
    Full_Adder FA_2422(s2422, c2422, in2422_1, in2422_2, s1223[0]);
    wire[0:0] s2423, in2423_1, in2423_2;
    wire c2423;
    assign in2423_1 = {c1848};
    assign in2423_2 = {c1849};
    Full_Adder FA_2423(s2423, c2423, in2423_1, in2423_2, c1847);
    wire[0:0] s2424, in2424_1, in2424_2;
    wire c2424;
    assign in2424_1 = {c1851};
    assign in2424_2 = {c1852};
    Full_Adder FA_2424(s2424, c2424, in2424_1, in2424_2, c1850);
    wire[0:0] s2425, in2425_1, in2425_2;
    wire c2425;
    assign in2425_1 = {c1854};
    assign in2425_2 = {s1855[0]};
    Full_Adder FA_2425(s2425, c2425, in2425_1, in2425_2, c1853);
    wire[0:0] s2426, in2426_1, in2426_2;
    wire c2426;
    assign in2426_1 = {s1857[0]};
    assign in2426_2 = {s1858[0]};
    Full_Adder FA_2426(s2426, c2426, in2426_1, in2426_2, s1856[0]);
    wire[0:0] s2427, in2427_1, in2427_2;
    wire c2427;
    assign in2427_1 = {s1860[0]};
    assign in2427_2 = {s1861[0]};
    Full_Adder FA_2427(s2427, c2427, in2427_1, in2427_2, s1859[0]);
    wire[0:0] s2428, in2428_1, in2428_2;
    wire c2428;
    assign in2428_1 = {s1232[0]};
    assign in2428_2 = {c1855};
    Full_Adder FA_2428(s2428, c2428, in2428_1, in2428_2, s1231[0]);
    wire[0:0] s2429, in2429_1, in2429_2;
    wire c2429;
    assign in2429_1 = {c1857};
    assign in2429_2 = {c1858};
    Full_Adder FA_2429(s2429, c2429, in2429_1, in2429_2, c1856);
    wire[0:0] s2430, in2430_1, in2430_2;
    wire c2430;
    assign in2430_1 = {c1860};
    assign in2430_2 = {c1861};
    Full_Adder FA_2430(s2430, c2430, in2430_1, in2430_2, c1859);
    wire[0:0] s2431, in2431_1, in2431_2;
    wire c2431;
    assign in2431_1 = {c1863};
    assign in2431_2 = {s1864[0]};
    Full_Adder FA_2431(s2431, c2431, in2431_1, in2431_2, c1862);
    wire[0:0] s2432, in2432_1, in2432_2;
    wire c2432;
    assign in2432_1 = {s1866[0]};
    assign in2432_2 = {s1867[0]};
    Full_Adder FA_2432(s2432, c2432, in2432_1, in2432_2, s1865[0]);
    wire[0:0] s2433, in2433_1, in2433_2;
    wire c2433;
    assign in2433_1 = {s1869[0]};
    assign in2433_2 = {s1870[0]};
    Full_Adder FA_2433(s2433, c2433, in2433_1, in2433_2, s1868[0]);
    wire[0:0] s2434, in2434_1, in2434_2;
    wire c2434;
    assign in2434_1 = {s1239[0]};
    assign in2434_2 = {c1864};
    Full_Adder FA_2434(s2434, c2434, in2434_1, in2434_2, s1238[0]);
    wire[0:0] s2435, in2435_1, in2435_2;
    wire c2435;
    assign in2435_1 = {c1866};
    assign in2435_2 = {c1867};
    Full_Adder FA_2435(s2435, c2435, in2435_1, in2435_2, c1865);
    wire[0:0] s2436, in2436_1, in2436_2;
    wire c2436;
    assign in2436_1 = {c1869};
    assign in2436_2 = {c1870};
    Full_Adder FA_2436(s2436, c2436, in2436_1, in2436_2, c1868);
    wire[0:0] s2437, in2437_1, in2437_2;
    wire c2437;
    assign in2437_1 = {c1872};
    assign in2437_2 = {s1873[0]};
    Full_Adder FA_2437(s2437, c2437, in2437_1, in2437_2, c1871);
    wire[0:0] s2438, in2438_1, in2438_2;
    wire c2438;
    assign in2438_1 = {s1875[0]};
    assign in2438_2 = {s1876[0]};
    Full_Adder FA_2438(s2438, c2438, in2438_1, in2438_2, s1874[0]);
    wire[0:0] s2439, in2439_1, in2439_2;
    wire c2439;
    assign in2439_1 = {s1878[0]};
    assign in2439_2 = {s1879[0]};
    Full_Adder FA_2439(s2439, c2439, in2439_1, in2439_2, s1877[0]);
    wire[0:0] s2440, in2440_1, in2440_2;
    wire c2440;
    assign in2440_1 = {s1245[0]};
    assign in2440_2 = {c1873};
    Full_Adder FA_2440(s2440, c2440, in2440_1, in2440_2, s1244[0]);
    wire[0:0] s2441, in2441_1, in2441_2;
    wire c2441;
    assign in2441_1 = {c1875};
    assign in2441_2 = {c1876};
    Full_Adder FA_2441(s2441, c2441, in2441_1, in2441_2, c1874);
    wire[0:0] s2442, in2442_1, in2442_2;
    wire c2442;
    assign in2442_1 = {c1878};
    assign in2442_2 = {c1879};
    Full_Adder FA_2442(s2442, c2442, in2442_1, in2442_2, c1877);
    wire[0:0] s2443, in2443_1, in2443_2;
    wire c2443;
    assign in2443_1 = {c1881};
    assign in2443_2 = {s1882[0]};
    Full_Adder FA_2443(s2443, c2443, in2443_1, in2443_2, c1880);
    wire[0:0] s2444, in2444_1, in2444_2;
    wire c2444;
    assign in2444_1 = {s1884[0]};
    assign in2444_2 = {s1885[0]};
    Full_Adder FA_2444(s2444, c2444, in2444_1, in2444_2, s1883[0]);
    wire[0:0] s2445, in2445_1, in2445_2;
    wire c2445;
    assign in2445_1 = {s1887[0]};
    assign in2445_2 = {s1888[0]};
    Full_Adder FA_2445(s2445, c2445, in2445_1, in2445_2, s1886[0]);
    wire[0:0] s2446, in2446_1, in2446_2;
    wire c2446;
    assign in2446_1 = {s1250[0]};
    assign in2446_2 = {c1882};
    Full_Adder FA_2446(s2446, c2446, in2446_1, in2446_2, s1249[0]);
    wire[0:0] s2447, in2447_1, in2447_2;
    wire c2447;
    assign in2447_1 = {c1884};
    assign in2447_2 = {c1885};
    Full_Adder FA_2447(s2447, c2447, in2447_1, in2447_2, c1883);
    wire[0:0] s2448, in2448_1, in2448_2;
    wire c2448;
    assign in2448_1 = {c1887};
    assign in2448_2 = {c1888};
    Full_Adder FA_2448(s2448, c2448, in2448_1, in2448_2, c1886);
    wire[0:0] s2449, in2449_1, in2449_2;
    wire c2449;
    assign in2449_1 = {c1890};
    assign in2449_2 = {s1891[0]};
    Full_Adder FA_2449(s2449, c2449, in2449_1, in2449_2, c1889);
    wire[0:0] s2450, in2450_1, in2450_2;
    wire c2450;
    assign in2450_1 = {s1893[0]};
    assign in2450_2 = {s1894[0]};
    Full_Adder FA_2450(s2450, c2450, in2450_1, in2450_2, s1892[0]);
    wire[0:0] s2451, in2451_1, in2451_2;
    wire c2451;
    assign in2451_1 = {s1896[0]};
    assign in2451_2 = {s1897[0]};
    Full_Adder FA_2451(s2451, c2451, in2451_1, in2451_2, s1895[0]);
    wire[0:0] s2452, in2452_1, in2452_2;
    wire c2452;
    assign in2452_1 = {s1254[0]};
    assign in2452_2 = {c1891};
    Full_Adder FA_2452(s2452, c2452, in2452_1, in2452_2, s1253[0]);
    wire[0:0] s2453, in2453_1, in2453_2;
    wire c2453;
    assign in2453_1 = {c1893};
    assign in2453_2 = {c1894};
    Full_Adder FA_2453(s2453, c2453, in2453_1, in2453_2, c1892);
    wire[0:0] s2454, in2454_1, in2454_2;
    wire c2454;
    assign in2454_1 = {c1896};
    assign in2454_2 = {c1897};
    Full_Adder FA_2454(s2454, c2454, in2454_1, in2454_2, c1895);
    wire[0:0] s2455, in2455_1, in2455_2;
    wire c2455;
    assign in2455_1 = {c1899};
    assign in2455_2 = {s1900[0]};
    Full_Adder FA_2455(s2455, c2455, in2455_1, in2455_2, c1898);
    wire[0:0] s2456, in2456_1, in2456_2;
    wire c2456;
    assign in2456_1 = {s1902[0]};
    assign in2456_2 = {s1903[0]};
    Full_Adder FA_2456(s2456, c2456, in2456_1, in2456_2, s1901[0]);
    wire[0:0] s2457, in2457_1, in2457_2;
    wire c2457;
    assign in2457_1 = {s1905[0]};
    assign in2457_2 = {s1906[0]};
    Full_Adder FA_2457(s2457, c2457, in2457_1, in2457_2, s1904[0]);
    wire[0:0] s2458, in2458_1, in2458_2;
    wire c2458;
    assign in2458_1 = {s1257[0]};
    assign in2458_2 = {c1900};
    Full_Adder FA_2458(s2458, c2458, in2458_1, in2458_2, s1256[0]);
    wire[0:0] s2459, in2459_1, in2459_2;
    wire c2459;
    assign in2459_1 = {c1902};
    assign in2459_2 = {c1903};
    Full_Adder FA_2459(s2459, c2459, in2459_1, in2459_2, c1901);
    wire[0:0] s2460, in2460_1, in2460_2;
    wire c2460;
    assign in2460_1 = {c1905};
    assign in2460_2 = {c1906};
    Full_Adder FA_2460(s2460, c2460, in2460_1, in2460_2, c1904);
    wire[0:0] s2461, in2461_1, in2461_2;
    wire c2461;
    assign in2461_1 = {c1908};
    assign in2461_2 = {s1909[0]};
    Full_Adder FA_2461(s2461, c2461, in2461_1, in2461_2, c1907);
    wire[0:0] s2462, in2462_1, in2462_2;
    wire c2462;
    assign in2462_1 = {s1911[0]};
    assign in2462_2 = {s1912[0]};
    Full_Adder FA_2462(s2462, c2462, in2462_1, in2462_2, s1910[0]);
    wire[0:0] s2463, in2463_1, in2463_2;
    wire c2463;
    assign in2463_1 = {s1914[0]};
    assign in2463_2 = {s1915[0]};
    Full_Adder FA_2463(s2463, c2463, in2463_1, in2463_2, s1913[0]);
    wire[0:0] s2464, in2464_1, in2464_2;
    wire c2464;
    assign in2464_1 = {s1259[0]};
    assign in2464_2 = {c1909};
    Full_Adder FA_2464(s2464, c2464, in2464_1, in2464_2, s1258[0]);
    wire[0:0] s2465, in2465_1, in2465_2;
    wire c2465;
    assign in2465_1 = {c1911};
    assign in2465_2 = {c1912};
    Full_Adder FA_2465(s2465, c2465, in2465_1, in2465_2, c1910);
    wire[0:0] s2466, in2466_1, in2466_2;
    wire c2466;
    assign in2466_1 = {c1914};
    assign in2466_2 = {c1915};
    Full_Adder FA_2466(s2466, c2466, in2466_1, in2466_2, c1913);
    wire[0:0] s2467, in2467_1, in2467_2;
    wire c2467;
    assign in2467_1 = {c1917};
    assign in2467_2 = {s1918[0]};
    Full_Adder FA_2467(s2467, c2467, in2467_1, in2467_2, c1916);
    wire[0:0] s2468, in2468_1, in2468_2;
    wire c2468;
    assign in2468_1 = {s1920[0]};
    assign in2468_2 = {s1921[0]};
    Full_Adder FA_2468(s2468, c2468, in2468_1, in2468_2, s1919[0]);
    wire[0:0] s2469, in2469_1, in2469_2;
    wire c2469;
    assign in2469_1 = {s1923[0]};
    assign in2469_2 = {s1924[0]};
    Full_Adder FA_2469(s2469, c2469, in2469_1, in2469_2, s1922[0]);
    wire[0:0] s2470, in2470_1, in2470_2;
    wire c2470;
    assign in2470_1 = {s1260[0]};
    assign in2470_2 = {c1918};
    Full_Adder FA_2470(s2470, c2470, in2470_1, in2470_2, c1259);
    wire[0:0] s2471, in2471_1, in2471_2;
    wire c2471;
    assign in2471_1 = {c1920};
    assign in2471_2 = {c1921};
    Full_Adder FA_2471(s2471, c2471, in2471_1, in2471_2, c1919);
    wire[0:0] s2472, in2472_1, in2472_2;
    wire c2472;
    assign in2472_1 = {c1923};
    assign in2472_2 = {c1924};
    Full_Adder FA_2472(s2472, c2472, in2472_1, in2472_2, c1922);
    wire[0:0] s2473, in2473_1, in2473_2;
    wire c2473;
    assign in2473_1 = {c1926};
    assign in2473_2 = {s1927[0]};
    Full_Adder FA_2473(s2473, c2473, in2473_1, in2473_2, c1925);
    wire[0:0] s2474, in2474_1, in2474_2;
    wire c2474;
    assign in2474_1 = {s1929[0]};
    assign in2474_2 = {s1930[0]};
    Full_Adder FA_2474(s2474, c2474, in2474_1, in2474_2, s1928[0]);
    wire[0:0] s2475, in2475_1, in2475_2;
    wire c2475;
    assign in2475_1 = {s1932[0]};
    assign in2475_2 = {s1933[0]};
    Full_Adder FA_2475(s2475, c2475, in2475_1, in2475_2, s1931[0]);
    wire[0:0] s2476, in2476_1, in2476_2;
    wire c2476;
    assign in2476_1 = {c1260};
    assign in2476_2 = {c1927};
    Full_Adder FA_2476(s2476, c2476, in2476_1, in2476_2, pp63[36]);
    wire[0:0] s2477, in2477_1, in2477_2;
    wire c2477;
    assign in2477_1 = {c1929};
    assign in2477_2 = {c1930};
    Full_Adder FA_2477(s2477, c2477, in2477_1, in2477_2, c1928);
    wire[0:0] s2478, in2478_1, in2478_2;
    wire c2478;
    assign in2478_1 = {c1932};
    assign in2478_2 = {c1933};
    Full_Adder FA_2478(s2478, c2478, in2478_1, in2478_2, c1931);
    wire[0:0] s2479, in2479_1, in2479_2;
    wire c2479;
    assign in2479_1 = {c1935};
    assign in2479_2 = {s1936[0]};
    Full_Adder FA_2479(s2479, c2479, in2479_1, in2479_2, c1934);
    wire[0:0] s2480, in2480_1, in2480_2;
    wire c2480;
    assign in2480_1 = {s1938[0]};
    assign in2480_2 = {s1939[0]};
    Full_Adder FA_2480(s2480, c2480, in2480_1, in2480_2, s1937[0]);
    wire[0:0] s2481, in2481_1, in2481_2;
    wire c2481;
    assign in2481_1 = {s1941[0]};
    assign in2481_2 = {s1942[0]};
    Full_Adder FA_2481(s2481, c2481, in2481_1, in2481_2, s1940[0]);
    wire[0:0] s2482, in2482_1, in2482_2;
    wire c2482;
    assign in2482_1 = {pp62[38]};
    assign in2482_2 = {pp63[37]};
    Full_Adder FA_2482(s2482, c2482, in2482_1, in2482_2, pp61[39]);
    wire[0:0] s2483, in2483_1, in2483_2;
    wire c2483;
    assign in2483_1 = {c1937};
    assign in2483_2 = {c1938};
    Full_Adder FA_2483(s2483, c2483, in2483_1, in2483_2, c1936);
    wire[0:0] s2484, in2484_1, in2484_2;
    wire c2484;
    assign in2484_1 = {c1940};
    assign in2484_2 = {c1941};
    Full_Adder FA_2484(s2484, c2484, in2484_1, in2484_2, c1939);
    wire[0:0] s2485, in2485_1, in2485_2;
    wire c2485;
    assign in2485_1 = {c1943};
    assign in2485_2 = {c1944};
    Full_Adder FA_2485(s2485, c2485, in2485_1, in2485_2, c1942);
    wire[0:0] s2486, in2486_1, in2486_2;
    wire c2486;
    assign in2486_1 = {s1946[0]};
    assign in2486_2 = {s1947[0]};
    Full_Adder FA_2486(s2486, c2486, in2486_1, in2486_2, s1945[0]);
    wire[0:0] s2487, in2487_1, in2487_2;
    wire c2487;
    assign in2487_1 = {s1949[0]};
    assign in2487_2 = {s1950[0]};
    Full_Adder FA_2487(s2487, c2487, in2487_1, in2487_2, s1948[0]);
    wire[0:0] s2488, in2488_1, in2488_2;
    wire c2488;
    assign in2488_1 = {pp60[41]};
    assign in2488_2 = {pp61[40]};
    Full_Adder FA_2488(s2488, c2488, in2488_1, in2488_2, pp59[42]);
    wire[0:0] s2489, in2489_1, in2489_2;
    wire c2489;
    assign in2489_1 = {pp63[38]};
    assign in2489_2 = {c1945};
    Full_Adder FA_2489(s2489, c2489, in2489_1, in2489_2, pp62[39]);
    wire[0:0] s2490, in2490_1, in2490_2;
    wire c2490;
    assign in2490_1 = {c1947};
    assign in2490_2 = {c1948};
    Full_Adder FA_2490(s2490, c2490, in2490_1, in2490_2, c1946);
    wire[0:0] s2491, in2491_1, in2491_2;
    wire c2491;
    assign in2491_1 = {c1950};
    assign in2491_2 = {c1951};
    Full_Adder FA_2491(s2491, c2491, in2491_1, in2491_2, c1949);
    wire[0:0] s2492, in2492_1, in2492_2;
    wire c2492;
    assign in2492_1 = {s1953[0]};
    assign in2492_2 = {s1954[0]};
    Full_Adder FA_2492(s2492, c2492, in2492_1, in2492_2, c1952);
    wire[0:0] s2493, in2493_1, in2493_2;
    wire c2493;
    assign in2493_1 = {s1956[0]};
    assign in2493_2 = {s1957[0]};
    Full_Adder FA_2493(s2493, c2493, in2493_1, in2493_2, s1955[0]);
    wire[0:0] s2494, in2494_1, in2494_2;
    wire c2494;
    assign in2494_1 = {pp58[44]};
    assign in2494_2 = {pp59[43]};
    Full_Adder FA_2494(s2494, c2494, in2494_1, in2494_2, pp57[45]);
    wire[0:0] s2495, in2495_1, in2495_2;
    wire c2495;
    assign in2495_1 = {pp61[41]};
    assign in2495_2 = {pp62[40]};
    Full_Adder FA_2495(s2495, c2495, in2495_1, in2495_2, pp60[42]);
    wire[0:0] s2496, in2496_1, in2496_2;
    wire c2496;
    assign in2496_1 = {c1953};
    assign in2496_2 = {c1954};
    Full_Adder FA_2496(s2496, c2496, in2496_1, in2496_2, pp63[39]);
    wire[0:0] s2497, in2497_1, in2497_2;
    wire c2497;
    assign in2497_1 = {c1956};
    assign in2497_2 = {c1957};
    Full_Adder FA_2497(s2497, c2497, in2497_1, in2497_2, c1955);
    wire[0:0] s2498, in2498_1, in2498_2;
    wire c2498;
    assign in2498_1 = {c1959};
    assign in2498_2 = {s1960[0]};
    Full_Adder FA_2498(s2498, c2498, in2498_1, in2498_2, c1958);
    wire[0:0] s2499, in2499_1, in2499_2;
    wire c2499;
    assign in2499_1 = {s1962[0]};
    assign in2499_2 = {s1963[0]};
    Full_Adder FA_2499(s2499, c2499, in2499_1, in2499_2, s1961[0]);
    wire[0:0] s2500, in2500_1, in2500_2;
    wire c2500;
    assign in2500_1 = {pp56[47]};
    assign in2500_2 = {pp57[46]};
    Full_Adder FA_2500(s2500, c2500, in2500_1, in2500_2, pp55[48]);
    wire[0:0] s2501, in2501_1, in2501_2;
    wire c2501;
    assign in2501_1 = {pp59[44]};
    assign in2501_2 = {pp60[43]};
    Full_Adder FA_2501(s2501, c2501, in2501_1, in2501_2, pp58[45]);
    wire[0:0] s2502, in2502_1, in2502_2;
    wire c2502;
    assign in2502_1 = {pp62[41]};
    assign in2502_2 = {pp63[40]};
    Full_Adder FA_2502(s2502, c2502, in2502_1, in2502_2, pp61[42]);
    wire[0:0] s2503, in2503_1, in2503_2;
    wire c2503;
    assign in2503_1 = {c1961};
    assign in2503_2 = {c1962};
    Full_Adder FA_2503(s2503, c2503, in2503_1, in2503_2, c1960);
    wire[0:0] s2504, in2504_1, in2504_2;
    wire c2504;
    assign in2504_1 = {c1964};
    assign in2504_2 = {c1965};
    Full_Adder FA_2504(s2504, c2504, in2504_1, in2504_2, c1963);
    wire[0:0] s2505, in2505_1, in2505_2;
    wire c2505;
    assign in2505_1 = {s1967[0]};
    assign in2505_2 = {s1968[0]};
    Full_Adder FA_2505(s2505, c2505, in2505_1, in2505_2, s1966[0]);
    wire[0:0] s2506, in2506_1, in2506_2;
    wire c2506;
    assign in2506_1 = {pp54[50]};
    assign in2506_2 = {pp55[49]};
    Full_Adder FA_2506(s2506, c2506, in2506_1, in2506_2, pp53[51]);
    wire[0:0] s2507, in2507_1, in2507_2;
    wire c2507;
    assign in2507_1 = {pp57[47]};
    assign in2507_2 = {pp58[46]};
    Full_Adder FA_2507(s2507, c2507, in2507_1, in2507_2, pp56[48]);
    wire[0:0] s2508, in2508_1, in2508_2;
    wire c2508;
    assign in2508_1 = {pp60[44]};
    assign in2508_2 = {pp61[43]};
    Full_Adder FA_2508(s2508, c2508, in2508_1, in2508_2, pp59[45]);
    wire[0:0] s2509, in2509_1, in2509_2;
    wire c2509;
    assign in2509_1 = {pp63[41]};
    assign in2509_2 = {c1966};
    Full_Adder FA_2509(s2509, c2509, in2509_1, in2509_2, pp62[42]);
    wire[0:0] s2510, in2510_1, in2510_2;
    wire c2510;
    assign in2510_1 = {c1968};
    assign in2510_2 = {c1969};
    Full_Adder FA_2510(s2510, c2510, in2510_1, in2510_2, c1967);
    wire[0:0] s2511, in2511_1, in2511_2;
    wire c2511;
    assign in2511_1 = {s1971[0]};
    assign in2511_2 = {s1972[0]};
    Full_Adder FA_2511(s2511, c2511, in2511_1, in2511_2, c1970);
    wire[0:0] s2512, in2512_1, in2512_2;
    wire c2512;
    assign in2512_1 = {pp52[53]};
    assign in2512_2 = {pp53[52]};
    Full_Adder FA_2512(s2512, c2512, in2512_1, in2512_2, pp51[54]);
    wire[0:0] s2513, in2513_1, in2513_2;
    wire c2513;
    assign in2513_1 = {pp55[50]};
    assign in2513_2 = {pp56[49]};
    Full_Adder FA_2513(s2513, c2513, in2513_1, in2513_2, pp54[51]);
    wire[0:0] s2514, in2514_1, in2514_2;
    wire c2514;
    assign in2514_1 = {pp58[47]};
    assign in2514_2 = {pp59[46]};
    Full_Adder FA_2514(s2514, c2514, in2514_1, in2514_2, pp57[48]);
    wire[0:0] s2515, in2515_1, in2515_2;
    wire c2515;
    assign in2515_1 = {pp61[44]};
    assign in2515_2 = {pp62[43]};
    Full_Adder FA_2515(s2515, c2515, in2515_1, in2515_2, pp60[45]);
    wire[0:0] s2516, in2516_1, in2516_2;
    wire c2516;
    assign in2516_1 = {c1971};
    assign in2516_2 = {c1972};
    Full_Adder FA_2516(s2516, c2516, in2516_1, in2516_2, pp63[42]);
    wire[0:0] s2517, in2517_1, in2517_2;
    wire c2517;
    assign in2517_1 = {c1974};
    assign in2517_2 = {s1975[0]};
    Full_Adder FA_2517(s2517, c2517, in2517_1, in2517_2, c1973);
    wire[0:0] s2518, in2518_1, in2518_2;
    wire c2518;
    assign in2518_1 = {pp50[56]};
    assign in2518_2 = {pp51[55]};
    Full_Adder FA_2518(s2518, c2518, in2518_1, in2518_2, pp49[57]);
    wire[0:0] s2519, in2519_1, in2519_2;
    wire c2519;
    assign in2519_1 = {pp53[53]};
    assign in2519_2 = {pp54[52]};
    Full_Adder FA_2519(s2519, c2519, in2519_1, in2519_2, pp52[54]);
    wire[0:0] s2520, in2520_1, in2520_2;
    wire c2520;
    assign in2520_1 = {pp56[50]};
    assign in2520_2 = {pp57[49]};
    Full_Adder FA_2520(s2520, c2520, in2520_1, in2520_2, pp55[51]);
    wire[0:0] s2521, in2521_1, in2521_2;
    wire c2521;
    assign in2521_1 = {pp59[47]};
    assign in2521_2 = {pp60[46]};
    Full_Adder FA_2521(s2521, c2521, in2521_1, in2521_2, pp58[48]);
    wire[0:0] s2522, in2522_1, in2522_2;
    wire c2522;
    assign in2522_1 = {pp62[44]};
    assign in2522_2 = {pp63[43]};
    Full_Adder FA_2522(s2522, c2522, in2522_1, in2522_2, pp61[45]);
    wire[0:0] s2523, in2523_1, in2523_2;
    wire c2523;
    assign in2523_1 = {c1976};
    assign in2523_2 = {c1977};
    Full_Adder FA_2523(s2523, c2523, in2523_1, in2523_2, c1975);
    wire[0:0] s2524, in2524_1, in2524_2;
    wire c2524;
    assign in2524_1 = {pp48[59]};
    assign in2524_2 = {pp49[58]};
    Full_Adder FA_2524(s2524, c2524, in2524_1, in2524_2, pp47[60]);
    wire[0:0] s2525, in2525_1, in2525_2;
    wire c2525;
    assign in2525_1 = {pp51[56]};
    assign in2525_2 = {pp52[55]};
    Full_Adder FA_2525(s2525, c2525, in2525_1, in2525_2, pp50[57]);
    wire[0:0] s2526, in2526_1, in2526_2;
    wire c2526;
    assign in2526_1 = {pp54[53]};
    assign in2526_2 = {pp55[52]};
    Full_Adder FA_2526(s2526, c2526, in2526_1, in2526_2, pp53[54]);
    wire[0:0] s2527, in2527_1, in2527_2;
    wire c2527;
    assign in2527_1 = {pp57[50]};
    assign in2527_2 = {pp58[49]};
    Full_Adder FA_2527(s2527, c2527, in2527_1, in2527_2, pp56[51]);
    wire[0:0] s2528, in2528_1, in2528_2;
    wire c2528;
    assign in2528_1 = {pp60[47]};
    assign in2528_2 = {pp61[46]};
    Full_Adder FA_2528(s2528, c2528, in2528_1, in2528_2, pp59[48]);
    wire[0:0] s2529, in2529_1, in2529_2;
    wire c2529;
    assign in2529_1 = {pp63[44]};
    assign in2529_2 = {c1978};
    Full_Adder FA_2529(s2529, c2529, in2529_1, in2529_2, pp62[45]);
    wire[0:0] s2530, in2530_1, in2530_2;
    wire c2530;
    assign in2530_1 = {pp46[62]};
    assign in2530_2 = {pp47[61]};
    Full_Adder FA_2530(s2530, c2530, in2530_1, in2530_2, pp45[63]);
    wire[0:0] s2531, in2531_1, in2531_2;
    wire c2531;
    assign in2531_1 = {pp49[59]};
    assign in2531_2 = {pp50[58]};
    Full_Adder FA_2531(s2531, c2531, in2531_1, in2531_2, pp48[60]);
    wire[0:0] s2532, in2532_1, in2532_2;
    wire c2532;
    assign in2532_1 = {pp52[56]};
    assign in2532_2 = {pp53[55]};
    Full_Adder FA_2532(s2532, c2532, in2532_1, in2532_2, pp51[57]);
    wire[0:0] s2533, in2533_1, in2533_2;
    wire c2533;
    assign in2533_1 = {pp55[53]};
    assign in2533_2 = {pp56[52]};
    Full_Adder FA_2533(s2533, c2533, in2533_1, in2533_2, pp54[54]);
    wire[0:0] s2534, in2534_1, in2534_2;
    wire c2534;
    assign in2534_1 = {pp58[50]};
    assign in2534_2 = {pp59[49]};
    Full_Adder FA_2534(s2534, c2534, in2534_1, in2534_2, pp57[51]);
    wire[0:0] s2535, in2535_1, in2535_2;
    wire c2535;
    assign in2535_1 = {pp61[47]};
    assign in2535_2 = {pp62[46]};
    Full_Adder FA_2535(s2535, c2535, in2535_1, in2535_2, pp60[48]);
    wire[0:0] s2536, in2536_1, in2536_2;
    wire c2536;
    assign in2536_1 = {pp47[62]};
    assign in2536_2 = {pp48[61]};
    Full_Adder FA_2536(s2536, c2536, in2536_1, in2536_2, pp46[63]);
    wire[0:0] s2537, in2537_1, in2537_2;
    wire c2537;
    assign in2537_1 = {pp50[59]};
    assign in2537_2 = {pp51[58]};
    Full_Adder FA_2537(s2537, c2537, in2537_1, in2537_2, pp49[60]);
    wire[0:0] s2538, in2538_1, in2538_2;
    wire c2538;
    assign in2538_1 = {pp53[56]};
    assign in2538_2 = {pp54[55]};
    Full_Adder FA_2538(s2538, c2538, in2538_1, in2538_2, pp52[57]);
    wire[0:0] s2539, in2539_1, in2539_2;
    wire c2539;
    assign in2539_1 = {pp56[53]};
    assign in2539_2 = {pp57[52]};
    Full_Adder FA_2539(s2539, c2539, in2539_1, in2539_2, pp55[54]);
    wire[0:0] s2540, in2540_1, in2540_2;
    wire c2540;
    assign in2540_1 = {pp59[50]};
    assign in2540_2 = {pp60[49]};
    Full_Adder FA_2540(s2540, c2540, in2540_1, in2540_2, pp58[51]);
    wire[0:0] s2541, in2541_1, in2541_2;
    wire c2541;
    assign in2541_1 = {pp48[62]};
    assign in2541_2 = {pp49[61]};
    Full_Adder FA_2541(s2541, c2541, in2541_1, in2541_2, pp47[63]);
    wire[0:0] s2542, in2542_1, in2542_2;
    wire c2542;
    assign in2542_1 = {pp51[59]};
    assign in2542_2 = {pp52[58]};
    Full_Adder FA_2542(s2542, c2542, in2542_1, in2542_2, pp50[60]);
    wire[0:0] s2543, in2543_1, in2543_2;
    wire c2543;
    assign in2543_1 = {pp54[56]};
    assign in2543_2 = {pp55[55]};
    Full_Adder FA_2543(s2543, c2543, in2543_1, in2543_2, pp53[57]);
    wire[0:0] s2544, in2544_1, in2544_2;
    wire c2544;
    assign in2544_1 = {pp57[53]};
    assign in2544_2 = {pp58[52]};
    Full_Adder FA_2544(s2544, c2544, in2544_1, in2544_2, pp56[54]);
    wire[0:0] s2545, in2545_1, in2545_2;
    wire c2545;
    assign in2545_1 = {pp49[62]};
    assign in2545_2 = {pp50[61]};
    Full_Adder FA_2545(s2545, c2545, in2545_1, in2545_2, pp48[63]);
    wire[0:0] s2546, in2546_1, in2546_2;
    wire c2546;
    assign in2546_1 = {pp52[59]};
    assign in2546_2 = {pp53[58]};
    Full_Adder FA_2546(s2546, c2546, in2546_1, in2546_2, pp51[60]);
    wire[0:0] s2547, in2547_1, in2547_2;
    wire c2547;
    assign in2547_1 = {pp55[56]};
    assign in2547_2 = {pp56[55]};
    Full_Adder FA_2547(s2547, c2547, in2547_1, in2547_2, pp54[57]);
    wire[0:0] s2548, in2548_1, in2548_2;
    wire c2548;
    assign in2548_1 = {pp50[62]};
    assign in2548_2 = {pp51[61]};
    Full_Adder FA_2548(s2548, c2548, in2548_1, in2548_2, pp49[63]);
    wire[0:0] s2549, in2549_1, in2549_2;
    wire c2549;
    assign in2549_1 = {pp53[59]};
    assign in2549_2 = {pp54[58]};
    Full_Adder FA_2549(s2549, c2549, in2549_1, in2549_2, pp52[60]);
    wire[0:0] s2550, in2550_1, in2550_2;
    wire c2550;
    assign in2550_1 = {pp51[62]};
    assign in2550_2 = {pp52[61]};
    Full_Adder FA_2550(s2550, c2550, in2550_1, in2550_2, pp50[63]);

    /*Stage 5*/
    wire[0:0] s2551, in2551_1, in2551_2;
    wire c2551;
    assign in2551_1 = {pp0[10]};
    assign in2551_2 = {pp1[9]};
    Half_Adder HA_2551(s2551, c2551, in2551_1, in2551_2);
    wire[0:0] s2552, in2552_1, in2552_2;
    wire c2552;
    assign in2552_1 = {pp1[10]};
    assign in2552_2 = {pp2[9]};
    Full_Adder FA_2552(s2552, c2552, in2552_1, in2552_2, pp0[11]);
    wire[0:0] s2553, in2553_1, in2553_2;
    wire c2553;
    assign in2553_1 = {pp3[8]};
    assign in2553_2 = {pp4[7]};
    Half_Adder HA_2553(s2553, c2553, in2553_1, in2553_2);
    wire[0:0] s2554, in2554_1, in2554_2;
    wire c2554;
    assign in2554_1 = {pp1[11]};
    assign in2554_2 = {pp2[10]};
    Full_Adder FA_2554(s2554, c2554, in2554_1, in2554_2, pp0[12]);
    wire[0:0] s2555, in2555_1, in2555_2;
    wire c2555;
    assign in2555_1 = {pp4[8]};
    assign in2555_2 = {pp5[7]};
    Full_Adder FA_2555(s2555, c2555, in2555_1, in2555_2, pp3[9]);
    wire[0:0] s2556, in2556_1, in2556_2;
    wire c2556;
    assign in2556_1 = {pp6[6]};
    assign in2556_2 = {pp7[5]};
    Half_Adder HA_2556(s2556, c2556, in2556_1, in2556_2);
    wire[0:0] s2557, in2557_1, in2557_2;
    wire c2557;
    assign in2557_1 = {pp1[12]};
    assign in2557_2 = {pp2[11]};
    Full_Adder FA_2557(s2557, c2557, in2557_1, in2557_2, pp0[13]);
    wire[0:0] s2558, in2558_1, in2558_2;
    wire c2558;
    assign in2558_1 = {pp4[9]};
    assign in2558_2 = {pp5[8]};
    Full_Adder FA_2558(s2558, c2558, in2558_1, in2558_2, pp3[10]);
    wire[0:0] s2559, in2559_1, in2559_2;
    wire c2559;
    assign in2559_1 = {pp7[6]};
    assign in2559_2 = {pp8[5]};
    Full_Adder FA_2559(s2559, c2559, in2559_1, in2559_2, pp6[7]);
    wire[0:0] s2560, in2560_1, in2560_2;
    wire c2560;
    assign in2560_1 = {pp9[4]};
    assign in2560_2 = {pp10[3]};
    Half_Adder HA_2560(s2560, c2560, in2560_1, in2560_2);
    wire[0:0] s2561, in2561_1, in2561_2;
    wire c2561;
    assign in2561_1 = {pp3[11]};
    assign in2561_2 = {pp4[10]};
    Full_Adder FA_2561(s2561, c2561, in2561_1, in2561_2, pp2[12]);
    wire[0:0] s2562, in2562_1, in2562_2;
    wire c2562;
    assign in2562_1 = {pp6[8]};
    assign in2562_2 = {pp7[7]};
    Full_Adder FA_2562(s2562, c2562, in2562_1, in2562_2, pp5[9]);
    wire[0:0] s2563, in2563_1, in2563_2;
    wire c2563;
    assign in2563_1 = {pp9[5]};
    assign in2563_2 = {pp10[4]};
    Full_Adder FA_2563(s2563, c2563, in2563_1, in2563_2, pp8[6]);
    wire[0:0] s2564, in2564_1, in2564_2;
    wire c2564;
    assign in2564_1 = {pp12[2]};
    assign in2564_2 = {pp13[1]};
    Full_Adder FA_2564(s2564, c2564, in2564_1, in2564_2, pp11[3]);
    wire[0:0] s2565, in2565_1, in2565_2;
    wire c2565;
    assign in2565_1 = {pp6[9]};
    assign in2565_2 = {pp7[8]};
    Full_Adder FA_2565(s2565, c2565, in2565_1, in2565_2, pp5[10]);
    wire[0:0] s2566, in2566_1, in2566_2;
    wire c2566;
    assign in2566_1 = {pp9[6]};
    assign in2566_2 = {pp10[5]};
    Full_Adder FA_2566(s2566, c2566, in2566_1, in2566_2, pp8[7]);
    wire[0:0] s2567, in2567_1, in2567_2;
    wire c2567;
    assign in2567_1 = {pp12[3]};
    assign in2567_2 = {pp13[2]};
    Full_Adder FA_2567(s2567, c2567, in2567_1, in2567_2, pp11[4]);
    wire[0:0] s2568, in2568_1, in2568_2;
    wire c2568;
    assign in2568_1 = {pp15[0]};
    assign in2568_2 = {c1981};
    Full_Adder FA_2568(s2568, c2568, in2568_1, in2568_2, pp14[1]);
    wire[0:0] s2569, in2569_1, in2569_2;
    wire c2569;
    assign in2569_1 = {pp9[7]};
    assign in2569_2 = {pp10[6]};
    Full_Adder FA_2569(s2569, c2569, in2569_1, in2569_2, pp8[8]);
    wire[0:0] s2570, in2570_1, in2570_2;
    wire c2570;
    assign in2570_1 = {pp12[4]};
    assign in2570_2 = {pp13[3]};
    Full_Adder FA_2570(s2570, c2570, in2570_1, in2570_2, pp11[5]);
    wire[0:0] s2571, in2571_1, in2571_2;
    wire c2571;
    assign in2571_1 = {pp15[1]};
    assign in2571_2 = {pp16[0]};
    Full_Adder FA_2571(s2571, c2571, in2571_1, in2571_2, pp14[2]);
    wire[0:0] s2572, in2572_1, in2572_2;
    wire c2572;
    assign in2572_1 = {c1983};
    assign in2572_2 = {s1984[0]};
    Full_Adder FA_2572(s2572, c2572, in2572_1, in2572_2, c1982);
    wire[0:0] s2573, in2573_1, in2573_2;
    wire c2573;
    assign in2573_1 = {pp12[5]};
    assign in2573_2 = {pp13[4]};
    Full_Adder FA_2573(s2573, c2573, in2573_1, in2573_2, pp11[6]);
    wire[0:0] s2574, in2574_1, in2574_2;
    wire c2574;
    assign in2574_1 = {pp15[2]};
    assign in2574_2 = {pp16[1]};
    Full_Adder FA_2574(s2574, c2574, in2574_1, in2574_2, pp14[3]);
    wire[0:0] s2575, in2575_1, in2575_2;
    wire c2575;
    assign in2575_1 = {c1984};
    assign in2575_2 = {c1985};
    Full_Adder FA_2575(s2575, c2575, in2575_1, in2575_2, pp17[0]);
    wire[0:0] s2576, in2576_1, in2576_2;
    wire c2576;
    assign in2576_1 = {s1987[0]};
    assign in2576_2 = {s1988[0]};
    Full_Adder FA_2576(s2576, c2576, in2576_1, in2576_2, c1986);
    wire[0:0] s2577, in2577_1, in2577_2;
    wire c2577;
    assign in2577_1 = {pp15[3]};
    assign in2577_2 = {pp16[2]};
    Full_Adder FA_2577(s2577, c2577, in2577_1, in2577_2, pp14[4]);
    wire[0:0] s2578, in2578_1, in2578_2;
    wire c2578;
    assign in2578_1 = {pp18[0]};
    assign in2578_2 = {c1987};
    Full_Adder FA_2578(s2578, c2578, in2578_1, in2578_2, pp17[1]);
    wire[0:0] s2579, in2579_1, in2579_2;
    wire c2579;
    assign in2579_1 = {c1989};
    assign in2579_2 = {c1990};
    Full_Adder FA_2579(s2579, c2579, in2579_1, in2579_2, c1988);
    wire[0:0] s2580, in2580_1, in2580_2;
    wire c2580;
    assign in2580_1 = {s1992[0]};
    assign in2580_2 = {s1993[0]};
    Full_Adder FA_2580(s2580, c2580, in2580_1, in2580_2, s1991[0]);
    wire[0:0] s2581, in2581_1, in2581_2;
    wire c2581;
    assign in2581_1 = {pp18[1]};
    assign in2581_2 = {pp19[0]};
    Full_Adder FA_2581(s2581, c2581, in2581_1, in2581_2, pp17[2]);
    wire[0:0] s2582, in2582_1, in2582_2;
    wire c2582;
    assign in2582_1 = {c1992};
    assign in2582_2 = {c1993};
    Full_Adder FA_2582(s2582, c2582, in2582_1, in2582_2, c1991);
    wire[0:0] s2583, in2583_1, in2583_2;
    wire c2583;
    assign in2583_1 = {c1995};
    assign in2583_2 = {s1996[0]};
    Full_Adder FA_2583(s2583, c2583, in2583_1, in2583_2, c1994);
    wire[0:0] s2584, in2584_1, in2584_2;
    wire c2584;
    assign in2584_1 = {s1998[0]};
    assign in2584_2 = {s1999[0]};
    Full_Adder FA_2584(s2584, c2584, in2584_1, in2584_2, s1997[0]);
    wire[0:0] s2585, in2585_1, in2585_2;
    wire c2585;
    assign in2585_1 = {s1261[0]};
    assign in2585_2 = {c1996};
    Full_Adder FA_2585(s2585, c2585, in2585_1, in2585_2, pp20[0]);
    wire[0:0] s2586, in2586_1, in2586_2;
    wire c2586;
    assign in2586_1 = {c1998};
    assign in2586_2 = {c1999};
    Full_Adder FA_2586(s2586, c2586, in2586_1, in2586_2, c1997);
    wire[0:0] s2587, in2587_1, in2587_2;
    wire c2587;
    assign in2587_1 = {c2001};
    assign in2587_2 = {s2002[0]};
    Full_Adder FA_2587(s2587, c2587, in2587_1, in2587_2, c2000);
    wire[0:0] s2588, in2588_1, in2588_2;
    wire c2588;
    assign in2588_1 = {s2004[0]};
    assign in2588_2 = {s2005[0]};
    Full_Adder FA_2588(s2588, c2588, in2588_1, in2588_2, s2003[0]);
    wire[0:0] s2589, in2589_1, in2589_2;
    wire c2589;
    assign in2589_1 = {s1263[0]};
    assign in2589_2 = {c2002};
    Full_Adder FA_2589(s2589, c2589, in2589_1, in2589_2, s1262[0]);
    wire[0:0] s2590, in2590_1, in2590_2;
    wire c2590;
    assign in2590_1 = {c2004};
    assign in2590_2 = {c2005};
    Full_Adder FA_2590(s2590, c2590, in2590_1, in2590_2, c2003);
    wire[0:0] s2591, in2591_1, in2591_2;
    wire c2591;
    assign in2591_1 = {c2007};
    assign in2591_2 = {s2008[0]};
    Full_Adder FA_2591(s2591, c2591, in2591_1, in2591_2, c2006);
    wire[0:0] s2592, in2592_1, in2592_2;
    wire c2592;
    assign in2592_1 = {s2010[0]};
    assign in2592_2 = {s2011[0]};
    Full_Adder FA_2592(s2592, c2592, in2592_1, in2592_2, s2009[0]);
    wire[0:0] s2593, in2593_1, in2593_2;
    wire c2593;
    assign in2593_1 = {s1266[0]};
    assign in2593_2 = {c2008};
    Full_Adder FA_2593(s2593, c2593, in2593_1, in2593_2, s1265[0]);
    wire[0:0] s2594, in2594_1, in2594_2;
    wire c2594;
    assign in2594_1 = {c2010};
    assign in2594_2 = {c2011};
    Full_Adder FA_2594(s2594, c2594, in2594_1, in2594_2, c2009);
    wire[0:0] s2595, in2595_1, in2595_2;
    wire c2595;
    assign in2595_1 = {c2013};
    assign in2595_2 = {s2014[0]};
    Full_Adder FA_2595(s2595, c2595, in2595_1, in2595_2, c2012);
    wire[0:0] s2596, in2596_1, in2596_2;
    wire c2596;
    assign in2596_1 = {s2016[0]};
    assign in2596_2 = {s2017[0]};
    Full_Adder FA_2596(s2596, c2596, in2596_1, in2596_2, s2015[0]);
    wire[0:0] s2597, in2597_1, in2597_2;
    wire c2597;
    assign in2597_1 = {s1270[0]};
    assign in2597_2 = {c2014};
    Full_Adder FA_2597(s2597, c2597, in2597_1, in2597_2, s1269[0]);
    wire[0:0] s2598, in2598_1, in2598_2;
    wire c2598;
    assign in2598_1 = {c2016};
    assign in2598_2 = {c2017};
    Full_Adder FA_2598(s2598, c2598, in2598_1, in2598_2, c2015);
    wire[0:0] s2599, in2599_1, in2599_2;
    wire c2599;
    assign in2599_1 = {c2019};
    assign in2599_2 = {s2020[0]};
    Full_Adder FA_2599(s2599, c2599, in2599_1, in2599_2, c2018);
    wire[0:0] s2600, in2600_1, in2600_2;
    wire c2600;
    assign in2600_1 = {s2022[0]};
    assign in2600_2 = {s2023[0]};
    Full_Adder FA_2600(s2600, c2600, in2600_1, in2600_2, s2021[0]);
    wire[0:0] s2601, in2601_1, in2601_2;
    wire c2601;
    assign in2601_1 = {s1275[0]};
    assign in2601_2 = {c2020};
    Full_Adder FA_2601(s2601, c2601, in2601_1, in2601_2, s1274[0]);
    wire[0:0] s2602, in2602_1, in2602_2;
    wire c2602;
    assign in2602_1 = {c2022};
    assign in2602_2 = {c2023};
    Full_Adder FA_2602(s2602, c2602, in2602_1, in2602_2, c2021);
    wire[0:0] s2603, in2603_1, in2603_2;
    wire c2603;
    assign in2603_1 = {c2025};
    assign in2603_2 = {s2026[0]};
    Full_Adder FA_2603(s2603, c2603, in2603_1, in2603_2, c2024);
    wire[0:0] s2604, in2604_1, in2604_2;
    wire c2604;
    assign in2604_1 = {s2028[0]};
    assign in2604_2 = {s2029[0]};
    Full_Adder FA_2604(s2604, c2604, in2604_1, in2604_2, s2027[0]);
    wire[0:0] s2605, in2605_1, in2605_2;
    wire c2605;
    assign in2605_1 = {s1281[0]};
    assign in2605_2 = {c2026};
    Full_Adder FA_2605(s2605, c2605, in2605_1, in2605_2, s1280[0]);
    wire[0:0] s2606, in2606_1, in2606_2;
    wire c2606;
    assign in2606_1 = {c2028};
    assign in2606_2 = {c2029};
    Full_Adder FA_2606(s2606, c2606, in2606_1, in2606_2, c2027);
    wire[0:0] s2607, in2607_1, in2607_2;
    wire c2607;
    assign in2607_1 = {c2031};
    assign in2607_2 = {s2032[0]};
    Full_Adder FA_2607(s2607, c2607, in2607_1, in2607_2, c2030);
    wire[0:0] s2608, in2608_1, in2608_2;
    wire c2608;
    assign in2608_1 = {s2034[0]};
    assign in2608_2 = {s2035[0]};
    Full_Adder FA_2608(s2608, c2608, in2608_1, in2608_2, s2033[0]);
    wire[0:0] s2609, in2609_1, in2609_2;
    wire c2609;
    assign in2609_1 = {s1288[0]};
    assign in2609_2 = {c2032};
    Full_Adder FA_2609(s2609, c2609, in2609_1, in2609_2, s1287[0]);
    wire[0:0] s2610, in2610_1, in2610_2;
    wire c2610;
    assign in2610_1 = {c2034};
    assign in2610_2 = {c2035};
    Full_Adder FA_2610(s2610, c2610, in2610_1, in2610_2, c2033);
    wire[0:0] s2611, in2611_1, in2611_2;
    wire c2611;
    assign in2611_1 = {c2037};
    assign in2611_2 = {s2038[0]};
    Full_Adder FA_2611(s2611, c2611, in2611_1, in2611_2, c2036);
    wire[0:0] s2612, in2612_1, in2612_2;
    wire c2612;
    assign in2612_1 = {s2040[0]};
    assign in2612_2 = {s2041[0]};
    Full_Adder FA_2612(s2612, c2612, in2612_1, in2612_2, s2039[0]);
    wire[0:0] s2613, in2613_1, in2613_2;
    wire c2613;
    assign in2613_1 = {s1296[0]};
    assign in2613_2 = {c2038};
    Full_Adder FA_2613(s2613, c2613, in2613_1, in2613_2, s1295[0]);
    wire[0:0] s2614, in2614_1, in2614_2;
    wire c2614;
    assign in2614_1 = {c2040};
    assign in2614_2 = {c2041};
    Full_Adder FA_2614(s2614, c2614, in2614_1, in2614_2, c2039);
    wire[0:0] s2615, in2615_1, in2615_2;
    wire c2615;
    assign in2615_1 = {c2043};
    assign in2615_2 = {s2044[0]};
    Full_Adder FA_2615(s2615, c2615, in2615_1, in2615_2, c2042);
    wire[0:0] s2616, in2616_1, in2616_2;
    wire c2616;
    assign in2616_1 = {s2046[0]};
    assign in2616_2 = {s2047[0]};
    Full_Adder FA_2616(s2616, c2616, in2616_1, in2616_2, s2045[0]);
    wire[0:0] s2617, in2617_1, in2617_2;
    wire c2617;
    assign in2617_1 = {s1305[0]};
    assign in2617_2 = {c2044};
    Full_Adder FA_2617(s2617, c2617, in2617_1, in2617_2, s1304[0]);
    wire[0:0] s2618, in2618_1, in2618_2;
    wire c2618;
    assign in2618_1 = {c2046};
    assign in2618_2 = {c2047};
    Full_Adder FA_2618(s2618, c2618, in2618_1, in2618_2, c2045);
    wire[0:0] s2619, in2619_1, in2619_2;
    wire c2619;
    assign in2619_1 = {c2049};
    assign in2619_2 = {s2050[0]};
    Full_Adder FA_2619(s2619, c2619, in2619_1, in2619_2, c2048);
    wire[0:0] s2620, in2620_1, in2620_2;
    wire c2620;
    assign in2620_1 = {s2052[0]};
    assign in2620_2 = {s2053[0]};
    Full_Adder FA_2620(s2620, c2620, in2620_1, in2620_2, s2051[0]);
    wire[0:0] s2621, in2621_1, in2621_2;
    wire c2621;
    assign in2621_1 = {s1314[0]};
    assign in2621_2 = {c2050};
    Full_Adder FA_2621(s2621, c2621, in2621_1, in2621_2, s1313[0]);
    wire[0:0] s2622, in2622_1, in2622_2;
    wire c2622;
    assign in2622_1 = {c2052};
    assign in2622_2 = {c2053};
    Full_Adder FA_2622(s2622, c2622, in2622_1, in2622_2, c2051);
    wire[0:0] s2623, in2623_1, in2623_2;
    wire c2623;
    assign in2623_1 = {c2055};
    assign in2623_2 = {s2056[0]};
    Full_Adder FA_2623(s2623, c2623, in2623_1, in2623_2, c2054);
    wire[0:0] s2624, in2624_1, in2624_2;
    wire c2624;
    assign in2624_1 = {s2058[0]};
    assign in2624_2 = {s2059[0]};
    Full_Adder FA_2624(s2624, c2624, in2624_1, in2624_2, s2057[0]);
    wire[0:0] s2625, in2625_1, in2625_2;
    wire c2625;
    assign in2625_1 = {s1323[0]};
    assign in2625_2 = {c2056};
    Full_Adder FA_2625(s2625, c2625, in2625_1, in2625_2, s1322[0]);
    wire[0:0] s2626, in2626_1, in2626_2;
    wire c2626;
    assign in2626_1 = {c2058};
    assign in2626_2 = {c2059};
    Full_Adder FA_2626(s2626, c2626, in2626_1, in2626_2, c2057);
    wire[0:0] s2627, in2627_1, in2627_2;
    wire c2627;
    assign in2627_1 = {c2061};
    assign in2627_2 = {s2062[0]};
    Full_Adder FA_2627(s2627, c2627, in2627_1, in2627_2, c2060);
    wire[0:0] s2628, in2628_1, in2628_2;
    wire c2628;
    assign in2628_1 = {s2064[0]};
    assign in2628_2 = {s2065[0]};
    Full_Adder FA_2628(s2628, c2628, in2628_1, in2628_2, s2063[0]);
    wire[0:0] s2629, in2629_1, in2629_2;
    wire c2629;
    assign in2629_1 = {s1332[0]};
    assign in2629_2 = {c2062};
    Full_Adder FA_2629(s2629, c2629, in2629_1, in2629_2, s1331[0]);
    wire[0:0] s2630, in2630_1, in2630_2;
    wire c2630;
    assign in2630_1 = {c2064};
    assign in2630_2 = {c2065};
    Full_Adder FA_2630(s2630, c2630, in2630_1, in2630_2, c2063);
    wire[0:0] s2631, in2631_1, in2631_2;
    wire c2631;
    assign in2631_1 = {c2067};
    assign in2631_2 = {s2068[0]};
    Full_Adder FA_2631(s2631, c2631, in2631_1, in2631_2, c2066);
    wire[0:0] s2632, in2632_1, in2632_2;
    wire c2632;
    assign in2632_1 = {s2070[0]};
    assign in2632_2 = {s2071[0]};
    Full_Adder FA_2632(s2632, c2632, in2632_1, in2632_2, s2069[0]);
    wire[0:0] s2633, in2633_1, in2633_2;
    wire c2633;
    assign in2633_1 = {s1341[0]};
    assign in2633_2 = {c2068};
    Full_Adder FA_2633(s2633, c2633, in2633_1, in2633_2, s1340[0]);
    wire[0:0] s2634, in2634_1, in2634_2;
    wire c2634;
    assign in2634_1 = {c2070};
    assign in2634_2 = {c2071};
    Full_Adder FA_2634(s2634, c2634, in2634_1, in2634_2, c2069);
    wire[0:0] s2635, in2635_1, in2635_2;
    wire c2635;
    assign in2635_1 = {c2073};
    assign in2635_2 = {s2074[0]};
    Full_Adder FA_2635(s2635, c2635, in2635_1, in2635_2, c2072);
    wire[0:0] s2636, in2636_1, in2636_2;
    wire c2636;
    assign in2636_1 = {s2076[0]};
    assign in2636_2 = {s2077[0]};
    Full_Adder FA_2636(s2636, c2636, in2636_1, in2636_2, s2075[0]);
    wire[0:0] s2637, in2637_1, in2637_2;
    wire c2637;
    assign in2637_1 = {s1350[0]};
    assign in2637_2 = {c2074};
    Full_Adder FA_2637(s2637, c2637, in2637_1, in2637_2, s1349[0]);
    wire[0:0] s2638, in2638_1, in2638_2;
    wire c2638;
    assign in2638_1 = {c2076};
    assign in2638_2 = {c2077};
    Full_Adder FA_2638(s2638, c2638, in2638_1, in2638_2, c2075);
    wire[0:0] s2639, in2639_1, in2639_2;
    wire c2639;
    assign in2639_1 = {c2079};
    assign in2639_2 = {s2080[0]};
    Full_Adder FA_2639(s2639, c2639, in2639_1, in2639_2, c2078);
    wire[0:0] s2640, in2640_1, in2640_2;
    wire c2640;
    assign in2640_1 = {s2082[0]};
    assign in2640_2 = {s2083[0]};
    Full_Adder FA_2640(s2640, c2640, in2640_1, in2640_2, s2081[0]);
    wire[0:0] s2641, in2641_1, in2641_2;
    wire c2641;
    assign in2641_1 = {s1359[0]};
    assign in2641_2 = {c2080};
    Full_Adder FA_2641(s2641, c2641, in2641_1, in2641_2, s1358[0]);
    wire[0:0] s2642, in2642_1, in2642_2;
    wire c2642;
    assign in2642_1 = {c2082};
    assign in2642_2 = {c2083};
    Full_Adder FA_2642(s2642, c2642, in2642_1, in2642_2, c2081);
    wire[0:0] s2643, in2643_1, in2643_2;
    wire c2643;
    assign in2643_1 = {c2085};
    assign in2643_2 = {s2086[0]};
    Full_Adder FA_2643(s2643, c2643, in2643_1, in2643_2, c2084);
    wire[0:0] s2644, in2644_1, in2644_2;
    wire c2644;
    assign in2644_1 = {s2088[0]};
    assign in2644_2 = {s2089[0]};
    Full_Adder FA_2644(s2644, c2644, in2644_1, in2644_2, s2087[0]);
    wire[0:0] s2645, in2645_1, in2645_2;
    wire c2645;
    assign in2645_1 = {s1368[0]};
    assign in2645_2 = {c2086};
    Full_Adder FA_2645(s2645, c2645, in2645_1, in2645_2, s1367[0]);
    wire[0:0] s2646, in2646_1, in2646_2;
    wire c2646;
    assign in2646_1 = {c2088};
    assign in2646_2 = {c2089};
    Full_Adder FA_2646(s2646, c2646, in2646_1, in2646_2, c2087);
    wire[0:0] s2647, in2647_1, in2647_2;
    wire c2647;
    assign in2647_1 = {c2091};
    assign in2647_2 = {s2092[0]};
    Full_Adder FA_2647(s2647, c2647, in2647_1, in2647_2, c2090);
    wire[0:0] s2648, in2648_1, in2648_2;
    wire c2648;
    assign in2648_1 = {s2094[0]};
    assign in2648_2 = {s2095[0]};
    Full_Adder FA_2648(s2648, c2648, in2648_1, in2648_2, s2093[0]);
    wire[0:0] s2649, in2649_1, in2649_2;
    wire c2649;
    assign in2649_1 = {s1377[0]};
    assign in2649_2 = {c2092};
    Full_Adder FA_2649(s2649, c2649, in2649_1, in2649_2, s1376[0]);
    wire[0:0] s2650, in2650_1, in2650_2;
    wire c2650;
    assign in2650_1 = {c2094};
    assign in2650_2 = {c2095};
    Full_Adder FA_2650(s2650, c2650, in2650_1, in2650_2, c2093);
    wire[0:0] s2651, in2651_1, in2651_2;
    wire c2651;
    assign in2651_1 = {c2097};
    assign in2651_2 = {s2098[0]};
    Full_Adder FA_2651(s2651, c2651, in2651_1, in2651_2, c2096);
    wire[0:0] s2652, in2652_1, in2652_2;
    wire c2652;
    assign in2652_1 = {s2100[0]};
    assign in2652_2 = {s2101[0]};
    Full_Adder FA_2652(s2652, c2652, in2652_1, in2652_2, s2099[0]);
    wire[0:0] s2653, in2653_1, in2653_2;
    wire c2653;
    assign in2653_1 = {s1386[0]};
    assign in2653_2 = {c2098};
    Full_Adder FA_2653(s2653, c2653, in2653_1, in2653_2, s1385[0]);
    wire[0:0] s2654, in2654_1, in2654_2;
    wire c2654;
    assign in2654_1 = {c2100};
    assign in2654_2 = {c2101};
    Full_Adder FA_2654(s2654, c2654, in2654_1, in2654_2, c2099);
    wire[0:0] s2655, in2655_1, in2655_2;
    wire c2655;
    assign in2655_1 = {c2103};
    assign in2655_2 = {s2104[0]};
    Full_Adder FA_2655(s2655, c2655, in2655_1, in2655_2, c2102);
    wire[0:0] s2656, in2656_1, in2656_2;
    wire c2656;
    assign in2656_1 = {s2106[0]};
    assign in2656_2 = {s2107[0]};
    Full_Adder FA_2656(s2656, c2656, in2656_1, in2656_2, s2105[0]);
    wire[0:0] s2657, in2657_1, in2657_2;
    wire c2657;
    assign in2657_1 = {s1395[0]};
    assign in2657_2 = {c2104};
    Full_Adder FA_2657(s2657, c2657, in2657_1, in2657_2, s1394[0]);
    wire[0:0] s2658, in2658_1, in2658_2;
    wire c2658;
    assign in2658_1 = {c2106};
    assign in2658_2 = {c2107};
    Full_Adder FA_2658(s2658, c2658, in2658_1, in2658_2, c2105);
    wire[0:0] s2659, in2659_1, in2659_2;
    wire c2659;
    assign in2659_1 = {c2109};
    assign in2659_2 = {s2110[0]};
    Full_Adder FA_2659(s2659, c2659, in2659_1, in2659_2, c2108);
    wire[0:0] s2660, in2660_1, in2660_2;
    wire c2660;
    assign in2660_1 = {s2112[0]};
    assign in2660_2 = {s2113[0]};
    Full_Adder FA_2660(s2660, c2660, in2660_1, in2660_2, s2111[0]);
    wire[0:0] s2661, in2661_1, in2661_2;
    wire c2661;
    assign in2661_1 = {s1404[0]};
    assign in2661_2 = {c2110};
    Full_Adder FA_2661(s2661, c2661, in2661_1, in2661_2, s1403[0]);
    wire[0:0] s2662, in2662_1, in2662_2;
    wire c2662;
    assign in2662_1 = {c2112};
    assign in2662_2 = {c2113};
    Full_Adder FA_2662(s2662, c2662, in2662_1, in2662_2, c2111);
    wire[0:0] s2663, in2663_1, in2663_2;
    wire c2663;
    assign in2663_1 = {c2115};
    assign in2663_2 = {s2116[0]};
    Full_Adder FA_2663(s2663, c2663, in2663_1, in2663_2, c2114);
    wire[0:0] s2664, in2664_1, in2664_2;
    wire c2664;
    assign in2664_1 = {s2118[0]};
    assign in2664_2 = {s2119[0]};
    Full_Adder FA_2664(s2664, c2664, in2664_1, in2664_2, s2117[0]);
    wire[0:0] s2665, in2665_1, in2665_2;
    wire c2665;
    assign in2665_1 = {s1413[0]};
    assign in2665_2 = {c2116};
    Full_Adder FA_2665(s2665, c2665, in2665_1, in2665_2, s1412[0]);
    wire[0:0] s2666, in2666_1, in2666_2;
    wire c2666;
    assign in2666_1 = {c2118};
    assign in2666_2 = {c2119};
    Full_Adder FA_2666(s2666, c2666, in2666_1, in2666_2, c2117);
    wire[0:0] s2667, in2667_1, in2667_2;
    wire c2667;
    assign in2667_1 = {c2121};
    assign in2667_2 = {s2122[0]};
    Full_Adder FA_2667(s2667, c2667, in2667_1, in2667_2, c2120);
    wire[0:0] s2668, in2668_1, in2668_2;
    wire c2668;
    assign in2668_1 = {s2124[0]};
    assign in2668_2 = {s2125[0]};
    Full_Adder FA_2668(s2668, c2668, in2668_1, in2668_2, s2123[0]);
    wire[0:0] s2669, in2669_1, in2669_2;
    wire c2669;
    assign in2669_1 = {s1422[0]};
    assign in2669_2 = {c2122};
    Full_Adder FA_2669(s2669, c2669, in2669_1, in2669_2, s1421[0]);
    wire[0:0] s2670, in2670_1, in2670_2;
    wire c2670;
    assign in2670_1 = {c2124};
    assign in2670_2 = {c2125};
    Full_Adder FA_2670(s2670, c2670, in2670_1, in2670_2, c2123);
    wire[0:0] s2671, in2671_1, in2671_2;
    wire c2671;
    assign in2671_1 = {c2127};
    assign in2671_2 = {s2128[0]};
    Full_Adder FA_2671(s2671, c2671, in2671_1, in2671_2, c2126);
    wire[0:0] s2672, in2672_1, in2672_2;
    wire c2672;
    assign in2672_1 = {s2130[0]};
    assign in2672_2 = {s2131[0]};
    Full_Adder FA_2672(s2672, c2672, in2672_1, in2672_2, s2129[0]);
    wire[0:0] s2673, in2673_1, in2673_2;
    wire c2673;
    assign in2673_1 = {s1431[0]};
    assign in2673_2 = {c2128};
    Full_Adder FA_2673(s2673, c2673, in2673_1, in2673_2, s1430[0]);
    wire[0:0] s2674, in2674_1, in2674_2;
    wire c2674;
    assign in2674_1 = {c2130};
    assign in2674_2 = {c2131};
    Full_Adder FA_2674(s2674, c2674, in2674_1, in2674_2, c2129);
    wire[0:0] s2675, in2675_1, in2675_2;
    wire c2675;
    assign in2675_1 = {c2133};
    assign in2675_2 = {s2134[0]};
    Full_Adder FA_2675(s2675, c2675, in2675_1, in2675_2, c2132);
    wire[0:0] s2676, in2676_1, in2676_2;
    wire c2676;
    assign in2676_1 = {s2136[0]};
    assign in2676_2 = {s2137[0]};
    Full_Adder FA_2676(s2676, c2676, in2676_1, in2676_2, s2135[0]);
    wire[0:0] s2677, in2677_1, in2677_2;
    wire c2677;
    assign in2677_1 = {s1440[0]};
    assign in2677_2 = {c2134};
    Full_Adder FA_2677(s2677, c2677, in2677_1, in2677_2, s1439[0]);
    wire[0:0] s2678, in2678_1, in2678_2;
    wire c2678;
    assign in2678_1 = {c2136};
    assign in2678_2 = {c2137};
    Full_Adder FA_2678(s2678, c2678, in2678_1, in2678_2, c2135);
    wire[0:0] s2679, in2679_1, in2679_2;
    wire c2679;
    assign in2679_1 = {c2139};
    assign in2679_2 = {s2140[0]};
    Full_Adder FA_2679(s2679, c2679, in2679_1, in2679_2, c2138);
    wire[0:0] s2680, in2680_1, in2680_2;
    wire c2680;
    assign in2680_1 = {s2142[0]};
    assign in2680_2 = {s2143[0]};
    Full_Adder FA_2680(s2680, c2680, in2680_1, in2680_2, s2141[0]);
    wire[0:0] s2681, in2681_1, in2681_2;
    wire c2681;
    assign in2681_1 = {s1449[0]};
    assign in2681_2 = {c2140};
    Full_Adder FA_2681(s2681, c2681, in2681_1, in2681_2, s1448[0]);
    wire[0:0] s2682, in2682_1, in2682_2;
    wire c2682;
    assign in2682_1 = {c2142};
    assign in2682_2 = {c2143};
    Full_Adder FA_2682(s2682, c2682, in2682_1, in2682_2, c2141);
    wire[0:0] s2683, in2683_1, in2683_2;
    wire c2683;
    assign in2683_1 = {c2145};
    assign in2683_2 = {s2146[0]};
    Full_Adder FA_2683(s2683, c2683, in2683_1, in2683_2, c2144);
    wire[0:0] s2684, in2684_1, in2684_2;
    wire c2684;
    assign in2684_1 = {s2148[0]};
    assign in2684_2 = {s2149[0]};
    Full_Adder FA_2684(s2684, c2684, in2684_1, in2684_2, s2147[0]);
    wire[0:0] s2685, in2685_1, in2685_2;
    wire c2685;
    assign in2685_1 = {s1458[0]};
    assign in2685_2 = {c2146};
    Full_Adder FA_2685(s2685, c2685, in2685_1, in2685_2, s1457[0]);
    wire[0:0] s2686, in2686_1, in2686_2;
    wire c2686;
    assign in2686_1 = {c2148};
    assign in2686_2 = {c2149};
    Full_Adder FA_2686(s2686, c2686, in2686_1, in2686_2, c2147);
    wire[0:0] s2687, in2687_1, in2687_2;
    wire c2687;
    assign in2687_1 = {c2151};
    assign in2687_2 = {s2152[0]};
    Full_Adder FA_2687(s2687, c2687, in2687_1, in2687_2, c2150);
    wire[0:0] s2688, in2688_1, in2688_2;
    wire c2688;
    assign in2688_1 = {s2154[0]};
    assign in2688_2 = {s2155[0]};
    Full_Adder FA_2688(s2688, c2688, in2688_1, in2688_2, s2153[0]);
    wire[0:0] s2689, in2689_1, in2689_2;
    wire c2689;
    assign in2689_1 = {s1467[0]};
    assign in2689_2 = {c2152};
    Full_Adder FA_2689(s2689, c2689, in2689_1, in2689_2, s1466[0]);
    wire[0:0] s2690, in2690_1, in2690_2;
    wire c2690;
    assign in2690_1 = {c2154};
    assign in2690_2 = {c2155};
    Full_Adder FA_2690(s2690, c2690, in2690_1, in2690_2, c2153);
    wire[0:0] s2691, in2691_1, in2691_2;
    wire c2691;
    assign in2691_1 = {c2157};
    assign in2691_2 = {s2158[0]};
    Full_Adder FA_2691(s2691, c2691, in2691_1, in2691_2, c2156);
    wire[0:0] s2692, in2692_1, in2692_2;
    wire c2692;
    assign in2692_1 = {s2160[0]};
    assign in2692_2 = {s2161[0]};
    Full_Adder FA_2692(s2692, c2692, in2692_1, in2692_2, s2159[0]);
    wire[0:0] s2693, in2693_1, in2693_2;
    wire c2693;
    assign in2693_1 = {s1476[0]};
    assign in2693_2 = {c2158};
    Full_Adder FA_2693(s2693, c2693, in2693_1, in2693_2, s1475[0]);
    wire[0:0] s2694, in2694_1, in2694_2;
    wire c2694;
    assign in2694_1 = {c2160};
    assign in2694_2 = {c2161};
    Full_Adder FA_2694(s2694, c2694, in2694_1, in2694_2, c2159);
    wire[0:0] s2695, in2695_1, in2695_2;
    wire c2695;
    assign in2695_1 = {c2163};
    assign in2695_2 = {s2164[0]};
    Full_Adder FA_2695(s2695, c2695, in2695_1, in2695_2, c2162);
    wire[0:0] s2696, in2696_1, in2696_2;
    wire c2696;
    assign in2696_1 = {s2166[0]};
    assign in2696_2 = {s2167[0]};
    Full_Adder FA_2696(s2696, c2696, in2696_1, in2696_2, s2165[0]);
    wire[0:0] s2697, in2697_1, in2697_2;
    wire c2697;
    assign in2697_1 = {s1485[0]};
    assign in2697_2 = {c2164};
    Full_Adder FA_2697(s2697, c2697, in2697_1, in2697_2, s1484[0]);
    wire[0:0] s2698, in2698_1, in2698_2;
    wire c2698;
    assign in2698_1 = {c2166};
    assign in2698_2 = {c2167};
    Full_Adder FA_2698(s2698, c2698, in2698_1, in2698_2, c2165);
    wire[0:0] s2699, in2699_1, in2699_2;
    wire c2699;
    assign in2699_1 = {c2169};
    assign in2699_2 = {s2170[0]};
    Full_Adder FA_2699(s2699, c2699, in2699_1, in2699_2, c2168);
    wire[0:0] s2700, in2700_1, in2700_2;
    wire c2700;
    assign in2700_1 = {s2172[0]};
    assign in2700_2 = {s2173[0]};
    Full_Adder FA_2700(s2700, c2700, in2700_1, in2700_2, s2171[0]);
    wire[0:0] s2701, in2701_1, in2701_2;
    wire c2701;
    assign in2701_1 = {s1494[0]};
    assign in2701_2 = {c2170};
    Full_Adder FA_2701(s2701, c2701, in2701_1, in2701_2, s1493[0]);
    wire[0:0] s2702, in2702_1, in2702_2;
    wire c2702;
    assign in2702_1 = {c2172};
    assign in2702_2 = {c2173};
    Full_Adder FA_2702(s2702, c2702, in2702_1, in2702_2, c2171);
    wire[0:0] s2703, in2703_1, in2703_2;
    wire c2703;
    assign in2703_1 = {c2175};
    assign in2703_2 = {s2176[0]};
    Full_Adder FA_2703(s2703, c2703, in2703_1, in2703_2, c2174);
    wire[0:0] s2704, in2704_1, in2704_2;
    wire c2704;
    assign in2704_1 = {s2178[0]};
    assign in2704_2 = {s2179[0]};
    Full_Adder FA_2704(s2704, c2704, in2704_1, in2704_2, s2177[0]);
    wire[0:0] s2705, in2705_1, in2705_2;
    wire c2705;
    assign in2705_1 = {s1503[0]};
    assign in2705_2 = {c2176};
    Full_Adder FA_2705(s2705, c2705, in2705_1, in2705_2, s1502[0]);
    wire[0:0] s2706, in2706_1, in2706_2;
    wire c2706;
    assign in2706_1 = {c2178};
    assign in2706_2 = {c2179};
    Full_Adder FA_2706(s2706, c2706, in2706_1, in2706_2, c2177);
    wire[0:0] s2707, in2707_1, in2707_2;
    wire c2707;
    assign in2707_1 = {c2181};
    assign in2707_2 = {s2182[0]};
    Full_Adder FA_2707(s2707, c2707, in2707_1, in2707_2, c2180);
    wire[0:0] s2708, in2708_1, in2708_2;
    wire c2708;
    assign in2708_1 = {s2184[0]};
    assign in2708_2 = {s2185[0]};
    Full_Adder FA_2708(s2708, c2708, in2708_1, in2708_2, s2183[0]);
    wire[0:0] s2709, in2709_1, in2709_2;
    wire c2709;
    assign in2709_1 = {s1512[0]};
    assign in2709_2 = {c2182};
    Full_Adder FA_2709(s2709, c2709, in2709_1, in2709_2, s1511[0]);
    wire[0:0] s2710, in2710_1, in2710_2;
    wire c2710;
    assign in2710_1 = {c2184};
    assign in2710_2 = {c2185};
    Full_Adder FA_2710(s2710, c2710, in2710_1, in2710_2, c2183);
    wire[0:0] s2711, in2711_1, in2711_2;
    wire c2711;
    assign in2711_1 = {c2187};
    assign in2711_2 = {s2188[0]};
    Full_Adder FA_2711(s2711, c2711, in2711_1, in2711_2, c2186);
    wire[0:0] s2712, in2712_1, in2712_2;
    wire c2712;
    assign in2712_1 = {s2190[0]};
    assign in2712_2 = {s2191[0]};
    Full_Adder FA_2712(s2712, c2712, in2712_1, in2712_2, s2189[0]);
    wire[0:0] s2713, in2713_1, in2713_2;
    wire c2713;
    assign in2713_1 = {s1521[0]};
    assign in2713_2 = {c2188};
    Full_Adder FA_2713(s2713, c2713, in2713_1, in2713_2, s1520[0]);
    wire[0:0] s2714, in2714_1, in2714_2;
    wire c2714;
    assign in2714_1 = {c2190};
    assign in2714_2 = {c2191};
    Full_Adder FA_2714(s2714, c2714, in2714_1, in2714_2, c2189);
    wire[0:0] s2715, in2715_1, in2715_2;
    wire c2715;
    assign in2715_1 = {c2193};
    assign in2715_2 = {s2194[0]};
    Full_Adder FA_2715(s2715, c2715, in2715_1, in2715_2, c2192);
    wire[0:0] s2716, in2716_1, in2716_2;
    wire c2716;
    assign in2716_1 = {s2196[0]};
    assign in2716_2 = {s2197[0]};
    Full_Adder FA_2716(s2716, c2716, in2716_1, in2716_2, s2195[0]);
    wire[0:0] s2717, in2717_1, in2717_2;
    wire c2717;
    assign in2717_1 = {s1530[0]};
    assign in2717_2 = {c2194};
    Full_Adder FA_2717(s2717, c2717, in2717_1, in2717_2, s1529[0]);
    wire[0:0] s2718, in2718_1, in2718_2;
    wire c2718;
    assign in2718_1 = {c2196};
    assign in2718_2 = {c2197};
    Full_Adder FA_2718(s2718, c2718, in2718_1, in2718_2, c2195);
    wire[0:0] s2719, in2719_1, in2719_2;
    wire c2719;
    assign in2719_1 = {c2199};
    assign in2719_2 = {s2200[0]};
    Full_Adder FA_2719(s2719, c2719, in2719_1, in2719_2, c2198);
    wire[0:0] s2720, in2720_1, in2720_2;
    wire c2720;
    assign in2720_1 = {s2202[0]};
    assign in2720_2 = {s2203[0]};
    Full_Adder FA_2720(s2720, c2720, in2720_1, in2720_2, s2201[0]);
    wire[0:0] s2721, in2721_1, in2721_2;
    wire c2721;
    assign in2721_1 = {s1539[0]};
    assign in2721_2 = {c2200};
    Full_Adder FA_2721(s2721, c2721, in2721_1, in2721_2, s1538[0]);
    wire[0:0] s2722, in2722_1, in2722_2;
    wire c2722;
    assign in2722_1 = {c2202};
    assign in2722_2 = {c2203};
    Full_Adder FA_2722(s2722, c2722, in2722_1, in2722_2, c2201);
    wire[0:0] s2723, in2723_1, in2723_2;
    wire c2723;
    assign in2723_1 = {c2205};
    assign in2723_2 = {s2206[0]};
    Full_Adder FA_2723(s2723, c2723, in2723_1, in2723_2, c2204);
    wire[0:0] s2724, in2724_1, in2724_2;
    wire c2724;
    assign in2724_1 = {s2208[0]};
    assign in2724_2 = {s2209[0]};
    Full_Adder FA_2724(s2724, c2724, in2724_1, in2724_2, s2207[0]);
    wire[0:0] s2725, in2725_1, in2725_2;
    wire c2725;
    assign in2725_1 = {s1548[0]};
    assign in2725_2 = {c2206};
    Full_Adder FA_2725(s2725, c2725, in2725_1, in2725_2, s1547[0]);
    wire[0:0] s2726, in2726_1, in2726_2;
    wire c2726;
    assign in2726_1 = {c2208};
    assign in2726_2 = {c2209};
    Full_Adder FA_2726(s2726, c2726, in2726_1, in2726_2, c2207);
    wire[0:0] s2727, in2727_1, in2727_2;
    wire c2727;
    assign in2727_1 = {c2211};
    assign in2727_2 = {s2212[0]};
    Full_Adder FA_2727(s2727, c2727, in2727_1, in2727_2, c2210);
    wire[0:0] s2728, in2728_1, in2728_2;
    wire c2728;
    assign in2728_1 = {s2214[0]};
    assign in2728_2 = {s2215[0]};
    Full_Adder FA_2728(s2728, c2728, in2728_1, in2728_2, s2213[0]);
    wire[0:0] s2729, in2729_1, in2729_2;
    wire c2729;
    assign in2729_1 = {s1557[0]};
    assign in2729_2 = {c2212};
    Full_Adder FA_2729(s2729, c2729, in2729_1, in2729_2, s1556[0]);
    wire[0:0] s2730, in2730_1, in2730_2;
    wire c2730;
    assign in2730_1 = {c2214};
    assign in2730_2 = {c2215};
    Full_Adder FA_2730(s2730, c2730, in2730_1, in2730_2, c2213);
    wire[0:0] s2731, in2731_1, in2731_2;
    wire c2731;
    assign in2731_1 = {c2217};
    assign in2731_2 = {s2218[0]};
    Full_Adder FA_2731(s2731, c2731, in2731_1, in2731_2, c2216);
    wire[0:0] s2732, in2732_1, in2732_2;
    wire c2732;
    assign in2732_1 = {s2220[0]};
    assign in2732_2 = {s2221[0]};
    Full_Adder FA_2732(s2732, c2732, in2732_1, in2732_2, s2219[0]);
    wire[0:0] s2733, in2733_1, in2733_2;
    wire c2733;
    assign in2733_1 = {s1566[0]};
    assign in2733_2 = {c2218};
    Full_Adder FA_2733(s2733, c2733, in2733_1, in2733_2, s1565[0]);
    wire[0:0] s2734, in2734_1, in2734_2;
    wire c2734;
    assign in2734_1 = {c2220};
    assign in2734_2 = {c2221};
    Full_Adder FA_2734(s2734, c2734, in2734_1, in2734_2, c2219);
    wire[0:0] s2735, in2735_1, in2735_2;
    wire c2735;
    assign in2735_1 = {c2223};
    assign in2735_2 = {s2224[0]};
    Full_Adder FA_2735(s2735, c2735, in2735_1, in2735_2, c2222);
    wire[0:0] s2736, in2736_1, in2736_2;
    wire c2736;
    assign in2736_1 = {s2226[0]};
    assign in2736_2 = {s2227[0]};
    Full_Adder FA_2736(s2736, c2736, in2736_1, in2736_2, s2225[0]);
    wire[0:0] s2737, in2737_1, in2737_2;
    wire c2737;
    assign in2737_1 = {s1575[0]};
    assign in2737_2 = {c2224};
    Full_Adder FA_2737(s2737, c2737, in2737_1, in2737_2, s1574[0]);
    wire[0:0] s2738, in2738_1, in2738_2;
    wire c2738;
    assign in2738_1 = {c2226};
    assign in2738_2 = {c2227};
    Full_Adder FA_2738(s2738, c2738, in2738_1, in2738_2, c2225);
    wire[0:0] s2739, in2739_1, in2739_2;
    wire c2739;
    assign in2739_1 = {c2229};
    assign in2739_2 = {s2230[0]};
    Full_Adder FA_2739(s2739, c2739, in2739_1, in2739_2, c2228);
    wire[0:0] s2740, in2740_1, in2740_2;
    wire c2740;
    assign in2740_1 = {s2232[0]};
    assign in2740_2 = {s2233[0]};
    Full_Adder FA_2740(s2740, c2740, in2740_1, in2740_2, s2231[0]);
    wire[0:0] s2741, in2741_1, in2741_2;
    wire c2741;
    assign in2741_1 = {s1584[0]};
    assign in2741_2 = {c2230};
    Full_Adder FA_2741(s2741, c2741, in2741_1, in2741_2, s1583[0]);
    wire[0:0] s2742, in2742_1, in2742_2;
    wire c2742;
    assign in2742_1 = {c2232};
    assign in2742_2 = {c2233};
    Full_Adder FA_2742(s2742, c2742, in2742_1, in2742_2, c2231);
    wire[0:0] s2743, in2743_1, in2743_2;
    wire c2743;
    assign in2743_1 = {c2235};
    assign in2743_2 = {s2236[0]};
    Full_Adder FA_2743(s2743, c2743, in2743_1, in2743_2, c2234);
    wire[0:0] s2744, in2744_1, in2744_2;
    wire c2744;
    assign in2744_1 = {s2238[0]};
    assign in2744_2 = {s2239[0]};
    Full_Adder FA_2744(s2744, c2744, in2744_1, in2744_2, s2237[0]);
    wire[0:0] s2745, in2745_1, in2745_2;
    wire c2745;
    assign in2745_1 = {s1593[0]};
    assign in2745_2 = {c2236};
    Full_Adder FA_2745(s2745, c2745, in2745_1, in2745_2, s1592[0]);
    wire[0:0] s2746, in2746_1, in2746_2;
    wire c2746;
    assign in2746_1 = {c2238};
    assign in2746_2 = {c2239};
    Full_Adder FA_2746(s2746, c2746, in2746_1, in2746_2, c2237);
    wire[0:0] s2747, in2747_1, in2747_2;
    wire c2747;
    assign in2747_1 = {c2241};
    assign in2747_2 = {s2242[0]};
    Full_Adder FA_2747(s2747, c2747, in2747_1, in2747_2, c2240);
    wire[0:0] s2748, in2748_1, in2748_2;
    wire c2748;
    assign in2748_1 = {s2244[0]};
    assign in2748_2 = {s2245[0]};
    Full_Adder FA_2748(s2748, c2748, in2748_1, in2748_2, s2243[0]);
    wire[0:0] s2749, in2749_1, in2749_2;
    wire c2749;
    assign in2749_1 = {s1602[0]};
    assign in2749_2 = {c2242};
    Full_Adder FA_2749(s2749, c2749, in2749_1, in2749_2, s1601[0]);
    wire[0:0] s2750, in2750_1, in2750_2;
    wire c2750;
    assign in2750_1 = {c2244};
    assign in2750_2 = {c2245};
    Full_Adder FA_2750(s2750, c2750, in2750_1, in2750_2, c2243);
    wire[0:0] s2751, in2751_1, in2751_2;
    wire c2751;
    assign in2751_1 = {c2247};
    assign in2751_2 = {s2248[0]};
    Full_Adder FA_2751(s2751, c2751, in2751_1, in2751_2, c2246);
    wire[0:0] s2752, in2752_1, in2752_2;
    wire c2752;
    assign in2752_1 = {s2250[0]};
    assign in2752_2 = {s2251[0]};
    Full_Adder FA_2752(s2752, c2752, in2752_1, in2752_2, s2249[0]);
    wire[0:0] s2753, in2753_1, in2753_2;
    wire c2753;
    assign in2753_1 = {s1611[0]};
    assign in2753_2 = {c2248};
    Full_Adder FA_2753(s2753, c2753, in2753_1, in2753_2, s1610[0]);
    wire[0:0] s2754, in2754_1, in2754_2;
    wire c2754;
    assign in2754_1 = {c2250};
    assign in2754_2 = {c2251};
    Full_Adder FA_2754(s2754, c2754, in2754_1, in2754_2, c2249);
    wire[0:0] s2755, in2755_1, in2755_2;
    wire c2755;
    assign in2755_1 = {c2253};
    assign in2755_2 = {s2254[0]};
    Full_Adder FA_2755(s2755, c2755, in2755_1, in2755_2, c2252);
    wire[0:0] s2756, in2756_1, in2756_2;
    wire c2756;
    assign in2756_1 = {s2256[0]};
    assign in2756_2 = {s2257[0]};
    Full_Adder FA_2756(s2756, c2756, in2756_1, in2756_2, s2255[0]);
    wire[0:0] s2757, in2757_1, in2757_2;
    wire c2757;
    assign in2757_1 = {s1620[0]};
    assign in2757_2 = {c2254};
    Full_Adder FA_2757(s2757, c2757, in2757_1, in2757_2, s1619[0]);
    wire[0:0] s2758, in2758_1, in2758_2;
    wire c2758;
    assign in2758_1 = {c2256};
    assign in2758_2 = {c2257};
    Full_Adder FA_2758(s2758, c2758, in2758_1, in2758_2, c2255);
    wire[0:0] s2759, in2759_1, in2759_2;
    wire c2759;
    assign in2759_1 = {c2259};
    assign in2759_2 = {s2260[0]};
    Full_Adder FA_2759(s2759, c2759, in2759_1, in2759_2, c2258);
    wire[0:0] s2760, in2760_1, in2760_2;
    wire c2760;
    assign in2760_1 = {s2262[0]};
    assign in2760_2 = {s2263[0]};
    Full_Adder FA_2760(s2760, c2760, in2760_1, in2760_2, s2261[0]);
    wire[0:0] s2761, in2761_1, in2761_2;
    wire c2761;
    assign in2761_1 = {s1629[0]};
    assign in2761_2 = {c2260};
    Full_Adder FA_2761(s2761, c2761, in2761_1, in2761_2, s1628[0]);
    wire[0:0] s2762, in2762_1, in2762_2;
    wire c2762;
    assign in2762_1 = {c2262};
    assign in2762_2 = {c2263};
    Full_Adder FA_2762(s2762, c2762, in2762_1, in2762_2, c2261);
    wire[0:0] s2763, in2763_1, in2763_2;
    wire c2763;
    assign in2763_1 = {c2265};
    assign in2763_2 = {s2266[0]};
    Full_Adder FA_2763(s2763, c2763, in2763_1, in2763_2, c2264);
    wire[0:0] s2764, in2764_1, in2764_2;
    wire c2764;
    assign in2764_1 = {s2268[0]};
    assign in2764_2 = {s2269[0]};
    Full_Adder FA_2764(s2764, c2764, in2764_1, in2764_2, s2267[0]);
    wire[0:0] s2765, in2765_1, in2765_2;
    wire c2765;
    assign in2765_1 = {s1638[0]};
    assign in2765_2 = {c2266};
    Full_Adder FA_2765(s2765, c2765, in2765_1, in2765_2, s1637[0]);
    wire[0:0] s2766, in2766_1, in2766_2;
    wire c2766;
    assign in2766_1 = {c2268};
    assign in2766_2 = {c2269};
    Full_Adder FA_2766(s2766, c2766, in2766_1, in2766_2, c2267);
    wire[0:0] s2767, in2767_1, in2767_2;
    wire c2767;
    assign in2767_1 = {c2271};
    assign in2767_2 = {s2272[0]};
    Full_Adder FA_2767(s2767, c2767, in2767_1, in2767_2, c2270);
    wire[0:0] s2768, in2768_1, in2768_2;
    wire c2768;
    assign in2768_1 = {s2274[0]};
    assign in2768_2 = {s2275[0]};
    Full_Adder FA_2768(s2768, c2768, in2768_1, in2768_2, s2273[0]);
    wire[0:0] s2769, in2769_1, in2769_2;
    wire c2769;
    assign in2769_1 = {s1647[0]};
    assign in2769_2 = {c2272};
    Full_Adder FA_2769(s2769, c2769, in2769_1, in2769_2, s1646[0]);
    wire[0:0] s2770, in2770_1, in2770_2;
    wire c2770;
    assign in2770_1 = {c2274};
    assign in2770_2 = {c2275};
    Full_Adder FA_2770(s2770, c2770, in2770_1, in2770_2, c2273);
    wire[0:0] s2771, in2771_1, in2771_2;
    wire c2771;
    assign in2771_1 = {c2277};
    assign in2771_2 = {s2278[0]};
    Full_Adder FA_2771(s2771, c2771, in2771_1, in2771_2, c2276);
    wire[0:0] s2772, in2772_1, in2772_2;
    wire c2772;
    assign in2772_1 = {s2280[0]};
    assign in2772_2 = {s2281[0]};
    Full_Adder FA_2772(s2772, c2772, in2772_1, in2772_2, s2279[0]);
    wire[0:0] s2773, in2773_1, in2773_2;
    wire c2773;
    assign in2773_1 = {s1656[0]};
    assign in2773_2 = {c2278};
    Full_Adder FA_2773(s2773, c2773, in2773_1, in2773_2, s1655[0]);
    wire[0:0] s2774, in2774_1, in2774_2;
    wire c2774;
    assign in2774_1 = {c2280};
    assign in2774_2 = {c2281};
    Full_Adder FA_2774(s2774, c2774, in2774_1, in2774_2, c2279);
    wire[0:0] s2775, in2775_1, in2775_2;
    wire c2775;
    assign in2775_1 = {c2283};
    assign in2775_2 = {s2284[0]};
    Full_Adder FA_2775(s2775, c2775, in2775_1, in2775_2, c2282);
    wire[0:0] s2776, in2776_1, in2776_2;
    wire c2776;
    assign in2776_1 = {s2286[0]};
    assign in2776_2 = {s2287[0]};
    Full_Adder FA_2776(s2776, c2776, in2776_1, in2776_2, s2285[0]);
    wire[0:0] s2777, in2777_1, in2777_2;
    wire c2777;
    assign in2777_1 = {s1665[0]};
    assign in2777_2 = {c2284};
    Full_Adder FA_2777(s2777, c2777, in2777_1, in2777_2, s1664[0]);
    wire[0:0] s2778, in2778_1, in2778_2;
    wire c2778;
    assign in2778_1 = {c2286};
    assign in2778_2 = {c2287};
    Full_Adder FA_2778(s2778, c2778, in2778_1, in2778_2, c2285);
    wire[0:0] s2779, in2779_1, in2779_2;
    wire c2779;
    assign in2779_1 = {c2289};
    assign in2779_2 = {s2290[0]};
    Full_Adder FA_2779(s2779, c2779, in2779_1, in2779_2, c2288);
    wire[0:0] s2780, in2780_1, in2780_2;
    wire c2780;
    assign in2780_1 = {s2292[0]};
    assign in2780_2 = {s2293[0]};
    Full_Adder FA_2780(s2780, c2780, in2780_1, in2780_2, s2291[0]);
    wire[0:0] s2781, in2781_1, in2781_2;
    wire c2781;
    assign in2781_1 = {s1674[0]};
    assign in2781_2 = {c2290};
    Full_Adder FA_2781(s2781, c2781, in2781_1, in2781_2, s1673[0]);
    wire[0:0] s2782, in2782_1, in2782_2;
    wire c2782;
    assign in2782_1 = {c2292};
    assign in2782_2 = {c2293};
    Full_Adder FA_2782(s2782, c2782, in2782_1, in2782_2, c2291);
    wire[0:0] s2783, in2783_1, in2783_2;
    wire c2783;
    assign in2783_1 = {c2295};
    assign in2783_2 = {s2296[0]};
    Full_Adder FA_2783(s2783, c2783, in2783_1, in2783_2, c2294);
    wire[0:0] s2784, in2784_1, in2784_2;
    wire c2784;
    assign in2784_1 = {s2298[0]};
    assign in2784_2 = {s2299[0]};
    Full_Adder FA_2784(s2784, c2784, in2784_1, in2784_2, s2297[0]);
    wire[0:0] s2785, in2785_1, in2785_2;
    wire c2785;
    assign in2785_1 = {s1683[0]};
    assign in2785_2 = {c2296};
    Full_Adder FA_2785(s2785, c2785, in2785_1, in2785_2, s1682[0]);
    wire[0:0] s2786, in2786_1, in2786_2;
    wire c2786;
    assign in2786_1 = {c2298};
    assign in2786_2 = {c2299};
    Full_Adder FA_2786(s2786, c2786, in2786_1, in2786_2, c2297);
    wire[0:0] s2787, in2787_1, in2787_2;
    wire c2787;
    assign in2787_1 = {c2301};
    assign in2787_2 = {s2302[0]};
    Full_Adder FA_2787(s2787, c2787, in2787_1, in2787_2, c2300);
    wire[0:0] s2788, in2788_1, in2788_2;
    wire c2788;
    assign in2788_1 = {s2304[0]};
    assign in2788_2 = {s2305[0]};
    Full_Adder FA_2788(s2788, c2788, in2788_1, in2788_2, s2303[0]);
    wire[0:0] s2789, in2789_1, in2789_2;
    wire c2789;
    assign in2789_1 = {s1692[0]};
    assign in2789_2 = {c2302};
    Full_Adder FA_2789(s2789, c2789, in2789_1, in2789_2, s1691[0]);
    wire[0:0] s2790, in2790_1, in2790_2;
    wire c2790;
    assign in2790_1 = {c2304};
    assign in2790_2 = {c2305};
    Full_Adder FA_2790(s2790, c2790, in2790_1, in2790_2, c2303);
    wire[0:0] s2791, in2791_1, in2791_2;
    wire c2791;
    assign in2791_1 = {c2307};
    assign in2791_2 = {s2308[0]};
    Full_Adder FA_2791(s2791, c2791, in2791_1, in2791_2, c2306);
    wire[0:0] s2792, in2792_1, in2792_2;
    wire c2792;
    assign in2792_1 = {s2310[0]};
    assign in2792_2 = {s2311[0]};
    Full_Adder FA_2792(s2792, c2792, in2792_1, in2792_2, s2309[0]);
    wire[0:0] s2793, in2793_1, in2793_2;
    wire c2793;
    assign in2793_1 = {s1701[0]};
    assign in2793_2 = {c2308};
    Full_Adder FA_2793(s2793, c2793, in2793_1, in2793_2, s1700[0]);
    wire[0:0] s2794, in2794_1, in2794_2;
    wire c2794;
    assign in2794_1 = {c2310};
    assign in2794_2 = {c2311};
    Full_Adder FA_2794(s2794, c2794, in2794_1, in2794_2, c2309);
    wire[0:0] s2795, in2795_1, in2795_2;
    wire c2795;
    assign in2795_1 = {c2313};
    assign in2795_2 = {s2314[0]};
    Full_Adder FA_2795(s2795, c2795, in2795_1, in2795_2, c2312);
    wire[0:0] s2796, in2796_1, in2796_2;
    wire c2796;
    assign in2796_1 = {s2316[0]};
    assign in2796_2 = {s2317[0]};
    Full_Adder FA_2796(s2796, c2796, in2796_1, in2796_2, s2315[0]);
    wire[0:0] s2797, in2797_1, in2797_2;
    wire c2797;
    assign in2797_1 = {s1710[0]};
    assign in2797_2 = {c2314};
    Full_Adder FA_2797(s2797, c2797, in2797_1, in2797_2, s1709[0]);
    wire[0:0] s2798, in2798_1, in2798_2;
    wire c2798;
    assign in2798_1 = {c2316};
    assign in2798_2 = {c2317};
    Full_Adder FA_2798(s2798, c2798, in2798_1, in2798_2, c2315);
    wire[0:0] s2799, in2799_1, in2799_2;
    wire c2799;
    assign in2799_1 = {c2319};
    assign in2799_2 = {s2320[0]};
    Full_Adder FA_2799(s2799, c2799, in2799_1, in2799_2, c2318);
    wire[0:0] s2800, in2800_1, in2800_2;
    wire c2800;
    assign in2800_1 = {s2322[0]};
    assign in2800_2 = {s2323[0]};
    Full_Adder FA_2800(s2800, c2800, in2800_1, in2800_2, s2321[0]);
    wire[0:0] s2801, in2801_1, in2801_2;
    wire c2801;
    assign in2801_1 = {s1719[0]};
    assign in2801_2 = {c2320};
    Full_Adder FA_2801(s2801, c2801, in2801_1, in2801_2, s1718[0]);
    wire[0:0] s2802, in2802_1, in2802_2;
    wire c2802;
    assign in2802_1 = {c2322};
    assign in2802_2 = {c2323};
    Full_Adder FA_2802(s2802, c2802, in2802_1, in2802_2, c2321);
    wire[0:0] s2803, in2803_1, in2803_2;
    wire c2803;
    assign in2803_1 = {c2325};
    assign in2803_2 = {s2326[0]};
    Full_Adder FA_2803(s2803, c2803, in2803_1, in2803_2, c2324);
    wire[0:0] s2804, in2804_1, in2804_2;
    wire c2804;
    assign in2804_1 = {s2328[0]};
    assign in2804_2 = {s2329[0]};
    Full_Adder FA_2804(s2804, c2804, in2804_1, in2804_2, s2327[0]);
    wire[0:0] s2805, in2805_1, in2805_2;
    wire c2805;
    assign in2805_1 = {s1728[0]};
    assign in2805_2 = {c2326};
    Full_Adder FA_2805(s2805, c2805, in2805_1, in2805_2, s1727[0]);
    wire[0:0] s2806, in2806_1, in2806_2;
    wire c2806;
    assign in2806_1 = {c2328};
    assign in2806_2 = {c2329};
    Full_Adder FA_2806(s2806, c2806, in2806_1, in2806_2, c2327);
    wire[0:0] s2807, in2807_1, in2807_2;
    wire c2807;
    assign in2807_1 = {c2331};
    assign in2807_2 = {s2332[0]};
    Full_Adder FA_2807(s2807, c2807, in2807_1, in2807_2, c2330);
    wire[0:0] s2808, in2808_1, in2808_2;
    wire c2808;
    assign in2808_1 = {s2334[0]};
    assign in2808_2 = {s2335[0]};
    Full_Adder FA_2808(s2808, c2808, in2808_1, in2808_2, s2333[0]);
    wire[0:0] s2809, in2809_1, in2809_2;
    wire c2809;
    assign in2809_1 = {s1737[0]};
    assign in2809_2 = {c2332};
    Full_Adder FA_2809(s2809, c2809, in2809_1, in2809_2, s1736[0]);
    wire[0:0] s2810, in2810_1, in2810_2;
    wire c2810;
    assign in2810_1 = {c2334};
    assign in2810_2 = {c2335};
    Full_Adder FA_2810(s2810, c2810, in2810_1, in2810_2, c2333);
    wire[0:0] s2811, in2811_1, in2811_2;
    wire c2811;
    assign in2811_1 = {c2337};
    assign in2811_2 = {s2338[0]};
    Full_Adder FA_2811(s2811, c2811, in2811_1, in2811_2, c2336);
    wire[0:0] s2812, in2812_1, in2812_2;
    wire c2812;
    assign in2812_1 = {s2340[0]};
    assign in2812_2 = {s2341[0]};
    Full_Adder FA_2812(s2812, c2812, in2812_1, in2812_2, s2339[0]);
    wire[0:0] s2813, in2813_1, in2813_2;
    wire c2813;
    assign in2813_1 = {s1746[0]};
    assign in2813_2 = {c2338};
    Full_Adder FA_2813(s2813, c2813, in2813_1, in2813_2, s1745[0]);
    wire[0:0] s2814, in2814_1, in2814_2;
    wire c2814;
    assign in2814_1 = {c2340};
    assign in2814_2 = {c2341};
    Full_Adder FA_2814(s2814, c2814, in2814_1, in2814_2, c2339);
    wire[0:0] s2815, in2815_1, in2815_2;
    wire c2815;
    assign in2815_1 = {c2343};
    assign in2815_2 = {s2344[0]};
    Full_Adder FA_2815(s2815, c2815, in2815_1, in2815_2, c2342);
    wire[0:0] s2816, in2816_1, in2816_2;
    wire c2816;
    assign in2816_1 = {s2346[0]};
    assign in2816_2 = {s2347[0]};
    Full_Adder FA_2816(s2816, c2816, in2816_1, in2816_2, s2345[0]);
    wire[0:0] s2817, in2817_1, in2817_2;
    wire c2817;
    assign in2817_1 = {s1755[0]};
    assign in2817_2 = {c2344};
    Full_Adder FA_2817(s2817, c2817, in2817_1, in2817_2, s1754[0]);
    wire[0:0] s2818, in2818_1, in2818_2;
    wire c2818;
    assign in2818_1 = {c2346};
    assign in2818_2 = {c2347};
    Full_Adder FA_2818(s2818, c2818, in2818_1, in2818_2, c2345);
    wire[0:0] s2819, in2819_1, in2819_2;
    wire c2819;
    assign in2819_1 = {c2349};
    assign in2819_2 = {s2350[0]};
    Full_Adder FA_2819(s2819, c2819, in2819_1, in2819_2, c2348);
    wire[0:0] s2820, in2820_1, in2820_2;
    wire c2820;
    assign in2820_1 = {s2352[0]};
    assign in2820_2 = {s2353[0]};
    Full_Adder FA_2820(s2820, c2820, in2820_1, in2820_2, s2351[0]);
    wire[0:0] s2821, in2821_1, in2821_2;
    wire c2821;
    assign in2821_1 = {s1764[0]};
    assign in2821_2 = {c2350};
    Full_Adder FA_2821(s2821, c2821, in2821_1, in2821_2, s1763[0]);
    wire[0:0] s2822, in2822_1, in2822_2;
    wire c2822;
    assign in2822_1 = {c2352};
    assign in2822_2 = {c2353};
    Full_Adder FA_2822(s2822, c2822, in2822_1, in2822_2, c2351);
    wire[0:0] s2823, in2823_1, in2823_2;
    wire c2823;
    assign in2823_1 = {c2355};
    assign in2823_2 = {s2356[0]};
    Full_Adder FA_2823(s2823, c2823, in2823_1, in2823_2, c2354);
    wire[0:0] s2824, in2824_1, in2824_2;
    wire c2824;
    assign in2824_1 = {s2358[0]};
    assign in2824_2 = {s2359[0]};
    Full_Adder FA_2824(s2824, c2824, in2824_1, in2824_2, s2357[0]);
    wire[0:0] s2825, in2825_1, in2825_2;
    wire c2825;
    assign in2825_1 = {s1773[0]};
    assign in2825_2 = {c2356};
    Full_Adder FA_2825(s2825, c2825, in2825_1, in2825_2, s1772[0]);
    wire[0:0] s2826, in2826_1, in2826_2;
    wire c2826;
    assign in2826_1 = {c2358};
    assign in2826_2 = {c2359};
    Full_Adder FA_2826(s2826, c2826, in2826_1, in2826_2, c2357);
    wire[0:0] s2827, in2827_1, in2827_2;
    wire c2827;
    assign in2827_1 = {c2361};
    assign in2827_2 = {s2362[0]};
    Full_Adder FA_2827(s2827, c2827, in2827_1, in2827_2, c2360);
    wire[0:0] s2828, in2828_1, in2828_2;
    wire c2828;
    assign in2828_1 = {s2364[0]};
    assign in2828_2 = {s2365[0]};
    Full_Adder FA_2828(s2828, c2828, in2828_1, in2828_2, s2363[0]);
    wire[0:0] s2829, in2829_1, in2829_2;
    wire c2829;
    assign in2829_1 = {s1782[0]};
    assign in2829_2 = {c2362};
    Full_Adder FA_2829(s2829, c2829, in2829_1, in2829_2, s1781[0]);
    wire[0:0] s2830, in2830_1, in2830_2;
    wire c2830;
    assign in2830_1 = {c2364};
    assign in2830_2 = {c2365};
    Full_Adder FA_2830(s2830, c2830, in2830_1, in2830_2, c2363);
    wire[0:0] s2831, in2831_1, in2831_2;
    wire c2831;
    assign in2831_1 = {c2367};
    assign in2831_2 = {s2368[0]};
    Full_Adder FA_2831(s2831, c2831, in2831_1, in2831_2, c2366);
    wire[0:0] s2832, in2832_1, in2832_2;
    wire c2832;
    assign in2832_1 = {s2370[0]};
    assign in2832_2 = {s2371[0]};
    Full_Adder FA_2832(s2832, c2832, in2832_1, in2832_2, s2369[0]);
    wire[0:0] s2833, in2833_1, in2833_2;
    wire c2833;
    assign in2833_1 = {s1791[0]};
    assign in2833_2 = {c2368};
    Full_Adder FA_2833(s2833, c2833, in2833_1, in2833_2, s1790[0]);
    wire[0:0] s2834, in2834_1, in2834_2;
    wire c2834;
    assign in2834_1 = {c2370};
    assign in2834_2 = {c2371};
    Full_Adder FA_2834(s2834, c2834, in2834_1, in2834_2, c2369);
    wire[0:0] s2835, in2835_1, in2835_2;
    wire c2835;
    assign in2835_1 = {c2373};
    assign in2835_2 = {s2374[0]};
    Full_Adder FA_2835(s2835, c2835, in2835_1, in2835_2, c2372);
    wire[0:0] s2836, in2836_1, in2836_2;
    wire c2836;
    assign in2836_1 = {s2376[0]};
    assign in2836_2 = {s2377[0]};
    Full_Adder FA_2836(s2836, c2836, in2836_1, in2836_2, s2375[0]);
    wire[0:0] s2837, in2837_1, in2837_2;
    wire c2837;
    assign in2837_1 = {s1800[0]};
    assign in2837_2 = {c2374};
    Full_Adder FA_2837(s2837, c2837, in2837_1, in2837_2, s1799[0]);
    wire[0:0] s2838, in2838_1, in2838_2;
    wire c2838;
    assign in2838_1 = {c2376};
    assign in2838_2 = {c2377};
    Full_Adder FA_2838(s2838, c2838, in2838_1, in2838_2, c2375);
    wire[0:0] s2839, in2839_1, in2839_2;
    wire c2839;
    assign in2839_1 = {c2379};
    assign in2839_2 = {s2380[0]};
    Full_Adder FA_2839(s2839, c2839, in2839_1, in2839_2, c2378);
    wire[0:0] s2840, in2840_1, in2840_2;
    wire c2840;
    assign in2840_1 = {s2382[0]};
    assign in2840_2 = {s2383[0]};
    Full_Adder FA_2840(s2840, c2840, in2840_1, in2840_2, s2381[0]);
    wire[0:0] s2841, in2841_1, in2841_2;
    wire c2841;
    assign in2841_1 = {s1809[0]};
    assign in2841_2 = {c2380};
    Full_Adder FA_2841(s2841, c2841, in2841_1, in2841_2, s1808[0]);
    wire[0:0] s2842, in2842_1, in2842_2;
    wire c2842;
    assign in2842_1 = {c2382};
    assign in2842_2 = {c2383};
    Full_Adder FA_2842(s2842, c2842, in2842_1, in2842_2, c2381);
    wire[0:0] s2843, in2843_1, in2843_2;
    wire c2843;
    assign in2843_1 = {c2385};
    assign in2843_2 = {s2386[0]};
    Full_Adder FA_2843(s2843, c2843, in2843_1, in2843_2, c2384);
    wire[0:0] s2844, in2844_1, in2844_2;
    wire c2844;
    assign in2844_1 = {s2388[0]};
    assign in2844_2 = {s2389[0]};
    Full_Adder FA_2844(s2844, c2844, in2844_1, in2844_2, s2387[0]);
    wire[0:0] s2845, in2845_1, in2845_2;
    wire c2845;
    assign in2845_1 = {s1818[0]};
    assign in2845_2 = {c2386};
    Full_Adder FA_2845(s2845, c2845, in2845_1, in2845_2, s1817[0]);
    wire[0:0] s2846, in2846_1, in2846_2;
    wire c2846;
    assign in2846_1 = {c2388};
    assign in2846_2 = {c2389};
    Full_Adder FA_2846(s2846, c2846, in2846_1, in2846_2, c2387);
    wire[0:0] s2847, in2847_1, in2847_2;
    wire c2847;
    assign in2847_1 = {c2391};
    assign in2847_2 = {s2392[0]};
    Full_Adder FA_2847(s2847, c2847, in2847_1, in2847_2, c2390);
    wire[0:0] s2848, in2848_1, in2848_2;
    wire c2848;
    assign in2848_1 = {s2394[0]};
    assign in2848_2 = {s2395[0]};
    Full_Adder FA_2848(s2848, c2848, in2848_1, in2848_2, s2393[0]);
    wire[0:0] s2849, in2849_1, in2849_2;
    wire c2849;
    assign in2849_1 = {s1827[0]};
    assign in2849_2 = {c2392};
    Full_Adder FA_2849(s2849, c2849, in2849_1, in2849_2, s1826[0]);
    wire[0:0] s2850, in2850_1, in2850_2;
    wire c2850;
    assign in2850_1 = {c2394};
    assign in2850_2 = {c2395};
    Full_Adder FA_2850(s2850, c2850, in2850_1, in2850_2, c2393);
    wire[0:0] s2851, in2851_1, in2851_2;
    wire c2851;
    assign in2851_1 = {c2397};
    assign in2851_2 = {s2398[0]};
    Full_Adder FA_2851(s2851, c2851, in2851_1, in2851_2, c2396);
    wire[0:0] s2852, in2852_1, in2852_2;
    wire c2852;
    assign in2852_1 = {s2400[0]};
    assign in2852_2 = {s2401[0]};
    Full_Adder FA_2852(s2852, c2852, in2852_1, in2852_2, s2399[0]);
    wire[0:0] s2853, in2853_1, in2853_2;
    wire c2853;
    assign in2853_1 = {s1836[0]};
    assign in2853_2 = {c2398};
    Full_Adder FA_2853(s2853, c2853, in2853_1, in2853_2, s1835[0]);
    wire[0:0] s2854, in2854_1, in2854_2;
    wire c2854;
    assign in2854_1 = {c2400};
    assign in2854_2 = {c2401};
    Full_Adder FA_2854(s2854, c2854, in2854_1, in2854_2, c2399);
    wire[0:0] s2855, in2855_1, in2855_2;
    wire c2855;
    assign in2855_1 = {c2403};
    assign in2855_2 = {s2404[0]};
    Full_Adder FA_2855(s2855, c2855, in2855_1, in2855_2, c2402);
    wire[0:0] s2856, in2856_1, in2856_2;
    wire c2856;
    assign in2856_1 = {s2406[0]};
    assign in2856_2 = {s2407[0]};
    Full_Adder FA_2856(s2856, c2856, in2856_1, in2856_2, s2405[0]);
    wire[0:0] s2857, in2857_1, in2857_2;
    wire c2857;
    assign in2857_1 = {s1845[0]};
    assign in2857_2 = {c2404};
    Full_Adder FA_2857(s2857, c2857, in2857_1, in2857_2, s1844[0]);
    wire[0:0] s2858, in2858_1, in2858_2;
    wire c2858;
    assign in2858_1 = {c2406};
    assign in2858_2 = {c2407};
    Full_Adder FA_2858(s2858, c2858, in2858_1, in2858_2, c2405);
    wire[0:0] s2859, in2859_1, in2859_2;
    wire c2859;
    assign in2859_1 = {c2409};
    assign in2859_2 = {s2410[0]};
    Full_Adder FA_2859(s2859, c2859, in2859_1, in2859_2, c2408);
    wire[0:0] s2860, in2860_1, in2860_2;
    wire c2860;
    assign in2860_1 = {s2412[0]};
    assign in2860_2 = {s2413[0]};
    Full_Adder FA_2860(s2860, c2860, in2860_1, in2860_2, s2411[0]);
    wire[0:0] s2861, in2861_1, in2861_2;
    wire c2861;
    assign in2861_1 = {s1854[0]};
    assign in2861_2 = {c2410};
    Full_Adder FA_2861(s2861, c2861, in2861_1, in2861_2, s1853[0]);
    wire[0:0] s2862, in2862_1, in2862_2;
    wire c2862;
    assign in2862_1 = {c2412};
    assign in2862_2 = {c2413};
    Full_Adder FA_2862(s2862, c2862, in2862_1, in2862_2, c2411);
    wire[0:0] s2863, in2863_1, in2863_2;
    wire c2863;
    assign in2863_1 = {c2415};
    assign in2863_2 = {s2416[0]};
    Full_Adder FA_2863(s2863, c2863, in2863_1, in2863_2, c2414);
    wire[0:0] s2864, in2864_1, in2864_2;
    wire c2864;
    assign in2864_1 = {s2418[0]};
    assign in2864_2 = {s2419[0]};
    Full_Adder FA_2864(s2864, c2864, in2864_1, in2864_2, s2417[0]);
    wire[0:0] s2865, in2865_1, in2865_2;
    wire c2865;
    assign in2865_1 = {s1863[0]};
    assign in2865_2 = {c2416};
    Full_Adder FA_2865(s2865, c2865, in2865_1, in2865_2, s1862[0]);
    wire[0:0] s2866, in2866_1, in2866_2;
    wire c2866;
    assign in2866_1 = {c2418};
    assign in2866_2 = {c2419};
    Full_Adder FA_2866(s2866, c2866, in2866_1, in2866_2, c2417);
    wire[0:0] s2867, in2867_1, in2867_2;
    wire c2867;
    assign in2867_1 = {c2421};
    assign in2867_2 = {s2422[0]};
    Full_Adder FA_2867(s2867, c2867, in2867_1, in2867_2, c2420);
    wire[0:0] s2868, in2868_1, in2868_2;
    wire c2868;
    assign in2868_1 = {s2424[0]};
    assign in2868_2 = {s2425[0]};
    Full_Adder FA_2868(s2868, c2868, in2868_1, in2868_2, s2423[0]);
    wire[0:0] s2869, in2869_1, in2869_2;
    wire c2869;
    assign in2869_1 = {s1872[0]};
    assign in2869_2 = {c2422};
    Full_Adder FA_2869(s2869, c2869, in2869_1, in2869_2, s1871[0]);
    wire[0:0] s2870, in2870_1, in2870_2;
    wire c2870;
    assign in2870_1 = {c2424};
    assign in2870_2 = {c2425};
    Full_Adder FA_2870(s2870, c2870, in2870_1, in2870_2, c2423);
    wire[0:0] s2871, in2871_1, in2871_2;
    wire c2871;
    assign in2871_1 = {c2427};
    assign in2871_2 = {s2428[0]};
    Full_Adder FA_2871(s2871, c2871, in2871_1, in2871_2, c2426);
    wire[0:0] s2872, in2872_1, in2872_2;
    wire c2872;
    assign in2872_1 = {s2430[0]};
    assign in2872_2 = {s2431[0]};
    Full_Adder FA_2872(s2872, c2872, in2872_1, in2872_2, s2429[0]);
    wire[0:0] s2873, in2873_1, in2873_2;
    wire c2873;
    assign in2873_1 = {s1881[0]};
    assign in2873_2 = {c2428};
    Full_Adder FA_2873(s2873, c2873, in2873_1, in2873_2, s1880[0]);
    wire[0:0] s2874, in2874_1, in2874_2;
    wire c2874;
    assign in2874_1 = {c2430};
    assign in2874_2 = {c2431};
    Full_Adder FA_2874(s2874, c2874, in2874_1, in2874_2, c2429);
    wire[0:0] s2875, in2875_1, in2875_2;
    wire c2875;
    assign in2875_1 = {c2433};
    assign in2875_2 = {s2434[0]};
    Full_Adder FA_2875(s2875, c2875, in2875_1, in2875_2, c2432);
    wire[0:0] s2876, in2876_1, in2876_2;
    wire c2876;
    assign in2876_1 = {s2436[0]};
    assign in2876_2 = {s2437[0]};
    Full_Adder FA_2876(s2876, c2876, in2876_1, in2876_2, s2435[0]);
    wire[0:0] s2877, in2877_1, in2877_2;
    wire c2877;
    assign in2877_1 = {s1890[0]};
    assign in2877_2 = {c2434};
    Full_Adder FA_2877(s2877, c2877, in2877_1, in2877_2, s1889[0]);
    wire[0:0] s2878, in2878_1, in2878_2;
    wire c2878;
    assign in2878_1 = {c2436};
    assign in2878_2 = {c2437};
    Full_Adder FA_2878(s2878, c2878, in2878_1, in2878_2, c2435);
    wire[0:0] s2879, in2879_1, in2879_2;
    wire c2879;
    assign in2879_1 = {c2439};
    assign in2879_2 = {s2440[0]};
    Full_Adder FA_2879(s2879, c2879, in2879_1, in2879_2, c2438);
    wire[0:0] s2880, in2880_1, in2880_2;
    wire c2880;
    assign in2880_1 = {s2442[0]};
    assign in2880_2 = {s2443[0]};
    Full_Adder FA_2880(s2880, c2880, in2880_1, in2880_2, s2441[0]);
    wire[0:0] s2881, in2881_1, in2881_2;
    wire c2881;
    assign in2881_1 = {s1899[0]};
    assign in2881_2 = {c2440};
    Full_Adder FA_2881(s2881, c2881, in2881_1, in2881_2, s1898[0]);
    wire[0:0] s2882, in2882_1, in2882_2;
    wire c2882;
    assign in2882_1 = {c2442};
    assign in2882_2 = {c2443};
    Full_Adder FA_2882(s2882, c2882, in2882_1, in2882_2, c2441);
    wire[0:0] s2883, in2883_1, in2883_2;
    wire c2883;
    assign in2883_1 = {c2445};
    assign in2883_2 = {s2446[0]};
    Full_Adder FA_2883(s2883, c2883, in2883_1, in2883_2, c2444);
    wire[0:0] s2884, in2884_1, in2884_2;
    wire c2884;
    assign in2884_1 = {s2448[0]};
    assign in2884_2 = {s2449[0]};
    Full_Adder FA_2884(s2884, c2884, in2884_1, in2884_2, s2447[0]);
    wire[0:0] s2885, in2885_1, in2885_2;
    wire c2885;
    assign in2885_1 = {s1908[0]};
    assign in2885_2 = {c2446};
    Full_Adder FA_2885(s2885, c2885, in2885_1, in2885_2, s1907[0]);
    wire[0:0] s2886, in2886_1, in2886_2;
    wire c2886;
    assign in2886_1 = {c2448};
    assign in2886_2 = {c2449};
    Full_Adder FA_2886(s2886, c2886, in2886_1, in2886_2, c2447);
    wire[0:0] s2887, in2887_1, in2887_2;
    wire c2887;
    assign in2887_1 = {c2451};
    assign in2887_2 = {s2452[0]};
    Full_Adder FA_2887(s2887, c2887, in2887_1, in2887_2, c2450);
    wire[0:0] s2888, in2888_1, in2888_2;
    wire c2888;
    assign in2888_1 = {s2454[0]};
    assign in2888_2 = {s2455[0]};
    Full_Adder FA_2888(s2888, c2888, in2888_1, in2888_2, s2453[0]);
    wire[0:0] s2889, in2889_1, in2889_2;
    wire c2889;
    assign in2889_1 = {s1917[0]};
    assign in2889_2 = {c2452};
    Full_Adder FA_2889(s2889, c2889, in2889_1, in2889_2, s1916[0]);
    wire[0:0] s2890, in2890_1, in2890_2;
    wire c2890;
    assign in2890_1 = {c2454};
    assign in2890_2 = {c2455};
    Full_Adder FA_2890(s2890, c2890, in2890_1, in2890_2, c2453);
    wire[0:0] s2891, in2891_1, in2891_2;
    wire c2891;
    assign in2891_1 = {c2457};
    assign in2891_2 = {s2458[0]};
    Full_Adder FA_2891(s2891, c2891, in2891_1, in2891_2, c2456);
    wire[0:0] s2892, in2892_1, in2892_2;
    wire c2892;
    assign in2892_1 = {s2460[0]};
    assign in2892_2 = {s2461[0]};
    Full_Adder FA_2892(s2892, c2892, in2892_1, in2892_2, s2459[0]);
    wire[0:0] s2893, in2893_1, in2893_2;
    wire c2893;
    assign in2893_1 = {s1926[0]};
    assign in2893_2 = {c2458};
    Full_Adder FA_2893(s2893, c2893, in2893_1, in2893_2, s1925[0]);
    wire[0:0] s2894, in2894_1, in2894_2;
    wire c2894;
    assign in2894_1 = {c2460};
    assign in2894_2 = {c2461};
    Full_Adder FA_2894(s2894, c2894, in2894_1, in2894_2, c2459);
    wire[0:0] s2895, in2895_1, in2895_2;
    wire c2895;
    assign in2895_1 = {c2463};
    assign in2895_2 = {s2464[0]};
    Full_Adder FA_2895(s2895, c2895, in2895_1, in2895_2, c2462);
    wire[0:0] s2896, in2896_1, in2896_2;
    wire c2896;
    assign in2896_1 = {s2466[0]};
    assign in2896_2 = {s2467[0]};
    Full_Adder FA_2896(s2896, c2896, in2896_1, in2896_2, s2465[0]);
    wire[0:0] s2897, in2897_1, in2897_2;
    wire c2897;
    assign in2897_1 = {s1935[0]};
    assign in2897_2 = {c2464};
    Full_Adder FA_2897(s2897, c2897, in2897_1, in2897_2, s1934[0]);
    wire[0:0] s2898, in2898_1, in2898_2;
    wire c2898;
    assign in2898_1 = {c2466};
    assign in2898_2 = {c2467};
    Full_Adder FA_2898(s2898, c2898, in2898_1, in2898_2, c2465);
    wire[0:0] s2899, in2899_1, in2899_2;
    wire c2899;
    assign in2899_1 = {c2469};
    assign in2899_2 = {s2470[0]};
    Full_Adder FA_2899(s2899, c2899, in2899_1, in2899_2, c2468);
    wire[0:0] s2900, in2900_1, in2900_2;
    wire c2900;
    assign in2900_1 = {s2472[0]};
    assign in2900_2 = {s2473[0]};
    Full_Adder FA_2900(s2900, c2900, in2900_1, in2900_2, s2471[0]);
    wire[0:0] s2901, in2901_1, in2901_2;
    wire c2901;
    assign in2901_1 = {s1944[0]};
    assign in2901_2 = {c2470};
    Full_Adder FA_2901(s2901, c2901, in2901_1, in2901_2, s1943[0]);
    wire[0:0] s2902, in2902_1, in2902_2;
    wire c2902;
    assign in2902_1 = {c2472};
    assign in2902_2 = {c2473};
    Full_Adder FA_2902(s2902, c2902, in2902_1, in2902_2, c2471);
    wire[0:0] s2903, in2903_1, in2903_2;
    wire c2903;
    assign in2903_1 = {c2475};
    assign in2903_2 = {s2476[0]};
    Full_Adder FA_2903(s2903, c2903, in2903_1, in2903_2, c2474);
    wire[0:0] s2904, in2904_1, in2904_2;
    wire c2904;
    assign in2904_1 = {s2478[0]};
    assign in2904_2 = {s2479[0]};
    Full_Adder FA_2904(s2904, c2904, in2904_1, in2904_2, s2477[0]);
    wire[0:0] s2905, in2905_1, in2905_2;
    wire c2905;
    assign in2905_1 = {s1952[0]};
    assign in2905_2 = {c2476};
    Full_Adder FA_2905(s2905, c2905, in2905_1, in2905_2, s1951[0]);
    wire[0:0] s2906, in2906_1, in2906_2;
    wire c2906;
    assign in2906_1 = {c2478};
    assign in2906_2 = {c2479};
    Full_Adder FA_2906(s2906, c2906, in2906_1, in2906_2, c2477);
    wire[0:0] s2907, in2907_1, in2907_2;
    wire c2907;
    assign in2907_1 = {c2481};
    assign in2907_2 = {s2482[0]};
    Full_Adder FA_2907(s2907, c2907, in2907_1, in2907_2, c2480);
    wire[0:0] s2908, in2908_1, in2908_2;
    wire c2908;
    assign in2908_1 = {s2484[0]};
    assign in2908_2 = {s2485[0]};
    Full_Adder FA_2908(s2908, c2908, in2908_1, in2908_2, s2483[0]);
    wire[0:0] s2909, in2909_1, in2909_2;
    wire c2909;
    assign in2909_1 = {s1959[0]};
    assign in2909_2 = {c2482};
    Full_Adder FA_2909(s2909, c2909, in2909_1, in2909_2, s1958[0]);
    wire[0:0] s2910, in2910_1, in2910_2;
    wire c2910;
    assign in2910_1 = {c2484};
    assign in2910_2 = {c2485};
    Full_Adder FA_2910(s2910, c2910, in2910_1, in2910_2, c2483);
    wire[0:0] s2911, in2911_1, in2911_2;
    wire c2911;
    assign in2911_1 = {c2487};
    assign in2911_2 = {s2488[0]};
    Full_Adder FA_2911(s2911, c2911, in2911_1, in2911_2, c2486);
    wire[0:0] s2912, in2912_1, in2912_2;
    wire c2912;
    assign in2912_1 = {s2490[0]};
    assign in2912_2 = {s2491[0]};
    Full_Adder FA_2912(s2912, c2912, in2912_1, in2912_2, s2489[0]);
    wire[0:0] s2913, in2913_1, in2913_2;
    wire c2913;
    assign in2913_1 = {s1965[0]};
    assign in2913_2 = {c2488};
    Full_Adder FA_2913(s2913, c2913, in2913_1, in2913_2, s1964[0]);
    wire[0:0] s2914, in2914_1, in2914_2;
    wire c2914;
    assign in2914_1 = {c2490};
    assign in2914_2 = {c2491};
    Full_Adder FA_2914(s2914, c2914, in2914_1, in2914_2, c2489);
    wire[0:0] s2915, in2915_1, in2915_2;
    wire c2915;
    assign in2915_1 = {c2493};
    assign in2915_2 = {s2494[0]};
    Full_Adder FA_2915(s2915, c2915, in2915_1, in2915_2, c2492);
    wire[0:0] s2916, in2916_1, in2916_2;
    wire c2916;
    assign in2916_1 = {s2496[0]};
    assign in2916_2 = {s2497[0]};
    Full_Adder FA_2916(s2916, c2916, in2916_1, in2916_2, s2495[0]);
    wire[0:0] s2917, in2917_1, in2917_2;
    wire c2917;
    assign in2917_1 = {s1970[0]};
    assign in2917_2 = {c2494};
    Full_Adder FA_2917(s2917, c2917, in2917_1, in2917_2, s1969[0]);
    wire[0:0] s2918, in2918_1, in2918_2;
    wire c2918;
    assign in2918_1 = {c2496};
    assign in2918_2 = {c2497};
    Full_Adder FA_2918(s2918, c2918, in2918_1, in2918_2, c2495);
    wire[0:0] s2919, in2919_1, in2919_2;
    wire c2919;
    assign in2919_1 = {c2499};
    assign in2919_2 = {s2500[0]};
    Full_Adder FA_2919(s2919, c2919, in2919_1, in2919_2, c2498);
    wire[0:0] s2920, in2920_1, in2920_2;
    wire c2920;
    assign in2920_1 = {s2502[0]};
    assign in2920_2 = {s2503[0]};
    Full_Adder FA_2920(s2920, c2920, in2920_1, in2920_2, s2501[0]);
    wire[0:0] s2921, in2921_1, in2921_2;
    wire c2921;
    assign in2921_1 = {s1974[0]};
    assign in2921_2 = {c2500};
    Full_Adder FA_2921(s2921, c2921, in2921_1, in2921_2, s1973[0]);
    wire[0:0] s2922, in2922_1, in2922_2;
    wire c2922;
    assign in2922_1 = {c2502};
    assign in2922_2 = {c2503};
    Full_Adder FA_2922(s2922, c2922, in2922_1, in2922_2, c2501);
    wire[0:0] s2923, in2923_1, in2923_2;
    wire c2923;
    assign in2923_1 = {c2505};
    assign in2923_2 = {s2506[0]};
    Full_Adder FA_2923(s2923, c2923, in2923_1, in2923_2, c2504);
    wire[0:0] s2924, in2924_1, in2924_2;
    wire c2924;
    assign in2924_1 = {s2508[0]};
    assign in2924_2 = {s2509[0]};
    Full_Adder FA_2924(s2924, c2924, in2924_1, in2924_2, s2507[0]);
    wire[0:0] s2925, in2925_1, in2925_2;
    wire c2925;
    assign in2925_1 = {s1977[0]};
    assign in2925_2 = {c2506};
    Full_Adder FA_2925(s2925, c2925, in2925_1, in2925_2, s1976[0]);
    wire[0:0] s2926, in2926_1, in2926_2;
    wire c2926;
    assign in2926_1 = {c2508};
    assign in2926_2 = {c2509};
    Full_Adder FA_2926(s2926, c2926, in2926_1, in2926_2, c2507);
    wire[0:0] s2927, in2927_1, in2927_2;
    wire c2927;
    assign in2927_1 = {c2511};
    assign in2927_2 = {s2512[0]};
    Full_Adder FA_2927(s2927, c2927, in2927_1, in2927_2, c2510);
    wire[0:0] s2928, in2928_1, in2928_2;
    wire c2928;
    assign in2928_1 = {s2514[0]};
    assign in2928_2 = {s2515[0]};
    Full_Adder FA_2928(s2928, c2928, in2928_1, in2928_2, s2513[0]);
    wire[0:0] s2929, in2929_1, in2929_2;
    wire c2929;
    assign in2929_1 = {s1979[0]};
    assign in2929_2 = {c2512};
    Full_Adder FA_2929(s2929, c2929, in2929_1, in2929_2, s1978[0]);
    wire[0:0] s2930, in2930_1, in2930_2;
    wire c2930;
    assign in2930_1 = {c2514};
    assign in2930_2 = {c2515};
    Full_Adder FA_2930(s2930, c2930, in2930_1, in2930_2, c2513);
    wire[0:0] s2931, in2931_1, in2931_2;
    wire c2931;
    assign in2931_1 = {c2517};
    assign in2931_2 = {s2518[0]};
    Full_Adder FA_2931(s2931, c2931, in2931_1, in2931_2, c2516);
    wire[0:0] s2932, in2932_1, in2932_2;
    wire c2932;
    assign in2932_1 = {s2520[0]};
    assign in2932_2 = {s2521[0]};
    Full_Adder FA_2932(s2932, c2932, in2932_1, in2932_2, s2519[0]);
    wire[0:0] s2933, in2933_1, in2933_2;
    wire c2933;
    assign in2933_1 = {s1980[0]};
    assign in2933_2 = {c2518};
    Full_Adder FA_2933(s2933, c2933, in2933_1, in2933_2, c1979);
    wire[0:0] s2934, in2934_1, in2934_2;
    wire c2934;
    assign in2934_1 = {c2520};
    assign in2934_2 = {c2521};
    Full_Adder FA_2934(s2934, c2934, in2934_1, in2934_2, c2519);
    wire[0:0] s2935, in2935_1, in2935_2;
    wire c2935;
    assign in2935_1 = {c2523};
    assign in2935_2 = {s2524[0]};
    Full_Adder FA_2935(s2935, c2935, in2935_1, in2935_2, c2522);
    wire[0:0] s2936, in2936_1, in2936_2;
    wire c2936;
    assign in2936_1 = {s2526[0]};
    assign in2936_2 = {s2527[0]};
    Full_Adder FA_2936(s2936, c2936, in2936_1, in2936_2, s2525[0]);
    wire[0:0] s2937, in2937_1, in2937_2;
    wire c2937;
    assign in2937_1 = {c1980};
    assign in2937_2 = {c2524};
    Full_Adder FA_2937(s2937, c2937, in2937_1, in2937_2, pp63[45]);
    wire[0:0] s2938, in2938_1, in2938_2;
    wire c2938;
    assign in2938_1 = {c2526};
    assign in2938_2 = {c2527};
    Full_Adder FA_2938(s2938, c2938, in2938_1, in2938_2, c2525);
    wire[0:0] s2939, in2939_1, in2939_2;
    wire c2939;
    assign in2939_1 = {c2529};
    assign in2939_2 = {s2530[0]};
    Full_Adder FA_2939(s2939, c2939, in2939_1, in2939_2, c2528);
    wire[0:0] s2940, in2940_1, in2940_2;
    wire c2940;
    assign in2940_1 = {s2532[0]};
    assign in2940_2 = {s2533[0]};
    Full_Adder FA_2940(s2940, c2940, in2940_1, in2940_2, s2531[0]);
    wire[0:0] s2941, in2941_1, in2941_2;
    wire c2941;
    assign in2941_1 = {pp62[47]};
    assign in2941_2 = {pp63[46]};
    Full_Adder FA_2941(s2941, c2941, in2941_1, in2941_2, pp61[48]);
    wire[0:0] s2942, in2942_1, in2942_2;
    wire c2942;
    assign in2942_1 = {c2531};
    assign in2942_2 = {c2532};
    Full_Adder FA_2942(s2942, c2942, in2942_1, in2942_2, c2530);
    wire[0:0] s2943, in2943_1, in2943_2;
    wire c2943;
    assign in2943_1 = {c2534};
    assign in2943_2 = {c2535};
    Full_Adder FA_2943(s2943, c2943, in2943_1, in2943_2, c2533);
    wire[0:0] s2944, in2944_1, in2944_2;
    wire c2944;
    assign in2944_1 = {s2537[0]};
    assign in2944_2 = {s2538[0]};
    Full_Adder FA_2944(s2944, c2944, in2944_1, in2944_2, s2536[0]);
    wire[0:0] s2945, in2945_1, in2945_2;
    wire c2945;
    assign in2945_1 = {pp60[50]};
    assign in2945_2 = {pp61[49]};
    Full_Adder FA_2945(s2945, c2945, in2945_1, in2945_2, pp59[51]);
    wire[0:0] s2946, in2946_1, in2946_2;
    wire c2946;
    assign in2946_1 = {pp63[47]};
    assign in2946_2 = {c2536};
    Full_Adder FA_2946(s2946, c2946, in2946_1, in2946_2, pp62[48]);
    wire[0:0] s2947, in2947_1, in2947_2;
    wire c2947;
    assign in2947_1 = {c2538};
    assign in2947_2 = {c2539};
    Full_Adder FA_2947(s2947, c2947, in2947_1, in2947_2, c2537);
    wire[0:0] s2948, in2948_1, in2948_2;
    wire c2948;
    assign in2948_1 = {s2541[0]};
    assign in2948_2 = {s2542[0]};
    Full_Adder FA_2948(s2948, c2948, in2948_1, in2948_2, c2540);
    wire[0:0] s2949, in2949_1, in2949_2;
    wire c2949;
    assign in2949_1 = {pp58[53]};
    assign in2949_2 = {pp59[52]};
    Full_Adder FA_2949(s2949, c2949, in2949_1, in2949_2, pp57[54]);
    wire[0:0] s2950, in2950_1, in2950_2;
    wire c2950;
    assign in2950_1 = {pp61[50]};
    assign in2950_2 = {pp62[49]};
    Full_Adder FA_2950(s2950, c2950, in2950_1, in2950_2, pp60[51]);
    wire[0:0] s2951, in2951_1, in2951_2;
    wire c2951;
    assign in2951_1 = {c2541};
    assign in2951_2 = {c2542};
    Full_Adder FA_2951(s2951, c2951, in2951_1, in2951_2, pp63[48]);
    wire[0:0] s2952, in2952_1, in2952_2;
    wire c2952;
    assign in2952_1 = {c2544};
    assign in2952_2 = {s2545[0]};
    Full_Adder FA_2952(s2952, c2952, in2952_1, in2952_2, c2543);
    wire[0:0] s2953, in2953_1, in2953_2;
    wire c2953;
    assign in2953_1 = {pp56[56]};
    assign in2953_2 = {pp57[55]};
    Full_Adder FA_2953(s2953, c2953, in2953_1, in2953_2, pp55[57]);
    wire[0:0] s2954, in2954_1, in2954_2;
    wire c2954;
    assign in2954_1 = {pp59[53]};
    assign in2954_2 = {pp60[52]};
    Full_Adder FA_2954(s2954, c2954, in2954_1, in2954_2, pp58[54]);
    wire[0:0] s2955, in2955_1, in2955_2;
    wire c2955;
    assign in2955_1 = {pp62[50]};
    assign in2955_2 = {pp63[49]};
    Full_Adder FA_2955(s2955, c2955, in2955_1, in2955_2, pp61[51]);
    wire[0:0] s2956, in2956_1, in2956_2;
    wire c2956;
    assign in2956_1 = {c2546};
    assign in2956_2 = {c2547};
    Full_Adder FA_2956(s2956, c2956, in2956_1, in2956_2, c2545);
    wire[0:0] s2957, in2957_1, in2957_2;
    wire c2957;
    assign in2957_1 = {pp54[59]};
    assign in2957_2 = {pp55[58]};
    Full_Adder FA_2957(s2957, c2957, in2957_1, in2957_2, pp53[60]);
    wire[0:0] s2958, in2958_1, in2958_2;
    wire c2958;
    assign in2958_1 = {pp57[56]};
    assign in2958_2 = {pp58[55]};
    Full_Adder FA_2958(s2958, c2958, in2958_1, in2958_2, pp56[57]);
    wire[0:0] s2959, in2959_1, in2959_2;
    wire c2959;
    assign in2959_1 = {pp60[53]};
    assign in2959_2 = {pp61[52]};
    Full_Adder FA_2959(s2959, c2959, in2959_1, in2959_2, pp59[54]);
    wire[0:0] s2960, in2960_1, in2960_2;
    wire c2960;
    assign in2960_1 = {pp63[50]};
    assign in2960_2 = {c2548};
    Full_Adder FA_2960(s2960, c2960, in2960_1, in2960_2, pp62[51]);
    wire[0:0] s2961, in2961_1, in2961_2;
    wire c2961;
    assign in2961_1 = {pp52[62]};
    assign in2961_2 = {pp53[61]};
    Full_Adder FA_2961(s2961, c2961, in2961_1, in2961_2, pp51[63]);
    wire[0:0] s2962, in2962_1, in2962_2;
    wire c2962;
    assign in2962_1 = {pp55[59]};
    assign in2962_2 = {pp56[58]};
    Full_Adder FA_2962(s2962, c2962, in2962_1, in2962_2, pp54[60]);
    wire[0:0] s2963, in2963_1, in2963_2;
    wire c2963;
    assign in2963_1 = {pp58[56]};
    assign in2963_2 = {pp59[55]};
    Full_Adder FA_2963(s2963, c2963, in2963_1, in2963_2, pp57[57]);
    wire[0:0] s2964, in2964_1, in2964_2;
    wire c2964;
    assign in2964_1 = {pp61[53]};
    assign in2964_2 = {pp62[52]};
    Full_Adder FA_2964(s2964, c2964, in2964_1, in2964_2, pp60[54]);
    wire[0:0] s2965, in2965_1, in2965_2;
    wire c2965;
    assign in2965_1 = {pp53[62]};
    assign in2965_2 = {pp54[61]};
    Full_Adder FA_2965(s2965, c2965, in2965_1, in2965_2, pp52[63]);
    wire[0:0] s2966, in2966_1, in2966_2;
    wire c2966;
    assign in2966_1 = {pp56[59]};
    assign in2966_2 = {pp57[58]};
    Full_Adder FA_2966(s2966, c2966, in2966_1, in2966_2, pp55[60]);
    wire[0:0] s2967, in2967_1, in2967_2;
    wire c2967;
    assign in2967_1 = {pp59[56]};
    assign in2967_2 = {pp60[55]};
    Full_Adder FA_2967(s2967, c2967, in2967_1, in2967_2, pp58[57]);
    wire[0:0] s2968, in2968_1, in2968_2;
    wire c2968;
    assign in2968_1 = {pp54[62]};
    assign in2968_2 = {pp55[61]};
    Full_Adder FA_2968(s2968, c2968, in2968_1, in2968_2, pp53[63]);
    wire[0:0] s2969, in2969_1, in2969_2;
    wire c2969;
    assign in2969_1 = {pp57[59]};
    assign in2969_2 = {pp58[58]};
    Full_Adder FA_2969(s2969, c2969, in2969_1, in2969_2, pp56[60]);
    wire[0:0] s2970, in2970_1, in2970_2;
    wire c2970;
    assign in2970_1 = {pp55[62]};
    assign in2970_2 = {pp56[61]};
    Full_Adder FA_2970(s2970, c2970, in2970_1, in2970_2, pp54[63]);

    /*Stage 6*/
    wire[0:0] s2971, in2971_1, in2971_2;
    wire c2971;
    assign in2971_1 = {pp0[7]};
    assign in2971_2 = {pp1[6]};
    Half_Adder HA_2971(s2971, c2971, in2971_1, in2971_2);
    wire[0:0] s2972, in2972_1, in2972_2;
    wire c2972;
    assign in2972_1 = {pp1[7]};
    assign in2972_2 = {pp2[6]};
    Full_Adder FA_2972(s2972, c2972, in2972_1, in2972_2, pp0[8]);
    wire[0:0] s2973, in2973_1, in2973_2;
    wire c2973;
    assign in2973_1 = {pp3[5]};
    assign in2973_2 = {pp4[4]};
    Half_Adder HA_2973(s2973, c2973, in2973_1, in2973_2);
    wire[0:0] s2974, in2974_1, in2974_2;
    wire c2974;
    assign in2974_1 = {pp1[8]};
    assign in2974_2 = {pp2[7]};
    Full_Adder FA_2974(s2974, c2974, in2974_1, in2974_2, pp0[9]);
    wire[0:0] s2975, in2975_1, in2975_2;
    wire c2975;
    assign in2975_1 = {pp4[5]};
    assign in2975_2 = {pp5[4]};
    Full_Adder FA_2975(s2975, c2975, in2975_1, in2975_2, pp3[6]);
    wire[0:0] s2976, in2976_1, in2976_2;
    wire c2976;
    assign in2976_1 = {pp6[3]};
    assign in2976_2 = {pp7[2]};
    Half_Adder HA_2976(s2976, c2976, in2976_1, in2976_2);
    wire[0:0] s2977, in2977_1, in2977_2;
    wire c2977;
    assign in2977_1 = {pp3[7]};
    assign in2977_2 = {pp4[6]};
    Full_Adder FA_2977(s2977, c2977, in2977_1, in2977_2, pp2[8]);
    wire[0:0] s2978, in2978_1, in2978_2;
    wire c2978;
    assign in2978_1 = {pp6[4]};
    assign in2978_2 = {pp7[3]};
    Full_Adder FA_2978(s2978, c2978, in2978_1, in2978_2, pp5[5]);
    wire[0:0] s2979, in2979_1, in2979_2;
    wire c2979;
    assign in2979_1 = {pp9[1]};
    assign in2979_2 = {pp10[0]};
    Full_Adder FA_2979(s2979, c2979, in2979_1, in2979_2, pp8[2]);
    wire[0:0] s2980, in2980_1, in2980_2;
    wire c2980;
    assign in2980_1 = {pp6[5]};
    assign in2980_2 = {pp7[4]};
    Full_Adder FA_2980(s2980, c2980, in2980_1, in2980_2, pp5[6]);
    wire[0:0] s2981, in2981_1, in2981_2;
    wire c2981;
    assign in2981_1 = {pp9[2]};
    assign in2981_2 = {pp10[1]};
    Full_Adder FA_2981(s2981, c2981, in2981_1, in2981_2, pp8[3]);
    wire[0:0] s2982, in2982_1, in2982_2;
    wire c2982;
    assign in2982_1 = {c2551};
    assign in2982_2 = {s2552[0]};
    Full_Adder FA_2982(s2982, c2982, in2982_1, in2982_2, pp11[0]);
    wire[0:0] s2983, in2983_1, in2983_2;
    wire c2983;
    assign in2983_1 = {pp9[3]};
    assign in2983_2 = {pp10[2]};
    Full_Adder FA_2983(s2983, c2983, in2983_1, in2983_2, pp8[4]);
    wire[0:0] s2984, in2984_1, in2984_2;
    wire c2984;
    assign in2984_1 = {pp12[0]};
    assign in2984_2 = {c2552};
    Full_Adder FA_2984(s2984, c2984, in2984_1, in2984_2, pp11[1]);
    wire[0:0] s2985, in2985_1, in2985_2;
    wire c2985;
    assign in2985_1 = {s2554[0]};
    assign in2985_2 = {s2555[0]};
    Full_Adder FA_2985(s2985, c2985, in2985_1, in2985_2, c2553);
    wire[0:0] s2986, in2986_1, in2986_2;
    wire c2986;
    assign in2986_1 = {pp12[1]};
    assign in2986_2 = {pp13[0]};
    Full_Adder FA_2986(s2986, c2986, in2986_1, in2986_2, pp11[2]);
    wire[0:0] s2987, in2987_1, in2987_2;
    wire c2987;
    assign in2987_1 = {c2555};
    assign in2987_2 = {c2556};
    Full_Adder FA_2987(s2987, c2987, in2987_1, in2987_2, c2554);
    wire[0:0] s2988, in2988_1, in2988_2;
    wire c2988;
    assign in2988_1 = {s2558[0]};
    assign in2988_2 = {s2559[0]};
    Full_Adder FA_2988(s2988, c2988, in2988_1, in2988_2, s2557[0]);
    wire[0:0] s2989, in2989_1, in2989_2;
    wire c2989;
    assign in2989_1 = {s1981[0]};
    assign in2989_2 = {c2557};
    Full_Adder FA_2989(s2989, c2989, in2989_1, in2989_2, pp14[0]);
    wire[0:0] s2990, in2990_1, in2990_2;
    wire c2990;
    assign in2990_1 = {c2559};
    assign in2990_2 = {c2560};
    Full_Adder FA_2990(s2990, c2990, in2990_1, in2990_2, c2558);
    wire[0:0] s2991, in2991_1, in2991_2;
    wire c2991;
    assign in2991_1 = {s2562[0]};
    assign in2991_2 = {s2563[0]};
    Full_Adder FA_2991(s2991, c2991, in2991_1, in2991_2, s2561[0]);
    wire[0:0] s2992, in2992_1, in2992_2;
    wire c2992;
    assign in2992_1 = {s1983[0]};
    assign in2992_2 = {c2561};
    Full_Adder FA_2992(s2992, c2992, in2992_1, in2992_2, s1982[0]);
    wire[0:0] s2993, in2993_1, in2993_2;
    wire c2993;
    assign in2993_1 = {c2563};
    assign in2993_2 = {c2564};
    Full_Adder FA_2993(s2993, c2993, in2993_1, in2993_2, c2562);
    wire[0:0] s2994, in2994_1, in2994_2;
    wire c2994;
    assign in2994_1 = {s2566[0]};
    assign in2994_2 = {s2567[0]};
    Full_Adder FA_2994(s2994, c2994, in2994_1, in2994_2, s2565[0]);
    wire[0:0] s2995, in2995_1, in2995_2;
    wire c2995;
    assign in2995_1 = {s1986[0]};
    assign in2995_2 = {c2565};
    Full_Adder FA_2995(s2995, c2995, in2995_1, in2995_2, s1985[0]);
    wire[0:0] s2996, in2996_1, in2996_2;
    wire c2996;
    assign in2996_1 = {c2567};
    assign in2996_2 = {c2568};
    Full_Adder FA_2996(s2996, c2996, in2996_1, in2996_2, c2566);
    wire[0:0] s2997, in2997_1, in2997_2;
    wire c2997;
    assign in2997_1 = {s2570[0]};
    assign in2997_2 = {s2571[0]};
    Full_Adder FA_2997(s2997, c2997, in2997_1, in2997_2, s2569[0]);
    wire[0:0] s2998, in2998_1, in2998_2;
    wire c2998;
    assign in2998_1 = {s1990[0]};
    assign in2998_2 = {c2569};
    Full_Adder FA_2998(s2998, c2998, in2998_1, in2998_2, s1989[0]);
    wire[0:0] s2999, in2999_1, in2999_2;
    wire c2999;
    assign in2999_1 = {c2571};
    assign in2999_2 = {c2572};
    Full_Adder FA_2999(s2999, c2999, in2999_1, in2999_2, c2570);
    wire[0:0] s3000, in3000_1, in3000_2;
    wire c3000;
    assign in3000_1 = {s2574[0]};
    assign in3000_2 = {s2575[0]};
    Full_Adder FA_3000(s3000, c3000, in3000_1, in3000_2, s2573[0]);
    wire[0:0] s3001, in3001_1, in3001_2;
    wire c3001;
    assign in3001_1 = {s1995[0]};
    assign in3001_2 = {c2573};
    Full_Adder FA_3001(s3001, c3001, in3001_1, in3001_2, s1994[0]);
    wire[0:0] s3002, in3002_1, in3002_2;
    wire c3002;
    assign in3002_1 = {c2575};
    assign in3002_2 = {c2576};
    Full_Adder FA_3002(s3002, c3002, in3002_1, in3002_2, c2574);
    wire[0:0] s3003, in3003_1, in3003_2;
    wire c3003;
    assign in3003_1 = {s2578[0]};
    assign in3003_2 = {s2579[0]};
    Full_Adder FA_3003(s3003, c3003, in3003_1, in3003_2, s2577[0]);
    wire[0:0] s3004, in3004_1, in3004_2;
    wire c3004;
    assign in3004_1 = {s2001[0]};
    assign in3004_2 = {c2577};
    Full_Adder FA_3004(s3004, c3004, in3004_1, in3004_2, s2000[0]);
    wire[0:0] s3005, in3005_1, in3005_2;
    wire c3005;
    assign in3005_1 = {c2579};
    assign in3005_2 = {c2580};
    Full_Adder FA_3005(s3005, c3005, in3005_1, in3005_2, c2578);
    wire[0:0] s3006, in3006_1, in3006_2;
    wire c3006;
    assign in3006_1 = {s2582[0]};
    assign in3006_2 = {s2583[0]};
    Full_Adder FA_3006(s3006, c3006, in3006_1, in3006_2, s2581[0]);
    wire[0:0] s3007, in3007_1, in3007_2;
    wire c3007;
    assign in3007_1 = {s2007[0]};
    assign in3007_2 = {c2581};
    Full_Adder FA_3007(s3007, c3007, in3007_1, in3007_2, s2006[0]);
    wire[0:0] s3008, in3008_1, in3008_2;
    wire c3008;
    assign in3008_1 = {c2583};
    assign in3008_2 = {c2584};
    Full_Adder FA_3008(s3008, c3008, in3008_1, in3008_2, c2582);
    wire[0:0] s3009, in3009_1, in3009_2;
    wire c3009;
    assign in3009_1 = {s2586[0]};
    assign in3009_2 = {s2587[0]};
    Full_Adder FA_3009(s3009, c3009, in3009_1, in3009_2, s2585[0]);
    wire[0:0] s3010, in3010_1, in3010_2;
    wire c3010;
    assign in3010_1 = {s2013[0]};
    assign in3010_2 = {c2585};
    Full_Adder FA_3010(s3010, c3010, in3010_1, in3010_2, s2012[0]);
    wire[0:0] s3011, in3011_1, in3011_2;
    wire c3011;
    assign in3011_1 = {c2587};
    assign in3011_2 = {c2588};
    Full_Adder FA_3011(s3011, c3011, in3011_1, in3011_2, c2586);
    wire[0:0] s3012, in3012_1, in3012_2;
    wire c3012;
    assign in3012_1 = {s2590[0]};
    assign in3012_2 = {s2591[0]};
    Full_Adder FA_3012(s3012, c3012, in3012_1, in3012_2, s2589[0]);
    wire[0:0] s3013, in3013_1, in3013_2;
    wire c3013;
    assign in3013_1 = {s2019[0]};
    assign in3013_2 = {c2589};
    Full_Adder FA_3013(s3013, c3013, in3013_1, in3013_2, s2018[0]);
    wire[0:0] s3014, in3014_1, in3014_2;
    wire c3014;
    assign in3014_1 = {c2591};
    assign in3014_2 = {c2592};
    Full_Adder FA_3014(s3014, c3014, in3014_1, in3014_2, c2590);
    wire[0:0] s3015, in3015_1, in3015_2;
    wire c3015;
    assign in3015_1 = {s2594[0]};
    assign in3015_2 = {s2595[0]};
    Full_Adder FA_3015(s3015, c3015, in3015_1, in3015_2, s2593[0]);
    wire[0:0] s3016, in3016_1, in3016_2;
    wire c3016;
    assign in3016_1 = {s2025[0]};
    assign in3016_2 = {c2593};
    Full_Adder FA_3016(s3016, c3016, in3016_1, in3016_2, s2024[0]);
    wire[0:0] s3017, in3017_1, in3017_2;
    wire c3017;
    assign in3017_1 = {c2595};
    assign in3017_2 = {c2596};
    Full_Adder FA_3017(s3017, c3017, in3017_1, in3017_2, c2594);
    wire[0:0] s3018, in3018_1, in3018_2;
    wire c3018;
    assign in3018_1 = {s2598[0]};
    assign in3018_2 = {s2599[0]};
    Full_Adder FA_3018(s3018, c3018, in3018_1, in3018_2, s2597[0]);
    wire[0:0] s3019, in3019_1, in3019_2;
    wire c3019;
    assign in3019_1 = {s2031[0]};
    assign in3019_2 = {c2597};
    Full_Adder FA_3019(s3019, c3019, in3019_1, in3019_2, s2030[0]);
    wire[0:0] s3020, in3020_1, in3020_2;
    wire c3020;
    assign in3020_1 = {c2599};
    assign in3020_2 = {c2600};
    Full_Adder FA_3020(s3020, c3020, in3020_1, in3020_2, c2598);
    wire[0:0] s3021, in3021_1, in3021_2;
    wire c3021;
    assign in3021_1 = {s2602[0]};
    assign in3021_2 = {s2603[0]};
    Full_Adder FA_3021(s3021, c3021, in3021_1, in3021_2, s2601[0]);
    wire[0:0] s3022, in3022_1, in3022_2;
    wire c3022;
    assign in3022_1 = {s2037[0]};
    assign in3022_2 = {c2601};
    Full_Adder FA_3022(s3022, c3022, in3022_1, in3022_2, s2036[0]);
    wire[0:0] s3023, in3023_1, in3023_2;
    wire c3023;
    assign in3023_1 = {c2603};
    assign in3023_2 = {c2604};
    Full_Adder FA_3023(s3023, c3023, in3023_1, in3023_2, c2602);
    wire[0:0] s3024, in3024_1, in3024_2;
    wire c3024;
    assign in3024_1 = {s2606[0]};
    assign in3024_2 = {s2607[0]};
    Full_Adder FA_3024(s3024, c3024, in3024_1, in3024_2, s2605[0]);
    wire[0:0] s3025, in3025_1, in3025_2;
    wire c3025;
    assign in3025_1 = {s2043[0]};
    assign in3025_2 = {c2605};
    Full_Adder FA_3025(s3025, c3025, in3025_1, in3025_2, s2042[0]);
    wire[0:0] s3026, in3026_1, in3026_2;
    wire c3026;
    assign in3026_1 = {c2607};
    assign in3026_2 = {c2608};
    Full_Adder FA_3026(s3026, c3026, in3026_1, in3026_2, c2606);
    wire[0:0] s3027, in3027_1, in3027_2;
    wire c3027;
    assign in3027_1 = {s2610[0]};
    assign in3027_2 = {s2611[0]};
    Full_Adder FA_3027(s3027, c3027, in3027_1, in3027_2, s2609[0]);
    wire[0:0] s3028, in3028_1, in3028_2;
    wire c3028;
    assign in3028_1 = {s2049[0]};
    assign in3028_2 = {c2609};
    Full_Adder FA_3028(s3028, c3028, in3028_1, in3028_2, s2048[0]);
    wire[0:0] s3029, in3029_1, in3029_2;
    wire c3029;
    assign in3029_1 = {c2611};
    assign in3029_2 = {c2612};
    Full_Adder FA_3029(s3029, c3029, in3029_1, in3029_2, c2610);
    wire[0:0] s3030, in3030_1, in3030_2;
    wire c3030;
    assign in3030_1 = {s2614[0]};
    assign in3030_2 = {s2615[0]};
    Full_Adder FA_3030(s3030, c3030, in3030_1, in3030_2, s2613[0]);
    wire[0:0] s3031, in3031_1, in3031_2;
    wire c3031;
    assign in3031_1 = {s2055[0]};
    assign in3031_2 = {c2613};
    Full_Adder FA_3031(s3031, c3031, in3031_1, in3031_2, s2054[0]);
    wire[0:0] s3032, in3032_1, in3032_2;
    wire c3032;
    assign in3032_1 = {c2615};
    assign in3032_2 = {c2616};
    Full_Adder FA_3032(s3032, c3032, in3032_1, in3032_2, c2614);
    wire[0:0] s3033, in3033_1, in3033_2;
    wire c3033;
    assign in3033_1 = {s2618[0]};
    assign in3033_2 = {s2619[0]};
    Full_Adder FA_3033(s3033, c3033, in3033_1, in3033_2, s2617[0]);
    wire[0:0] s3034, in3034_1, in3034_2;
    wire c3034;
    assign in3034_1 = {s2061[0]};
    assign in3034_2 = {c2617};
    Full_Adder FA_3034(s3034, c3034, in3034_1, in3034_2, s2060[0]);
    wire[0:0] s3035, in3035_1, in3035_2;
    wire c3035;
    assign in3035_1 = {c2619};
    assign in3035_2 = {c2620};
    Full_Adder FA_3035(s3035, c3035, in3035_1, in3035_2, c2618);
    wire[0:0] s3036, in3036_1, in3036_2;
    wire c3036;
    assign in3036_1 = {s2622[0]};
    assign in3036_2 = {s2623[0]};
    Full_Adder FA_3036(s3036, c3036, in3036_1, in3036_2, s2621[0]);
    wire[0:0] s3037, in3037_1, in3037_2;
    wire c3037;
    assign in3037_1 = {s2067[0]};
    assign in3037_2 = {c2621};
    Full_Adder FA_3037(s3037, c3037, in3037_1, in3037_2, s2066[0]);
    wire[0:0] s3038, in3038_1, in3038_2;
    wire c3038;
    assign in3038_1 = {c2623};
    assign in3038_2 = {c2624};
    Full_Adder FA_3038(s3038, c3038, in3038_1, in3038_2, c2622);
    wire[0:0] s3039, in3039_1, in3039_2;
    wire c3039;
    assign in3039_1 = {s2626[0]};
    assign in3039_2 = {s2627[0]};
    Full_Adder FA_3039(s3039, c3039, in3039_1, in3039_2, s2625[0]);
    wire[0:0] s3040, in3040_1, in3040_2;
    wire c3040;
    assign in3040_1 = {s2073[0]};
    assign in3040_2 = {c2625};
    Full_Adder FA_3040(s3040, c3040, in3040_1, in3040_2, s2072[0]);
    wire[0:0] s3041, in3041_1, in3041_2;
    wire c3041;
    assign in3041_1 = {c2627};
    assign in3041_2 = {c2628};
    Full_Adder FA_3041(s3041, c3041, in3041_1, in3041_2, c2626);
    wire[0:0] s3042, in3042_1, in3042_2;
    wire c3042;
    assign in3042_1 = {s2630[0]};
    assign in3042_2 = {s2631[0]};
    Full_Adder FA_3042(s3042, c3042, in3042_1, in3042_2, s2629[0]);
    wire[0:0] s3043, in3043_1, in3043_2;
    wire c3043;
    assign in3043_1 = {s2079[0]};
    assign in3043_2 = {c2629};
    Full_Adder FA_3043(s3043, c3043, in3043_1, in3043_2, s2078[0]);
    wire[0:0] s3044, in3044_1, in3044_2;
    wire c3044;
    assign in3044_1 = {c2631};
    assign in3044_2 = {c2632};
    Full_Adder FA_3044(s3044, c3044, in3044_1, in3044_2, c2630);
    wire[0:0] s3045, in3045_1, in3045_2;
    wire c3045;
    assign in3045_1 = {s2634[0]};
    assign in3045_2 = {s2635[0]};
    Full_Adder FA_3045(s3045, c3045, in3045_1, in3045_2, s2633[0]);
    wire[0:0] s3046, in3046_1, in3046_2;
    wire c3046;
    assign in3046_1 = {s2085[0]};
    assign in3046_2 = {c2633};
    Full_Adder FA_3046(s3046, c3046, in3046_1, in3046_2, s2084[0]);
    wire[0:0] s3047, in3047_1, in3047_2;
    wire c3047;
    assign in3047_1 = {c2635};
    assign in3047_2 = {c2636};
    Full_Adder FA_3047(s3047, c3047, in3047_1, in3047_2, c2634);
    wire[0:0] s3048, in3048_1, in3048_2;
    wire c3048;
    assign in3048_1 = {s2638[0]};
    assign in3048_2 = {s2639[0]};
    Full_Adder FA_3048(s3048, c3048, in3048_1, in3048_2, s2637[0]);
    wire[0:0] s3049, in3049_1, in3049_2;
    wire c3049;
    assign in3049_1 = {s2091[0]};
    assign in3049_2 = {c2637};
    Full_Adder FA_3049(s3049, c3049, in3049_1, in3049_2, s2090[0]);
    wire[0:0] s3050, in3050_1, in3050_2;
    wire c3050;
    assign in3050_1 = {c2639};
    assign in3050_2 = {c2640};
    Full_Adder FA_3050(s3050, c3050, in3050_1, in3050_2, c2638);
    wire[0:0] s3051, in3051_1, in3051_2;
    wire c3051;
    assign in3051_1 = {s2642[0]};
    assign in3051_2 = {s2643[0]};
    Full_Adder FA_3051(s3051, c3051, in3051_1, in3051_2, s2641[0]);
    wire[0:0] s3052, in3052_1, in3052_2;
    wire c3052;
    assign in3052_1 = {s2097[0]};
    assign in3052_2 = {c2641};
    Full_Adder FA_3052(s3052, c3052, in3052_1, in3052_2, s2096[0]);
    wire[0:0] s3053, in3053_1, in3053_2;
    wire c3053;
    assign in3053_1 = {c2643};
    assign in3053_2 = {c2644};
    Full_Adder FA_3053(s3053, c3053, in3053_1, in3053_2, c2642);
    wire[0:0] s3054, in3054_1, in3054_2;
    wire c3054;
    assign in3054_1 = {s2646[0]};
    assign in3054_2 = {s2647[0]};
    Full_Adder FA_3054(s3054, c3054, in3054_1, in3054_2, s2645[0]);
    wire[0:0] s3055, in3055_1, in3055_2;
    wire c3055;
    assign in3055_1 = {s2103[0]};
    assign in3055_2 = {c2645};
    Full_Adder FA_3055(s3055, c3055, in3055_1, in3055_2, s2102[0]);
    wire[0:0] s3056, in3056_1, in3056_2;
    wire c3056;
    assign in3056_1 = {c2647};
    assign in3056_2 = {c2648};
    Full_Adder FA_3056(s3056, c3056, in3056_1, in3056_2, c2646);
    wire[0:0] s3057, in3057_1, in3057_2;
    wire c3057;
    assign in3057_1 = {s2650[0]};
    assign in3057_2 = {s2651[0]};
    Full_Adder FA_3057(s3057, c3057, in3057_1, in3057_2, s2649[0]);
    wire[0:0] s3058, in3058_1, in3058_2;
    wire c3058;
    assign in3058_1 = {s2109[0]};
    assign in3058_2 = {c2649};
    Full_Adder FA_3058(s3058, c3058, in3058_1, in3058_2, s2108[0]);
    wire[0:0] s3059, in3059_1, in3059_2;
    wire c3059;
    assign in3059_1 = {c2651};
    assign in3059_2 = {c2652};
    Full_Adder FA_3059(s3059, c3059, in3059_1, in3059_2, c2650);
    wire[0:0] s3060, in3060_1, in3060_2;
    wire c3060;
    assign in3060_1 = {s2654[0]};
    assign in3060_2 = {s2655[0]};
    Full_Adder FA_3060(s3060, c3060, in3060_1, in3060_2, s2653[0]);
    wire[0:0] s3061, in3061_1, in3061_2;
    wire c3061;
    assign in3061_1 = {s2115[0]};
    assign in3061_2 = {c2653};
    Full_Adder FA_3061(s3061, c3061, in3061_1, in3061_2, s2114[0]);
    wire[0:0] s3062, in3062_1, in3062_2;
    wire c3062;
    assign in3062_1 = {c2655};
    assign in3062_2 = {c2656};
    Full_Adder FA_3062(s3062, c3062, in3062_1, in3062_2, c2654);
    wire[0:0] s3063, in3063_1, in3063_2;
    wire c3063;
    assign in3063_1 = {s2658[0]};
    assign in3063_2 = {s2659[0]};
    Full_Adder FA_3063(s3063, c3063, in3063_1, in3063_2, s2657[0]);
    wire[0:0] s3064, in3064_1, in3064_2;
    wire c3064;
    assign in3064_1 = {s2121[0]};
    assign in3064_2 = {c2657};
    Full_Adder FA_3064(s3064, c3064, in3064_1, in3064_2, s2120[0]);
    wire[0:0] s3065, in3065_1, in3065_2;
    wire c3065;
    assign in3065_1 = {c2659};
    assign in3065_2 = {c2660};
    Full_Adder FA_3065(s3065, c3065, in3065_1, in3065_2, c2658);
    wire[0:0] s3066, in3066_1, in3066_2;
    wire c3066;
    assign in3066_1 = {s2662[0]};
    assign in3066_2 = {s2663[0]};
    Full_Adder FA_3066(s3066, c3066, in3066_1, in3066_2, s2661[0]);
    wire[0:0] s3067, in3067_1, in3067_2;
    wire c3067;
    assign in3067_1 = {s2127[0]};
    assign in3067_2 = {c2661};
    Full_Adder FA_3067(s3067, c3067, in3067_1, in3067_2, s2126[0]);
    wire[0:0] s3068, in3068_1, in3068_2;
    wire c3068;
    assign in3068_1 = {c2663};
    assign in3068_2 = {c2664};
    Full_Adder FA_3068(s3068, c3068, in3068_1, in3068_2, c2662);
    wire[0:0] s3069, in3069_1, in3069_2;
    wire c3069;
    assign in3069_1 = {s2666[0]};
    assign in3069_2 = {s2667[0]};
    Full_Adder FA_3069(s3069, c3069, in3069_1, in3069_2, s2665[0]);
    wire[0:0] s3070, in3070_1, in3070_2;
    wire c3070;
    assign in3070_1 = {s2133[0]};
    assign in3070_2 = {c2665};
    Full_Adder FA_3070(s3070, c3070, in3070_1, in3070_2, s2132[0]);
    wire[0:0] s3071, in3071_1, in3071_2;
    wire c3071;
    assign in3071_1 = {c2667};
    assign in3071_2 = {c2668};
    Full_Adder FA_3071(s3071, c3071, in3071_1, in3071_2, c2666);
    wire[0:0] s3072, in3072_1, in3072_2;
    wire c3072;
    assign in3072_1 = {s2670[0]};
    assign in3072_2 = {s2671[0]};
    Full_Adder FA_3072(s3072, c3072, in3072_1, in3072_2, s2669[0]);
    wire[0:0] s3073, in3073_1, in3073_2;
    wire c3073;
    assign in3073_1 = {s2139[0]};
    assign in3073_2 = {c2669};
    Full_Adder FA_3073(s3073, c3073, in3073_1, in3073_2, s2138[0]);
    wire[0:0] s3074, in3074_1, in3074_2;
    wire c3074;
    assign in3074_1 = {c2671};
    assign in3074_2 = {c2672};
    Full_Adder FA_3074(s3074, c3074, in3074_1, in3074_2, c2670);
    wire[0:0] s3075, in3075_1, in3075_2;
    wire c3075;
    assign in3075_1 = {s2674[0]};
    assign in3075_2 = {s2675[0]};
    Full_Adder FA_3075(s3075, c3075, in3075_1, in3075_2, s2673[0]);
    wire[0:0] s3076, in3076_1, in3076_2;
    wire c3076;
    assign in3076_1 = {s2145[0]};
    assign in3076_2 = {c2673};
    Full_Adder FA_3076(s3076, c3076, in3076_1, in3076_2, s2144[0]);
    wire[0:0] s3077, in3077_1, in3077_2;
    wire c3077;
    assign in3077_1 = {c2675};
    assign in3077_2 = {c2676};
    Full_Adder FA_3077(s3077, c3077, in3077_1, in3077_2, c2674);
    wire[0:0] s3078, in3078_1, in3078_2;
    wire c3078;
    assign in3078_1 = {s2678[0]};
    assign in3078_2 = {s2679[0]};
    Full_Adder FA_3078(s3078, c3078, in3078_1, in3078_2, s2677[0]);
    wire[0:0] s3079, in3079_1, in3079_2;
    wire c3079;
    assign in3079_1 = {s2151[0]};
    assign in3079_2 = {c2677};
    Full_Adder FA_3079(s3079, c3079, in3079_1, in3079_2, s2150[0]);
    wire[0:0] s3080, in3080_1, in3080_2;
    wire c3080;
    assign in3080_1 = {c2679};
    assign in3080_2 = {c2680};
    Full_Adder FA_3080(s3080, c3080, in3080_1, in3080_2, c2678);
    wire[0:0] s3081, in3081_1, in3081_2;
    wire c3081;
    assign in3081_1 = {s2682[0]};
    assign in3081_2 = {s2683[0]};
    Full_Adder FA_3081(s3081, c3081, in3081_1, in3081_2, s2681[0]);
    wire[0:0] s3082, in3082_1, in3082_2;
    wire c3082;
    assign in3082_1 = {s2157[0]};
    assign in3082_2 = {c2681};
    Full_Adder FA_3082(s3082, c3082, in3082_1, in3082_2, s2156[0]);
    wire[0:0] s3083, in3083_1, in3083_2;
    wire c3083;
    assign in3083_1 = {c2683};
    assign in3083_2 = {c2684};
    Full_Adder FA_3083(s3083, c3083, in3083_1, in3083_2, c2682);
    wire[0:0] s3084, in3084_1, in3084_2;
    wire c3084;
    assign in3084_1 = {s2686[0]};
    assign in3084_2 = {s2687[0]};
    Full_Adder FA_3084(s3084, c3084, in3084_1, in3084_2, s2685[0]);
    wire[0:0] s3085, in3085_1, in3085_2;
    wire c3085;
    assign in3085_1 = {s2163[0]};
    assign in3085_2 = {c2685};
    Full_Adder FA_3085(s3085, c3085, in3085_1, in3085_2, s2162[0]);
    wire[0:0] s3086, in3086_1, in3086_2;
    wire c3086;
    assign in3086_1 = {c2687};
    assign in3086_2 = {c2688};
    Full_Adder FA_3086(s3086, c3086, in3086_1, in3086_2, c2686);
    wire[0:0] s3087, in3087_1, in3087_2;
    wire c3087;
    assign in3087_1 = {s2690[0]};
    assign in3087_2 = {s2691[0]};
    Full_Adder FA_3087(s3087, c3087, in3087_1, in3087_2, s2689[0]);
    wire[0:0] s3088, in3088_1, in3088_2;
    wire c3088;
    assign in3088_1 = {s2169[0]};
    assign in3088_2 = {c2689};
    Full_Adder FA_3088(s3088, c3088, in3088_1, in3088_2, s2168[0]);
    wire[0:0] s3089, in3089_1, in3089_2;
    wire c3089;
    assign in3089_1 = {c2691};
    assign in3089_2 = {c2692};
    Full_Adder FA_3089(s3089, c3089, in3089_1, in3089_2, c2690);
    wire[0:0] s3090, in3090_1, in3090_2;
    wire c3090;
    assign in3090_1 = {s2694[0]};
    assign in3090_2 = {s2695[0]};
    Full_Adder FA_3090(s3090, c3090, in3090_1, in3090_2, s2693[0]);
    wire[0:0] s3091, in3091_1, in3091_2;
    wire c3091;
    assign in3091_1 = {s2175[0]};
    assign in3091_2 = {c2693};
    Full_Adder FA_3091(s3091, c3091, in3091_1, in3091_2, s2174[0]);
    wire[0:0] s3092, in3092_1, in3092_2;
    wire c3092;
    assign in3092_1 = {c2695};
    assign in3092_2 = {c2696};
    Full_Adder FA_3092(s3092, c3092, in3092_1, in3092_2, c2694);
    wire[0:0] s3093, in3093_1, in3093_2;
    wire c3093;
    assign in3093_1 = {s2698[0]};
    assign in3093_2 = {s2699[0]};
    Full_Adder FA_3093(s3093, c3093, in3093_1, in3093_2, s2697[0]);
    wire[0:0] s3094, in3094_1, in3094_2;
    wire c3094;
    assign in3094_1 = {s2181[0]};
    assign in3094_2 = {c2697};
    Full_Adder FA_3094(s3094, c3094, in3094_1, in3094_2, s2180[0]);
    wire[0:0] s3095, in3095_1, in3095_2;
    wire c3095;
    assign in3095_1 = {c2699};
    assign in3095_2 = {c2700};
    Full_Adder FA_3095(s3095, c3095, in3095_1, in3095_2, c2698);
    wire[0:0] s3096, in3096_1, in3096_2;
    wire c3096;
    assign in3096_1 = {s2702[0]};
    assign in3096_2 = {s2703[0]};
    Full_Adder FA_3096(s3096, c3096, in3096_1, in3096_2, s2701[0]);
    wire[0:0] s3097, in3097_1, in3097_2;
    wire c3097;
    assign in3097_1 = {s2187[0]};
    assign in3097_2 = {c2701};
    Full_Adder FA_3097(s3097, c3097, in3097_1, in3097_2, s2186[0]);
    wire[0:0] s3098, in3098_1, in3098_2;
    wire c3098;
    assign in3098_1 = {c2703};
    assign in3098_2 = {c2704};
    Full_Adder FA_3098(s3098, c3098, in3098_1, in3098_2, c2702);
    wire[0:0] s3099, in3099_1, in3099_2;
    wire c3099;
    assign in3099_1 = {s2706[0]};
    assign in3099_2 = {s2707[0]};
    Full_Adder FA_3099(s3099, c3099, in3099_1, in3099_2, s2705[0]);
    wire[0:0] s3100, in3100_1, in3100_2;
    wire c3100;
    assign in3100_1 = {s2193[0]};
    assign in3100_2 = {c2705};
    Full_Adder FA_3100(s3100, c3100, in3100_1, in3100_2, s2192[0]);
    wire[0:0] s3101, in3101_1, in3101_2;
    wire c3101;
    assign in3101_1 = {c2707};
    assign in3101_2 = {c2708};
    Full_Adder FA_3101(s3101, c3101, in3101_1, in3101_2, c2706);
    wire[0:0] s3102, in3102_1, in3102_2;
    wire c3102;
    assign in3102_1 = {s2710[0]};
    assign in3102_2 = {s2711[0]};
    Full_Adder FA_3102(s3102, c3102, in3102_1, in3102_2, s2709[0]);
    wire[0:0] s3103, in3103_1, in3103_2;
    wire c3103;
    assign in3103_1 = {s2199[0]};
    assign in3103_2 = {c2709};
    Full_Adder FA_3103(s3103, c3103, in3103_1, in3103_2, s2198[0]);
    wire[0:0] s3104, in3104_1, in3104_2;
    wire c3104;
    assign in3104_1 = {c2711};
    assign in3104_2 = {c2712};
    Full_Adder FA_3104(s3104, c3104, in3104_1, in3104_2, c2710);
    wire[0:0] s3105, in3105_1, in3105_2;
    wire c3105;
    assign in3105_1 = {s2714[0]};
    assign in3105_2 = {s2715[0]};
    Full_Adder FA_3105(s3105, c3105, in3105_1, in3105_2, s2713[0]);
    wire[0:0] s3106, in3106_1, in3106_2;
    wire c3106;
    assign in3106_1 = {s2205[0]};
    assign in3106_2 = {c2713};
    Full_Adder FA_3106(s3106, c3106, in3106_1, in3106_2, s2204[0]);
    wire[0:0] s3107, in3107_1, in3107_2;
    wire c3107;
    assign in3107_1 = {c2715};
    assign in3107_2 = {c2716};
    Full_Adder FA_3107(s3107, c3107, in3107_1, in3107_2, c2714);
    wire[0:0] s3108, in3108_1, in3108_2;
    wire c3108;
    assign in3108_1 = {s2718[0]};
    assign in3108_2 = {s2719[0]};
    Full_Adder FA_3108(s3108, c3108, in3108_1, in3108_2, s2717[0]);
    wire[0:0] s3109, in3109_1, in3109_2;
    wire c3109;
    assign in3109_1 = {s2211[0]};
    assign in3109_2 = {c2717};
    Full_Adder FA_3109(s3109, c3109, in3109_1, in3109_2, s2210[0]);
    wire[0:0] s3110, in3110_1, in3110_2;
    wire c3110;
    assign in3110_1 = {c2719};
    assign in3110_2 = {c2720};
    Full_Adder FA_3110(s3110, c3110, in3110_1, in3110_2, c2718);
    wire[0:0] s3111, in3111_1, in3111_2;
    wire c3111;
    assign in3111_1 = {s2722[0]};
    assign in3111_2 = {s2723[0]};
    Full_Adder FA_3111(s3111, c3111, in3111_1, in3111_2, s2721[0]);
    wire[0:0] s3112, in3112_1, in3112_2;
    wire c3112;
    assign in3112_1 = {s2217[0]};
    assign in3112_2 = {c2721};
    Full_Adder FA_3112(s3112, c3112, in3112_1, in3112_2, s2216[0]);
    wire[0:0] s3113, in3113_1, in3113_2;
    wire c3113;
    assign in3113_1 = {c2723};
    assign in3113_2 = {c2724};
    Full_Adder FA_3113(s3113, c3113, in3113_1, in3113_2, c2722);
    wire[0:0] s3114, in3114_1, in3114_2;
    wire c3114;
    assign in3114_1 = {s2726[0]};
    assign in3114_2 = {s2727[0]};
    Full_Adder FA_3114(s3114, c3114, in3114_1, in3114_2, s2725[0]);
    wire[0:0] s3115, in3115_1, in3115_2;
    wire c3115;
    assign in3115_1 = {s2223[0]};
    assign in3115_2 = {c2725};
    Full_Adder FA_3115(s3115, c3115, in3115_1, in3115_2, s2222[0]);
    wire[0:0] s3116, in3116_1, in3116_2;
    wire c3116;
    assign in3116_1 = {c2727};
    assign in3116_2 = {c2728};
    Full_Adder FA_3116(s3116, c3116, in3116_1, in3116_2, c2726);
    wire[0:0] s3117, in3117_1, in3117_2;
    wire c3117;
    assign in3117_1 = {s2730[0]};
    assign in3117_2 = {s2731[0]};
    Full_Adder FA_3117(s3117, c3117, in3117_1, in3117_2, s2729[0]);
    wire[0:0] s3118, in3118_1, in3118_2;
    wire c3118;
    assign in3118_1 = {s2229[0]};
    assign in3118_2 = {c2729};
    Full_Adder FA_3118(s3118, c3118, in3118_1, in3118_2, s2228[0]);
    wire[0:0] s3119, in3119_1, in3119_2;
    wire c3119;
    assign in3119_1 = {c2731};
    assign in3119_2 = {c2732};
    Full_Adder FA_3119(s3119, c3119, in3119_1, in3119_2, c2730);
    wire[0:0] s3120, in3120_1, in3120_2;
    wire c3120;
    assign in3120_1 = {s2734[0]};
    assign in3120_2 = {s2735[0]};
    Full_Adder FA_3120(s3120, c3120, in3120_1, in3120_2, s2733[0]);
    wire[0:0] s3121, in3121_1, in3121_2;
    wire c3121;
    assign in3121_1 = {s2235[0]};
    assign in3121_2 = {c2733};
    Full_Adder FA_3121(s3121, c3121, in3121_1, in3121_2, s2234[0]);
    wire[0:0] s3122, in3122_1, in3122_2;
    wire c3122;
    assign in3122_1 = {c2735};
    assign in3122_2 = {c2736};
    Full_Adder FA_3122(s3122, c3122, in3122_1, in3122_2, c2734);
    wire[0:0] s3123, in3123_1, in3123_2;
    wire c3123;
    assign in3123_1 = {s2738[0]};
    assign in3123_2 = {s2739[0]};
    Full_Adder FA_3123(s3123, c3123, in3123_1, in3123_2, s2737[0]);
    wire[0:0] s3124, in3124_1, in3124_2;
    wire c3124;
    assign in3124_1 = {s2241[0]};
    assign in3124_2 = {c2737};
    Full_Adder FA_3124(s3124, c3124, in3124_1, in3124_2, s2240[0]);
    wire[0:0] s3125, in3125_1, in3125_2;
    wire c3125;
    assign in3125_1 = {c2739};
    assign in3125_2 = {c2740};
    Full_Adder FA_3125(s3125, c3125, in3125_1, in3125_2, c2738);
    wire[0:0] s3126, in3126_1, in3126_2;
    wire c3126;
    assign in3126_1 = {s2742[0]};
    assign in3126_2 = {s2743[0]};
    Full_Adder FA_3126(s3126, c3126, in3126_1, in3126_2, s2741[0]);
    wire[0:0] s3127, in3127_1, in3127_2;
    wire c3127;
    assign in3127_1 = {s2247[0]};
    assign in3127_2 = {c2741};
    Full_Adder FA_3127(s3127, c3127, in3127_1, in3127_2, s2246[0]);
    wire[0:0] s3128, in3128_1, in3128_2;
    wire c3128;
    assign in3128_1 = {c2743};
    assign in3128_2 = {c2744};
    Full_Adder FA_3128(s3128, c3128, in3128_1, in3128_2, c2742);
    wire[0:0] s3129, in3129_1, in3129_2;
    wire c3129;
    assign in3129_1 = {s2746[0]};
    assign in3129_2 = {s2747[0]};
    Full_Adder FA_3129(s3129, c3129, in3129_1, in3129_2, s2745[0]);
    wire[0:0] s3130, in3130_1, in3130_2;
    wire c3130;
    assign in3130_1 = {s2253[0]};
    assign in3130_2 = {c2745};
    Full_Adder FA_3130(s3130, c3130, in3130_1, in3130_2, s2252[0]);
    wire[0:0] s3131, in3131_1, in3131_2;
    wire c3131;
    assign in3131_1 = {c2747};
    assign in3131_2 = {c2748};
    Full_Adder FA_3131(s3131, c3131, in3131_1, in3131_2, c2746);
    wire[0:0] s3132, in3132_1, in3132_2;
    wire c3132;
    assign in3132_1 = {s2750[0]};
    assign in3132_2 = {s2751[0]};
    Full_Adder FA_3132(s3132, c3132, in3132_1, in3132_2, s2749[0]);
    wire[0:0] s3133, in3133_1, in3133_2;
    wire c3133;
    assign in3133_1 = {s2259[0]};
    assign in3133_2 = {c2749};
    Full_Adder FA_3133(s3133, c3133, in3133_1, in3133_2, s2258[0]);
    wire[0:0] s3134, in3134_1, in3134_2;
    wire c3134;
    assign in3134_1 = {c2751};
    assign in3134_2 = {c2752};
    Full_Adder FA_3134(s3134, c3134, in3134_1, in3134_2, c2750);
    wire[0:0] s3135, in3135_1, in3135_2;
    wire c3135;
    assign in3135_1 = {s2754[0]};
    assign in3135_2 = {s2755[0]};
    Full_Adder FA_3135(s3135, c3135, in3135_1, in3135_2, s2753[0]);
    wire[0:0] s3136, in3136_1, in3136_2;
    wire c3136;
    assign in3136_1 = {s2265[0]};
    assign in3136_2 = {c2753};
    Full_Adder FA_3136(s3136, c3136, in3136_1, in3136_2, s2264[0]);
    wire[0:0] s3137, in3137_1, in3137_2;
    wire c3137;
    assign in3137_1 = {c2755};
    assign in3137_2 = {c2756};
    Full_Adder FA_3137(s3137, c3137, in3137_1, in3137_2, c2754);
    wire[0:0] s3138, in3138_1, in3138_2;
    wire c3138;
    assign in3138_1 = {s2758[0]};
    assign in3138_2 = {s2759[0]};
    Full_Adder FA_3138(s3138, c3138, in3138_1, in3138_2, s2757[0]);
    wire[0:0] s3139, in3139_1, in3139_2;
    wire c3139;
    assign in3139_1 = {s2271[0]};
    assign in3139_2 = {c2757};
    Full_Adder FA_3139(s3139, c3139, in3139_1, in3139_2, s2270[0]);
    wire[0:0] s3140, in3140_1, in3140_2;
    wire c3140;
    assign in3140_1 = {c2759};
    assign in3140_2 = {c2760};
    Full_Adder FA_3140(s3140, c3140, in3140_1, in3140_2, c2758);
    wire[0:0] s3141, in3141_1, in3141_2;
    wire c3141;
    assign in3141_1 = {s2762[0]};
    assign in3141_2 = {s2763[0]};
    Full_Adder FA_3141(s3141, c3141, in3141_1, in3141_2, s2761[0]);
    wire[0:0] s3142, in3142_1, in3142_2;
    wire c3142;
    assign in3142_1 = {s2277[0]};
    assign in3142_2 = {c2761};
    Full_Adder FA_3142(s3142, c3142, in3142_1, in3142_2, s2276[0]);
    wire[0:0] s3143, in3143_1, in3143_2;
    wire c3143;
    assign in3143_1 = {c2763};
    assign in3143_2 = {c2764};
    Full_Adder FA_3143(s3143, c3143, in3143_1, in3143_2, c2762);
    wire[0:0] s3144, in3144_1, in3144_2;
    wire c3144;
    assign in3144_1 = {s2766[0]};
    assign in3144_2 = {s2767[0]};
    Full_Adder FA_3144(s3144, c3144, in3144_1, in3144_2, s2765[0]);
    wire[0:0] s3145, in3145_1, in3145_2;
    wire c3145;
    assign in3145_1 = {s2283[0]};
    assign in3145_2 = {c2765};
    Full_Adder FA_3145(s3145, c3145, in3145_1, in3145_2, s2282[0]);
    wire[0:0] s3146, in3146_1, in3146_2;
    wire c3146;
    assign in3146_1 = {c2767};
    assign in3146_2 = {c2768};
    Full_Adder FA_3146(s3146, c3146, in3146_1, in3146_2, c2766);
    wire[0:0] s3147, in3147_1, in3147_2;
    wire c3147;
    assign in3147_1 = {s2770[0]};
    assign in3147_2 = {s2771[0]};
    Full_Adder FA_3147(s3147, c3147, in3147_1, in3147_2, s2769[0]);
    wire[0:0] s3148, in3148_1, in3148_2;
    wire c3148;
    assign in3148_1 = {s2289[0]};
    assign in3148_2 = {c2769};
    Full_Adder FA_3148(s3148, c3148, in3148_1, in3148_2, s2288[0]);
    wire[0:0] s3149, in3149_1, in3149_2;
    wire c3149;
    assign in3149_1 = {c2771};
    assign in3149_2 = {c2772};
    Full_Adder FA_3149(s3149, c3149, in3149_1, in3149_2, c2770);
    wire[0:0] s3150, in3150_1, in3150_2;
    wire c3150;
    assign in3150_1 = {s2774[0]};
    assign in3150_2 = {s2775[0]};
    Full_Adder FA_3150(s3150, c3150, in3150_1, in3150_2, s2773[0]);
    wire[0:0] s3151, in3151_1, in3151_2;
    wire c3151;
    assign in3151_1 = {s2295[0]};
    assign in3151_2 = {c2773};
    Full_Adder FA_3151(s3151, c3151, in3151_1, in3151_2, s2294[0]);
    wire[0:0] s3152, in3152_1, in3152_2;
    wire c3152;
    assign in3152_1 = {c2775};
    assign in3152_2 = {c2776};
    Full_Adder FA_3152(s3152, c3152, in3152_1, in3152_2, c2774);
    wire[0:0] s3153, in3153_1, in3153_2;
    wire c3153;
    assign in3153_1 = {s2778[0]};
    assign in3153_2 = {s2779[0]};
    Full_Adder FA_3153(s3153, c3153, in3153_1, in3153_2, s2777[0]);
    wire[0:0] s3154, in3154_1, in3154_2;
    wire c3154;
    assign in3154_1 = {s2301[0]};
    assign in3154_2 = {c2777};
    Full_Adder FA_3154(s3154, c3154, in3154_1, in3154_2, s2300[0]);
    wire[0:0] s3155, in3155_1, in3155_2;
    wire c3155;
    assign in3155_1 = {c2779};
    assign in3155_2 = {c2780};
    Full_Adder FA_3155(s3155, c3155, in3155_1, in3155_2, c2778);
    wire[0:0] s3156, in3156_1, in3156_2;
    wire c3156;
    assign in3156_1 = {s2782[0]};
    assign in3156_2 = {s2783[0]};
    Full_Adder FA_3156(s3156, c3156, in3156_1, in3156_2, s2781[0]);
    wire[0:0] s3157, in3157_1, in3157_2;
    wire c3157;
    assign in3157_1 = {s2307[0]};
    assign in3157_2 = {c2781};
    Full_Adder FA_3157(s3157, c3157, in3157_1, in3157_2, s2306[0]);
    wire[0:0] s3158, in3158_1, in3158_2;
    wire c3158;
    assign in3158_1 = {c2783};
    assign in3158_2 = {c2784};
    Full_Adder FA_3158(s3158, c3158, in3158_1, in3158_2, c2782);
    wire[0:0] s3159, in3159_1, in3159_2;
    wire c3159;
    assign in3159_1 = {s2786[0]};
    assign in3159_2 = {s2787[0]};
    Full_Adder FA_3159(s3159, c3159, in3159_1, in3159_2, s2785[0]);
    wire[0:0] s3160, in3160_1, in3160_2;
    wire c3160;
    assign in3160_1 = {s2313[0]};
    assign in3160_2 = {c2785};
    Full_Adder FA_3160(s3160, c3160, in3160_1, in3160_2, s2312[0]);
    wire[0:0] s3161, in3161_1, in3161_2;
    wire c3161;
    assign in3161_1 = {c2787};
    assign in3161_2 = {c2788};
    Full_Adder FA_3161(s3161, c3161, in3161_1, in3161_2, c2786);
    wire[0:0] s3162, in3162_1, in3162_2;
    wire c3162;
    assign in3162_1 = {s2790[0]};
    assign in3162_2 = {s2791[0]};
    Full_Adder FA_3162(s3162, c3162, in3162_1, in3162_2, s2789[0]);
    wire[0:0] s3163, in3163_1, in3163_2;
    wire c3163;
    assign in3163_1 = {s2319[0]};
    assign in3163_2 = {c2789};
    Full_Adder FA_3163(s3163, c3163, in3163_1, in3163_2, s2318[0]);
    wire[0:0] s3164, in3164_1, in3164_2;
    wire c3164;
    assign in3164_1 = {c2791};
    assign in3164_2 = {c2792};
    Full_Adder FA_3164(s3164, c3164, in3164_1, in3164_2, c2790);
    wire[0:0] s3165, in3165_1, in3165_2;
    wire c3165;
    assign in3165_1 = {s2794[0]};
    assign in3165_2 = {s2795[0]};
    Full_Adder FA_3165(s3165, c3165, in3165_1, in3165_2, s2793[0]);
    wire[0:0] s3166, in3166_1, in3166_2;
    wire c3166;
    assign in3166_1 = {s2325[0]};
    assign in3166_2 = {c2793};
    Full_Adder FA_3166(s3166, c3166, in3166_1, in3166_2, s2324[0]);
    wire[0:0] s3167, in3167_1, in3167_2;
    wire c3167;
    assign in3167_1 = {c2795};
    assign in3167_2 = {c2796};
    Full_Adder FA_3167(s3167, c3167, in3167_1, in3167_2, c2794);
    wire[0:0] s3168, in3168_1, in3168_2;
    wire c3168;
    assign in3168_1 = {s2798[0]};
    assign in3168_2 = {s2799[0]};
    Full_Adder FA_3168(s3168, c3168, in3168_1, in3168_2, s2797[0]);
    wire[0:0] s3169, in3169_1, in3169_2;
    wire c3169;
    assign in3169_1 = {s2331[0]};
    assign in3169_2 = {c2797};
    Full_Adder FA_3169(s3169, c3169, in3169_1, in3169_2, s2330[0]);
    wire[0:0] s3170, in3170_1, in3170_2;
    wire c3170;
    assign in3170_1 = {c2799};
    assign in3170_2 = {c2800};
    Full_Adder FA_3170(s3170, c3170, in3170_1, in3170_2, c2798);
    wire[0:0] s3171, in3171_1, in3171_2;
    wire c3171;
    assign in3171_1 = {s2802[0]};
    assign in3171_2 = {s2803[0]};
    Full_Adder FA_3171(s3171, c3171, in3171_1, in3171_2, s2801[0]);
    wire[0:0] s3172, in3172_1, in3172_2;
    wire c3172;
    assign in3172_1 = {s2337[0]};
    assign in3172_2 = {c2801};
    Full_Adder FA_3172(s3172, c3172, in3172_1, in3172_2, s2336[0]);
    wire[0:0] s3173, in3173_1, in3173_2;
    wire c3173;
    assign in3173_1 = {c2803};
    assign in3173_2 = {c2804};
    Full_Adder FA_3173(s3173, c3173, in3173_1, in3173_2, c2802);
    wire[0:0] s3174, in3174_1, in3174_2;
    wire c3174;
    assign in3174_1 = {s2806[0]};
    assign in3174_2 = {s2807[0]};
    Full_Adder FA_3174(s3174, c3174, in3174_1, in3174_2, s2805[0]);
    wire[0:0] s3175, in3175_1, in3175_2;
    wire c3175;
    assign in3175_1 = {s2343[0]};
    assign in3175_2 = {c2805};
    Full_Adder FA_3175(s3175, c3175, in3175_1, in3175_2, s2342[0]);
    wire[0:0] s3176, in3176_1, in3176_2;
    wire c3176;
    assign in3176_1 = {c2807};
    assign in3176_2 = {c2808};
    Full_Adder FA_3176(s3176, c3176, in3176_1, in3176_2, c2806);
    wire[0:0] s3177, in3177_1, in3177_2;
    wire c3177;
    assign in3177_1 = {s2810[0]};
    assign in3177_2 = {s2811[0]};
    Full_Adder FA_3177(s3177, c3177, in3177_1, in3177_2, s2809[0]);
    wire[0:0] s3178, in3178_1, in3178_2;
    wire c3178;
    assign in3178_1 = {s2349[0]};
    assign in3178_2 = {c2809};
    Full_Adder FA_3178(s3178, c3178, in3178_1, in3178_2, s2348[0]);
    wire[0:0] s3179, in3179_1, in3179_2;
    wire c3179;
    assign in3179_1 = {c2811};
    assign in3179_2 = {c2812};
    Full_Adder FA_3179(s3179, c3179, in3179_1, in3179_2, c2810);
    wire[0:0] s3180, in3180_1, in3180_2;
    wire c3180;
    assign in3180_1 = {s2814[0]};
    assign in3180_2 = {s2815[0]};
    Full_Adder FA_3180(s3180, c3180, in3180_1, in3180_2, s2813[0]);
    wire[0:0] s3181, in3181_1, in3181_2;
    wire c3181;
    assign in3181_1 = {s2355[0]};
    assign in3181_2 = {c2813};
    Full_Adder FA_3181(s3181, c3181, in3181_1, in3181_2, s2354[0]);
    wire[0:0] s3182, in3182_1, in3182_2;
    wire c3182;
    assign in3182_1 = {c2815};
    assign in3182_2 = {c2816};
    Full_Adder FA_3182(s3182, c3182, in3182_1, in3182_2, c2814);
    wire[0:0] s3183, in3183_1, in3183_2;
    wire c3183;
    assign in3183_1 = {s2818[0]};
    assign in3183_2 = {s2819[0]};
    Full_Adder FA_3183(s3183, c3183, in3183_1, in3183_2, s2817[0]);
    wire[0:0] s3184, in3184_1, in3184_2;
    wire c3184;
    assign in3184_1 = {s2361[0]};
    assign in3184_2 = {c2817};
    Full_Adder FA_3184(s3184, c3184, in3184_1, in3184_2, s2360[0]);
    wire[0:0] s3185, in3185_1, in3185_2;
    wire c3185;
    assign in3185_1 = {c2819};
    assign in3185_2 = {c2820};
    Full_Adder FA_3185(s3185, c3185, in3185_1, in3185_2, c2818);
    wire[0:0] s3186, in3186_1, in3186_2;
    wire c3186;
    assign in3186_1 = {s2822[0]};
    assign in3186_2 = {s2823[0]};
    Full_Adder FA_3186(s3186, c3186, in3186_1, in3186_2, s2821[0]);
    wire[0:0] s3187, in3187_1, in3187_2;
    wire c3187;
    assign in3187_1 = {s2367[0]};
    assign in3187_2 = {c2821};
    Full_Adder FA_3187(s3187, c3187, in3187_1, in3187_2, s2366[0]);
    wire[0:0] s3188, in3188_1, in3188_2;
    wire c3188;
    assign in3188_1 = {c2823};
    assign in3188_2 = {c2824};
    Full_Adder FA_3188(s3188, c3188, in3188_1, in3188_2, c2822);
    wire[0:0] s3189, in3189_1, in3189_2;
    wire c3189;
    assign in3189_1 = {s2826[0]};
    assign in3189_2 = {s2827[0]};
    Full_Adder FA_3189(s3189, c3189, in3189_1, in3189_2, s2825[0]);
    wire[0:0] s3190, in3190_1, in3190_2;
    wire c3190;
    assign in3190_1 = {s2373[0]};
    assign in3190_2 = {c2825};
    Full_Adder FA_3190(s3190, c3190, in3190_1, in3190_2, s2372[0]);
    wire[0:0] s3191, in3191_1, in3191_2;
    wire c3191;
    assign in3191_1 = {c2827};
    assign in3191_2 = {c2828};
    Full_Adder FA_3191(s3191, c3191, in3191_1, in3191_2, c2826);
    wire[0:0] s3192, in3192_1, in3192_2;
    wire c3192;
    assign in3192_1 = {s2830[0]};
    assign in3192_2 = {s2831[0]};
    Full_Adder FA_3192(s3192, c3192, in3192_1, in3192_2, s2829[0]);
    wire[0:0] s3193, in3193_1, in3193_2;
    wire c3193;
    assign in3193_1 = {s2379[0]};
    assign in3193_2 = {c2829};
    Full_Adder FA_3193(s3193, c3193, in3193_1, in3193_2, s2378[0]);
    wire[0:0] s3194, in3194_1, in3194_2;
    wire c3194;
    assign in3194_1 = {c2831};
    assign in3194_2 = {c2832};
    Full_Adder FA_3194(s3194, c3194, in3194_1, in3194_2, c2830);
    wire[0:0] s3195, in3195_1, in3195_2;
    wire c3195;
    assign in3195_1 = {s2834[0]};
    assign in3195_2 = {s2835[0]};
    Full_Adder FA_3195(s3195, c3195, in3195_1, in3195_2, s2833[0]);
    wire[0:0] s3196, in3196_1, in3196_2;
    wire c3196;
    assign in3196_1 = {s2385[0]};
    assign in3196_2 = {c2833};
    Full_Adder FA_3196(s3196, c3196, in3196_1, in3196_2, s2384[0]);
    wire[0:0] s3197, in3197_1, in3197_2;
    wire c3197;
    assign in3197_1 = {c2835};
    assign in3197_2 = {c2836};
    Full_Adder FA_3197(s3197, c3197, in3197_1, in3197_2, c2834);
    wire[0:0] s3198, in3198_1, in3198_2;
    wire c3198;
    assign in3198_1 = {s2838[0]};
    assign in3198_2 = {s2839[0]};
    Full_Adder FA_3198(s3198, c3198, in3198_1, in3198_2, s2837[0]);
    wire[0:0] s3199, in3199_1, in3199_2;
    wire c3199;
    assign in3199_1 = {s2391[0]};
    assign in3199_2 = {c2837};
    Full_Adder FA_3199(s3199, c3199, in3199_1, in3199_2, s2390[0]);
    wire[0:0] s3200, in3200_1, in3200_2;
    wire c3200;
    assign in3200_1 = {c2839};
    assign in3200_2 = {c2840};
    Full_Adder FA_3200(s3200, c3200, in3200_1, in3200_2, c2838);
    wire[0:0] s3201, in3201_1, in3201_2;
    wire c3201;
    assign in3201_1 = {s2842[0]};
    assign in3201_2 = {s2843[0]};
    Full_Adder FA_3201(s3201, c3201, in3201_1, in3201_2, s2841[0]);
    wire[0:0] s3202, in3202_1, in3202_2;
    wire c3202;
    assign in3202_1 = {s2397[0]};
    assign in3202_2 = {c2841};
    Full_Adder FA_3202(s3202, c3202, in3202_1, in3202_2, s2396[0]);
    wire[0:0] s3203, in3203_1, in3203_2;
    wire c3203;
    assign in3203_1 = {c2843};
    assign in3203_2 = {c2844};
    Full_Adder FA_3203(s3203, c3203, in3203_1, in3203_2, c2842);
    wire[0:0] s3204, in3204_1, in3204_2;
    wire c3204;
    assign in3204_1 = {s2846[0]};
    assign in3204_2 = {s2847[0]};
    Full_Adder FA_3204(s3204, c3204, in3204_1, in3204_2, s2845[0]);
    wire[0:0] s3205, in3205_1, in3205_2;
    wire c3205;
    assign in3205_1 = {s2403[0]};
    assign in3205_2 = {c2845};
    Full_Adder FA_3205(s3205, c3205, in3205_1, in3205_2, s2402[0]);
    wire[0:0] s3206, in3206_1, in3206_2;
    wire c3206;
    assign in3206_1 = {c2847};
    assign in3206_2 = {c2848};
    Full_Adder FA_3206(s3206, c3206, in3206_1, in3206_2, c2846);
    wire[0:0] s3207, in3207_1, in3207_2;
    wire c3207;
    assign in3207_1 = {s2850[0]};
    assign in3207_2 = {s2851[0]};
    Full_Adder FA_3207(s3207, c3207, in3207_1, in3207_2, s2849[0]);
    wire[0:0] s3208, in3208_1, in3208_2;
    wire c3208;
    assign in3208_1 = {s2409[0]};
    assign in3208_2 = {c2849};
    Full_Adder FA_3208(s3208, c3208, in3208_1, in3208_2, s2408[0]);
    wire[0:0] s3209, in3209_1, in3209_2;
    wire c3209;
    assign in3209_1 = {c2851};
    assign in3209_2 = {c2852};
    Full_Adder FA_3209(s3209, c3209, in3209_1, in3209_2, c2850);
    wire[0:0] s3210, in3210_1, in3210_2;
    wire c3210;
    assign in3210_1 = {s2854[0]};
    assign in3210_2 = {s2855[0]};
    Full_Adder FA_3210(s3210, c3210, in3210_1, in3210_2, s2853[0]);
    wire[0:0] s3211, in3211_1, in3211_2;
    wire c3211;
    assign in3211_1 = {s2415[0]};
    assign in3211_2 = {c2853};
    Full_Adder FA_3211(s3211, c3211, in3211_1, in3211_2, s2414[0]);
    wire[0:0] s3212, in3212_1, in3212_2;
    wire c3212;
    assign in3212_1 = {c2855};
    assign in3212_2 = {c2856};
    Full_Adder FA_3212(s3212, c3212, in3212_1, in3212_2, c2854);
    wire[0:0] s3213, in3213_1, in3213_2;
    wire c3213;
    assign in3213_1 = {s2858[0]};
    assign in3213_2 = {s2859[0]};
    Full_Adder FA_3213(s3213, c3213, in3213_1, in3213_2, s2857[0]);
    wire[0:0] s3214, in3214_1, in3214_2;
    wire c3214;
    assign in3214_1 = {s2421[0]};
    assign in3214_2 = {c2857};
    Full_Adder FA_3214(s3214, c3214, in3214_1, in3214_2, s2420[0]);
    wire[0:0] s3215, in3215_1, in3215_2;
    wire c3215;
    assign in3215_1 = {c2859};
    assign in3215_2 = {c2860};
    Full_Adder FA_3215(s3215, c3215, in3215_1, in3215_2, c2858);
    wire[0:0] s3216, in3216_1, in3216_2;
    wire c3216;
    assign in3216_1 = {s2862[0]};
    assign in3216_2 = {s2863[0]};
    Full_Adder FA_3216(s3216, c3216, in3216_1, in3216_2, s2861[0]);
    wire[0:0] s3217, in3217_1, in3217_2;
    wire c3217;
    assign in3217_1 = {s2427[0]};
    assign in3217_2 = {c2861};
    Full_Adder FA_3217(s3217, c3217, in3217_1, in3217_2, s2426[0]);
    wire[0:0] s3218, in3218_1, in3218_2;
    wire c3218;
    assign in3218_1 = {c2863};
    assign in3218_2 = {c2864};
    Full_Adder FA_3218(s3218, c3218, in3218_1, in3218_2, c2862);
    wire[0:0] s3219, in3219_1, in3219_2;
    wire c3219;
    assign in3219_1 = {s2866[0]};
    assign in3219_2 = {s2867[0]};
    Full_Adder FA_3219(s3219, c3219, in3219_1, in3219_2, s2865[0]);
    wire[0:0] s3220, in3220_1, in3220_2;
    wire c3220;
    assign in3220_1 = {s2433[0]};
    assign in3220_2 = {c2865};
    Full_Adder FA_3220(s3220, c3220, in3220_1, in3220_2, s2432[0]);
    wire[0:0] s3221, in3221_1, in3221_2;
    wire c3221;
    assign in3221_1 = {c2867};
    assign in3221_2 = {c2868};
    Full_Adder FA_3221(s3221, c3221, in3221_1, in3221_2, c2866);
    wire[0:0] s3222, in3222_1, in3222_2;
    wire c3222;
    assign in3222_1 = {s2870[0]};
    assign in3222_2 = {s2871[0]};
    Full_Adder FA_3222(s3222, c3222, in3222_1, in3222_2, s2869[0]);
    wire[0:0] s3223, in3223_1, in3223_2;
    wire c3223;
    assign in3223_1 = {s2439[0]};
    assign in3223_2 = {c2869};
    Full_Adder FA_3223(s3223, c3223, in3223_1, in3223_2, s2438[0]);
    wire[0:0] s3224, in3224_1, in3224_2;
    wire c3224;
    assign in3224_1 = {c2871};
    assign in3224_2 = {c2872};
    Full_Adder FA_3224(s3224, c3224, in3224_1, in3224_2, c2870);
    wire[0:0] s3225, in3225_1, in3225_2;
    wire c3225;
    assign in3225_1 = {s2874[0]};
    assign in3225_2 = {s2875[0]};
    Full_Adder FA_3225(s3225, c3225, in3225_1, in3225_2, s2873[0]);
    wire[0:0] s3226, in3226_1, in3226_2;
    wire c3226;
    assign in3226_1 = {s2445[0]};
    assign in3226_2 = {c2873};
    Full_Adder FA_3226(s3226, c3226, in3226_1, in3226_2, s2444[0]);
    wire[0:0] s3227, in3227_1, in3227_2;
    wire c3227;
    assign in3227_1 = {c2875};
    assign in3227_2 = {c2876};
    Full_Adder FA_3227(s3227, c3227, in3227_1, in3227_2, c2874);
    wire[0:0] s3228, in3228_1, in3228_2;
    wire c3228;
    assign in3228_1 = {s2878[0]};
    assign in3228_2 = {s2879[0]};
    Full_Adder FA_3228(s3228, c3228, in3228_1, in3228_2, s2877[0]);
    wire[0:0] s3229, in3229_1, in3229_2;
    wire c3229;
    assign in3229_1 = {s2451[0]};
    assign in3229_2 = {c2877};
    Full_Adder FA_3229(s3229, c3229, in3229_1, in3229_2, s2450[0]);
    wire[0:0] s3230, in3230_1, in3230_2;
    wire c3230;
    assign in3230_1 = {c2879};
    assign in3230_2 = {c2880};
    Full_Adder FA_3230(s3230, c3230, in3230_1, in3230_2, c2878);
    wire[0:0] s3231, in3231_1, in3231_2;
    wire c3231;
    assign in3231_1 = {s2882[0]};
    assign in3231_2 = {s2883[0]};
    Full_Adder FA_3231(s3231, c3231, in3231_1, in3231_2, s2881[0]);
    wire[0:0] s3232, in3232_1, in3232_2;
    wire c3232;
    assign in3232_1 = {s2457[0]};
    assign in3232_2 = {c2881};
    Full_Adder FA_3232(s3232, c3232, in3232_1, in3232_2, s2456[0]);
    wire[0:0] s3233, in3233_1, in3233_2;
    wire c3233;
    assign in3233_1 = {c2883};
    assign in3233_2 = {c2884};
    Full_Adder FA_3233(s3233, c3233, in3233_1, in3233_2, c2882);
    wire[0:0] s3234, in3234_1, in3234_2;
    wire c3234;
    assign in3234_1 = {s2886[0]};
    assign in3234_2 = {s2887[0]};
    Full_Adder FA_3234(s3234, c3234, in3234_1, in3234_2, s2885[0]);
    wire[0:0] s3235, in3235_1, in3235_2;
    wire c3235;
    assign in3235_1 = {s2463[0]};
    assign in3235_2 = {c2885};
    Full_Adder FA_3235(s3235, c3235, in3235_1, in3235_2, s2462[0]);
    wire[0:0] s3236, in3236_1, in3236_2;
    wire c3236;
    assign in3236_1 = {c2887};
    assign in3236_2 = {c2888};
    Full_Adder FA_3236(s3236, c3236, in3236_1, in3236_2, c2886);
    wire[0:0] s3237, in3237_1, in3237_2;
    wire c3237;
    assign in3237_1 = {s2890[0]};
    assign in3237_2 = {s2891[0]};
    Full_Adder FA_3237(s3237, c3237, in3237_1, in3237_2, s2889[0]);
    wire[0:0] s3238, in3238_1, in3238_2;
    wire c3238;
    assign in3238_1 = {s2469[0]};
    assign in3238_2 = {c2889};
    Full_Adder FA_3238(s3238, c3238, in3238_1, in3238_2, s2468[0]);
    wire[0:0] s3239, in3239_1, in3239_2;
    wire c3239;
    assign in3239_1 = {c2891};
    assign in3239_2 = {c2892};
    Full_Adder FA_3239(s3239, c3239, in3239_1, in3239_2, c2890);
    wire[0:0] s3240, in3240_1, in3240_2;
    wire c3240;
    assign in3240_1 = {s2894[0]};
    assign in3240_2 = {s2895[0]};
    Full_Adder FA_3240(s3240, c3240, in3240_1, in3240_2, s2893[0]);
    wire[0:0] s3241, in3241_1, in3241_2;
    wire c3241;
    assign in3241_1 = {s2475[0]};
    assign in3241_2 = {c2893};
    Full_Adder FA_3241(s3241, c3241, in3241_1, in3241_2, s2474[0]);
    wire[0:0] s3242, in3242_1, in3242_2;
    wire c3242;
    assign in3242_1 = {c2895};
    assign in3242_2 = {c2896};
    Full_Adder FA_3242(s3242, c3242, in3242_1, in3242_2, c2894);
    wire[0:0] s3243, in3243_1, in3243_2;
    wire c3243;
    assign in3243_1 = {s2898[0]};
    assign in3243_2 = {s2899[0]};
    Full_Adder FA_3243(s3243, c3243, in3243_1, in3243_2, s2897[0]);
    wire[0:0] s3244, in3244_1, in3244_2;
    wire c3244;
    assign in3244_1 = {s2481[0]};
    assign in3244_2 = {c2897};
    Full_Adder FA_3244(s3244, c3244, in3244_1, in3244_2, s2480[0]);
    wire[0:0] s3245, in3245_1, in3245_2;
    wire c3245;
    assign in3245_1 = {c2899};
    assign in3245_2 = {c2900};
    Full_Adder FA_3245(s3245, c3245, in3245_1, in3245_2, c2898);
    wire[0:0] s3246, in3246_1, in3246_2;
    wire c3246;
    assign in3246_1 = {s2902[0]};
    assign in3246_2 = {s2903[0]};
    Full_Adder FA_3246(s3246, c3246, in3246_1, in3246_2, s2901[0]);
    wire[0:0] s3247, in3247_1, in3247_2;
    wire c3247;
    assign in3247_1 = {s2487[0]};
    assign in3247_2 = {c2901};
    Full_Adder FA_3247(s3247, c3247, in3247_1, in3247_2, s2486[0]);
    wire[0:0] s3248, in3248_1, in3248_2;
    wire c3248;
    assign in3248_1 = {c2903};
    assign in3248_2 = {c2904};
    Full_Adder FA_3248(s3248, c3248, in3248_1, in3248_2, c2902);
    wire[0:0] s3249, in3249_1, in3249_2;
    wire c3249;
    assign in3249_1 = {s2906[0]};
    assign in3249_2 = {s2907[0]};
    Full_Adder FA_3249(s3249, c3249, in3249_1, in3249_2, s2905[0]);
    wire[0:0] s3250, in3250_1, in3250_2;
    wire c3250;
    assign in3250_1 = {s2493[0]};
    assign in3250_2 = {c2905};
    Full_Adder FA_3250(s3250, c3250, in3250_1, in3250_2, s2492[0]);
    wire[0:0] s3251, in3251_1, in3251_2;
    wire c3251;
    assign in3251_1 = {c2907};
    assign in3251_2 = {c2908};
    Full_Adder FA_3251(s3251, c3251, in3251_1, in3251_2, c2906);
    wire[0:0] s3252, in3252_1, in3252_2;
    wire c3252;
    assign in3252_1 = {s2910[0]};
    assign in3252_2 = {s2911[0]};
    Full_Adder FA_3252(s3252, c3252, in3252_1, in3252_2, s2909[0]);
    wire[0:0] s3253, in3253_1, in3253_2;
    wire c3253;
    assign in3253_1 = {s2499[0]};
    assign in3253_2 = {c2909};
    Full_Adder FA_3253(s3253, c3253, in3253_1, in3253_2, s2498[0]);
    wire[0:0] s3254, in3254_1, in3254_2;
    wire c3254;
    assign in3254_1 = {c2911};
    assign in3254_2 = {c2912};
    Full_Adder FA_3254(s3254, c3254, in3254_1, in3254_2, c2910);
    wire[0:0] s3255, in3255_1, in3255_2;
    wire c3255;
    assign in3255_1 = {s2914[0]};
    assign in3255_2 = {s2915[0]};
    Full_Adder FA_3255(s3255, c3255, in3255_1, in3255_2, s2913[0]);
    wire[0:0] s3256, in3256_1, in3256_2;
    wire c3256;
    assign in3256_1 = {s2505[0]};
    assign in3256_2 = {c2913};
    Full_Adder FA_3256(s3256, c3256, in3256_1, in3256_2, s2504[0]);
    wire[0:0] s3257, in3257_1, in3257_2;
    wire c3257;
    assign in3257_1 = {c2915};
    assign in3257_2 = {c2916};
    Full_Adder FA_3257(s3257, c3257, in3257_1, in3257_2, c2914);
    wire[0:0] s3258, in3258_1, in3258_2;
    wire c3258;
    assign in3258_1 = {s2918[0]};
    assign in3258_2 = {s2919[0]};
    Full_Adder FA_3258(s3258, c3258, in3258_1, in3258_2, s2917[0]);
    wire[0:0] s3259, in3259_1, in3259_2;
    wire c3259;
    assign in3259_1 = {s2511[0]};
    assign in3259_2 = {c2917};
    Full_Adder FA_3259(s3259, c3259, in3259_1, in3259_2, s2510[0]);
    wire[0:0] s3260, in3260_1, in3260_2;
    wire c3260;
    assign in3260_1 = {c2919};
    assign in3260_2 = {c2920};
    Full_Adder FA_3260(s3260, c3260, in3260_1, in3260_2, c2918);
    wire[0:0] s3261, in3261_1, in3261_2;
    wire c3261;
    assign in3261_1 = {s2922[0]};
    assign in3261_2 = {s2923[0]};
    Full_Adder FA_3261(s3261, c3261, in3261_1, in3261_2, s2921[0]);
    wire[0:0] s3262, in3262_1, in3262_2;
    wire c3262;
    assign in3262_1 = {s2517[0]};
    assign in3262_2 = {c2921};
    Full_Adder FA_3262(s3262, c3262, in3262_1, in3262_2, s2516[0]);
    wire[0:0] s3263, in3263_1, in3263_2;
    wire c3263;
    assign in3263_1 = {c2923};
    assign in3263_2 = {c2924};
    Full_Adder FA_3263(s3263, c3263, in3263_1, in3263_2, c2922);
    wire[0:0] s3264, in3264_1, in3264_2;
    wire c3264;
    assign in3264_1 = {s2926[0]};
    assign in3264_2 = {s2927[0]};
    Full_Adder FA_3264(s3264, c3264, in3264_1, in3264_2, s2925[0]);
    wire[0:0] s3265, in3265_1, in3265_2;
    wire c3265;
    assign in3265_1 = {s2523[0]};
    assign in3265_2 = {c2925};
    Full_Adder FA_3265(s3265, c3265, in3265_1, in3265_2, s2522[0]);
    wire[0:0] s3266, in3266_1, in3266_2;
    wire c3266;
    assign in3266_1 = {c2927};
    assign in3266_2 = {c2928};
    Full_Adder FA_3266(s3266, c3266, in3266_1, in3266_2, c2926);
    wire[0:0] s3267, in3267_1, in3267_2;
    wire c3267;
    assign in3267_1 = {s2930[0]};
    assign in3267_2 = {s2931[0]};
    Full_Adder FA_3267(s3267, c3267, in3267_1, in3267_2, s2929[0]);
    wire[0:0] s3268, in3268_1, in3268_2;
    wire c3268;
    assign in3268_1 = {s2529[0]};
    assign in3268_2 = {c2929};
    Full_Adder FA_3268(s3268, c3268, in3268_1, in3268_2, s2528[0]);
    wire[0:0] s3269, in3269_1, in3269_2;
    wire c3269;
    assign in3269_1 = {c2931};
    assign in3269_2 = {c2932};
    Full_Adder FA_3269(s3269, c3269, in3269_1, in3269_2, c2930);
    wire[0:0] s3270, in3270_1, in3270_2;
    wire c3270;
    assign in3270_1 = {s2934[0]};
    assign in3270_2 = {s2935[0]};
    Full_Adder FA_3270(s3270, c3270, in3270_1, in3270_2, s2933[0]);
    wire[0:0] s3271, in3271_1, in3271_2;
    wire c3271;
    assign in3271_1 = {s2535[0]};
    assign in3271_2 = {c2933};
    Full_Adder FA_3271(s3271, c3271, in3271_1, in3271_2, s2534[0]);
    wire[0:0] s3272, in3272_1, in3272_2;
    wire c3272;
    assign in3272_1 = {c2935};
    assign in3272_2 = {c2936};
    Full_Adder FA_3272(s3272, c3272, in3272_1, in3272_2, c2934);
    wire[0:0] s3273, in3273_1, in3273_2;
    wire c3273;
    assign in3273_1 = {s2938[0]};
    assign in3273_2 = {s2939[0]};
    Full_Adder FA_3273(s3273, c3273, in3273_1, in3273_2, s2937[0]);
    wire[0:0] s3274, in3274_1, in3274_2;
    wire c3274;
    assign in3274_1 = {s2540[0]};
    assign in3274_2 = {c2937};
    Full_Adder FA_3274(s3274, c3274, in3274_1, in3274_2, s2539[0]);
    wire[0:0] s3275, in3275_1, in3275_2;
    wire c3275;
    assign in3275_1 = {c2939};
    assign in3275_2 = {c2940};
    Full_Adder FA_3275(s3275, c3275, in3275_1, in3275_2, c2938);
    wire[0:0] s3276, in3276_1, in3276_2;
    wire c3276;
    assign in3276_1 = {s2942[0]};
    assign in3276_2 = {s2943[0]};
    Full_Adder FA_3276(s3276, c3276, in3276_1, in3276_2, s2941[0]);
    wire[0:0] s3277, in3277_1, in3277_2;
    wire c3277;
    assign in3277_1 = {s2544[0]};
    assign in3277_2 = {c2941};
    Full_Adder FA_3277(s3277, c3277, in3277_1, in3277_2, s2543[0]);
    wire[0:0] s3278, in3278_1, in3278_2;
    wire c3278;
    assign in3278_1 = {c2943};
    assign in3278_2 = {c2944};
    Full_Adder FA_3278(s3278, c3278, in3278_1, in3278_2, c2942);
    wire[0:0] s3279, in3279_1, in3279_2;
    wire c3279;
    assign in3279_1 = {s2946[0]};
    assign in3279_2 = {s2947[0]};
    Full_Adder FA_3279(s3279, c3279, in3279_1, in3279_2, s2945[0]);
    wire[0:0] s3280, in3280_1, in3280_2;
    wire c3280;
    assign in3280_1 = {s2547[0]};
    assign in3280_2 = {c2945};
    Full_Adder FA_3280(s3280, c3280, in3280_1, in3280_2, s2546[0]);
    wire[0:0] s3281, in3281_1, in3281_2;
    wire c3281;
    assign in3281_1 = {c2947};
    assign in3281_2 = {c2948};
    Full_Adder FA_3281(s3281, c3281, in3281_1, in3281_2, c2946);
    wire[0:0] s3282, in3282_1, in3282_2;
    wire c3282;
    assign in3282_1 = {s2950[0]};
    assign in3282_2 = {s2951[0]};
    Full_Adder FA_3282(s3282, c3282, in3282_1, in3282_2, s2949[0]);
    wire[0:0] s3283, in3283_1, in3283_2;
    wire c3283;
    assign in3283_1 = {s2549[0]};
    assign in3283_2 = {c2949};
    Full_Adder FA_3283(s3283, c3283, in3283_1, in3283_2, s2548[0]);
    wire[0:0] s3284, in3284_1, in3284_2;
    wire c3284;
    assign in3284_1 = {c2951};
    assign in3284_2 = {c2952};
    Full_Adder FA_3284(s3284, c3284, in3284_1, in3284_2, c2950);
    wire[0:0] s3285, in3285_1, in3285_2;
    wire c3285;
    assign in3285_1 = {s2954[0]};
    assign in3285_2 = {s2955[0]};
    Full_Adder FA_3285(s3285, c3285, in3285_1, in3285_2, s2953[0]);
    wire[0:0] s3286, in3286_1, in3286_2;
    wire c3286;
    assign in3286_1 = {s2550[0]};
    assign in3286_2 = {c2953};
    Full_Adder FA_3286(s3286, c3286, in3286_1, in3286_2, c2549);
    wire[0:0] s3287, in3287_1, in3287_2;
    wire c3287;
    assign in3287_1 = {c2955};
    assign in3287_2 = {c2956};
    Full_Adder FA_3287(s3287, c3287, in3287_1, in3287_2, c2954);
    wire[0:0] s3288, in3288_1, in3288_2;
    wire c3288;
    assign in3288_1 = {s2958[0]};
    assign in3288_2 = {s2959[0]};
    Full_Adder FA_3288(s3288, c3288, in3288_1, in3288_2, s2957[0]);
    wire[0:0] s3289, in3289_1, in3289_2;
    wire c3289;
    assign in3289_1 = {c2550};
    assign in3289_2 = {c2957};
    Full_Adder FA_3289(s3289, c3289, in3289_1, in3289_2, pp63[51]);
    wire[0:0] s3290, in3290_1, in3290_2;
    wire c3290;
    assign in3290_1 = {c2959};
    assign in3290_2 = {c2960};
    Full_Adder FA_3290(s3290, c3290, in3290_1, in3290_2, c2958);
    wire[0:0] s3291, in3291_1, in3291_2;
    wire c3291;
    assign in3291_1 = {s2962[0]};
    assign in3291_2 = {s2963[0]};
    Full_Adder FA_3291(s3291, c3291, in3291_1, in3291_2, s2961[0]);
    wire[0:0] s3292, in3292_1, in3292_2;
    wire c3292;
    assign in3292_1 = {pp62[53]};
    assign in3292_2 = {pp63[52]};
    Full_Adder FA_3292(s3292, c3292, in3292_1, in3292_2, pp61[54]);
    wire[0:0] s3293, in3293_1, in3293_2;
    wire c3293;
    assign in3293_1 = {c2962};
    assign in3293_2 = {c2963};
    Full_Adder FA_3293(s3293, c3293, in3293_1, in3293_2, c2961);
    wire[0:0] s3294, in3294_1, in3294_2;
    wire c3294;
    assign in3294_1 = {s2965[0]};
    assign in3294_2 = {s2966[0]};
    Full_Adder FA_3294(s3294, c3294, in3294_1, in3294_2, c2964);
    wire[0:0] s3295, in3295_1, in3295_2;
    wire c3295;
    assign in3295_1 = {pp60[56]};
    assign in3295_2 = {pp61[55]};
    Full_Adder FA_3295(s3295, c3295, in3295_1, in3295_2, pp59[57]);
    wire[0:0] s3296, in3296_1, in3296_2;
    wire c3296;
    assign in3296_1 = {pp63[53]};
    assign in3296_2 = {c2965};
    Full_Adder FA_3296(s3296, c3296, in3296_1, in3296_2, pp62[54]);
    wire[0:0] s3297, in3297_1, in3297_2;
    wire c3297;
    assign in3297_1 = {c2967};
    assign in3297_2 = {s2968[0]};
    Full_Adder FA_3297(s3297, c3297, in3297_1, in3297_2, c2966);
    wire[0:0] s3298, in3298_1, in3298_2;
    wire c3298;
    assign in3298_1 = {pp58[59]};
    assign in3298_2 = {pp59[58]};
    Full_Adder FA_3298(s3298, c3298, in3298_1, in3298_2, pp57[60]);
    wire[0:0] s3299, in3299_1, in3299_2;
    wire c3299;
    assign in3299_1 = {pp61[56]};
    assign in3299_2 = {pp62[55]};
    Full_Adder FA_3299(s3299, c3299, in3299_1, in3299_2, pp60[57]);
    wire[0:0] s3300, in3300_1, in3300_2;
    wire c3300;
    assign in3300_1 = {c2968};
    assign in3300_2 = {c2969};
    Full_Adder FA_3300(s3300, c3300, in3300_1, in3300_2, pp63[54]);
    wire[0:0] s3301, in3301_1, in3301_2;
    wire c3301;
    assign in3301_1 = {pp56[62]};
    assign in3301_2 = {pp57[61]};
    Full_Adder FA_3301(s3301, c3301, in3301_1, in3301_2, pp55[63]);
    wire[0:0] s3302, in3302_1, in3302_2;
    wire c3302;
    assign in3302_1 = {pp59[59]};
    assign in3302_2 = {pp60[58]};
    Full_Adder FA_3302(s3302, c3302, in3302_1, in3302_2, pp58[60]);
    wire[0:0] s3303, in3303_1, in3303_2;
    wire c3303;
    assign in3303_1 = {pp62[56]};
    assign in3303_2 = {pp63[55]};
    Full_Adder FA_3303(s3303, c3303, in3303_1, in3303_2, pp61[57]);
    wire[0:0] s3304, in3304_1, in3304_2;
    wire c3304;
    assign in3304_1 = {pp57[62]};
    assign in3304_2 = {pp58[61]};
    Full_Adder FA_3304(s3304, c3304, in3304_1, in3304_2, pp56[63]);
    wire[0:0] s3305, in3305_1, in3305_2;
    wire c3305;
    assign in3305_1 = {pp60[59]};
    assign in3305_2 = {pp61[58]};
    Full_Adder FA_3305(s3305, c3305, in3305_1, in3305_2, pp59[60]);
    wire[0:0] s3306, in3306_1, in3306_2;
    wire c3306;
    assign in3306_1 = {pp58[62]};
    assign in3306_2 = {pp59[61]};
    Full_Adder FA_3306(s3306, c3306, in3306_1, in3306_2, pp57[63]);

    /*Stage 7*/
    wire[0:0] s3307, in3307_1, in3307_2;
    wire c3307;
    assign in3307_1 = {pp0[5]};
    assign in3307_2 = {pp1[4]};
    Half_Adder HA_3307(s3307, c3307, in3307_1, in3307_2);
    wire[0:0] s3308, in3308_1, in3308_2;
    wire c3308;
    assign in3308_1 = {pp1[5]};
    assign in3308_2 = {pp2[4]};
    Full_Adder FA_3308(s3308, c3308, in3308_1, in3308_2, pp0[6]);
    wire[0:0] s3309, in3309_1, in3309_2;
    wire c3309;
    assign in3309_1 = {pp3[3]};
    assign in3309_2 = {pp4[2]};
    Half_Adder HA_3309(s3309, c3309, in3309_1, in3309_2);
    wire[0:0] s3310, in3310_1, in3310_2;
    wire c3310;
    assign in3310_1 = {pp3[4]};
    assign in3310_2 = {pp4[3]};
    Full_Adder FA_3310(s3310, c3310, in3310_1, in3310_2, pp2[5]);
    wire[0:0] s3311, in3311_1, in3311_2;
    wire c3311;
    assign in3311_1 = {pp6[1]};
    assign in3311_2 = {pp7[0]};
    Full_Adder FA_3311(s3311, c3311, in3311_1, in3311_2, pp5[2]);
    wire[0:0] s3312, in3312_1, in3312_2;
    wire c3312;
    assign in3312_1 = {pp6[2]};
    assign in3312_2 = {pp7[1]};
    Full_Adder FA_3312(s3312, c3312, in3312_1, in3312_2, pp5[3]);
    wire[0:0] s3313, in3313_1, in3313_2;
    wire c3313;
    assign in3313_1 = {c2971};
    assign in3313_2 = {s2972[0]};
    Full_Adder FA_3313(s3313, c3313, in3313_1, in3313_2, pp8[0]);
    wire[0:0] s3314, in3314_1, in3314_2;
    wire c3314;
    assign in3314_1 = {pp9[0]};
    assign in3314_2 = {c2972};
    Full_Adder FA_3314(s3314, c3314, in3314_1, in3314_2, pp8[1]);
    wire[0:0] s3315, in3315_1, in3315_2;
    wire c3315;
    assign in3315_1 = {s2974[0]};
    assign in3315_2 = {s2975[0]};
    Full_Adder FA_3315(s3315, c3315, in3315_1, in3315_2, c2973);
    wire[0:0] s3316, in3316_1, in3316_2;
    wire c3316;
    assign in3316_1 = {c2974};
    assign in3316_2 = {c2975};
    Full_Adder FA_3316(s3316, c3316, in3316_1, in3316_2, s2551[0]);
    wire[0:0] s3317, in3317_1, in3317_2;
    wire c3317;
    assign in3317_1 = {s2977[0]};
    assign in3317_2 = {s2978[0]};
    Full_Adder FA_3317(s3317, c3317, in3317_1, in3317_2, c2976);
    wire[0:0] s3318, in3318_1, in3318_2;
    wire c3318;
    assign in3318_1 = {c2977};
    assign in3318_2 = {c2978};
    Full_Adder FA_3318(s3318, c3318, in3318_1, in3318_2, s2553[0]);
    wire[0:0] s3319, in3319_1, in3319_2;
    wire c3319;
    assign in3319_1 = {s2980[0]};
    assign in3319_2 = {s2981[0]};
    Full_Adder FA_3319(s3319, c3319, in3319_1, in3319_2, c2979);
    wire[0:0] s3320, in3320_1, in3320_2;
    wire c3320;
    assign in3320_1 = {c2980};
    assign in3320_2 = {c2981};
    Full_Adder FA_3320(s3320, c3320, in3320_1, in3320_2, s2556[0]);
    wire[0:0] s3321, in3321_1, in3321_2;
    wire c3321;
    assign in3321_1 = {s2983[0]};
    assign in3321_2 = {s2984[0]};
    Full_Adder FA_3321(s3321, c3321, in3321_1, in3321_2, c2982);
    wire[0:0] s3322, in3322_1, in3322_2;
    wire c3322;
    assign in3322_1 = {c2983};
    assign in3322_2 = {c2984};
    Full_Adder FA_3322(s3322, c3322, in3322_1, in3322_2, s2560[0]);
    wire[0:0] s3323, in3323_1, in3323_2;
    wire c3323;
    assign in3323_1 = {s2986[0]};
    assign in3323_2 = {s2987[0]};
    Full_Adder FA_3323(s3323, c3323, in3323_1, in3323_2, c2985);
    wire[0:0] s3324, in3324_1, in3324_2;
    wire c3324;
    assign in3324_1 = {c2986};
    assign in3324_2 = {c2987};
    Full_Adder FA_3324(s3324, c3324, in3324_1, in3324_2, s2564[0]);
    wire[0:0] s3325, in3325_1, in3325_2;
    wire c3325;
    assign in3325_1 = {s2989[0]};
    assign in3325_2 = {s2990[0]};
    Full_Adder FA_3325(s3325, c3325, in3325_1, in3325_2, c2988);
    wire[0:0] s3326, in3326_1, in3326_2;
    wire c3326;
    assign in3326_1 = {c2989};
    assign in3326_2 = {c2990};
    Full_Adder FA_3326(s3326, c3326, in3326_1, in3326_2, s2568[0]);
    wire[0:0] s3327, in3327_1, in3327_2;
    wire c3327;
    assign in3327_1 = {s2992[0]};
    assign in3327_2 = {s2993[0]};
    Full_Adder FA_3327(s3327, c3327, in3327_1, in3327_2, c2991);
    wire[0:0] s3328, in3328_1, in3328_2;
    wire c3328;
    assign in3328_1 = {c2992};
    assign in3328_2 = {c2993};
    Full_Adder FA_3328(s3328, c3328, in3328_1, in3328_2, s2572[0]);
    wire[0:0] s3329, in3329_1, in3329_2;
    wire c3329;
    assign in3329_1 = {s2995[0]};
    assign in3329_2 = {s2996[0]};
    Full_Adder FA_3329(s3329, c3329, in3329_1, in3329_2, c2994);
    wire[0:0] s3330, in3330_1, in3330_2;
    wire c3330;
    assign in3330_1 = {c2995};
    assign in3330_2 = {c2996};
    Full_Adder FA_3330(s3330, c3330, in3330_1, in3330_2, s2576[0]);
    wire[0:0] s3331, in3331_1, in3331_2;
    wire c3331;
    assign in3331_1 = {s2998[0]};
    assign in3331_2 = {s2999[0]};
    Full_Adder FA_3331(s3331, c3331, in3331_1, in3331_2, c2997);
    wire[0:0] s3332, in3332_1, in3332_2;
    wire c3332;
    assign in3332_1 = {c2998};
    assign in3332_2 = {c2999};
    Full_Adder FA_3332(s3332, c3332, in3332_1, in3332_2, s2580[0]);
    wire[0:0] s3333, in3333_1, in3333_2;
    wire c3333;
    assign in3333_1 = {s3001[0]};
    assign in3333_2 = {s3002[0]};
    Full_Adder FA_3333(s3333, c3333, in3333_1, in3333_2, c3000);
    wire[0:0] s3334, in3334_1, in3334_2;
    wire c3334;
    assign in3334_1 = {c3001};
    assign in3334_2 = {c3002};
    Full_Adder FA_3334(s3334, c3334, in3334_1, in3334_2, s2584[0]);
    wire[0:0] s3335, in3335_1, in3335_2;
    wire c3335;
    assign in3335_1 = {s3004[0]};
    assign in3335_2 = {s3005[0]};
    Full_Adder FA_3335(s3335, c3335, in3335_1, in3335_2, c3003);
    wire[0:0] s3336, in3336_1, in3336_2;
    wire c3336;
    assign in3336_1 = {c3004};
    assign in3336_2 = {c3005};
    Full_Adder FA_3336(s3336, c3336, in3336_1, in3336_2, s2588[0]);
    wire[0:0] s3337, in3337_1, in3337_2;
    wire c3337;
    assign in3337_1 = {s3007[0]};
    assign in3337_2 = {s3008[0]};
    Full_Adder FA_3337(s3337, c3337, in3337_1, in3337_2, c3006);
    wire[0:0] s3338, in3338_1, in3338_2;
    wire c3338;
    assign in3338_1 = {c3007};
    assign in3338_2 = {c3008};
    Full_Adder FA_3338(s3338, c3338, in3338_1, in3338_2, s2592[0]);
    wire[0:0] s3339, in3339_1, in3339_2;
    wire c3339;
    assign in3339_1 = {s3010[0]};
    assign in3339_2 = {s3011[0]};
    Full_Adder FA_3339(s3339, c3339, in3339_1, in3339_2, c3009);
    wire[0:0] s3340, in3340_1, in3340_2;
    wire c3340;
    assign in3340_1 = {c3010};
    assign in3340_2 = {c3011};
    Full_Adder FA_3340(s3340, c3340, in3340_1, in3340_2, s2596[0]);
    wire[0:0] s3341, in3341_1, in3341_2;
    wire c3341;
    assign in3341_1 = {s3013[0]};
    assign in3341_2 = {s3014[0]};
    Full_Adder FA_3341(s3341, c3341, in3341_1, in3341_2, c3012);
    wire[0:0] s3342, in3342_1, in3342_2;
    wire c3342;
    assign in3342_1 = {c3013};
    assign in3342_2 = {c3014};
    Full_Adder FA_3342(s3342, c3342, in3342_1, in3342_2, s2600[0]);
    wire[0:0] s3343, in3343_1, in3343_2;
    wire c3343;
    assign in3343_1 = {s3016[0]};
    assign in3343_2 = {s3017[0]};
    Full_Adder FA_3343(s3343, c3343, in3343_1, in3343_2, c3015);
    wire[0:0] s3344, in3344_1, in3344_2;
    wire c3344;
    assign in3344_1 = {c3016};
    assign in3344_2 = {c3017};
    Full_Adder FA_3344(s3344, c3344, in3344_1, in3344_2, s2604[0]);
    wire[0:0] s3345, in3345_1, in3345_2;
    wire c3345;
    assign in3345_1 = {s3019[0]};
    assign in3345_2 = {s3020[0]};
    Full_Adder FA_3345(s3345, c3345, in3345_1, in3345_2, c3018);
    wire[0:0] s3346, in3346_1, in3346_2;
    wire c3346;
    assign in3346_1 = {c3019};
    assign in3346_2 = {c3020};
    Full_Adder FA_3346(s3346, c3346, in3346_1, in3346_2, s2608[0]);
    wire[0:0] s3347, in3347_1, in3347_2;
    wire c3347;
    assign in3347_1 = {s3022[0]};
    assign in3347_2 = {s3023[0]};
    Full_Adder FA_3347(s3347, c3347, in3347_1, in3347_2, c3021);
    wire[0:0] s3348, in3348_1, in3348_2;
    wire c3348;
    assign in3348_1 = {c3022};
    assign in3348_2 = {c3023};
    Full_Adder FA_3348(s3348, c3348, in3348_1, in3348_2, s2612[0]);
    wire[0:0] s3349, in3349_1, in3349_2;
    wire c3349;
    assign in3349_1 = {s3025[0]};
    assign in3349_2 = {s3026[0]};
    Full_Adder FA_3349(s3349, c3349, in3349_1, in3349_2, c3024);
    wire[0:0] s3350, in3350_1, in3350_2;
    wire c3350;
    assign in3350_1 = {c3025};
    assign in3350_2 = {c3026};
    Full_Adder FA_3350(s3350, c3350, in3350_1, in3350_2, s2616[0]);
    wire[0:0] s3351, in3351_1, in3351_2;
    wire c3351;
    assign in3351_1 = {s3028[0]};
    assign in3351_2 = {s3029[0]};
    Full_Adder FA_3351(s3351, c3351, in3351_1, in3351_2, c3027);
    wire[0:0] s3352, in3352_1, in3352_2;
    wire c3352;
    assign in3352_1 = {c3028};
    assign in3352_2 = {c3029};
    Full_Adder FA_3352(s3352, c3352, in3352_1, in3352_2, s2620[0]);
    wire[0:0] s3353, in3353_1, in3353_2;
    wire c3353;
    assign in3353_1 = {s3031[0]};
    assign in3353_2 = {s3032[0]};
    Full_Adder FA_3353(s3353, c3353, in3353_1, in3353_2, c3030);
    wire[0:0] s3354, in3354_1, in3354_2;
    wire c3354;
    assign in3354_1 = {c3031};
    assign in3354_2 = {c3032};
    Full_Adder FA_3354(s3354, c3354, in3354_1, in3354_2, s2624[0]);
    wire[0:0] s3355, in3355_1, in3355_2;
    wire c3355;
    assign in3355_1 = {s3034[0]};
    assign in3355_2 = {s3035[0]};
    Full_Adder FA_3355(s3355, c3355, in3355_1, in3355_2, c3033);
    wire[0:0] s3356, in3356_1, in3356_2;
    wire c3356;
    assign in3356_1 = {c3034};
    assign in3356_2 = {c3035};
    Full_Adder FA_3356(s3356, c3356, in3356_1, in3356_2, s2628[0]);
    wire[0:0] s3357, in3357_1, in3357_2;
    wire c3357;
    assign in3357_1 = {s3037[0]};
    assign in3357_2 = {s3038[0]};
    Full_Adder FA_3357(s3357, c3357, in3357_1, in3357_2, c3036);
    wire[0:0] s3358, in3358_1, in3358_2;
    wire c3358;
    assign in3358_1 = {c3037};
    assign in3358_2 = {c3038};
    Full_Adder FA_3358(s3358, c3358, in3358_1, in3358_2, s2632[0]);
    wire[0:0] s3359, in3359_1, in3359_2;
    wire c3359;
    assign in3359_1 = {s3040[0]};
    assign in3359_2 = {s3041[0]};
    Full_Adder FA_3359(s3359, c3359, in3359_1, in3359_2, c3039);
    wire[0:0] s3360, in3360_1, in3360_2;
    wire c3360;
    assign in3360_1 = {c3040};
    assign in3360_2 = {c3041};
    Full_Adder FA_3360(s3360, c3360, in3360_1, in3360_2, s2636[0]);
    wire[0:0] s3361, in3361_1, in3361_2;
    wire c3361;
    assign in3361_1 = {s3043[0]};
    assign in3361_2 = {s3044[0]};
    Full_Adder FA_3361(s3361, c3361, in3361_1, in3361_2, c3042);
    wire[0:0] s3362, in3362_1, in3362_2;
    wire c3362;
    assign in3362_1 = {c3043};
    assign in3362_2 = {c3044};
    Full_Adder FA_3362(s3362, c3362, in3362_1, in3362_2, s2640[0]);
    wire[0:0] s3363, in3363_1, in3363_2;
    wire c3363;
    assign in3363_1 = {s3046[0]};
    assign in3363_2 = {s3047[0]};
    Full_Adder FA_3363(s3363, c3363, in3363_1, in3363_2, c3045);
    wire[0:0] s3364, in3364_1, in3364_2;
    wire c3364;
    assign in3364_1 = {c3046};
    assign in3364_2 = {c3047};
    Full_Adder FA_3364(s3364, c3364, in3364_1, in3364_2, s2644[0]);
    wire[0:0] s3365, in3365_1, in3365_2;
    wire c3365;
    assign in3365_1 = {s3049[0]};
    assign in3365_2 = {s3050[0]};
    Full_Adder FA_3365(s3365, c3365, in3365_1, in3365_2, c3048);
    wire[0:0] s3366, in3366_1, in3366_2;
    wire c3366;
    assign in3366_1 = {c3049};
    assign in3366_2 = {c3050};
    Full_Adder FA_3366(s3366, c3366, in3366_1, in3366_2, s2648[0]);
    wire[0:0] s3367, in3367_1, in3367_2;
    wire c3367;
    assign in3367_1 = {s3052[0]};
    assign in3367_2 = {s3053[0]};
    Full_Adder FA_3367(s3367, c3367, in3367_1, in3367_2, c3051);
    wire[0:0] s3368, in3368_1, in3368_2;
    wire c3368;
    assign in3368_1 = {c3052};
    assign in3368_2 = {c3053};
    Full_Adder FA_3368(s3368, c3368, in3368_1, in3368_2, s2652[0]);
    wire[0:0] s3369, in3369_1, in3369_2;
    wire c3369;
    assign in3369_1 = {s3055[0]};
    assign in3369_2 = {s3056[0]};
    Full_Adder FA_3369(s3369, c3369, in3369_1, in3369_2, c3054);
    wire[0:0] s3370, in3370_1, in3370_2;
    wire c3370;
    assign in3370_1 = {c3055};
    assign in3370_2 = {c3056};
    Full_Adder FA_3370(s3370, c3370, in3370_1, in3370_2, s2656[0]);
    wire[0:0] s3371, in3371_1, in3371_2;
    wire c3371;
    assign in3371_1 = {s3058[0]};
    assign in3371_2 = {s3059[0]};
    Full_Adder FA_3371(s3371, c3371, in3371_1, in3371_2, c3057);
    wire[0:0] s3372, in3372_1, in3372_2;
    wire c3372;
    assign in3372_1 = {c3058};
    assign in3372_2 = {c3059};
    Full_Adder FA_3372(s3372, c3372, in3372_1, in3372_2, s2660[0]);
    wire[0:0] s3373, in3373_1, in3373_2;
    wire c3373;
    assign in3373_1 = {s3061[0]};
    assign in3373_2 = {s3062[0]};
    Full_Adder FA_3373(s3373, c3373, in3373_1, in3373_2, c3060);
    wire[0:0] s3374, in3374_1, in3374_2;
    wire c3374;
    assign in3374_1 = {c3061};
    assign in3374_2 = {c3062};
    Full_Adder FA_3374(s3374, c3374, in3374_1, in3374_2, s2664[0]);
    wire[0:0] s3375, in3375_1, in3375_2;
    wire c3375;
    assign in3375_1 = {s3064[0]};
    assign in3375_2 = {s3065[0]};
    Full_Adder FA_3375(s3375, c3375, in3375_1, in3375_2, c3063);
    wire[0:0] s3376, in3376_1, in3376_2;
    wire c3376;
    assign in3376_1 = {c3064};
    assign in3376_2 = {c3065};
    Full_Adder FA_3376(s3376, c3376, in3376_1, in3376_2, s2668[0]);
    wire[0:0] s3377, in3377_1, in3377_2;
    wire c3377;
    assign in3377_1 = {s3067[0]};
    assign in3377_2 = {s3068[0]};
    Full_Adder FA_3377(s3377, c3377, in3377_1, in3377_2, c3066);
    wire[0:0] s3378, in3378_1, in3378_2;
    wire c3378;
    assign in3378_1 = {c3067};
    assign in3378_2 = {c3068};
    Full_Adder FA_3378(s3378, c3378, in3378_1, in3378_2, s2672[0]);
    wire[0:0] s3379, in3379_1, in3379_2;
    wire c3379;
    assign in3379_1 = {s3070[0]};
    assign in3379_2 = {s3071[0]};
    Full_Adder FA_3379(s3379, c3379, in3379_1, in3379_2, c3069);
    wire[0:0] s3380, in3380_1, in3380_2;
    wire c3380;
    assign in3380_1 = {c3070};
    assign in3380_2 = {c3071};
    Full_Adder FA_3380(s3380, c3380, in3380_1, in3380_2, s2676[0]);
    wire[0:0] s3381, in3381_1, in3381_2;
    wire c3381;
    assign in3381_1 = {s3073[0]};
    assign in3381_2 = {s3074[0]};
    Full_Adder FA_3381(s3381, c3381, in3381_1, in3381_2, c3072);
    wire[0:0] s3382, in3382_1, in3382_2;
    wire c3382;
    assign in3382_1 = {c3073};
    assign in3382_2 = {c3074};
    Full_Adder FA_3382(s3382, c3382, in3382_1, in3382_2, s2680[0]);
    wire[0:0] s3383, in3383_1, in3383_2;
    wire c3383;
    assign in3383_1 = {s3076[0]};
    assign in3383_2 = {s3077[0]};
    Full_Adder FA_3383(s3383, c3383, in3383_1, in3383_2, c3075);
    wire[0:0] s3384, in3384_1, in3384_2;
    wire c3384;
    assign in3384_1 = {c3076};
    assign in3384_2 = {c3077};
    Full_Adder FA_3384(s3384, c3384, in3384_1, in3384_2, s2684[0]);
    wire[0:0] s3385, in3385_1, in3385_2;
    wire c3385;
    assign in3385_1 = {s3079[0]};
    assign in3385_2 = {s3080[0]};
    Full_Adder FA_3385(s3385, c3385, in3385_1, in3385_2, c3078);
    wire[0:0] s3386, in3386_1, in3386_2;
    wire c3386;
    assign in3386_1 = {c3079};
    assign in3386_2 = {c3080};
    Full_Adder FA_3386(s3386, c3386, in3386_1, in3386_2, s2688[0]);
    wire[0:0] s3387, in3387_1, in3387_2;
    wire c3387;
    assign in3387_1 = {s3082[0]};
    assign in3387_2 = {s3083[0]};
    Full_Adder FA_3387(s3387, c3387, in3387_1, in3387_2, c3081);
    wire[0:0] s3388, in3388_1, in3388_2;
    wire c3388;
    assign in3388_1 = {c3082};
    assign in3388_2 = {c3083};
    Full_Adder FA_3388(s3388, c3388, in3388_1, in3388_2, s2692[0]);
    wire[0:0] s3389, in3389_1, in3389_2;
    wire c3389;
    assign in3389_1 = {s3085[0]};
    assign in3389_2 = {s3086[0]};
    Full_Adder FA_3389(s3389, c3389, in3389_1, in3389_2, c3084);
    wire[0:0] s3390, in3390_1, in3390_2;
    wire c3390;
    assign in3390_1 = {c3085};
    assign in3390_2 = {c3086};
    Full_Adder FA_3390(s3390, c3390, in3390_1, in3390_2, s2696[0]);
    wire[0:0] s3391, in3391_1, in3391_2;
    wire c3391;
    assign in3391_1 = {s3088[0]};
    assign in3391_2 = {s3089[0]};
    Full_Adder FA_3391(s3391, c3391, in3391_1, in3391_2, c3087);
    wire[0:0] s3392, in3392_1, in3392_2;
    wire c3392;
    assign in3392_1 = {c3088};
    assign in3392_2 = {c3089};
    Full_Adder FA_3392(s3392, c3392, in3392_1, in3392_2, s2700[0]);
    wire[0:0] s3393, in3393_1, in3393_2;
    wire c3393;
    assign in3393_1 = {s3091[0]};
    assign in3393_2 = {s3092[0]};
    Full_Adder FA_3393(s3393, c3393, in3393_1, in3393_2, c3090);
    wire[0:0] s3394, in3394_1, in3394_2;
    wire c3394;
    assign in3394_1 = {c3091};
    assign in3394_2 = {c3092};
    Full_Adder FA_3394(s3394, c3394, in3394_1, in3394_2, s2704[0]);
    wire[0:0] s3395, in3395_1, in3395_2;
    wire c3395;
    assign in3395_1 = {s3094[0]};
    assign in3395_2 = {s3095[0]};
    Full_Adder FA_3395(s3395, c3395, in3395_1, in3395_2, c3093);
    wire[0:0] s3396, in3396_1, in3396_2;
    wire c3396;
    assign in3396_1 = {c3094};
    assign in3396_2 = {c3095};
    Full_Adder FA_3396(s3396, c3396, in3396_1, in3396_2, s2708[0]);
    wire[0:0] s3397, in3397_1, in3397_2;
    wire c3397;
    assign in3397_1 = {s3097[0]};
    assign in3397_2 = {s3098[0]};
    Full_Adder FA_3397(s3397, c3397, in3397_1, in3397_2, c3096);
    wire[0:0] s3398, in3398_1, in3398_2;
    wire c3398;
    assign in3398_1 = {c3097};
    assign in3398_2 = {c3098};
    Full_Adder FA_3398(s3398, c3398, in3398_1, in3398_2, s2712[0]);
    wire[0:0] s3399, in3399_1, in3399_2;
    wire c3399;
    assign in3399_1 = {s3100[0]};
    assign in3399_2 = {s3101[0]};
    Full_Adder FA_3399(s3399, c3399, in3399_1, in3399_2, c3099);
    wire[0:0] s3400, in3400_1, in3400_2;
    wire c3400;
    assign in3400_1 = {c3100};
    assign in3400_2 = {c3101};
    Full_Adder FA_3400(s3400, c3400, in3400_1, in3400_2, s2716[0]);
    wire[0:0] s3401, in3401_1, in3401_2;
    wire c3401;
    assign in3401_1 = {s3103[0]};
    assign in3401_2 = {s3104[0]};
    Full_Adder FA_3401(s3401, c3401, in3401_1, in3401_2, c3102);
    wire[0:0] s3402, in3402_1, in3402_2;
    wire c3402;
    assign in3402_1 = {c3103};
    assign in3402_2 = {c3104};
    Full_Adder FA_3402(s3402, c3402, in3402_1, in3402_2, s2720[0]);
    wire[0:0] s3403, in3403_1, in3403_2;
    wire c3403;
    assign in3403_1 = {s3106[0]};
    assign in3403_2 = {s3107[0]};
    Full_Adder FA_3403(s3403, c3403, in3403_1, in3403_2, c3105);
    wire[0:0] s3404, in3404_1, in3404_2;
    wire c3404;
    assign in3404_1 = {c3106};
    assign in3404_2 = {c3107};
    Full_Adder FA_3404(s3404, c3404, in3404_1, in3404_2, s2724[0]);
    wire[0:0] s3405, in3405_1, in3405_2;
    wire c3405;
    assign in3405_1 = {s3109[0]};
    assign in3405_2 = {s3110[0]};
    Full_Adder FA_3405(s3405, c3405, in3405_1, in3405_2, c3108);
    wire[0:0] s3406, in3406_1, in3406_2;
    wire c3406;
    assign in3406_1 = {c3109};
    assign in3406_2 = {c3110};
    Full_Adder FA_3406(s3406, c3406, in3406_1, in3406_2, s2728[0]);
    wire[0:0] s3407, in3407_1, in3407_2;
    wire c3407;
    assign in3407_1 = {s3112[0]};
    assign in3407_2 = {s3113[0]};
    Full_Adder FA_3407(s3407, c3407, in3407_1, in3407_2, c3111);
    wire[0:0] s3408, in3408_1, in3408_2;
    wire c3408;
    assign in3408_1 = {c3112};
    assign in3408_2 = {c3113};
    Full_Adder FA_3408(s3408, c3408, in3408_1, in3408_2, s2732[0]);
    wire[0:0] s3409, in3409_1, in3409_2;
    wire c3409;
    assign in3409_1 = {s3115[0]};
    assign in3409_2 = {s3116[0]};
    Full_Adder FA_3409(s3409, c3409, in3409_1, in3409_2, c3114);
    wire[0:0] s3410, in3410_1, in3410_2;
    wire c3410;
    assign in3410_1 = {c3115};
    assign in3410_2 = {c3116};
    Full_Adder FA_3410(s3410, c3410, in3410_1, in3410_2, s2736[0]);
    wire[0:0] s3411, in3411_1, in3411_2;
    wire c3411;
    assign in3411_1 = {s3118[0]};
    assign in3411_2 = {s3119[0]};
    Full_Adder FA_3411(s3411, c3411, in3411_1, in3411_2, c3117);
    wire[0:0] s3412, in3412_1, in3412_2;
    wire c3412;
    assign in3412_1 = {c3118};
    assign in3412_2 = {c3119};
    Full_Adder FA_3412(s3412, c3412, in3412_1, in3412_2, s2740[0]);
    wire[0:0] s3413, in3413_1, in3413_2;
    wire c3413;
    assign in3413_1 = {s3121[0]};
    assign in3413_2 = {s3122[0]};
    Full_Adder FA_3413(s3413, c3413, in3413_1, in3413_2, c3120);
    wire[0:0] s3414, in3414_1, in3414_2;
    wire c3414;
    assign in3414_1 = {c3121};
    assign in3414_2 = {c3122};
    Full_Adder FA_3414(s3414, c3414, in3414_1, in3414_2, s2744[0]);
    wire[0:0] s3415, in3415_1, in3415_2;
    wire c3415;
    assign in3415_1 = {s3124[0]};
    assign in3415_2 = {s3125[0]};
    Full_Adder FA_3415(s3415, c3415, in3415_1, in3415_2, c3123);
    wire[0:0] s3416, in3416_1, in3416_2;
    wire c3416;
    assign in3416_1 = {c3124};
    assign in3416_2 = {c3125};
    Full_Adder FA_3416(s3416, c3416, in3416_1, in3416_2, s2748[0]);
    wire[0:0] s3417, in3417_1, in3417_2;
    wire c3417;
    assign in3417_1 = {s3127[0]};
    assign in3417_2 = {s3128[0]};
    Full_Adder FA_3417(s3417, c3417, in3417_1, in3417_2, c3126);
    wire[0:0] s3418, in3418_1, in3418_2;
    wire c3418;
    assign in3418_1 = {c3127};
    assign in3418_2 = {c3128};
    Full_Adder FA_3418(s3418, c3418, in3418_1, in3418_2, s2752[0]);
    wire[0:0] s3419, in3419_1, in3419_2;
    wire c3419;
    assign in3419_1 = {s3130[0]};
    assign in3419_2 = {s3131[0]};
    Full_Adder FA_3419(s3419, c3419, in3419_1, in3419_2, c3129);
    wire[0:0] s3420, in3420_1, in3420_2;
    wire c3420;
    assign in3420_1 = {c3130};
    assign in3420_2 = {c3131};
    Full_Adder FA_3420(s3420, c3420, in3420_1, in3420_2, s2756[0]);
    wire[0:0] s3421, in3421_1, in3421_2;
    wire c3421;
    assign in3421_1 = {s3133[0]};
    assign in3421_2 = {s3134[0]};
    Full_Adder FA_3421(s3421, c3421, in3421_1, in3421_2, c3132);
    wire[0:0] s3422, in3422_1, in3422_2;
    wire c3422;
    assign in3422_1 = {c3133};
    assign in3422_2 = {c3134};
    Full_Adder FA_3422(s3422, c3422, in3422_1, in3422_2, s2760[0]);
    wire[0:0] s3423, in3423_1, in3423_2;
    wire c3423;
    assign in3423_1 = {s3136[0]};
    assign in3423_2 = {s3137[0]};
    Full_Adder FA_3423(s3423, c3423, in3423_1, in3423_2, c3135);
    wire[0:0] s3424, in3424_1, in3424_2;
    wire c3424;
    assign in3424_1 = {c3136};
    assign in3424_2 = {c3137};
    Full_Adder FA_3424(s3424, c3424, in3424_1, in3424_2, s2764[0]);
    wire[0:0] s3425, in3425_1, in3425_2;
    wire c3425;
    assign in3425_1 = {s3139[0]};
    assign in3425_2 = {s3140[0]};
    Full_Adder FA_3425(s3425, c3425, in3425_1, in3425_2, c3138);
    wire[0:0] s3426, in3426_1, in3426_2;
    wire c3426;
    assign in3426_1 = {c3139};
    assign in3426_2 = {c3140};
    Full_Adder FA_3426(s3426, c3426, in3426_1, in3426_2, s2768[0]);
    wire[0:0] s3427, in3427_1, in3427_2;
    wire c3427;
    assign in3427_1 = {s3142[0]};
    assign in3427_2 = {s3143[0]};
    Full_Adder FA_3427(s3427, c3427, in3427_1, in3427_2, c3141);
    wire[0:0] s3428, in3428_1, in3428_2;
    wire c3428;
    assign in3428_1 = {c3142};
    assign in3428_2 = {c3143};
    Full_Adder FA_3428(s3428, c3428, in3428_1, in3428_2, s2772[0]);
    wire[0:0] s3429, in3429_1, in3429_2;
    wire c3429;
    assign in3429_1 = {s3145[0]};
    assign in3429_2 = {s3146[0]};
    Full_Adder FA_3429(s3429, c3429, in3429_1, in3429_2, c3144);
    wire[0:0] s3430, in3430_1, in3430_2;
    wire c3430;
    assign in3430_1 = {c3145};
    assign in3430_2 = {c3146};
    Full_Adder FA_3430(s3430, c3430, in3430_1, in3430_2, s2776[0]);
    wire[0:0] s3431, in3431_1, in3431_2;
    wire c3431;
    assign in3431_1 = {s3148[0]};
    assign in3431_2 = {s3149[0]};
    Full_Adder FA_3431(s3431, c3431, in3431_1, in3431_2, c3147);
    wire[0:0] s3432, in3432_1, in3432_2;
    wire c3432;
    assign in3432_1 = {c3148};
    assign in3432_2 = {c3149};
    Full_Adder FA_3432(s3432, c3432, in3432_1, in3432_2, s2780[0]);
    wire[0:0] s3433, in3433_1, in3433_2;
    wire c3433;
    assign in3433_1 = {s3151[0]};
    assign in3433_2 = {s3152[0]};
    Full_Adder FA_3433(s3433, c3433, in3433_1, in3433_2, c3150);
    wire[0:0] s3434, in3434_1, in3434_2;
    wire c3434;
    assign in3434_1 = {c3151};
    assign in3434_2 = {c3152};
    Full_Adder FA_3434(s3434, c3434, in3434_1, in3434_2, s2784[0]);
    wire[0:0] s3435, in3435_1, in3435_2;
    wire c3435;
    assign in3435_1 = {s3154[0]};
    assign in3435_2 = {s3155[0]};
    Full_Adder FA_3435(s3435, c3435, in3435_1, in3435_2, c3153);
    wire[0:0] s3436, in3436_1, in3436_2;
    wire c3436;
    assign in3436_1 = {c3154};
    assign in3436_2 = {c3155};
    Full_Adder FA_3436(s3436, c3436, in3436_1, in3436_2, s2788[0]);
    wire[0:0] s3437, in3437_1, in3437_2;
    wire c3437;
    assign in3437_1 = {s3157[0]};
    assign in3437_2 = {s3158[0]};
    Full_Adder FA_3437(s3437, c3437, in3437_1, in3437_2, c3156);
    wire[0:0] s3438, in3438_1, in3438_2;
    wire c3438;
    assign in3438_1 = {c3157};
    assign in3438_2 = {c3158};
    Full_Adder FA_3438(s3438, c3438, in3438_1, in3438_2, s2792[0]);
    wire[0:0] s3439, in3439_1, in3439_2;
    wire c3439;
    assign in3439_1 = {s3160[0]};
    assign in3439_2 = {s3161[0]};
    Full_Adder FA_3439(s3439, c3439, in3439_1, in3439_2, c3159);
    wire[0:0] s3440, in3440_1, in3440_2;
    wire c3440;
    assign in3440_1 = {c3160};
    assign in3440_2 = {c3161};
    Full_Adder FA_3440(s3440, c3440, in3440_1, in3440_2, s2796[0]);
    wire[0:0] s3441, in3441_1, in3441_2;
    wire c3441;
    assign in3441_1 = {s3163[0]};
    assign in3441_2 = {s3164[0]};
    Full_Adder FA_3441(s3441, c3441, in3441_1, in3441_2, c3162);
    wire[0:0] s3442, in3442_1, in3442_2;
    wire c3442;
    assign in3442_1 = {c3163};
    assign in3442_2 = {c3164};
    Full_Adder FA_3442(s3442, c3442, in3442_1, in3442_2, s2800[0]);
    wire[0:0] s3443, in3443_1, in3443_2;
    wire c3443;
    assign in3443_1 = {s3166[0]};
    assign in3443_2 = {s3167[0]};
    Full_Adder FA_3443(s3443, c3443, in3443_1, in3443_2, c3165);
    wire[0:0] s3444, in3444_1, in3444_2;
    wire c3444;
    assign in3444_1 = {c3166};
    assign in3444_2 = {c3167};
    Full_Adder FA_3444(s3444, c3444, in3444_1, in3444_2, s2804[0]);
    wire[0:0] s3445, in3445_1, in3445_2;
    wire c3445;
    assign in3445_1 = {s3169[0]};
    assign in3445_2 = {s3170[0]};
    Full_Adder FA_3445(s3445, c3445, in3445_1, in3445_2, c3168);
    wire[0:0] s3446, in3446_1, in3446_2;
    wire c3446;
    assign in3446_1 = {c3169};
    assign in3446_2 = {c3170};
    Full_Adder FA_3446(s3446, c3446, in3446_1, in3446_2, s2808[0]);
    wire[0:0] s3447, in3447_1, in3447_2;
    wire c3447;
    assign in3447_1 = {s3172[0]};
    assign in3447_2 = {s3173[0]};
    Full_Adder FA_3447(s3447, c3447, in3447_1, in3447_2, c3171);
    wire[0:0] s3448, in3448_1, in3448_2;
    wire c3448;
    assign in3448_1 = {c3172};
    assign in3448_2 = {c3173};
    Full_Adder FA_3448(s3448, c3448, in3448_1, in3448_2, s2812[0]);
    wire[0:0] s3449, in3449_1, in3449_2;
    wire c3449;
    assign in3449_1 = {s3175[0]};
    assign in3449_2 = {s3176[0]};
    Full_Adder FA_3449(s3449, c3449, in3449_1, in3449_2, c3174);
    wire[0:0] s3450, in3450_1, in3450_2;
    wire c3450;
    assign in3450_1 = {c3175};
    assign in3450_2 = {c3176};
    Full_Adder FA_3450(s3450, c3450, in3450_1, in3450_2, s2816[0]);
    wire[0:0] s3451, in3451_1, in3451_2;
    wire c3451;
    assign in3451_1 = {s3178[0]};
    assign in3451_2 = {s3179[0]};
    Full_Adder FA_3451(s3451, c3451, in3451_1, in3451_2, c3177);
    wire[0:0] s3452, in3452_1, in3452_2;
    wire c3452;
    assign in3452_1 = {c3178};
    assign in3452_2 = {c3179};
    Full_Adder FA_3452(s3452, c3452, in3452_1, in3452_2, s2820[0]);
    wire[0:0] s3453, in3453_1, in3453_2;
    wire c3453;
    assign in3453_1 = {s3181[0]};
    assign in3453_2 = {s3182[0]};
    Full_Adder FA_3453(s3453, c3453, in3453_1, in3453_2, c3180);
    wire[0:0] s3454, in3454_1, in3454_2;
    wire c3454;
    assign in3454_1 = {c3181};
    assign in3454_2 = {c3182};
    Full_Adder FA_3454(s3454, c3454, in3454_1, in3454_2, s2824[0]);
    wire[0:0] s3455, in3455_1, in3455_2;
    wire c3455;
    assign in3455_1 = {s3184[0]};
    assign in3455_2 = {s3185[0]};
    Full_Adder FA_3455(s3455, c3455, in3455_1, in3455_2, c3183);
    wire[0:0] s3456, in3456_1, in3456_2;
    wire c3456;
    assign in3456_1 = {c3184};
    assign in3456_2 = {c3185};
    Full_Adder FA_3456(s3456, c3456, in3456_1, in3456_2, s2828[0]);
    wire[0:0] s3457, in3457_1, in3457_2;
    wire c3457;
    assign in3457_1 = {s3187[0]};
    assign in3457_2 = {s3188[0]};
    Full_Adder FA_3457(s3457, c3457, in3457_1, in3457_2, c3186);
    wire[0:0] s3458, in3458_1, in3458_2;
    wire c3458;
    assign in3458_1 = {c3187};
    assign in3458_2 = {c3188};
    Full_Adder FA_3458(s3458, c3458, in3458_1, in3458_2, s2832[0]);
    wire[0:0] s3459, in3459_1, in3459_2;
    wire c3459;
    assign in3459_1 = {s3190[0]};
    assign in3459_2 = {s3191[0]};
    Full_Adder FA_3459(s3459, c3459, in3459_1, in3459_2, c3189);
    wire[0:0] s3460, in3460_1, in3460_2;
    wire c3460;
    assign in3460_1 = {c3190};
    assign in3460_2 = {c3191};
    Full_Adder FA_3460(s3460, c3460, in3460_1, in3460_2, s2836[0]);
    wire[0:0] s3461, in3461_1, in3461_2;
    wire c3461;
    assign in3461_1 = {s3193[0]};
    assign in3461_2 = {s3194[0]};
    Full_Adder FA_3461(s3461, c3461, in3461_1, in3461_2, c3192);
    wire[0:0] s3462, in3462_1, in3462_2;
    wire c3462;
    assign in3462_1 = {c3193};
    assign in3462_2 = {c3194};
    Full_Adder FA_3462(s3462, c3462, in3462_1, in3462_2, s2840[0]);
    wire[0:0] s3463, in3463_1, in3463_2;
    wire c3463;
    assign in3463_1 = {s3196[0]};
    assign in3463_2 = {s3197[0]};
    Full_Adder FA_3463(s3463, c3463, in3463_1, in3463_2, c3195);
    wire[0:0] s3464, in3464_1, in3464_2;
    wire c3464;
    assign in3464_1 = {c3196};
    assign in3464_2 = {c3197};
    Full_Adder FA_3464(s3464, c3464, in3464_1, in3464_2, s2844[0]);
    wire[0:0] s3465, in3465_1, in3465_2;
    wire c3465;
    assign in3465_1 = {s3199[0]};
    assign in3465_2 = {s3200[0]};
    Full_Adder FA_3465(s3465, c3465, in3465_1, in3465_2, c3198);
    wire[0:0] s3466, in3466_1, in3466_2;
    wire c3466;
    assign in3466_1 = {c3199};
    assign in3466_2 = {c3200};
    Full_Adder FA_3466(s3466, c3466, in3466_1, in3466_2, s2848[0]);
    wire[0:0] s3467, in3467_1, in3467_2;
    wire c3467;
    assign in3467_1 = {s3202[0]};
    assign in3467_2 = {s3203[0]};
    Full_Adder FA_3467(s3467, c3467, in3467_1, in3467_2, c3201);
    wire[0:0] s3468, in3468_1, in3468_2;
    wire c3468;
    assign in3468_1 = {c3202};
    assign in3468_2 = {c3203};
    Full_Adder FA_3468(s3468, c3468, in3468_1, in3468_2, s2852[0]);
    wire[0:0] s3469, in3469_1, in3469_2;
    wire c3469;
    assign in3469_1 = {s3205[0]};
    assign in3469_2 = {s3206[0]};
    Full_Adder FA_3469(s3469, c3469, in3469_1, in3469_2, c3204);
    wire[0:0] s3470, in3470_1, in3470_2;
    wire c3470;
    assign in3470_1 = {c3205};
    assign in3470_2 = {c3206};
    Full_Adder FA_3470(s3470, c3470, in3470_1, in3470_2, s2856[0]);
    wire[0:0] s3471, in3471_1, in3471_2;
    wire c3471;
    assign in3471_1 = {s3208[0]};
    assign in3471_2 = {s3209[0]};
    Full_Adder FA_3471(s3471, c3471, in3471_1, in3471_2, c3207);
    wire[0:0] s3472, in3472_1, in3472_2;
    wire c3472;
    assign in3472_1 = {c3208};
    assign in3472_2 = {c3209};
    Full_Adder FA_3472(s3472, c3472, in3472_1, in3472_2, s2860[0]);
    wire[0:0] s3473, in3473_1, in3473_2;
    wire c3473;
    assign in3473_1 = {s3211[0]};
    assign in3473_2 = {s3212[0]};
    Full_Adder FA_3473(s3473, c3473, in3473_1, in3473_2, c3210);
    wire[0:0] s3474, in3474_1, in3474_2;
    wire c3474;
    assign in3474_1 = {c3211};
    assign in3474_2 = {c3212};
    Full_Adder FA_3474(s3474, c3474, in3474_1, in3474_2, s2864[0]);
    wire[0:0] s3475, in3475_1, in3475_2;
    wire c3475;
    assign in3475_1 = {s3214[0]};
    assign in3475_2 = {s3215[0]};
    Full_Adder FA_3475(s3475, c3475, in3475_1, in3475_2, c3213);
    wire[0:0] s3476, in3476_1, in3476_2;
    wire c3476;
    assign in3476_1 = {c3214};
    assign in3476_2 = {c3215};
    Full_Adder FA_3476(s3476, c3476, in3476_1, in3476_2, s2868[0]);
    wire[0:0] s3477, in3477_1, in3477_2;
    wire c3477;
    assign in3477_1 = {s3217[0]};
    assign in3477_2 = {s3218[0]};
    Full_Adder FA_3477(s3477, c3477, in3477_1, in3477_2, c3216);
    wire[0:0] s3478, in3478_1, in3478_2;
    wire c3478;
    assign in3478_1 = {c3217};
    assign in3478_2 = {c3218};
    Full_Adder FA_3478(s3478, c3478, in3478_1, in3478_2, s2872[0]);
    wire[0:0] s3479, in3479_1, in3479_2;
    wire c3479;
    assign in3479_1 = {s3220[0]};
    assign in3479_2 = {s3221[0]};
    Full_Adder FA_3479(s3479, c3479, in3479_1, in3479_2, c3219);
    wire[0:0] s3480, in3480_1, in3480_2;
    wire c3480;
    assign in3480_1 = {c3220};
    assign in3480_2 = {c3221};
    Full_Adder FA_3480(s3480, c3480, in3480_1, in3480_2, s2876[0]);
    wire[0:0] s3481, in3481_1, in3481_2;
    wire c3481;
    assign in3481_1 = {s3223[0]};
    assign in3481_2 = {s3224[0]};
    Full_Adder FA_3481(s3481, c3481, in3481_1, in3481_2, c3222);
    wire[0:0] s3482, in3482_1, in3482_2;
    wire c3482;
    assign in3482_1 = {c3223};
    assign in3482_2 = {c3224};
    Full_Adder FA_3482(s3482, c3482, in3482_1, in3482_2, s2880[0]);
    wire[0:0] s3483, in3483_1, in3483_2;
    wire c3483;
    assign in3483_1 = {s3226[0]};
    assign in3483_2 = {s3227[0]};
    Full_Adder FA_3483(s3483, c3483, in3483_1, in3483_2, c3225);
    wire[0:0] s3484, in3484_1, in3484_2;
    wire c3484;
    assign in3484_1 = {c3226};
    assign in3484_2 = {c3227};
    Full_Adder FA_3484(s3484, c3484, in3484_1, in3484_2, s2884[0]);
    wire[0:0] s3485, in3485_1, in3485_2;
    wire c3485;
    assign in3485_1 = {s3229[0]};
    assign in3485_2 = {s3230[0]};
    Full_Adder FA_3485(s3485, c3485, in3485_1, in3485_2, c3228);
    wire[0:0] s3486, in3486_1, in3486_2;
    wire c3486;
    assign in3486_1 = {c3229};
    assign in3486_2 = {c3230};
    Full_Adder FA_3486(s3486, c3486, in3486_1, in3486_2, s2888[0]);
    wire[0:0] s3487, in3487_1, in3487_2;
    wire c3487;
    assign in3487_1 = {s3232[0]};
    assign in3487_2 = {s3233[0]};
    Full_Adder FA_3487(s3487, c3487, in3487_1, in3487_2, c3231);
    wire[0:0] s3488, in3488_1, in3488_2;
    wire c3488;
    assign in3488_1 = {c3232};
    assign in3488_2 = {c3233};
    Full_Adder FA_3488(s3488, c3488, in3488_1, in3488_2, s2892[0]);
    wire[0:0] s3489, in3489_1, in3489_2;
    wire c3489;
    assign in3489_1 = {s3235[0]};
    assign in3489_2 = {s3236[0]};
    Full_Adder FA_3489(s3489, c3489, in3489_1, in3489_2, c3234);
    wire[0:0] s3490, in3490_1, in3490_2;
    wire c3490;
    assign in3490_1 = {c3235};
    assign in3490_2 = {c3236};
    Full_Adder FA_3490(s3490, c3490, in3490_1, in3490_2, s2896[0]);
    wire[0:0] s3491, in3491_1, in3491_2;
    wire c3491;
    assign in3491_1 = {s3238[0]};
    assign in3491_2 = {s3239[0]};
    Full_Adder FA_3491(s3491, c3491, in3491_1, in3491_2, c3237);
    wire[0:0] s3492, in3492_1, in3492_2;
    wire c3492;
    assign in3492_1 = {c3238};
    assign in3492_2 = {c3239};
    Full_Adder FA_3492(s3492, c3492, in3492_1, in3492_2, s2900[0]);
    wire[0:0] s3493, in3493_1, in3493_2;
    wire c3493;
    assign in3493_1 = {s3241[0]};
    assign in3493_2 = {s3242[0]};
    Full_Adder FA_3493(s3493, c3493, in3493_1, in3493_2, c3240);
    wire[0:0] s3494, in3494_1, in3494_2;
    wire c3494;
    assign in3494_1 = {c3241};
    assign in3494_2 = {c3242};
    Full_Adder FA_3494(s3494, c3494, in3494_1, in3494_2, s2904[0]);
    wire[0:0] s3495, in3495_1, in3495_2;
    wire c3495;
    assign in3495_1 = {s3244[0]};
    assign in3495_2 = {s3245[0]};
    Full_Adder FA_3495(s3495, c3495, in3495_1, in3495_2, c3243);
    wire[0:0] s3496, in3496_1, in3496_2;
    wire c3496;
    assign in3496_1 = {c3244};
    assign in3496_2 = {c3245};
    Full_Adder FA_3496(s3496, c3496, in3496_1, in3496_2, s2908[0]);
    wire[0:0] s3497, in3497_1, in3497_2;
    wire c3497;
    assign in3497_1 = {s3247[0]};
    assign in3497_2 = {s3248[0]};
    Full_Adder FA_3497(s3497, c3497, in3497_1, in3497_2, c3246);
    wire[0:0] s3498, in3498_1, in3498_2;
    wire c3498;
    assign in3498_1 = {c3247};
    assign in3498_2 = {c3248};
    Full_Adder FA_3498(s3498, c3498, in3498_1, in3498_2, s2912[0]);
    wire[0:0] s3499, in3499_1, in3499_2;
    wire c3499;
    assign in3499_1 = {s3250[0]};
    assign in3499_2 = {s3251[0]};
    Full_Adder FA_3499(s3499, c3499, in3499_1, in3499_2, c3249);
    wire[0:0] s3500, in3500_1, in3500_2;
    wire c3500;
    assign in3500_1 = {c3250};
    assign in3500_2 = {c3251};
    Full_Adder FA_3500(s3500, c3500, in3500_1, in3500_2, s2916[0]);
    wire[0:0] s3501, in3501_1, in3501_2;
    wire c3501;
    assign in3501_1 = {s3253[0]};
    assign in3501_2 = {s3254[0]};
    Full_Adder FA_3501(s3501, c3501, in3501_1, in3501_2, c3252);
    wire[0:0] s3502, in3502_1, in3502_2;
    wire c3502;
    assign in3502_1 = {c3253};
    assign in3502_2 = {c3254};
    Full_Adder FA_3502(s3502, c3502, in3502_1, in3502_2, s2920[0]);
    wire[0:0] s3503, in3503_1, in3503_2;
    wire c3503;
    assign in3503_1 = {s3256[0]};
    assign in3503_2 = {s3257[0]};
    Full_Adder FA_3503(s3503, c3503, in3503_1, in3503_2, c3255);
    wire[0:0] s3504, in3504_1, in3504_2;
    wire c3504;
    assign in3504_1 = {c3256};
    assign in3504_2 = {c3257};
    Full_Adder FA_3504(s3504, c3504, in3504_1, in3504_2, s2924[0]);
    wire[0:0] s3505, in3505_1, in3505_2;
    wire c3505;
    assign in3505_1 = {s3259[0]};
    assign in3505_2 = {s3260[0]};
    Full_Adder FA_3505(s3505, c3505, in3505_1, in3505_2, c3258);
    wire[0:0] s3506, in3506_1, in3506_2;
    wire c3506;
    assign in3506_1 = {c3259};
    assign in3506_2 = {c3260};
    Full_Adder FA_3506(s3506, c3506, in3506_1, in3506_2, s2928[0]);
    wire[0:0] s3507, in3507_1, in3507_2;
    wire c3507;
    assign in3507_1 = {s3262[0]};
    assign in3507_2 = {s3263[0]};
    Full_Adder FA_3507(s3507, c3507, in3507_1, in3507_2, c3261);
    wire[0:0] s3508, in3508_1, in3508_2;
    wire c3508;
    assign in3508_1 = {c3262};
    assign in3508_2 = {c3263};
    Full_Adder FA_3508(s3508, c3508, in3508_1, in3508_2, s2932[0]);
    wire[0:0] s3509, in3509_1, in3509_2;
    wire c3509;
    assign in3509_1 = {s3265[0]};
    assign in3509_2 = {s3266[0]};
    Full_Adder FA_3509(s3509, c3509, in3509_1, in3509_2, c3264);
    wire[0:0] s3510, in3510_1, in3510_2;
    wire c3510;
    assign in3510_1 = {c3265};
    assign in3510_2 = {c3266};
    Full_Adder FA_3510(s3510, c3510, in3510_1, in3510_2, s2936[0]);
    wire[0:0] s3511, in3511_1, in3511_2;
    wire c3511;
    assign in3511_1 = {s3268[0]};
    assign in3511_2 = {s3269[0]};
    Full_Adder FA_3511(s3511, c3511, in3511_1, in3511_2, c3267);
    wire[0:0] s3512, in3512_1, in3512_2;
    wire c3512;
    assign in3512_1 = {c3268};
    assign in3512_2 = {c3269};
    Full_Adder FA_3512(s3512, c3512, in3512_1, in3512_2, s2940[0]);
    wire[0:0] s3513, in3513_1, in3513_2;
    wire c3513;
    assign in3513_1 = {s3271[0]};
    assign in3513_2 = {s3272[0]};
    Full_Adder FA_3513(s3513, c3513, in3513_1, in3513_2, c3270);
    wire[0:0] s3514, in3514_1, in3514_2;
    wire c3514;
    assign in3514_1 = {c3271};
    assign in3514_2 = {c3272};
    Full_Adder FA_3514(s3514, c3514, in3514_1, in3514_2, s2944[0]);
    wire[0:0] s3515, in3515_1, in3515_2;
    wire c3515;
    assign in3515_1 = {s3274[0]};
    assign in3515_2 = {s3275[0]};
    Full_Adder FA_3515(s3515, c3515, in3515_1, in3515_2, c3273);
    wire[0:0] s3516, in3516_1, in3516_2;
    wire c3516;
    assign in3516_1 = {c3274};
    assign in3516_2 = {c3275};
    Full_Adder FA_3516(s3516, c3516, in3516_1, in3516_2, s2948[0]);
    wire[0:0] s3517, in3517_1, in3517_2;
    wire c3517;
    assign in3517_1 = {s3277[0]};
    assign in3517_2 = {s3278[0]};
    Full_Adder FA_3517(s3517, c3517, in3517_1, in3517_2, c3276);
    wire[0:0] s3518, in3518_1, in3518_2;
    wire c3518;
    assign in3518_1 = {c3277};
    assign in3518_2 = {c3278};
    Full_Adder FA_3518(s3518, c3518, in3518_1, in3518_2, s2952[0]);
    wire[0:0] s3519, in3519_1, in3519_2;
    wire c3519;
    assign in3519_1 = {s3280[0]};
    assign in3519_2 = {s3281[0]};
    Full_Adder FA_3519(s3519, c3519, in3519_1, in3519_2, c3279);
    wire[0:0] s3520, in3520_1, in3520_2;
    wire c3520;
    assign in3520_1 = {c3280};
    assign in3520_2 = {c3281};
    Full_Adder FA_3520(s3520, c3520, in3520_1, in3520_2, s2956[0]);
    wire[0:0] s3521, in3521_1, in3521_2;
    wire c3521;
    assign in3521_1 = {s3283[0]};
    assign in3521_2 = {s3284[0]};
    Full_Adder FA_3521(s3521, c3521, in3521_1, in3521_2, c3282);
    wire[0:0] s3522, in3522_1, in3522_2;
    wire c3522;
    assign in3522_1 = {c3283};
    assign in3522_2 = {c3284};
    Full_Adder FA_3522(s3522, c3522, in3522_1, in3522_2, s2960[0]);
    wire[0:0] s3523, in3523_1, in3523_2;
    wire c3523;
    assign in3523_1 = {s3286[0]};
    assign in3523_2 = {s3287[0]};
    Full_Adder FA_3523(s3523, c3523, in3523_1, in3523_2, c3285);
    wire[0:0] s3524, in3524_1, in3524_2;
    wire c3524;
    assign in3524_1 = {c3286};
    assign in3524_2 = {c3287};
    Full_Adder FA_3524(s3524, c3524, in3524_1, in3524_2, s2964[0]);
    wire[0:0] s3525, in3525_1, in3525_2;
    wire c3525;
    assign in3525_1 = {s3289[0]};
    assign in3525_2 = {s3290[0]};
    Full_Adder FA_3525(s3525, c3525, in3525_1, in3525_2, c3288);
    wire[0:0] s3526, in3526_1, in3526_2;
    wire c3526;
    assign in3526_1 = {c3289};
    assign in3526_2 = {c3290};
    Full_Adder FA_3526(s3526, c3526, in3526_1, in3526_2, s2967[0]);
    wire[0:0] s3527, in3527_1, in3527_2;
    wire c3527;
    assign in3527_1 = {s3292[0]};
    assign in3527_2 = {s3293[0]};
    Full_Adder FA_3527(s3527, c3527, in3527_1, in3527_2, c3291);
    wire[0:0] s3528, in3528_1, in3528_2;
    wire c3528;
    assign in3528_1 = {c3292};
    assign in3528_2 = {c3293};
    Full_Adder FA_3528(s3528, c3528, in3528_1, in3528_2, s2969[0]);
    wire[0:0] s3529, in3529_1, in3529_2;
    wire c3529;
    assign in3529_1 = {s3295[0]};
    assign in3529_2 = {s3296[0]};
    Full_Adder FA_3529(s3529, c3529, in3529_1, in3529_2, c3294);
    wire[0:0] s3530, in3530_1, in3530_2;
    wire c3530;
    assign in3530_1 = {c3295};
    assign in3530_2 = {c3296};
    Full_Adder FA_3530(s3530, c3530, in3530_1, in3530_2, s2970[0]);
    wire[0:0] s3531, in3531_1, in3531_2;
    wire c3531;
    assign in3531_1 = {s3298[0]};
    assign in3531_2 = {s3299[0]};
    Full_Adder FA_3531(s3531, c3531, in3531_1, in3531_2, c3297);
    wire[0:0] s3532, in3532_1, in3532_2;
    wire c3532;
    assign in3532_1 = {c3298};
    assign in3532_2 = {c3299};
    Full_Adder FA_3532(s3532, c3532, in3532_1, in3532_2, c2970);
    wire[0:0] s3533, in3533_1, in3533_2;
    wire c3533;
    assign in3533_1 = {s3301[0]};
    assign in3533_2 = {s3302[0]};
    Full_Adder FA_3533(s3533, c3533, in3533_1, in3533_2, c3300);
    wire[0:0] s3534, in3534_1, in3534_2;
    wire c3534;
    assign in3534_1 = {pp63[56]};
    assign in3534_2 = {c3301};
    Full_Adder FA_3534(s3534, c3534, in3534_1, in3534_2, pp62[57]);
    wire[0:0] s3535, in3535_1, in3535_2;
    wire c3535;
    assign in3535_1 = {c3303};
    assign in3535_2 = {s3304[0]};
    Full_Adder FA_3535(s3535, c3535, in3535_1, in3535_2, c3302);
    wire[0:0] s3536, in3536_1, in3536_2;
    wire c3536;
    assign in3536_1 = {pp61[59]};
    assign in3536_2 = {pp62[58]};
    Full_Adder FA_3536(s3536, c3536, in3536_1, in3536_2, pp60[60]);
    wire[0:0] s3537, in3537_1, in3537_2;
    wire c3537;
    assign in3537_1 = {c3304};
    assign in3537_2 = {c3305};
    Full_Adder FA_3537(s3537, c3537, in3537_1, in3537_2, pp63[57]);
    wire[0:0] s3538, in3538_1, in3538_2;
    wire c3538;
    assign in3538_1 = {pp59[62]};
    assign in3538_2 = {pp60[61]};
    Full_Adder FA_3538(s3538, c3538, in3538_1, in3538_2, pp58[63]);
    wire[0:0] s3539, in3539_1, in3539_2;
    wire c3539;
    assign in3539_1 = {pp62[59]};
    assign in3539_2 = {pp63[58]};
    Full_Adder FA_3539(s3539, c3539, in3539_1, in3539_2, pp61[60]);
    wire[0:0] s3540, in3540_1, in3540_2;
    wire c3540;
    assign in3540_1 = {pp60[62]};
    assign in3540_2 = {pp61[61]};
    Full_Adder FA_3540(s3540, c3540, in3540_1, in3540_2, pp59[63]);

    /*Stage 8*/
    wire[0:0] s3541, in3541_1, in3541_2;
    wire c3541;
    assign in3541_1 = {pp0[4]};
    assign in3541_2 = {pp1[3]};
    Half_Adder HA_3541(s3541, c3541, in3541_1, in3541_2);
    wire[0:0] s3542, in3542_1, in3542_2;
    wire c3542;
    assign in3542_1 = {pp3[2]};
    assign in3542_2 = {pp4[1]};
    Full_Adder FA_3542(s3542, c3542, in3542_1, in3542_2, pp2[3]);
    wire[0:0] s3543, in3543_1, in3543_2;
    wire c3543;
    assign in3543_1 = {pp6[0]};
    assign in3543_2 = {c3307};
    Full_Adder FA_3543(s3543, c3543, in3543_1, in3543_2, pp5[1]);
    wire[0:0] s3544, in3544_1, in3544_2;
    wire c3544;
    assign in3544_1 = {c3308};
    assign in3544_2 = {c3309};
    Full_Adder FA_3544(s3544, c3544, in3544_1, in3544_2, s2971[0]);
    wire[0:0] s3545, in3545_1, in3545_2;
    wire c3545;
    assign in3545_1 = {c3310};
    assign in3545_2 = {c3311};
    Full_Adder FA_3545(s3545, c3545, in3545_1, in3545_2, s2973[0]);
    wire[0:0] s3546, in3546_1, in3546_2;
    wire c3546;
    assign in3546_1 = {c3312};
    assign in3546_2 = {c3313};
    Full_Adder FA_3546(s3546, c3546, in3546_1, in3546_2, s2976[0]);
    wire[0:0] s3547, in3547_1, in3547_2;
    wire c3547;
    assign in3547_1 = {c3314};
    assign in3547_2 = {c3315};
    Full_Adder FA_3547(s3547, c3547, in3547_1, in3547_2, s2979[0]);
    wire[0:0] s3548, in3548_1, in3548_2;
    wire c3548;
    assign in3548_1 = {c3316};
    assign in3548_2 = {c3317};
    Full_Adder FA_3548(s3548, c3548, in3548_1, in3548_2, s2982[0]);
    wire[0:0] s3549, in3549_1, in3549_2;
    wire c3549;
    assign in3549_1 = {c3318};
    assign in3549_2 = {c3319};
    Full_Adder FA_3549(s3549, c3549, in3549_1, in3549_2, s2985[0]);
    wire[0:0] s3550, in3550_1, in3550_2;
    wire c3550;
    assign in3550_1 = {c3320};
    assign in3550_2 = {c3321};
    Full_Adder FA_3550(s3550, c3550, in3550_1, in3550_2, s2988[0]);
    wire[0:0] s3551, in3551_1, in3551_2;
    wire c3551;
    assign in3551_1 = {c3322};
    assign in3551_2 = {c3323};
    Full_Adder FA_3551(s3551, c3551, in3551_1, in3551_2, s2991[0]);
    wire[0:0] s3552, in3552_1, in3552_2;
    wire c3552;
    assign in3552_1 = {c3324};
    assign in3552_2 = {c3325};
    Full_Adder FA_3552(s3552, c3552, in3552_1, in3552_2, s2994[0]);
    wire[0:0] s3553, in3553_1, in3553_2;
    wire c3553;
    assign in3553_1 = {c3326};
    assign in3553_2 = {c3327};
    Full_Adder FA_3553(s3553, c3553, in3553_1, in3553_2, s2997[0]);
    wire[0:0] s3554, in3554_1, in3554_2;
    wire c3554;
    assign in3554_1 = {c3328};
    assign in3554_2 = {c3329};
    Full_Adder FA_3554(s3554, c3554, in3554_1, in3554_2, s3000[0]);
    wire[0:0] s3555, in3555_1, in3555_2;
    wire c3555;
    assign in3555_1 = {c3330};
    assign in3555_2 = {c3331};
    Full_Adder FA_3555(s3555, c3555, in3555_1, in3555_2, s3003[0]);
    wire[0:0] s3556, in3556_1, in3556_2;
    wire c3556;
    assign in3556_1 = {c3332};
    assign in3556_2 = {c3333};
    Full_Adder FA_3556(s3556, c3556, in3556_1, in3556_2, s3006[0]);
    wire[0:0] s3557, in3557_1, in3557_2;
    wire c3557;
    assign in3557_1 = {c3334};
    assign in3557_2 = {c3335};
    Full_Adder FA_3557(s3557, c3557, in3557_1, in3557_2, s3009[0]);
    wire[0:0] s3558, in3558_1, in3558_2;
    wire c3558;
    assign in3558_1 = {c3336};
    assign in3558_2 = {c3337};
    Full_Adder FA_3558(s3558, c3558, in3558_1, in3558_2, s3012[0]);
    wire[0:0] s3559, in3559_1, in3559_2;
    wire c3559;
    assign in3559_1 = {c3338};
    assign in3559_2 = {c3339};
    Full_Adder FA_3559(s3559, c3559, in3559_1, in3559_2, s3015[0]);
    wire[0:0] s3560, in3560_1, in3560_2;
    wire c3560;
    assign in3560_1 = {c3340};
    assign in3560_2 = {c3341};
    Full_Adder FA_3560(s3560, c3560, in3560_1, in3560_2, s3018[0]);
    wire[0:0] s3561, in3561_1, in3561_2;
    wire c3561;
    assign in3561_1 = {c3342};
    assign in3561_2 = {c3343};
    Full_Adder FA_3561(s3561, c3561, in3561_1, in3561_2, s3021[0]);
    wire[0:0] s3562, in3562_1, in3562_2;
    wire c3562;
    assign in3562_1 = {c3344};
    assign in3562_2 = {c3345};
    Full_Adder FA_3562(s3562, c3562, in3562_1, in3562_2, s3024[0]);
    wire[0:0] s3563, in3563_1, in3563_2;
    wire c3563;
    assign in3563_1 = {c3346};
    assign in3563_2 = {c3347};
    Full_Adder FA_3563(s3563, c3563, in3563_1, in3563_2, s3027[0]);
    wire[0:0] s3564, in3564_1, in3564_2;
    wire c3564;
    assign in3564_1 = {c3348};
    assign in3564_2 = {c3349};
    Full_Adder FA_3564(s3564, c3564, in3564_1, in3564_2, s3030[0]);
    wire[0:0] s3565, in3565_1, in3565_2;
    wire c3565;
    assign in3565_1 = {c3350};
    assign in3565_2 = {c3351};
    Full_Adder FA_3565(s3565, c3565, in3565_1, in3565_2, s3033[0]);
    wire[0:0] s3566, in3566_1, in3566_2;
    wire c3566;
    assign in3566_1 = {c3352};
    assign in3566_2 = {c3353};
    Full_Adder FA_3566(s3566, c3566, in3566_1, in3566_2, s3036[0]);
    wire[0:0] s3567, in3567_1, in3567_2;
    wire c3567;
    assign in3567_1 = {c3354};
    assign in3567_2 = {c3355};
    Full_Adder FA_3567(s3567, c3567, in3567_1, in3567_2, s3039[0]);
    wire[0:0] s3568, in3568_1, in3568_2;
    wire c3568;
    assign in3568_1 = {c3356};
    assign in3568_2 = {c3357};
    Full_Adder FA_3568(s3568, c3568, in3568_1, in3568_2, s3042[0]);
    wire[0:0] s3569, in3569_1, in3569_2;
    wire c3569;
    assign in3569_1 = {c3358};
    assign in3569_2 = {c3359};
    Full_Adder FA_3569(s3569, c3569, in3569_1, in3569_2, s3045[0]);
    wire[0:0] s3570, in3570_1, in3570_2;
    wire c3570;
    assign in3570_1 = {c3360};
    assign in3570_2 = {c3361};
    Full_Adder FA_3570(s3570, c3570, in3570_1, in3570_2, s3048[0]);
    wire[0:0] s3571, in3571_1, in3571_2;
    wire c3571;
    assign in3571_1 = {c3362};
    assign in3571_2 = {c3363};
    Full_Adder FA_3571(s3571, c3571, in3571_1, in3571_2, s3051[0]);
    wire[0:0] s3572, in3572_1, in3572_2;
    wire c3572;
    assign in3572_1 = {c3364};
    assign in3572_2 = {c3365};
    Full_Adder FA_3572(s3572, c3572, in3572_1, in3572_2, s3054[0]);
    wire[0:0] s3573, in3573_1, in3573_2;
    wire c3573;
    assign in3573_1 = {c3366};
    assign in3573_2 = {c3367};
    Full_Adder FA_3573(s3573, c3573, in3573_1, in3573_2, s3057[0]);
    wire[0:0] s3574, in3574_1, in3574_2;
    wire c3574;
    assign in3574_1 = {c3368};
    assign in3574_2 = {c3369};
    Full_Adder FA_3574(s3574, c3574, in3574_1, in3574_2, s3060[0]);
    wire[0:0] s3575, in3575_1, in3575_2;
    wire c3575;
    assign in3575_1 = {c3370};
    assign in3575_2 = {c3371};
    Full_Adder FA_3575(s3575, c3575, in3575_1, in3575_2, s3063[0]);
    wire[0:0] s3576, in3576_1, in3576_2;
    wire c3576;
    assign in3576_1 = {c3372};
    assign in3576_2 = {c3373};
    Full_Adder FA_3576(s3576, c3576, in3576_1, in3576_2, s3066[0]);
    wire[0:0] s3577, in3577_1, in3577_2;
    wire c3577;
    assign in3577_1 = {c3374};
    assign in3577_2 = {c3375};
    Full_Adder FA_3577(s3577, c3577, in3577_1, in3577_2, s3069[0]);
    wire[0:0] s3578, in3578_1, in3578_2;
    wire c3578;
    assign in3578_1 = {c3376};
    assign in3578_2 = {c3377};
    Full_Adder FA_3578(s3578, c3578, in3578_1, in3578_2, s3072[0]);
    wire[0:0] s3579, in3579_1, in3579_2;
    wire c3579;
    assign in3579_1 = {c3378};
    assign in3579_2 = {c3379};
    Full_Adder FA_3579(s3579, c3579, in3579_1, in3579_2, s3075[0]);
    wire[0:0] s3580, in3580_1, in3580_2;
    wire c3580;
    assign in3580_1 = {c3380};
    assign in3580_2 = {c3381};
    Full_Adder FA_3580(s3580, c3580, in3580_1, in3580_2, s3078[0]);
    wire[0:0] s3581, in3581_1, in3581_2;
    wire c3581;
    assign in3581_1 = {c3382};
    assign in3581_2 = {c3383};
    Full_Adder FA_3581(s3581, c3581, in3581_1, in3581_2, s3081[0]);
    wire[0:0] s3582, in3582_1, in3582_2;
    wire c3582;
    assign in3582_1 = {c3384};
    assign in3582_2 = {c3385};
    Full_Adder FA_3582(s3582, c3582, in3582_1, in3582_2, s3084[0]);
    wire[0:0] s3583, in3583_1, in3583_2;
    wire c3583;
    assign in3583_1 = {c3386};
    assign in3583_2 = {c3387};
    Full_Adder FA_3583(s3583, c3583, in3583_1, in3583_2, s3087[0]);
    wire[0:0] s3584, in3584_1, in3584_2;
    wire c3584;
    assign in3584_1 = {c3388};
    assign in3584_2 = {c3389};
    Full_Adder FA_3584(s3584, c3584, in3584_1, in3584_2, s3090[0]);
    wire[0:0] s3585, in3585_1, in3585_2;
    wire c3585;
    assign in3585_1 = {c3390};
    assign in3585_2 = {c3391};
    Full_Adder FA_3585(s3585, c3585, in3585_1, in3585_2, s3093[0]);
    wire[0:0] s3586, in3586_1, in3586_2;
    wire c3586;
    assign in3586_1 = {c3392};
    assign in3586_2 = {c3393};
    Full_Adder FA_3586(s3586, c3586, in3586_1, in3586_2, s3096[0]);
    wire[0:0] s3587, in3587_1, in3587_2;
    wire c3587;
    assign in3587_1 = {c3394};
    assign in3587_2 = {c3395};
    Full_Adder FA_3587(s3587, c3587, in3587_1, in3587_2, s3099[0]);
    wire[0:0] s3588, in3588_1, in3588_2;
    wire c3588;
    assign in3588_1 = {c3396};
    assign in3588_2 = {c3397};
    Full_Adder FA_3588(s3588, c3588, in3588_1, in3588_2, s3102[0]);
    wire[0:0] s3589, in3589_1, in3589_2;
    wire c3589;
    assign in3589_1 = {c3398};
    assign in3589_2 = {c3399};
    Full_Adder FA_3589(s3589, c3589, in3589_1, in3589_2, s3105[0]);
    wire[0:0] s3590, in3590_1, in3590_2;
    wire c3590;
    assign in3590_1 = {c3400};
    assign in3590_2 = {c3401};
    Full_Adder FA_3590(s3590, c3590, in3590_1, in3590_2, s3108[0]);
    wire[0:0] s3591, in3591_1, in3591_2;
    wire c3591;
    assign in3591_1 = {c3402};
    assign in3591_2 = {c3403};
    Full_Adder FA_3591(s3591, c3591, in3591_1, in3591_2, s3111[0]);
    wire[0:0] s3592, in3592_1, in3592_2;
    wire c3592;
    assign in3592_1 = {c3404};
    assign in3592_2 = {c3405};
    Full_Adder FA_3592(s3592, c3592, in3592_1, in3592_2, s3114[0]);
    wire[0:0] s3593, in3593_1, in3593_2;
    wire c3593;
    assign in3593_1 = {c3406};
    assign in3593_2 = {c3407};
    Full_Adder FA_3593(s3593, c3593, in3593_1, in3593_2, s3117[0]);
    wire[0:0] s3594, in3594_1, in3594_2;
    wire c3594;
    assign in3594_1 = {c3408};
    assign in3594_2 = {c3409};
    Full_Adder FA_3594(s3594, c3594, in3594_1, in3594_2, s3120[0]);
    wire[0:0] s3595, in3595_1, in3595_2;
    wire c3595;
    assign in3595_1 = {c3410};
    assign in3595_2 = {c3411};
    Full_Adder FA_3595(s3595, c3595, in3595_1, in3595_2, s3123[0]);
    wire[0:0] s3596, in3596_1, in3596_2;
    wire c3596;
    assign in3596_1 = {c3412};
    assign in3596_2 = {c3413};
    Full_Adder FA_3596(s3596, c3596, in3596_1, in3596_2, s3126[0]);
    wire[0:0] s3597, in3597_1, in3597_2;
    wire c3597;
    assign in3597_1 = {c3414};
    assign in3597_2 = {c3415};
    Full_Adder FA_3597(s3597, c3597, in3597_1, in3597_2, s3129[0]);
    wire[0:0] s3598, in3598_1, in3598_2;
    wire c3598;
    assign in3598_1 = {c3416};
    assign in3598_2 = {c3417};
    Full_Adder FA_3598(s3598, c3598, in3598_1, in3598_2, s3132[0]);
    wire[0:0] s3599, in3599_1, in3599_2;
    wire c3599;
    assign in3599_1 = {c3418};
    assign in3599_2 = {c3419};
    Full_Adder FA_3599(s3599, c3599, in3599_1, in3599_2, s3135[0]);
    wire[0:0] s3600, in3600_1, in3600_2;
    wire c3600;
    assign in3600_1 = {c3420};
    assign in3600_2 = {c3421};
    Full_Adder FA_3600(s3600, c3600, in3600_1, in3600_2, s3138[0]);
    wire[0:0] s3601, in3601_1, in3601_2;
    wire c3601;
    assign in3601_1 = {c3422};
    assign in3601_2 = {c3423};
    Full_Adder FA_3601(s3601, c3601, in3601_1, in3601_2, s3141[0]);
    wire[0:0] s3602, in3602_1, in3602_2;
    wire c3602;
    assign in3602_1 = {c3424};
    assign in3602_2 = {c3425};
    Full_Adder FA_3602(s3602, c3602, in3602_1, in3602_2, s3144[0]);
    wire[0:0] s3603, in3603_1, in3603_2;
    wire c3603;
    assign in3603_1 = {c3426};
    assign in3603_2 = {c3427};
    Full_Adder FA_3603(s3603, c3603, in3603_1, in3603_2, s3147[0]);
    wire[0:0] s3604, in3604_1, in3604_2;
    wire c3604;
    assign in3604_1 = {c3428};
    assign in3604_2 = {c3429};
    Full_Adder FA_3604(s3604, c3604, in3604_1, in3604_2, s3150[0]);
    wire[0:0] s3605, in3605_1, in3605_2;
    wire c3605;
    assign in3605_1 = {c3430};
    assign in3605_2 = {c3431};
    Full_Adder FA_3605(s3605, c3605, in3605_1, in3605_2, s3153[0]);
    wire[0:0] s3606, in3606_1, in3606_2;
    wire c3606;
    assign in3606_1 = {c3432};
    assign in3606_2 = {c3433};
    Full_Adder FA_3606(s3606, c3606, in3606_1, in3606_2, s3156[0]);
    wire[0:0] s3607, in3607_1, in3607_2;
    wire c3607;
    assign in3607_1 = {c3434};
    assign in3607_2 = {c3435};
    Full_Adder FA_3607(s3607, c3607, in3607_1, in3607_2, s3159[0]);
    wire[0:0] s3608, in3608_1, in3608_2;
    wire c3608;
    assign in3608_1 = {c3436};
    assign in3608_2 = {c3437};
    Full_Adder FA_3608(s3608, c3608, in3608_1, in3608_2, s3162[0]);
    wire[0:0] s3609, in3609_1, in3609_2;
    wire c3609;
    assign in3609_1 = {c3438};
    assign in3609_2 = {c3439};
    Full_Adder FA_3609(s3609, c3609, in3609_1, in3609_2, s3165[0]);
    wire[0:0] s3610, in3610_1, in3610_2;
    wire c3610;
    assign in3610_1 = {c3440};
    assign in3610_2 = {c3441};
    Full_Adder FA_3610(s3610, c3610, in3610_1, in3610_2, s3168[0]);
    wire[0:0] s3611, in3611_1, in3611_2;
    wire c3611;
    assign in3611_1 = {c3442};
    assign in3611_2 = {c3443};
    Full_Adder FA_3611(s3611, c3611, in3611_1, in3611_2, s3171[0]);
    wire[0:0] s3612, in3612_1, in3612_2;
    wire c3612;
    assign in3612_1 = {c3444};
    assign in3612_2 = {c3445};
    Full_Adder FA_3612(s3612, c3612, in3612_1, in3612_2, s3174[0]);
    wire[0:0] s3613, in3613_1, in3613_2;
    wire c3613;
    assign in3613_1 = {c3446};
    assign in3613_2 = {c3447};
    Full_Adder FA_3613(s3613, c3613, in3613_1, in3613_2, s3177[0]);
    wire[0:0] s3614, in3614_1, in3614_2;
    wire c3614;
    assign in3614_1 = {c3448};
    assign in3614_2 = {c3449};
    Full_Adder FA_3614(s3614, c3614, in3614_1, in3614_2, s3180[0]);
    wire[0:0] s3615, in3615_1, in3615_2;
    wire c3615;
    assign in3615_1 = {c3450};
    assign in3615_2 = {c3451};
    Full_Adder FA_3615(s3615, c3615, in3615_1, in3615_2, s3183[0]);
    wire[0:0] s3616, in3616_1, in3616_2;
    wire c3616;
    assign in3616_1 = {c3452};
    assign in3616_2 = {c3453};
    Full_Adder FA_3616(s3616, c3616, in3616_1, in3616_2, s3186[0]);
    wire[0:0] s3617, in3617_1, in3617_2;
    wire c3617;
    assign in3617_1 = {c3454};
    assign in3617_2 = {c3455};
    Full_Adder FA_3617(s3617, c3617, in3617_1, in3617_2, s3189[0]);
    wire[0:0] s3618, in3618_1, in3618_2;
    wire c3618;
    assign in3618_1 = {c3456};
    assign in3618_2 = {c3457};
    Full_Adder FA_3618(s3618, c3618, in3618_1, in3618_2, s3192[0]);
    wire[0:0] s3619, in3619_1, in3619_2;
    wire c3619;
    assign in3619_1 = {c3458};
    assign in3619_2 = {c3459};
    Full_Adder FA_3619(s3619, c3619, in3619_1, in3619_2, s3195[0]);
    wire[0:0] s3620, in3620_1, in3620_2;
    wire c3620;
    assign in3620_1 = {c3460};
    assign in3620_2 = {c3461};
    Full_Adder FA_3620(s3620, c3620, in3620_1, in3620_2, s3198[0]);
    wire[0:0] s3621, in3621_1, in3621_2;
    wire c3621;
    assign in3621_1 = {c3462};
    assign in3621_2 = {c3463};
    Full_Adder FA_3621(s3621, c3621, in3621_1, in3621_2, s3201[0]);
    wire[0:0] s3622, in3622_1, in3622_2;
    wire c3622;
    assign in3622_1 = {c3464};
    assign in3622_2 = {c3465};
    Full_Adder FA_3622(s3622, c3622, in3622_1, in3622_2, s3204[0]);
    wire[0:0] s3623, in3623_1, in3623_2;
    wire c3623;
    assign in3623_1 = {c3466};
    assign in3623_2 = {c3467};
    Full_Adder FA_3623(s3623, c3623, in3623_1, in3623_2, s3207[0]);
    wire[0:0] s3624, in3624_1, in3624_2;
    wire c3624;
    assign in3624_1 = {c3468};
    assign in3624_2 = {c3469};
    Full_Adder FA_3624(s3624, c3624, in3624_1, in3624_2, s3210[0]);
    wire[0:0] s3625, in3625_1, in3625_2;
    wire c3625;
    assign in3625_1 = {c3470};
    assign in3625_2 = {c3471};
    Full_Adder FA_3625(s3625, c3625, in3625_1, in3625_2, s3213[0]);
    wire[0:0] s3626, in3626_1, in3626_2;
    wire c3626;
    assign in3626_1 = {c3472};
    assign in3626_2 = {c3473};
    Full_Adder FA_3626(s3626, c3626, in3626_1, in3626_2, s3216[0]);
    wire[0:0] s3627, in3627_1, in3627_2;
    wire c3627;
    assign in3627_1 = {c3474};
    assign in3627_2 = {c3475};
    Full_Adder FA_3627(s3627, c3627, in3627_1, in3627_2, s3219[0]);
    wire[0:0] s3628, in3628_1, in3628_2;
    wire c3628;
    assign in3628_1 = {c3476};
    assign in3628_2 = {c3477};
    Full_Adder FA_3628(s3628, c3628, in3628_1, in3628_2, s3222[0]);
    wire[0:0] s3629, in3629_1, in3629_2;
    wire c3629;
    assign in3629_1 = {c3478};
    assign in3629_2 = {c3479};
    Full_Adder FA_3629(s3629, c3629, in3629_1, in3629_2, s3225[0]);
    wire[0:0] s3630, in3630_1, in3630_2;
    wire c3630;
    assign in3630_1 = {c3480};
    assign in3630_2 = {c3481};
    Full_Adder FA_3630(s3630, c3630, in3630_1, in3630_2, s3228[0]);
    wire[0:0] s3631, in3631_1, in3631_2;
    wire c3631;
    assign in3631_1 = {c3482};
    assign in3631_2 = {c3483};
    Full_Adder FA_3631(s3631, c3631, in3631_1, in3631_2, s3231[0]);
    wire[0:0] s3632, in3632_1, in3632_2;
    wire c3632;
    assign in3632_1 = {c3484};
    assign in3632_2 = {c3485};
    Full_Adder FA_3632(s3632, c3632, in3632_1, in3632_2, s3234[0]);
    wire[0:0] s3633, in3633_1, in3633_2;
    wire c3633;
    assign in3633_1 = {c3486};
    assign in3633_2 = {c3487};
    Full_Adder FA_3633(s3633, c3633, in3633_1, in3633_2, s3237[0]);
    wire[0:0] s3634, in3634_1, in3634_2;
    wire c3634;
    assign in3634_1 = {c3488};
    assign in3634_2 = {c3489};
    Full_Adder FA_3634(s3634, c3634, in3634_1, in3634_2, s3240[0]);
    wire[0:0] s3635, in3635_1, in3635_2;
    wire c3635;
    assign in3635_1 = {c3490};
    assign in3635_2 = {c3491};
    Full_Adder FA_3635(s3635, c3635, in3635_1, in3635_2, s3243[0]);
    wire[0:0] s3636, in3636_1, in3636_2;
    wire c3636;
    assign in3636_1 = {c3492};
    assign in3636_2 = {c3493};
    Full_Adder FA_3636(s3636, c3636, in3636_1, in3636_2, s3246[0]);
    wire[0:0] s3637, in3637_1, in3637_2;
    wire c3637;
    assign in3637_1 = {c3494};
    assign in3637_2 = {c3495};
    Full_Adder FA_3637(s3637, c3637, in3637_1, in3637_2, s3249[0]);
    wire[0:0] s3638, in3638_1, in3638_2;
    wire c3638;
    assign in3638_1 = {c3496};
    assign in3638_2 = {c3497};
    Full_Adder FA_3638(s3638, c3638, in3638_1, in3638_2, s3252[0]);
    wire[0:0] s3639, in3639_1, in3639_2;
    wire c3639;
    assign in3639_1 = {c3498};
    assign in3639_2 = {c3499};
    Full_Adder FA_3639(s3639, c3639, in3639_1, in3639_2, s3255[0]);
    wire[0:0] s3640, in3640_1, in3640_2;
    wire c3640;
    assign in3640_1 = {c3500};
    assign in3640_2 = {c3501};
    Full_Adder FA_3640(s3640, c3640, in3640_1, in3640_2, s3258[0]);
    wire[0:0] s3641, in3641_1, in3641_2;
    wire c3641;
    assign in3641_1 = {c3502};
    assign in3641_2 = {c3503};
    Full_Adder FA_3641(s3641, c3641, in3641_1, in3641_2, s3261[0]);
    wire[0:0] s3642, in3642_1, in3642_2;
    wire c3642;
    assign in3642_1 = {c3504};
    assign in3642_2 = {c3505};
    Full_Adder FA_3642(s3642, c3642, in3642_1, in3642_2, s3264[0]);
    wire[0:0] s3643, in3643_1, in3643_2;
    wire c3643;
    assign in3643_1 = {c3506};
    assign in3643_2 = {c3507};
    Full_Adder FA_3643(s3643, c3643, in3643_1, in3643_2, s3267[0]);
    wire[0:0] s3644, in3644_1, in3644_2;
    wire c3644;
    assign in3644_1 = {c3508};
    assign in3644_2 = {c3509};
    Full_Adder FA_3644(s3644, c3644, in3644_1, in3644_2, s3270[0]);
    wire[0:0] s3645, in3645_1, in3645_2;
    wire c3645;
    assign in3645_1 = {c3510};
    assign in3645_2 = {c3511};
    Full_Adder FA_3645(s3645, c3645, in3645_1, in3645_2, s3273[0]);
    wire[0:0] s3646, in3646_1, in3646_2;
    wire c3646;
    assign in3646_1 = {c3512};
    assign in3646_2 = {c3513};
    Full_Adder FA_3646(s3646, c3646, in3646_1, in3646_2, s3276[0]);
    wire[0:0] s3647, in3647_1, in3647_2;
    wire c3647;
    assign in3647_1 = {c3514};
    assign in3647_2 = {c3515};
    Full_Adder FA_3647(s3647, c3647, in3647_1, in3647_2, s3279[0]);
    wire[0:0] s3648, in3648_1, in3648_2;
    wire c3648;
    assign in3648_1 = {c3516};
    assign in3648_2 = {c3517};
    Full_Adder FA_3648(s3648, c3648, in3648_1, in3648_2, s3282[0]);
    wire[0:0] s3649, in3649_1, in3649_2;
    wire c3649;
    assign in3649_1 = {c3518};
    assign in3649_2 = {c3519};
    Full_Adder FA_3649(s3649, c3649, in3649_1, in3649_2, s3285[0]);
    wire[0:0] s3650, in3650_1, in3650_2;
    wire c3650;
    assign in3650_1 = {c3520};
    assign in3650_2 = {c3521};
    Full_Adder FA_3650(s3650, c3650, in3650_1, in3650_2, s3288[0]);
    wire[0:0] s3651, in3651_1, in3651_2;
    wire c3651;
    assign in3651_1 = {c3522};
    assign in3651_2 = {c3523};
    Full_Adder FA_3651(s3651, c3651, in3651_1, in3651_2, s3291[0]);
    wire[0:0] s3652, in3652_1, in3652_2;
    wire c3652;
    assign in3652_1 = {c3524};
    assign in3652_2 = {c3525};
    Full_Adder FA_3652(s3652, c3652, in3652_1, in3652_2, s3294[0]);
    wire[0:0] s3653, in3653_1, in3653_2;
    wire c3653;
    assign in3653_1 = {c3526};
    assign in3653_2 = {c3527};
    Full_Adder FA_3653(s3653, c3653, in3653_1, in3653_2, s3297[0]);
    wire[0:0] s3654, in3654_1, in3654_2;
    wire c3654;
    assign in3654_1 = {c3528};
    assign in3654_2 = {c3529};
    Full_Adder FA_3654(s3654, c3654, in3654_1, in3654_2, s3300[0]);
    wire[0:0] s3655, in3655_1, in3655_2;
    wire c3655;
    assign in3655_1 = {c3530};
    assign in3655_2 = {c3531};
    Full_Adder FA_3655(s3655, c3655, in3655_1, in3655_2, s3303[0]);
    wire[0:0] s3656, in3656_1, in3656_2;
    wire c3656;
    assign in3656_1 = {c3532};
    assign in3656_2 = {c3533};
    Full_Adder FA_3656(s3656, c3656, in3656_1, in3656_2, s3305[0]);
    wire[0:0] s3657, in3657_1, in3657_2;
    wire c3657;
    assign in3657_1 = {c3534};
    assign in3657_2 = {c3535};
    Full_Adder FA_3657(s3657, c3657, in3657_1, in3657_2, s3306[0]);
    wire[0:0] s3658, in3658_1, in3658_2;
    wire c3658;
    assign in3658_1 = {c3536};
    assign in3658_2 = {c3537};
    Full_Adder FA_3658(s3658, c3658, in3658_1, in3658_2, c3306);
    wire[0:0] s3659, in3659_1, in3659_2;
    wire c3659;
    assign in3659_1 = {pp63[59]};
    assign in3659_2 = {c3538};
    Full_Adder FA_3659(s3659, c3659, in3659_1, in3659_2, pp62[60]);
    wire[0:0] s3660, in3660_1, in3660_2;
    wire c3660;
    assign in3660_1 = {pp61[62]};
    assign in3660_2 = {pp62[61]};
    Full_Adder FA_3660(s3660, c3660, in3660_1, in3660_2, pp60[63]);

    /*Stage 9*/
    wire[0:0] s3661, in3661_1, in3661_2;
    wire c3661;
    assign in3661_1 = {pp0[3]};
    assign in3661_2 = {pp1[2]};
    Half_Adder HA_3661(s3661, c3661, in3661_1, in3661_2);
    wire[0:0] s3662, in3662_1, in3662_2;
    wire c3662;
    assign in3662_1 = {pp3[1]};
    assign in3662_2 = {pp4[0]};
    Full_Adder FA_3662(s3662, c3662, in3662_1, in3662_2, pp2[2]);
    wire[0:0] s3663, in3663_1, in3663_2;
    wire c3663;
    assign in3663_1 = {s3307[0]};
    assign in3663_2 = {c3541};
    Full_Adder FA_3663(s3663, c3663, in3663_1, in3663_2, pp5[0]);
    wire[0:0] s3664, in3664_1, in3664_2;
    wire c3664;
    assign in3664_1 = {s3309[0]};
    assign in3664_2 = {c3542};
    Full_Adder FA_3664(s3664, c3664, in3664_1, in3664_2, s3308[0]);
    wire[0:0] s3665, in3665_1, in3665_2;
    wire c3665;
    assign in3665_1 = {s3311[0]};
    assign in3665_2 = {c3543};
    Full_Adder FA_3665(s3665, c3665, in3665_1, in3665_2, s3310[0]);
    wire[0:0] s3666, in3666_1, in3666_2;
    wire c3666;
    assign in3666_1 = {s3313[0]};
    assign in3666_2 = {c3544};
    Full_Adder FA_3666(s3666, c3666, in3666_1, in3666_2, s3312[0]);
    wire[0:0] s3667, in3667_1, in3667_2;
    wire c3667;
    assign in3667_1 = {s3315[0]};
    assign in3667_2 = {c3545};
    Full_Adder FA_3667(s3667, c3667, in3667_1, in3667_2, s3314[0]);
    wire[0:0] s3668, in3668_1, in3668_2;
    wire c3668;
    assign in3668_1 = {s3317[0]};
    assign in3668_2 = {c3546};
    Full_Adder FA_3668(s3668, c3668, in3668_1, in3668_2, s3316[0]);
    wire[0:0] s3669, in3669_1, in3669_2;
    wire c3669;
    assign in3669_1 = {s3319[0]};
    assign in3669_2 = {c3547};
    Full_Adder FA_3669(s3669, c3669, in3669_1, in3669_2, s3318[0]);
    wire[0:0] s3670, in3670_1, in3670_2;
    wire c3670;
    assign in3670_1 = {s3321[0]};
    assign in3670_2 = {c3548};
    Full_Adder FA_3670(s3670, c3670, in3670_1, in3670_2, s3320[0]);
    wire[0:0] s3671, in3671_1, in3671_2;
    wire c3671;
    assign in3671_1 = {s3323[0]};
    assign in3671_2 = {c3549};
    Full_Adder FA_3671(s3671, c3671, in3671_1, in3671_2, s3322[0]);
    wire[0:0] s3672, in3672_1, in3672_2;
    wire c3672;
    assign in3672_1 = {s3325[0]};
    assign in3672_2 = {c3550};
    Full_Adder FA_3672(s3672, c3672, in3672_1, in3672_2, s3324[0]);
    wire[0:0] s3673, in3673_1, in3673_2;
    wire c3673;
    assign in3673_1 = {s3327[0]};
    assign in3673_2 = {c3551};
    Full_Adder FA_3673(s3673, c3673, in3673_1, in3673_2, s3326[0]);
    wire[0:0] s3674, in3674_1, in3674_2;
    wire c3674;
    assign in3674_1 = {s3329[0]};
    assign in3674_2 = {c3552};
    Full_Adder FA_3674(s3674, c3674, in3674_1, in3674_2, s3328[0]);
    wire[0:0] s3675, in3675_1, in3675_2;
    wire c3675;
    assign in3675_1 = {s3331[0]};
    assign in3675_2 = {c3553};
    Full_Adder FA_3675(s3675, c3675, in3675_1, in3675_2, s3330[0]);
    wire[0:0] s3676, in3676_1, in3676_2;
    wire c3676;
    assign in3676_1 = {s3333[0]};
    assign in3676_2 = {c3554};
    Full_Adder FA_3676(s3676, c3676, in3676_1, in3676_2, s3332[0]);
    wire[0:0] s3677, in3677_1, in3677_2;
    wire c3677;
    assign in3677_1 = {s3335[0]};
    assign in3677_2 = {c3555};
    Full_Adder FA_3677(s3677, c3677, in3677_1, in3677_2, s3334[0]);
    wire[0:0] s3678, in3678_1, in3678_2;
    wire c3678;
    assign in3678_1 = {s3337[0]};
    assign in3678_2 = {c3556};
    Full_Adder FA_3678(s3678, c3678, in3678_1, in3678_2, s3336[0]);
    wire[0:0] s3679, in3679_1, in3679_2;
    wire c3679;
    assign in3679_1 = {s3339[0]};
    assign in3679_2 = {c3557};
    Full_Adder FA_3679(s3679, c3679, in3679_1, in3679_2, s3338[0]);
    wire[0:0] s3680, in3680_1, in3680_2;
    wire c3680;
    assign in3680_1 = {s3341[0]};
    assign in3680_2 = {c3558};
    Full_Adder FA_3680(s3680, c3680, in3680_1, in3680_2, s3340[0]);
    wire[0:0] s3681, in3681_1, in3681_2;
    wire c3681;
    assign in3681_1 = {s3343[0]};
    assign in3681_2 = {c3559};
    Full_Adder FA_3681(s3681, c3681, in3681_1, in3681_2, s3342[0]);
    wire[0:0] s3682, in3682_1, in3682_2;
    wire c3682;
    assign in3682_1 = {s3345[0]};
    assign in3682_2 = {c3560};
    Full_Adder FA_3682(s3682, c3682, in3682_1, in3682_2, s3344[0]);
    wire[0:0] s3683, in3683_1, in3683_2;
    wire c3683;
    assign in3683_1 = {s3347[0]};
    assign in3683_2 = {c3561};
    Full_Adder FA_3683(s3683, c3683, in3683_1, in3683_2, s3346[0]);
    wire[0:0] s3684, in3684_1, in3684_2;
    wire c3684;
    assign in3684_1 = {s3349[0]};
    assign in3684_2 = {c3562};
    Full_Adder FA_3684(s3684, c3684, in3684_1, in3684_2, s3348[0]);
    wire[0:0] s3685, in3685_1, in3685_2;
    wire c3685;
    assign in3685_1 = {s3351[0]};
    assign in3685_2 = {c3563};
    Full_Adder FA_3685(s3685, c3685, in3685_1, in3685_2, s3350[0]);
    wire[0:0] s3686, in3686_1, in3686_2;
    wire c3686;
    assign in3686_1 = {s3353[0]};
    assign in3686_2 = {c3564};
    Full_Adder FA_3686(s3686, c3686, in3686_1, in3686_2, s3352[0]);
    wire[0:0] s3687, in3687_1, in3687_2;
    wire c3687;
    assign in3687_1 = {s3355[0]};
    assign in3687_2 = {c3565};
    Full_Adder FA_3687(s3687, c3687, in3687_1, in3687_2, s3354[0]);
    wire[0:0] s3688, in3688_1, in3688_2;
    wire c3688;
    assign in3688_1 = {s3357[0]};
    assign in3688_2 = {c3566};
    Full_Adder FA_3688(s3688, c3688, in3688_1, in3688_2, s3356[0]);
    wire[0:0] s3689, in3689_1, in3689_2;
    wire c3689;
    assign in3689_1 = {s3359[0]};
    assign in3689_2 = {c3567};
    Full_Adder FA_3689(s3689, c3689, in3689_1, in3689_2, s3358[0]);
    wire[0:0] s3690, in3690_1, in3690_2;
    wire c3690;
    assign in3690_1 = {s3361[0]};
    assign in3690_2 = {c3568};
    Full_Adder FA_3690(s3690, c3690, in3690_1, in3690_2, s3360[0]);
    wire[0:0] s3691, in3691_1, in3691_2;
    wire c3691;
    assign in3691_1 = {s3363[0]};
    assign in3691_2 = {c3569};
    Full_Adder FA_3691(s3691, c3691, in3691_1, in3691_2, s3362[0]);
    wire[0:0] s3692, in3692_1, in3692_2;
    wire c3692;
    assign in3692_1 = {s3365[0]};
    assign in3692_2 = {c3570};
    Full_Adder FA_3692(s3692, c3692, in3692_1, in3692_2, s3364[0]);
    wire[0:0] s3693, in3693_1, in3693_2;
    wire c3693;
    assign in3693_1 = {s3367[0]};
    assign in3693_2 = {c3571};
    Full_Adder FA_3693(s3693, c3693, in3693_1, in3693_2, s3366[0]);
    wire[0:0] s3694, in3694_1, in3694_2;
    wire c3694;
    assign in3694_1 = {s3369[0]};
    assign in3694_2 = {c3572};
    Full_Adder FA_3694(s3694, c3694, in3694_1, in3694_2, s3368[0]);
    wire[0:0] s3695, in3695_1, in3695_2;
    wire c3695;
    assign in3695_1 = {s3371[0]};
    assign in3695_2 = {c3573};
    Full_Adder FA_3695(s3695, c3695, in3695_1, in3695_2, s3370[0]);
    wire[0:0] s3696, in3696_1, in3696_2;
    wire c3696;
    assign in3696_1 = {s3373[0]};
    assign in3696_2 = {c3574};
    Full_Adder FA_3696(s3696, c3696, in3696_1, in3696_2, s3372[0]);
    wire[0:0] s3697, in3697_1, in3697_2;
    wire c3697;
    assign in3697_1 = {s3375[0]};
    assign in3697_2 = {c3575};
    Full_Adder FA_3697(s3697, c3697, in3697_1, in3697_2, s3374[0]);
    wire[0:0] s3698, in3698_1, in3698_2;
    wire c3698;
    assign in3698_1 = {s3377[0]};
    assign in3698_2 = {c3576};
    Full_Adder FA_3698(s3698, c3698, in3698_1, in3698_2, s3376[0]);
    wire[0:0] s3699, in3699_1, in3699_2;
    wire c3699;
    assign in3699_1 = {s3379[0]};
    assign in3699_2 = {c3577};
    Full_Adder FA_3699(s3699, c3699, in3699_1, in3699_2, s3378[0]);
    wire[0:0] s3700, in3700_1, in3700_2;
    wire c3700;
    assign in3700_1 = {s3381[0]};
    assign in3700_2 = {c3578};
    Full_Adder FA_3700(s3700, c3700, in3700_1, in3700_2, s3380[0]);
    wire[0:0] s3701, in3701_1, in3701_2;
    wire c3701;
    assign in3701_1 = {s3383[0]};
    assign in3701_2 = {c3579};
    Full_Adder FA_3701(s3701, c3701, in3701_1, in3701_2, s3382[0]);
    wire[0:0] s3702, in3702_1, in3702_2;
    wire c3702;
    assign in3702_1 = {s3385[0]};
    assign in3702_2 = {c3580};
    Full_Adder FA_3702(s3702, c3702, in3702_1, in3702_2, s3384[0]);
    wire[0:0] s3703, in3703_1, in3703_2;
    wire c3703;
    assign in3703_1 = {s3387[0]};
    assign in3703_2 = {c3581};
    Full_Adder FA_3703(s3703, c3703, in3703_1, in3703_2, s3386[0]);
    wire[0:0] s3704, in3704_1, in3704_2;
    wire c3704;
    assign in3704_1 = {s3389[0]};
    assign in3704_2 = {c3582};
    Full_Adder FA_3704(s3704, c3704, in3704_1, in3704_2, s3388[0]);
    wire[0:0] s3705, in3705_1, in3705_2;
    wire c3705;
    assign in3705_1 = {s3391[0]};
    assign in3705_2 = {c3583};
    Full_Adder FA_3705(s3705, c3705, in3705_1, in3705_2, s3390[0]);
    wire[0:0] s3706, in3706_1, in3706_2;
    wire c3706;
    assign in3706_1 = {s3393[0]};
    assign in3706_2 = {c3584};
    Full_Adder FA_3706(s3706, c3706, in3706_1, in3706_2, s3392[0]);
    wire[0:0] s3707, in3707_1, in3707_2;
    wire c3707;
    assign in3707_1 = {s3395[0]};
    assign in3707_2 = {c3585};
    Full_Adder FA_3707(s3707, c3707, in3707_1, in3707_2, s3394[0]);
    wire[0:0] s3708, in3708_1, in3708_2;
    wire c3708;
    assign in3708_1 = {s3397[0]};
    assign in3708_2 = {c3586};
    Full_Adder FA_3708(s3708, c3708, in3708_1, in3708_2, s3396[0]);
    wire[0:0] s3709, in3709_1, in3709_2;
    wire c3709;
    assign in3709_1 = {s3399[0]};
    assign in3709_2 = {c3587};
    Full_Adder FA_3709(s3709, c3709, in3709_1, in3709_2, s3398[0]);
    wire[0:0] s3710, in3710_1, in3710_2;
    wire c3710;
    assign in3710_1 = {s3401[0]};
    assign in3710_2 = {c3588};
    Full_Adder FA_3710(s3710, c3710, in3710_1, in3710_2, s3400[0]);
    wire[0:0] s3711, in3711_1, in3711_2;
    wire c3711;
    assign in3711_1 = {s3403[0]};
    assign in3711_2 = {c3589};
    Full_Adder FA_3711(s3711, c3711, in3711_1, in3711_2, s3402[0]);
    wire[0:0] s3712, in3712_1, in3712_2;
    wire c3712;
    assign in3712_1 = {s3405[0]};
    assign in3712_2 = {c3590};
    Full_Adder FA_3712(s3712, c3712, in3712_1, in3712_2, s3404[0]);
    wire[0:0] s3713, in3713_1, in3713_2;
    wire c3713;
    assign in3713_1 = {s3407[0]};
    assign in3713_2 = {c3591};
    Full_Adder FA_3713(s3713, c3713, in3713_1, in3713_2, s3406[0]);
    wire[0:0] s3714, in3714_1, in3714_2;
    wire c3714;
    assign in3714_1 = {s3409[0]};
    assign in3714_2 = {c3592};
    Full_Adder FA_3714(s3714, c3714, in3714_1, in3714_2, s3408[0]);
    wire[0:0] s3715, in3715_1, in3715_2;
    wire c3715;
    assign in3715_1 = {s3411[0]};
    assign in3715_2 = {c3593};
    Full_Adder FA_3715(s3715, c3715, in3715_1, in3715_2, s3410[0]);
    wire[0:0] s3716, in3716_1, in3716_2;
    wire c3716;
    assign in3716_1 = {s3413[0]};
    assign in3716_2 = {c3594};
    Full_Adder FA_3716(s3716, c3716, in3716_1, in3716_2, s3412[0]);
    wire[0:0] s3717, in3717_1, in3717_2;
    wire c3717;
    assign in3717_1 = {s3415[0]};
    assign in3717_2 = {c3595};
    Full_Adder FA_3717(s3717, c3717, in3717_1, in3717_2, s3414[0]);
    wire[0:0] s3718, in3718_1, in3718_2;
    wire c3718;
    assign in3718_1 = {s3417[0]};
    assign in3718_2 = {c3596};
    Full_Adder FA_3718(s3718, c3718, in3718_1, in3718_2, s3416[0]);
    wire[0:0] s3719, in3719_1, in3719_2;
    wire c3719;
    assign in3719_1 = {s3419[0]};
    assign in3719_2 = {c3597};
    Full_Adder FA_3719(s3719, c3719, in3719_1, in3719_2, s3418[0]);
    wire[0:0] s3720, in3720_1, in3720_2;
    wire c3720;
    assign in3720_1 = {s3421[0]};
    assign in3720_2 = {c3598};
    Full_Adder FA_3720(s3720, c3720, in3720_1, in3720_2, s3420[0]);
    wire[0:0] s3721, in3721_1, in3721_2;
    wire c3721;
    assign in3721_1 = {s3423[0]};
    assign in3721_2 = {c3599};
    Full_Adder FA_3721(s3721, c3721, in3721_1, in3721_2, s3422[0]);
    wire[0:0] s3722, in3722_1, in3722_2;
    wire c3722;
    assign in3722_1 = {s3425[0]};
    assign in3722_2 = {c3600};
    Full_Adder FA_3722(s3722, c3722, in3722_1, in3722_2, s3424[0]);
    wire[0:0] s3723, in3723_1, in3723_2;
    wire c3723;
    assign in3723_1 = {s3427[0]};
    assign in3723_2 = {c3601};
    Full_Adder FA_3723(s3723, c3723, in3723_1, in3723_2, s3426[0]);
    wire[0:0] s3724, in3724_1, in3724_2;
    wire c3724;
    assign in3724_1 = {s3429[0]};
    assign in3724_2 = {c3602};
    Full_Adder FA_3724(s3724, c3724, in3724_1, in3724_2, s3428[0]);
    wire[0:0] s3725, in3725_1, in3725_2;
    wire c3725;
    assign in3725_1 = {s3431[0]};
    assign in3725_2 = {c3603};
    Full_Adder FA_3725(s3725, c3725, in3725_1, in3725_2, s3430[0]);
    wire[0:0] s3726, in3726_1, in3726_2;
    wire c3726;
    assign in3726_1 = {s3433[0]};
    assign in3726_2 = {c3604};
    Full_Adder FA_3726(s3726, c3726, in3726_1, in3726_2, s3432[0]);
    wire[0:0] s3727, in3727_1, in3727_2;
    wire c3727;
    assign in3727_1 = {s3435[0]};
    assign in3727_2 = {c3605};
    Full_Adder FA_3727(s3727, c3727, in3727_1, in3727_2, s3434[0]);
    wire[0:0] s3728, in3728_1, in3728_2;
    wire c3728;
    assign in3728_1 = {s3437[0]};
    assign in3728_2 = {c3606};
    Full_Adder FA_3728(s3728, c3728, in3728_1, in3728_2, s3436[0]);
    wire[0:0] s3729, in3729_1, in3729_2;
    wire c3729;
    assign in3729_1 = {s3439[0]};
    assign in3729_2 = {c3607};
    Full_Adder FA_3729(s3729, c3729, in3729_1, in3729_2, s3438[0]);
    wire[0:0] s3730, in3730_1, in3730_2;
    wire c3730;
    assign in3730_1 = {s3441[0]};
    assign in3730_2 = {c3608};
    Full_Adder FA_3730(s3730, c3730, in3730_1, in3730_2, s3440[0]);
    wire[0:0] s3731, in3731_1, in3731_2;
    wire c3731;
    assign in3731_1 = {s3443[0]};
    assign in3731_2 = {c3609};
    Full_Adder FA_3731(s3731, c3731, in3731_1, in3731_2, s3442[0]);
    wire[0:0] s3732, in3732_1, in3732_2;
    wire c3732;
    assign in3732_1 = {s3445[0]};
    assign in3732_2 = {c3610};
    Full_Adder FA_3732(s3732, c3732, in3732_1, in3732_2, s3444[0]);
    wire[0:0] s3733, in3733_1, in3733_2;
    wire c3733;
    assign in3733_1 = {s3447[0]};
    assign in3733_2 = {c3611};
    Full_Adder FA_3733(s3733, c3733, in3733_1, in3733_2, s3446[0]);
    wire[0:0] s3734, in3734_1, in3734_2;
    wire c3734;
    assign in3734_1 = {s3449[0]};
    assign in3734_2 = {c3612};
    Full_Adder FA_3734(s3734, c3734, in3734_1, in3734_2, s3448[0]);
    wire[0:0] s3735, in3735_1, in3735_2;
    wire c3735;
    assign in3735_1 = {s3451[0]};
    assign in3735_2 = {c3613};
    Full_Adder FA_3735(s3735, c3735, in3735_1, in3735_2, s3450[0]);
    wire[0:0] s3736, in3736_1, in3736_2;
    wire c3736;
    assign in3736_1 = {s3453[0]};
    assign in3736_2 = {c3614};
    Full_Adder FA_3736(s3736, c3736, in3736_1, in3736_2, s3452[0]);
    wire[0:0] s3737, in3737_1, in3737_2;
    wire c3737;
    assign in3737_1 = {s3455[0]};
    assign in3737_2 = {c3615};
    Full_Adder FA_3737(s3737, c3737, in3737_1, in3737_2, s3454[0]);
    wire[0:0] s3738, in3738_1, in3738_2;
    wire c3738;
    assign in3738_1 = {s3457[0]};
    assign in3738_2 = {c3616};
    Full_Adder FA_3738(s3738, c3738, in3738_1, in3738_2, s3456[0]);
    wire[0:0] s3739, in3739_1, in3739_2;
    wire c3739;
    assign in3739_1 = {s3459[0]};
    assign in3739_2 = {c3617};
    Full_Adder FA_3739(s3739, c3739, in3739_1, in3739_2, s3458[0]);
    wire[0:0] s3740, in3740_1, in3740_2;
    wire c3740;
    assign in3740_1 = {s3461[0]};
    assign in3740_2 = {c3618};
    Full_Adder FA_3740(s3740, c3740, in3740_1, in3740_2, s3460[0]);
    wire[0:0] s3741, in3741_1, in3741_2;
    wire c3741;
    assign in3741_1 = {s3463[0]};
    assign in3741_2 = {c3619};
    Full_Adder FA_3741(s3741, c3741, in3741_1, in3741_2, s3462[0]);
    wire[0:0] s3742, in3742_1, in3742_2;
    wire c3742;
    assign in3742_1 = {s3465[0]};
    assign in3742_2 = {c3620};
    Full_Adder FA_3742(s3742, c3742, in3742_1, in3742_2, s3464[0]);
    wire[0:0] s3743, in3743_1, in3743_2;
    wire c3743;
    assign in3743_1 = {s3467[0]};
    assign in3743_2 = {c3621};
    Full_Adder FA_3743(s3743, c3743, in3743_1, in3743_2, s3466[0]);
    wire[0:0] s3744, in3744_1, in3744_2;
    wire c3744;
    assign in3744_1 = {s3469[0]};
    assign in3744_2 = {c3622};
    Full_Adder FA_3744(s3744, c3744, in3744_1, in3744_2, s3468[0]);
    wire[0:0] s3745, in3745_1, in3745_2;
    wire c3745;
    assign in3745_1 = {s3471[0]};
    assign in3745_2 = {c3623};
    Full_Adder FA_3745(s3745, c3745, in3745_1, in3745_2, s3470[0]);
    wire[0:0] s3746, in3746_1, in3746_2;
    wire c3746;
    assign in3746_1 = {s3473[0]};
    assign in3746_2 = {c3624};
    Full_Adder FA_3746(s3746, c3746, in3746_1, in3746_2, s3472[0]);
    wire[0:0] s3747, in3747_1, in3747_2;
    wire c3747;
    assign in3747_1 = {s3475[0]};
    assign in3747_2 = {c3625};
    Full_Adder FA_3747(s3747, c3747, in3747_1, in3747_2, s3474[0]);
    wire[0:0] s3748, in3748_1, in3748_2;
    wire c3748;
    assign in3748_1 = {s3477[0]};
    assign in3748_2 = {c3626};
    Full_Adder FA_3748(s3748, c3748, in3748_1, in3748_2, s3476[0]);
    wire[0:0] s3749, in3749_1, in3749_2;
    wire c3749;
    assign in3749_1 = {s3479[0]};
    assign in3749_2 = {c3627};
    Full_Adder FA_3749(s3749, c3749, in3749_1, in3749_2, s3478[0]);
    wire[0:0] s3750, in3750_1, in3750_2;
    wire c3750;
    assign in3750_1 = {s3481[0]};
    assign in3750_2 = {c3628};
    Full_Adder FA_3750(s3750, c3750, in3750_1, in3750_2, s3480[0]);
    wire[0:0] s3751, in3751_1, in3751_2;
    wire c3751;
    assign in3751_1 = {s3483[0]};
    assign in3751_2 = {c3629};
    Full_Adder FA_3751(s3751, c3751, in3751_1, in3751_2, s3482[0]);
    wire[0:0] s3752, in3752_1, in3752_2;
    wire c3752;
    assign in3752_1 = {s3485[0]};
    assign in3752_2 = {c3630};
    Full_Adder FA_3752(s3752, c3752, in3752_1, in3752_2, s3484[0]);
    wire[0:0] s3753, in3753_1, in3753_2;
    wire c3753;
    assign in3753_1 = {s3487[0]};
    assign in3753_2 = {c3631};
    Full_Adder FA_3753(s3753, c3753, in3753_1, in3753_2, s3486[0]);
    wire[0:0] s3754, in3754_1, in3754_2;
    wire c3754;
    assign in3754_1 = {s3489[0]};
    assign in3754_2 = {c3632};
    Full_Adder FA_3754(s3754, c3754, in3754_1, in3754_2, s3488[0]);
    wire[0:0] s3755, in3755_1, in3755_2;
    wire c3755;
    assign in3755_1 = {s3491[0]};
    assign in3755_2 = {c3633};
    Full_Adder FA_3755(s3755, c3755, in3755_1, in3755_2, s3490[0]);
    wire[0:0] s3756, in3756_1, in3756_2;
    wire c3756;
    assign in3756_1 = {s3493[0]};
    assign in3756_2 = {c3634};
    Full_Adder FA_3756(s3756, c3756, in3756_1, in3756_2, s3492[0]);
    wire[0:0] s3757, in3757_1, in3757_2;
    wire c3757;
    assign in3757_1 = {s3495[0]};
    assign in3757_2 = {c3635};
    Full_Adder FA_3757(s3757, c3757, in3757_1, in3757_2, s3494[0]);
    wire[0:0] s3758, in3758_1, in3758_2;
    wire c3758;
    assign in3758_1 = {s3497[0]};
    assign in3758_2 = {c3636};
    Full_Adder FA_3758(s3758, c3758, in3758_1, in3758_2, s3496[0]);
    wire[0:0] s3759, in3759_1, in3759_2;
    wire c3759;
    assign in3759_1 = {s3499[0]};
    assign in3759_2 = {c3637};
    Full_Adder FA_3759(s3759, c3759, in3759_1, in3759_2, s3498[0]);
    wire[0:0] s3760, in3760_1, in3760_2;
    wire c3760;
    assign in3760_1 = {s3501[0]};
    assign in3760_2 = {c3638};
    Full_Adder FA_3760(s3760, c3760, in3760_1, in3760_2, s3500[0]);
    wire[0:0] s3761, in3761_1, in3761_2;
    wire c3761;
    assign in3761_1 = {s3503[0]};
    assign in3761_2 = {c3639};
    Full_Adder FA_3761(s3761, c3761, in3761_1, in3761_2, s3502[0]);
    wire[0:0] s3762, in3762_1, in3762_2;
    wire c3762;
    assign in3762_1 = {s3505[0]};
    assign in3762_2 = {c3640};
    Full_Adder FA_3762(s3762, c3762, in3762_1, in3762_2, s3504[0]);
    wire[0:0] s3763, in3763_1, in3763_2;
    wire c3763;
    assign in3763_1 = {s3507[0]};
    assign in3763_2 = {c3641};
    Full_Adder FA_3763(s3763, c3763, in3763_1, in3763_2, s3506[0]);
    wire[0:0] s3764, in3764_1, in3764_2;
    wire c3764;
    assign in3764_1 = {s3509[0]};
    assign in3764_2 = {c3642};
    Full_Adder FA_3764(s3764, c3764, in3764_1, in3764_2, s3508[0]);
    wire[0:0] s3765, in3765_1, in3765_2;
    wire c3765;
    assign in3765_1 = {s3511[0]};
    assign in3765_2 = {c3643};
    Full_Adder FA_3765(s3765, c3765, in3765_1, in3765_2, s3510[0]);
    wire[0:0] s3766, in3766_1, in3766_2;
    wire c3766;
    assign in3766_1 = {s3513[0]};
    assign in3766_2 = {c3644};
    Full_Adder FA_3766(s3766, c3766, in3766_1, in3766_2, s3512[0]);
    wire[0:0] s3767, in3767_1, in3767_2;
    wire c3767;
    assign in3767_1 = {s3515[0]};
    assign in3767_2 = {c3645};
    Full_Adder FA_3767(s3767, c3767, in3767_1, in3767_2, s3514[0]);
    wire[0:0] s3768, in3768_1, in3768_2;
    wire c3768;
    assign in3768_1 = {s3517[0]};
    assign in3768_2 = {c3646};
    Full_Adder FA_3768(s3768, c3768, in3768_1, in3768_2, s3516[0]);
    wire[0:0] s3769, in3769_1, in3769_2;
    wire c3769;
    assign in3769_1 = {s3519[0]};
    assign in3769_2 = {c3647};
    Full_Adder FA_3769(s3769, c3769, in3769_1, in3769_2, s3518[0]);
    wire[0:0] s3770, in3770_1, in3770_2;
    wire c3770;
    assign in3770_1 = {s3521[0]};
    assign in3770_2 = {c3648};
    Full_Adder FA_3770(s3770, c3770, in3770_1, in3770_2, s3520[0]);
    wire[0:0] s3771, in3771_1, in3771_2;
    wire c3771;
    assign in3771_1 = {s3523[0]};
    assign in3771_2 = {c3649};
    Full_Adder FA_3771(s3771, c3771, in3771_1, in3771_2, s3522[0]);
    wire[0:0] s3772, in3772_1, in3772_2;
    wire c3772;
    assign in3772_1 = {s3525[0]};
    assign in3772_2 = {c3650};
    Full_Adder FA_3772(s3772, c3772, in3772_1, in3772_2, s3524[0]);
    wire[0:0] s3773, in3773_1, in3773_2;
    wire c3773;
    assign in3773_1 = {s3527[0]};
    assign in3773_2 = {c3651};
    Full_Adder FA_3773(s3773, c3773, in3773_1, in3773_2, s3526[0]);
    wire[0:0] s3774, in3774_1, in3774_2;
    wire c3774;
    assign in3774_1 = {s3529[0]};
    assign in3774_2 = {c3652};
    Full_Adder FA_3774(s3774, c3774, in3774_1, in3774_2, s3528[0]);
    wire[0:0] s3775, in3775_1, in3775_2;
    wire c3775;
    assign in3775_1 = {s3531[0]};
    assign in3775_2 = {c3653};
    Full_Adder FA_3775(s3775, c3775, in3775_1, in3775_2, s3530[0]);
    wire[0:0] s3776, in3776_1, in3776_2;
    wire c3776;
    assign in3776_1 = {s3533[0]};
    assign in3776_2 = {c3654};
    Full_Adder FA_3776(s3776, c3776, in3776_1, in3776_2, s3532[0]);
    wire[0:0] s3777, in3777_1, in3777_2;
    wire c3777;
    assign in3777_1 = {s3535[0]};
    assign in3777_2 = {c3655};
    Full_Adder FA_3777(s3777, c3777, in3777_1, in3777_2, s3534[0]);
    wire[0:0] s3778, in3778_1, in3778_2;
    wire c3778;
    assign in3778_1 = {s3537[0]};
    assign in3778_2 = {c3656};
    Full_Adder FA_3778(s3778, c3778, in3778_1, in3778_2, s3536[0]);
    wire[0:0] s3779, in3779_1, in3779_2;
    wire c3779;
    assign in3779_1 = {s3539[0]};
    assign in3779_2 = {c3657};
    Full_Adder FA_3779(s3779, c3779, in3779_1, in3779_2, s3538[0]);
    wire[0:0] s3780, in3780_1, in3780_2;
    wire c3780;
    assign in3780_1 = {s3540[0]};
    assign in3780_2 = {c3658};
    Full_Adder FA_3780(s3780, c3780, in3780_1, in3780_2, c3539);
    wire[0:0] s3781, in3781_1, in3781_2;
    wire c3781;
    assign in3781_1 = {c3540};
    assign in3781_2 = {c3659};
    Full_Adder FA_3781(s3781, c3781, in3781_1, in3781_2, pp63[60]);
    wire[0:0] s3782, in3782_1, in3782_2;
    wire c3782;
    assign in3782_1 = {pp62[62]};
    assign in3782_2 = {pp63[61]};
    Full_Adder FA_3782(s3782, c3782, in3782_1, in3782_2, pp61[63]);

    /*Stage 10*/
    wire[0:0] s3783, in3783_1, in3783_2;
    wire c3783;
    assign in3783_1 = {pp0[2]};
    assign in3783_2 = {pp1[1]};
    Half_Adder HA_3783(s3783, c3783, in3783_1, in3783_2);
    wire[0:0] s3784, in3784_1, in3784_2;
    wire c3784;
    assign in3784_1 = {pp3[0]};
    assign in3784_2 = {s3661[0]};
    Full_Adder FA_3784(s3784, c3784, in3784_1, in3784_2, pp2[1]);
    wire[0:0] s3785, in3785_1, in3785_2;
    wire c3785;
    assign in3785_1 = {c3661};
    assign in3785_2 = {s3662[0]};
    Full_Adder FA_3785(s3785, c3785, in3785_1, in3785_2, s3541[0]);
    wire[0:0] s3786, in3786_1, in3786_2;
    wire c3786;
    assign in3786_1 = {c3662};
    assign in3786_2 = {s3663[0]};
    Full_Adder FA_3786(s3786, c3786, in3786_1, in3786_2, s3542[0]);
    wire[0:0] s3787, in3787_1, in3787_2;
    wire c3787;
    assign in3787_1 = {c3663};
    assign in3787_2 = {s3664[0]};
    Full_Adder FA_3787(s3787, c3787, in3787_1, in3787_2, s3543[0]);
    wire[0:0] s3788, in3788_1, in3788_2;
    wire c3788;
    assign in3788_1 = {c3664};
    assign in3788_2 = {s3665[0]};
    Full_Adder FA_3788(s3788, c3788, in3788_1, in3788_2, s3544[0]);
    wire[0:0] s3789, in3789_1, in3789_2;
    wire c3789;
    assign in3789_1 = {c3665};
    assign in3789_2 = {s3666[0]};
    Full_Adder FA_3789(s3789, c3789, in3789_1, in3789_2, s3545[0]);
    wire[0:0] s3790, in3790_1, in3790_2;
    wire c3790;
    assign in3790_1 = {c3666};
    assign in3790_2 = {s3667[0]};
    Full_Adder FA_3790(s3790, c3790, in3790_1, in3790_2, s3546[0]);
    wire[0:0] s3791, in3791_1, in3791_2;
    wire c3791;
    assign in3791_1 = {c3667};
    assign in3791_2 = {s3668[0]};
    Full_Adder FA_3791(s3791, c3791, in3791_1, in3791_2, s3547[0]);
    wire[0:0] s3792, in3792_1, in3792_2;
    wire c3792;
    assign in3792_1 = {c3668};
    assign in3792_2 = {s3669[0]};
    Full_Adder FA_3792(s3792, c3792, in3792_1, in3792_2, s3548[0]);
    wire[0:0] s3793, in3793_1, in3793_2;
    wire c3793;
    assign in3793_1 = {c3669};
    assign in3793_2 = {s3670[0]};
    Full_Adder FA_3793(s3793, c3793, in3793_1, in3793_2, s3549[0]);
    wire[0:0] s3794, in3794_1, in3794_2;
    wire c3794;
    assign in3794_1 = {c3670};
    assign in3794_2 = {s3671[0]};
    Full_Adder FA_3794(s3794, c3794, in3794_1, in3794_2, s3550[0]);
    wire[0:0] s3795, in3795_1, in3795_2;
    wire c3795;
    assign in3795_1 = {c3671};
    assign in3795_2 = {s3672[0]};
    Full_Adder FA_3795(s3795, c3795, in3795_1, in3795_2, s3551[0]);
    wire[0:0] s3796, in3796_1, in3796_2;
    wire c3796;
    assign in3796_1 = {c3672};
    assign in3796_2 = {s3673[0]};
    Full_Adder FA_3796(s3796, c3796, in3796_1, in3796_2, s3552[0]);
    wire[0:0] s3797, in3797_1, in3797_2;
    wire c3797;
    assign in3797_1 = {c3673};
    assign in3797_2 = {s3674[0]};
    Full_Adder FA_3797(s3797, c3797, in3797_1, in3797_2, s3553[0]);
    wire[0:0] s3798, in3798_1, in3798_2;
    wire c3798;
    assign in3798_1 = {c3674};
    assign in3798_2 = {s3675[0]};
    Full_Adder FA_3798(s3798, c3798, in3798_1, in3798_2, s3554[0]);
    wire[0:0] s3799, in3799_1, in3799_2;
    wire c3799;
    assign in3799_1 = {c3675};
    assign in3799_2 = {s3676[0]};
    Full_Adder FA_3799(s3799, c3799, in3799_1, in3799_2, s3555[0]);
    wire[0:0] s3800, in3800_1, in3800_2;
    wire c3800;
    assign in3800_1 = {c3676};
    assign in3800_2 = {s3677[0]};
    Full_Adder FA_3800(s3800, c3800, in3800_1, in3800_2, s3556[0]);
    wire[0:0] s3801, in3801_1, in3801_2;
    wire c3801;
    assign in3801_1 = {c3677};
    assign in3801_2 = {s3678[0]};
    Full_Adder FA_3801(s3801, c3801, in3801_1, in3801_2, s3557[0]);
    wire[0:0] s3802, in3802_1, in3802_2;
    wire c3802;
    assign in3802_1 = {c3678};
    assign in3802_2 = {s3679[0]};
    Full_Adder FA_3802(s3802, c3802, in3802_1, in3802_2, s3558[0]);
    wire[0:0] s3803, in3803_1, in3803_2;
    wire c3803;
    assign in3803_1 = {c3679};
    assign in3803_2 = {s3680[0]};
    Full_Adder FA_3803(s3803, c3803, in3803_1, in3803_2, s3559[0]);
    wire[0:0] s3804, in3804_1, in3804_2;
    wire c3804;
    assign in3804_1 = {c3680};
    assign in3804_2 = {s3681[0]};
    Full_Adder FA_3804(s3804, c3804, in3804_1, in3804_2, s3560[0]);
    wire[0:0] s3805, in3805_1, in3805_2;
    wire c3805;
    assign in3805_1 = {c3681};
    assign in3805_2 = {s3682[0]};
    Full_Adder FA_3805(s3805, c3805, in3805_1, in3805_2, s3561[0]);
    wire[0:0] s3806, in3806_1, in3806_2;
    wire c3806;
    assign in3806_1 = {c3682};
    assign in3806_2 = {s3683[0]};
    Full_Adder FA_3806(s3806, c3806, in3806_1, in3806_2, s3562[0]);
    wire[0:0] s3807, in3807_1, in3807_2;
    wire c3807;
    assign in3807_1 = {c3683};
    assign in3807_2 = {s3684[0]};
    Full_Adder FA_3807(s3807, c3807, in3807_1, in3807_2, s3563[0]);
    wire[0:0] s3808, in3808_1, in3808_2;
    wire c3808;
    assign in3808_1 = {c3684};
    assign in3808_2 = {s3685[0]};
    Full_Adder FA_3808(s3808, c3808, in3808_1, in3808_2, s3564[0]);
    wire[0:0] s3809, in3809_1, in3809_2;
    wire c3809;
    assign in3809_1 = {c3685};
    assign in3809_2 = {s3686[0]};
    Full_Adder FA_3809(s3809, c3809, in3809_1, in3809_2, s3565[0]);
    wire[0:0] s3810, in3810_1, in3810_2;
    wire c3810;
    assign in3810_1 = {c3686};
    assign in3810_2 = {s3687[0]};
    Full_Adder FA_3810(s3810, c3810, in3810_1, in3810_2, s3566[0]);
    wire[0:0] s3811, in3811_1, in3811_2;
    wire c3811;
    assign in3811_1 = {c3687};
    assign in3811_2 = {s3688[0]};
    Full_Adder FA_3811(s3811, c3811, in3811_1, in3811_2, s3567[0]);
    wire[0:0] s3812, in3812_1, in3812_2;
    wire c3812;
    assign in3812_1 = {c3688};
    assign in3812_2 = {s3689[0]};
    Full_Adder FA_3812(s3812, c3812, in3812_1, in3812_2, s3568[0]);
    wire[0:0] s3813, in3813_1, in3813_2;
    wire c3813;
    assign in3813_1 = {c3689};
    assign in3813_2 = {s3690[0]};
    Full_Adder FA_3813(s3813, c3813, in3813_1, in3813_2, s3569[0]);
    wire[0:0] s3814, in3814_1, in3814_2;
    wire c3814;
    assign in3814_1 = {c3690};
    assign in3814_2 = {s3691[0]};
    Full_Adder FA_3814(s3814, c3814, in3814_1, in3814_2, s3570[0]);
    wire[0:0] s3815, in3815_1, in3815_2;
    wire c3815;
    assign in3815_1 = {c3691};
    assign in3815_2 = {s3692[0]};
    Full_Adder FA_3815(s3815, c3815, in3815_1, in3815_2, s3571[0]);
    wire[0:0] s3816, in3816_1, in3816_2;
    wire c3816;
    assign in3816_1 = {c3692};
    assign in3816_2 = {s3693[0]};
    Full_Adder FA_3816(s3816, c3816, in3816_1, in3816_2, s3572[0]);
    wire[0:0] s3817, in3817_1, in3817_2;
    wire c3817;
    assign in3817_1 = {c3693};
    assign in3817_2 = {s3694[0]};
    Full_Adder FA_3817(s3817, c3817, in3817_1, in3817_2, s3573[0]);
    wire[0:0] s3818, in3818_1, in3818_2;
    wire c3818;
    assign in3818_1 = {c3694};
    assign in3818_2 = {s3695[0]};
    Full_Adder FA_3818(s3818, c3818, in3818_1, in3818_2, s3574[0]);
    wire[0:0] s3819, in3819_1, in3819_2;
    wire c3819;
    assign in3819_1 = {c3695};
    assign in3819_2 = {s3696[0]};
    Full_Adder FA_3819(s3819, c3819, in3819_1, in3819_2, s3575[0]);
    wire[0:0] s3820, in3820_1, in3820_2;
    wire c3820;
    assign in3820_1 = {c3696};
    assign in3820_2 = {s3697[0]};
    Full_Adder FA_3820(s3820, c3820, in3820_1, in3820_2, s3576[0]);
    wire[0:0] s3821, in3821_1, in3821_2;
    wire c3821;
    assign in3821_1 = {c3697};
    assign in3821_2 = {s3698[0]};
    Full_Adder FA_3821(s3821, c3821, in3821_1, in3821_2, s3577[0]);
    wire[0:0] s3822, in3822_1, in3822_2;
    wire c3822;
    assign in3822_1 = {c3698};
    assign in3822_2 = {s3699[0]};
    Full_Adder FA_3822(s3822, c3822, in3822_1, in3822_2, s3578[0]);
    wire[0:0] s3823, in3823_1, in3823_2;
    wire c3823;
    assign in3823_1 = {c3699};
    assign in3823_2 = {s3700[0]};
    Full_Adder FA_3823(s3823, c3823, in3823_1, in3823_2, s3579[0]);
    wire[0:0] s3824, in3824_1, in3824_2;
    wire c3824;
    assign in3824_1 = {c3700};
    assign in3824_2 = {s3701[0]};
    Full_Adder FA_3824(s3824, c3824, in3824_1, in3824_2, s3580[0]);
    wire[0:0] s3825, in3825_1, in3825_2;
    wire c3825;
    assign in3825_1 = {c3701};
    assign in3825_2 = {s3702[0]};
    Full_Adder FA_3825(s3825, c3825, in3825_1, in3825_2, s3581[0]);
    wire[0:0] s3826, in3826_1, in3826_2;
    wire c3826;
    assign in3826_1 = {c3702};
    assign in3826_2 = {s3703[0]};
    Full_Adder FA_3826(s3826, c3826, in3826_1, in3826_2, s3582[0]);
    wire[0:0] s3827, in3827_1, in3827_2;
    wire c3827;
    assign in3827_1 = {c3703};
    assign in3827_2 = {s3704[0]};
    Full_Adder FA_3827(s3827, c3827, in3827_1, in3827_2, s3583[0]);
    wire[0:0] s3828, in3828_1, in3828_2;
    wire c3828;
    assign in3828_1 = {c3704};
    assign in3828_2 = {s3705[0]};
    Full_Adder FA_3828(s3828, c3828, in3828_1, in3828_2, s3584[0]);
    wire[0:0] s3829, in3829_1, in3829_2;
    wire c3829;
    assign in3829_1 = {c3705};
    assign in3829_2 = {s3706[0]};
    Full_Adder FA_3829(s3829, c3829, in3829_1, in3829_2, s3585[0]);
    wire[0:0] s3830, in3830_1, in3830_2;
    wire c3830;
    assign in3830_1 = {c3706};
    assign in3830_2 = {s3707[0]};
    Full_Adder FA_3830(s3830, c3830, in3830_1, in3830_2, s3586[0]);
    wire[0:0] s3831, in3831_1, in3831_2;
    wire c3831;
    assign in3831_1 = {c3707};
    assign in3831_2 = {s3708[0]};
    Full_Adder FA_3831(s3831, c3831, in3831_1, in3831_2, s3587[0]);
    wire[0:0] s3832, in3832_1, in3832_2;
    wire c3832;
    assign in3832_1 = {c3708};
    assign in3832_2 = {s3709[0]};
    Full_Adder FA_3832(s3832, c3832, in3832_1, in3832_2, s3588[0]);
    wire[0:0] s3833, in3833_1, in3833_2;
    wire c3833;
    assign in3833_1 = {c3709};
    assign in3833_2 = {s3710[0]};
    Full_Adder FA_3833(s3833, c3833, in3833_1, in3833_2, s3589[0]);
    wire[0:0] s3834, in3834_1, in3834_2;
    wire c3834;
    assign in3834_1 = {c3710};
    assign in3834_2 = {s3711[0]};
    Full_Adder FA_3834(s3834, c3834, in3834_1, in3834_2, s3590[0]);
    wire[0:0] s3835, in3835_1, in3835_2;
    wire c3835;
    assign in3835_1 = {c3711};
    assign in3835_2 = {s3712[0]};
    Full_Adder FA_3835(s3835, c3835, in3835_1, in3835_2, s3591[0]);
    wire[0:0] s3836, in3836_1, in3836_2;
    wire c3836;
    assign in3836_1 = {c3712};
    assign in3836_2 = {s3713[0]};
    Full_Adder FA_3836(s3836, c3836, in3836_1, in3836_2, s3592[0]);
    wire[0:0] s3837, in3837_1, in3837_2;
    wire c3837;
    assign in3837_1 = {c3713};
    assign in3837_2 = {s3714[0]};
    Full_Adder FA_3837(s3837, c3837, in3837_1, in3837_2, s3593[0]);
    wire[0:0] s3838, in3838_1, in3838_2;
    wire c3838;
    assign in3838_1 = {c3714};
    assign in3838_2 = {s3715[0]};
    Full_Adder FA_3838(s3838, c3838, in3838_1, in3838_2, s3594[0]);
    wire[0:0] s3839, in3839_1, in3839_2;
    wire c3839;
    assign in3839_1 = {c3715};
    assign in3839_2 = {s3716[0]};
    Full_Adder FA_3839(s3839, c3839, in3839_1, in3839_2, s3595[0]);
    wire[0:0] s3840, in3840_1, in3840_2;
    wire c3840;
    assign in3840_1 = {c3716};
    assign in3840_2 = {s3717[0]};
    Full_Adder FA_3840(s3840, c3840, in3840_1, in3840_2, s3596[0]);
    wire[0:0] s3841, in3841_1, in3841_2;
    wire c3841;
    assign in3841_1 = {c3717};
    assign in3841_2 = {s3718[0]};
    Full_Adder FA_3841(s3841, c3841, in3841_1, in3841_2, s3597[0]);
    wire[0:0] s3842, in3842_1, in3842_2;
    wire c3842;
    assign in3842_1 = {c3718};
    assign in3842_2 = {s3719[0]};
    Full_Adder FA_3842(s3842, c3842, in3842_1, in3842_2, s3598[0]);
    wire[0:0] s3843, in3843_1, in3843_2;
    wire c3843;
    assign in3843_1 = {c3719};
    assign in3843_2 = {s3720[0]};
    Full_Adder FA_3843(s3843, c3843, in3843_1, in3843_2, s3599[0]);
    wire[0:0] s3844, in3844_1, in3844_2;
    wire c3844;
    assign in3844_1 = {c3720};
    assign in3844_2 = {s3721[0]};
    Full_Adder FA_3844(s3844, c3844, in3844_1, in3844_2, s3600[0]);
    wire[0:0] s3845, in3845_1, in3845_2;
    wire c3845;
    assign in3845_1 = {c3721};
    assign in3845_2 = {s3722[0]};
    Full_Adder FA_3845(s3845, c3845, in3845_1, in3845_2, s3601[0]);
    wire[0:0] s3846, in3846_1, in3846_2;
    wire c3846;
    assign in3846_1 = {c3722};
    assign in3846_2 = {s3723[0]};
    Full_Adder FA_3846(s3846, c3846, in3846_1, in3846_2, s3602[0]);
    wire[0:0] s3847, in3847_1, in3847_2;
    wire c3847;
    assign in3847_1 = {c3723};
    assign in3847_2 = {s3724[0]};
    Full_Adder FA_3847(s3847, c3847, in3847_1, in3847_2, s3603[0]);
    wire[0:0] s3848, in3848_1, in3848_2;
    wire c3848;
    assign in3848_1 = {c3724};
    assign in3848_2 = {s3725[0]};
    Full_Adder FA_3848(s3848, c3848, in3848_1, in3848_2, s3604[0]);
    wire[0:0] s3849, in3849_1, in3849_2;
    wire c3849;
    assign in3849_1 = {c3725};
    assign in3849_2 = {s3726[0]};
    Full_Adder FA_3849(s3849, c3849, in3849_1, in3849_2, s3605[0]);
    wire[0:0] s3850, in3850_1, in3850_2;
    wire c3850;
    assign in3850_1 = {c3726};
    assign in3850_2 = {s3727[0]};
    Full_Adder FA_3850(s3850, c3850, in3850_1, in3850_2, s3606[0]);
    wire[0:0] s3851, in3851_1, in3851_2;
    wire c3851;
    assign in3851_1 = {c3727};
    assign in3851_2 = {s3728[0]};
    Full_Adder FA_3851(s3851, c3851, in3851_1, in3851_2, s3607[0]);
    wire[0:0] s3852, in3852_1, in3852_2;
    wire c3852;
    assign in3852_1 = {c3728};
    assign in3852_2 = {s3729[0]};
    Full_Adder FA_3852(s3852, c3852, in3852_1, in3852_2, s3608[0]);
    wire[0:0] s3853, in3853_1, in3853_2;
    wire c3853;
    assign in3853_1 = {c3729};
    assign in3853_2 = {s3730[0]};
    Full_Adder FA_3853(s3853, c3853, in3853_1, in3853_2, s3609[0]);
    wire[0:0] s3854, in3854_1, in3854_2;
    wire c3854;
    assign in3854_1 = {c3730};
    assign in3854_2 = {s3731[0]};
    Full_Adder FA_3854(s3854, c3854, in3854_1, in3854_2, s3610[0]);
    wire[0:0] s3855, in3855_1, in3855_2;
    wire c3855;
    assign in3855_1 = {c3731};
    assign in3855_2 = {s3732[0]};
    Full_Adder FA_3855(s3855, c3855, in3855_1, in3855_2, s3611[0]);
    wire[0:0] s3856, in3856_1, in3856_2;
    wire c3856;
    assign in3856_1 = {c3732};
    assign in3856_2 = {s3733[0]};
    Full_Adder FA_3856(s3856, c3856, in3856_1, in3856_2, s3612[0]);
    wire[0:0] s3857, in3857_1, in3857_2;
    wire c3857;
    assign in3857_1 = {c3733};
    assign in3857_2 = {s3734[0]};
    Full_Adder FA_3857(s3857, c3857, in3857_1, in3857_2, s3613[0]);
    wire[0:0] s3858, in3858_1, in3858_2;
    wire c3858;
    assign in3858_1 = {c3734};
    assign in3858_2 = {s3735[0]};
    Full_Adder FA_3858(s3858, c3858, in3858_1, in3858_2, s3614[0]);
    wire[0:0] s3859, in3859_1, in3859_2;
    wire c3859;
    assign in3859_1 = {c3735};
    assign in3859_2 = {s3736[0]};
    Full_Adder FA_3859(s3859, c3859, in3859_1, in3859_2, s3615[0]);
    wire[0:0] s3860, in3860_1, in3860_2;
    wire c3860;
    assign in3860_1 = {c3736};
    assign in3860_2 = {s3737[0]};
    Full_Adder FA_3860(s3860, c3860, in3860_1, in3860_2, s3616[0]);
    wire[0:0] s3861, in3861_1, in3861_2;
    wire c3861;
    assign in3861_1 = {c3737};
    assign in3861_2 = {s3738[0]};
    Full_Adder FA_3861(s3861, c3861, in3861_1, in3861_2, s3617[0]);
    wire[0:0] s3862, in3862_1, in3862_2;
    wire c3862;
    assign in3862_1 = {c3738};
    assign in3862_2 = {s3739[0]};
    Full_Adder FA_3862(s3862, c3862, in3862_1, in3862_2, s3618[0]);
    wire[0:0] s3863, in3863_1, in3863_2;
    wire c3863;
    assign in3863_1 = {c3739};
    assign in3863_2 = {s3740[0]};
    Full_Adder FA_3863(s3863, c3863, in3863_1, in3863_2, s3619[0]);
    wire[0:0] s3864, in3864_1, in3864_2;
    wire c3864;
    assign in3864_1 = {c3740};
    assign in3864_2 = {s3741[0]};
    Full_Adder FA_3864(s3864, c3864, in3864_1, in3864_2, s3620[0]);
    wire[0:0] s3865, in3865_1, in3865_2;
    wire c3865;
    assign in3865_1 = {c3741};
    assign in3865_2 = {s3742[0]};
    Full_Adder FA_3865(s3865, c3865, in3865_1, in3865_2, s3621[0]);
    wire[0:0] s3866, in3866_1, in3866_2;
    wire c3866;
    assign in3866_1 = {c3742};
    assign in3866_2 = {s3743[0]};
    Full_Adder FA_3866(s3866, c3866, in3866_1, in3866_2, s3622[0]);
    wire[0:0] s3867, in3867_1, in3867_2;
    wire c3867;
    assign in3867_1 = {c3743};
    assign in3867_2 = {s3744[0]};
    Full_Adder FA_3867(s3867, c3867, in3867_1, in3867_2, s3623[0]);
    wire[0:0] s3868, in3868_1, in3868_2;
    wire c3868;
    assign in3868_1 = {c3744};
    assign in3868_2 = {s3745[0]};
    Full_Adder FA_3868(s3868, c3868, in3868_1, in3868_2, s3624[0]);
    wire[0:0] s3869, in3869_1, in3869_2;
    wire c3869;
    assign in3869_1 = {c3745};
    assign in3869_2 = {s3746[0]};
    Full_Adder FA_3869(s3869, c3869, in3869_1, in3869_2, s3625[0]);
    wire[0:0] s3870, in3870_1, in3870_2;
    wire c3870;
    assign in3870_1 = {c3746};
    assign in3870_2 = {s3747[0]};
    Full_Adder FA_3870(s3870, c3870, in3870_1, in3870_2, s3626[0]);
    wire[0:0] s3871, in3871_1, in3871_2;
    wire c3871;
    assign in3871_1 = {c3747};
    assign in3871_2 = {s3748[0]};
    Full_Adder FA_3871(s3871, c3871, in3871_1, in3871_2, s3627[0]);
    wire[0:0] s3872, in3872_1, in3872_2;
    wire c3872;
    assign in3872_1 = {c3748};
    assign in3872_2 = {s3749[0]};
    Full_Adder FA_3872(s3872, c3872, in3872_1, in3872_2, s3628[0]);
    wire[0:0] s3873, in3873_1, in3873_2;
    wire c3873;
    assign in3873_1 = {c3749};
    assign in3873_2 = {s3750[0]};
    Full_Adder FA_3873(s3873, c3873, in3873_1, in3873_2, s3629[0]);
    wire[0:0] s3874, in3874_1, in3874_2;
    wire c3874;
    assign in3874_1 = {c3750};
    assign in3874_2 = {s3751[0]};
    Full_Adder FA_3874(s3874, c3874, in3874_1, in3874_2, s3630[0]);
    wire[0:0] s3875, in3875_1, in3875_2;
    wire c3875;
    assign in3875_1 = {c3751};
    assign in3875_2 = {s3752[0]};
    Full_Adder FA_3875(s3875, c3875, in3875_1, in3875_2, s3631[0]);
    wire[0:0] s3876, in3876_1, in3876_2;
    wire c3876;
    assign in3876_1 = {c3752};
    assign in3876_2 = {s3753[0]};
    Full_Adder FA_3876(s3876, c3876, in3876_1, in3876_2, s3632[0]);
    wire[0:0] s3877, in3877_1, in3877_2;
    wire c3877;
    assign in3877_1 = {c3753};
    assign in3877_2 = {s3754[0]};
    Full_Adder FA_3877(s3877, c3877, in3877_1, in3877_2, s3633[0]);
    wire[0:0] s3878, in3878_1, in3878_2;
    wire c3878;
    assign in3878_1 = {c3754};
    assign in3878_2 = {s3755[0]};
    Full_Adder FA_3878(s3878, c3878, in3878_1, in3878_2, s3634[0]);
    wire[0:0] s3879, in3879_1, in3879_2;
    wire c3879;
    assign in3879_1 = {c3755};
    assign in3879_2 = {s3756[0]};
    Full_Adder FA_3879(s3879, c3879, in3879_1, in3879_2, s3635[0]);
    wire[0:0] s3880, in3880_1, in3880_2;
    wire c3880;
    assign in3880_1 = {c3756};
    assign in3880_2 = {s3757[0]};
    Full_Adder FA_3880(s3880, c3880, in3880_1, in3880_2, s3636[0]);
    wire[0:0] s3881, in3881_1, in3881_2;
    wire c3881;
    assign in3881_1 = {c3757};
    assign in3881_2 = {s3758[0]};
    Full_Adder FA_3881(s3881, c3881, in3881_1, in3881_2, s3637[0]);
    wire[0:0] s3882, in3882_1, in3882_2;
    wire c3882;
    assign in3882_1 = {c3758};
    assign in3882_2 = {s3759[0]};
    Full_Adder FA_3882(s3882, c3882, in3882_1, in3882_2, s3638[0]);
    wire[0:0] s3883, in3883_1, in3883_2;
    wire c3883;
    assign in3883_1 = {c3759};
    assign in3883_2 = {s3760[0]};
    Full_Adder FA_3883(s3883, c3883, in3883_1, in3883_2, s3639[0]);
    wire[0:0] s3884, in3884_1, in3884_2;
    wire c3884;
    assign in3884_1 = {c3760};
    assign in3884_2 = {s3761[0]};
    Full_Adder FA_3884(s3884, c3884, in3884_1, in3884_2, s3640[0]);
    wire[0:0] s3885, in3885_1, in3885_2;
    wire c3885;
    assign in3885_1 = {c3761};
    assign in3885_2 = {s3762[0]};
    Full_Adder FA_3885(s3885, c3885, in3885_1, in3885_2, s3641[0]);
    wire[0:0] s3886, in3886_1, in3886_2;
    wire c3886;
    assign in3886_1 = {c3762};
    assign in3886_2 = {s3763[0]};
    Full_Adder FA_3886(s3886, c3886, in3886_1, in3886_2, s3642[0]);
    wire[0:0] s3887, in3887_1, in3887_2;
    wire c3887;
    assign in3887_1 = {c3763};
    assign in3887_2 = {s3764[0]};
    Full_Adder FA_3887(s3887, c3887, in3887_1, in3887_2, s3643[0]);
    wire[0:0] s3888, in3888_1, in3888_2;
    wire c3888;
    assign in3888_1 = {c3764};
    assign in3888_2 = {s3765[0]};
    Full_Adder FA_3888(s3888, c3888, in3888_1, in3888_2, s3644[0]);
    wire[0:0] s3889, in3889_1, in3889_2;
    wire c3889;
    assign in3889_1 = {c3765};
    assign in3889_2 = {s3766[0]};
    Full_Adder FA_3889(s3889, c3889, in3889_1, in3889_2, s3645[0]);
    wire[0:0] s3890, in3890_1, in3890_2;
    wire c3890;
    assign in3890_1 = {c3766};
    assign in3890_2 = {s3767[0]};
    Full_Adder FA_3890(s3890, c3890, in3890_1, in3890_2, s3646[0]);
    wire[0:0] s3891, in3891_1, in3891_2;
    wire c3891;
    assign in3891_1 = {c3767};
    assign in3891_2 = {s3768[0]};
    Full_Adder FA_3891(s3891, c3891, in3891_1, in3891_2, s3647[0]);
    wire[0:0] s3892, in3892_1, in3892_2;
    wire c3892;
    assign in3892_1 = {c3768};
    assign in3892_2 = {s3769[0]};
    Full_Adder FA_3892(s3892, c3892, in3892_1, in3892_2, s3648[0]);
    wire[0:0] s3893, in3893_1, in3893_2;
    wire c3893;
    assign in3893_1 = {c3769};
    assign in3893_2 = {s3770[0]};
    Full_Adder FA_3893(s3893, c3893, in3893_1, in3893_2, s3649[0]);
    wire[0:0] s3894, in3894_1, in3894_2;
    wire c3894;
    assign in3894_1 = {c3770};
    assign in3894_2 = {s3771[0]};
    Full_Adder FA_3894(s3894, c3894, in3894_1, in3894_2, s3650[0]);
    wire[0:0] s3895, in3895_1, in3895_2;
    wire c3895;
    assign in3895_1 = {c3771};
    assign in3895_2 = {s3772[0]};
    Full_Adder FA_3895(s3895, c3895, in3895_1, in3895_2, s3651[0]);
    wire[0:0] s3896, in3896_1, in3896_2;
    wire c3896;
    assign in3896_1 = {c3772};
    assign in3896_2 = {s3773[0]};
    Full_Adder FA_3896(s3896, c3896, in3896_1, in3896_2, s3652[0]);
    wire[0:0] s3897, in3897_1, in3897_2;
    wire c3897;
    assign in3897_1 = {c3773};
    assign in3897_2 = {s3774[0]};
    Full_Adder FA_3897(s3897, c3897, in3897_1, in3897_2, s3653[0]);
    wire[0:0] s3898, in3898_1, in3898_2;
    wire c3898;
    assign in3898_1 = {c3774};
    assign in3898_2 = {s3775[0]};
    Full_Adder FA_3898(s3898, c3898, in3898_1, in3898_2, s3654[0]);
    wire[0:0] s3899, in3899_1, in3899_2;
    wire c3899;
    assign in3899_1 = {c3775};
    assign in3899_2 = {s3776[0]};
    Full_Adder FA_3899(s3899, c3899, in3899_1, in3899_2, s3655[0]);
    wire[0:0] s3900, in3900_1, in3900_2;
    wire c3900;
    assign in3900_1 = {c3776};
    assign in3900_2 = {s3777[0]};
    Full_Adder FA_3900(s3900, c3900, in3900_1, in3900_2, s3656[0]);
    wire[0:0] s3901, in3901_1, in3901_2;
    wire c3901;
    assign in3901_1 = {c3777};
    assign in3901_2 = {s3778[0]};
    Full_Adder FA_3901(s3901, c3901, in3901_1, in3901_2, s3657[0]);
    wire[0:0] s3902, in3902_1, in3902_2;
    wire c3902;
    assign in3902_1 = {c3778};
    assign in3902_2 = {s3779[0]};
    Full_Adder FA_3902(s3902, c3902, in3902_1, in3902_2, s3658[0]);
    wire[0:0] s3903, in3903_1, in3903_2;
    wire c3903;
    assign in3903_1 = {c3779};
    assign in3903_2 = {s3780[0]};
    Full_Adder FA_3903(s3903, c3903, in3903_1, in3903_2, s3659[0]);
    wire[0:0] s3904, in3904_1, in3904_2;
    wire c3904;
    assign in3904_1 = {c3780};
    assign in3904_2 = {s3781[0]};
    Full_Adder FA_3904(s3904, c3904, in3904_1, in3904_2, s3660[0]);
    wire[0:0] s3905, in3905_1, in3905_2;
    wire c3905;
    assign in3905_1 = {c3781};
    assign in3905_2 = {s3782[0]};
    Full_Adder FA_3905(s3905, c3905, in3905_1, in3905_2, c3660);
    wire[0:0] s3906, in3906_1, in3906_2;
    wire c3906;
    assign in3906_1 = {pp63[62]};
    assign in3906_2 = {c3782};
    Full_Adder FA_3906(s3906, c3906, in3906_1, in3906_2, pp62[63]);


    /*Final Stage 10*/
    wire[125:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],c3783,c3784,c3785,c3786,c3787,c3788,c3789,c3790,c3791,c3792,c3793,c3794,c3795,c3796,c3797,c3798,c3799,c3800,c3801,c3802,c3803,c3804,c3805,c3806,c3807,c3808,c3809,c3810,c3811,c3812,c3813,c3814,c3815,c3816,c3817,c3818,c3819,c3820,c3821,c3822,c3823,c3824,c3825,c3826,c3827,c3828,c3829,c3830,c3831,c3832,c3833,c3834,c3835,c3836,c3837,c3838,c3839,c3840,c3841,c3842,c3843,c3844,c3845,c3846,c3847,c3848,c3849,c3850,c3851,c3852,c3853,c3854,c3855,c3856,c3857,c3858,c3859,c3860,c3861,c3862,c3863,c3864,c3865,c3866,c3867,c3868,c3869,c3870,c3871,c3872,c3873,c3874,c3875,c3876,c3877,c3878,c3879,c3880,c3881,c3882,c3883,c3884,c3885,c3886,c3887,c3888,c3889,c3890,c3891,c3892,c3893,c3894,c3895,c3896,c3897,c3898,c3899,c3900,c3901,c3902,c3903,c3904,c3905,pp63[63]};
    assign in_2 = {pp1[0],s3783[0],s3784[0],s3785[0],s3786[0],s3787[0],s3788[0],s3789[0],s3790[0],s3791[0],s3792[0],s3793[0],s3794[0],s3795[0],s3796[0],s3797[0],s3798[0],s3799[0],s3800[0],s3801[0],s3802[0],s3803[0],s3804[0],s3805[0],s3806[0],s3807[0],s3808[0],s3809[0],s3810[0],s3811[0],s3812[0],s3813[0],s3814[0],s3815[0],s3816[0],s3817[0],s3818[0],s3819[0],s3820[0],s3821[0],s3822[0],s3823[0],s3824[0],s3825[0],s3826[0],s3827[0],s3828[0],s3829[0],s3830[0],s3831[0],s3832[0],s3833[0],s3834[0],s3835[0],s3836[0],s3837[0],s3838[0],s3839[0],s3840[0],s3841[0],s3842[0],s3843[0],s3844[0],s3845[0],s3846[0],s3847[0],s3848[0],s3849[0],s3850[0],s3851[0],s3852[0],s3853[0],s3854[0],s3855[0],s3856[0],s3857[0],s3858[0],s3859[0],s3860[0],s3861[0],s3862[0],s3863[0],s3864[0],s3865[0],s3866[0],s3867[0],s3868[0],s3869[0],s3870[0],s3871[0],s3872[0],s3873[0],s3874[0],s3875[0],s3876[0],s3877[0],s3878[0],s3879[0],s3880[0],s3881[0],s3882[0],s3883[0],s3884[0],s3885[0],s3886[0],s3887[0],s3888[0],s3889[0],s3890[0],s3891[0],s3892[0],s3893[0],s3894[0],s3895[0],s3896[0],s3897[0],s3898[0],s3899[0],s3900[0],s3901[0],s3902[0],s3903[0],s3904[0],s3905[0],s3906[0],c3906};
    CLA_126(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = c;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule

module CLA_126(output [125:0] sum, output cout, input [125:0] in1, input [125:0] in2);

    wire[125:0] G;
    wire[125:0] C;
    wire[125:0] P;

    assign G[0] = in1[125] & in2[125];
    assign P[0] = in1[125] ^ in2[125];
    assign G[1] = in1[124] & in2[124];
    assign P[1] = in1[124] ^ in2[124];
    assign G[2] = in1[123] & in2[123];
    assign P[2] = in1[123] ^ in2[123];
    assign G[3] = in1[122] & in2[122];
    assign P[3] = in1[122] ^ in2[122];
    assign G[4] = in1[121] & in2[121];
    assign P[4] = in1[121] ^ in2[121];
    assign G[5] = in1[120] & in2[120];
    assign P[5] = in1[120] ^ in2[120];
    assign G[6] = in1[119] & in2[119];
    assign P[6] = in1[119] ^ in2[119];
    assign G[7] = in1[118] & in2[118];
    assign P[7] = in1[118] ^ in2[118];
    assign G[8] = in1[117] & in2[117];
    assign P[8] = in1[117] ^ in2[117];
    assign G[9] = in1[116] & in2[116];
    assign P[9] = in1[116] ^ in2[116];
    assign G[10] = in1[115] & in2[115];
    assign P[10] = in1[115] ^ in2[115];
    assign G[11] = in1[114] & in2[114];
    assign P[11] = in1[114] ^ in2[114];
    assign G[12] = in1[113] & in2[113];
    assign P[12] = in1[113] ^ in2[113];
    assign G[13] = in1[112] & in2[112];
    assign P[13] = in1[112] ^ in2[112];
    assign G[14] = in1[111] & in2[111];
    assign P[14] = in1[111] ^ in2[111];
    assign G[15] = in1[110] & in2[110];
    assign P[15] = in1[110] ^ in2[110];
    assign G[16] = in1[109] & in2[109];
    assign P[16] = in1[109] ^ in2[109];
    assign G[17] = in1[108] & in2[108];
    assign P[17] = in1[108] ^ in2[108];
    assign G[18] = in1[107] & in2[107];
    assign P[18] = in1[107] ^ in2[107];
    assign G[19] = in1[106] & in2[106];
    assign P[19] = in1[106] ^ in2[106];
    assign G[20] = in1[105] & in2[105];
    assign P[20] = in1[105] ^ in2[105];
    assign G[21] = in1[104] & in2[104];
    assign P[21] = in1[104] ^ in2[104];
    assign G[22] = in1[103] & in2[103];
    assign P[22] = in1[103] ^ in2[103];
    assign G[23] = in1[102] & in2[102];
    assign P[23] = in1[102] ^ in2[102];
    assign G[24] = in1[101] & in2[101];
    assign P[24] = in1[101] ^ in2[101];
    assign G[25] = in1[100] & in2[100];
    assign P[25] = in1[100] ^ in2[100];
    assign G[26] = in1[99] & in2[99];
    assign P[26] = in1[99] ^ in2[99];
    assign G[27] = in1[98] & in2[98];
    assign P[27] = in1[98] ^ in2[98];
    assign G[28] = in1[97] & in2[97];
    assign P[28] = in1[97] ^ in2[97];
    assign G[29] = in1[96] & in2[96];
    assign P[29] = in1[96] ^ in2[96];
    assign G[30] = in1[95] & in2[95];
    assign P[30] = in1[95] ^ in2[95];
    assign G[31] = in1[94] & in2[94];
    assign P[31] = in1[94] ^ in2[94];
    assign G[32] = in1[93] & in2[93];
    assign P[32] = in1[93] ^ in2[93];
    assign G[33] = in1[92] & in2[92];
    assign P[33] = in1[92] ^ in2[92];
    assign G[34] = in1[91] & in2[91];
    assign P[34] = in1[91] ^ in2[91];
    assign G[35] = in1[90] & in2[90];
    assign P[35] = in1[90] ^ in2[90];
    assign G[36] = in1[89] & in2[89];
    assign P[36] = in1[89] ^ in2[89];
    assign G[37] = in1[88] & in2[88];
    assign P[37] = in1[88] ^ in2[88];
    assign G[38] = in1[87] & in2[87];
    assign P[38] = in1[87] ^ in2[87];
    assign G[39] = in1[86] & in2[86];
    assign P[39] = in1[86] ^ in2[86];
    assign G[40] = in1[85] & in2[85];
    assign P[40] = in1[85] ^ in2[85];
    assign G[41] = in1[84] & in2[84];
    assign P[41] = in1[84] ^ in2[84];
    assign G[42] = in1[83] & in2[83];
    assign P[42] = in1[83] ^ in2[83];
    assign G[43] = in1[82] & in2[82];
    assign P[43] = in1[82] ^ in2[82];
    assign G[44] = in1[81] & in2[81];
    assign P[44] = in1[81] ^ in2[81];
    assign G[45] = in1[80] & in2[80];
    assign P[45] = in1[80] ^ in2[80];
    assign G[46] = in1[79] & in2[79];
    assign P[46] = in1[79] ^ in2[79];
    assign G[47] = in1[78] & in2[78];
    assign P[47] = in1[78] ^ in2[78];
    assign G[48] = in1[77] & in2[77];
    assign P[48] = in1[77] ^ in2[77];
    assign G[49] = in1[76] & in2[76];
    assign P[49] = in1[76] ^ in2[76];
    assign G[50] = in1[75] & in2[75];
    assign P[50] = in1[75] ^ in2[75];
    assign G[51] = in1[74] & in2[74];
    assign P[51] = in1[74] ^ in2[74];
    assign G[52] = in1[73] & in2[73];
    assign P[52] = in1[73] ^ in2[73];
    assign G[53] = in1[72] & in2[72];
    assign P[53] = in1[72] ^ in2[72];
    assign G[54] = in1[71] & in2[71];
    assign P[54] = in1[71] ^ in2[71];
    assign G[55] = in1[70] & in2[70];
    assign P[55] = in1[70] ^ in2[70];
    assign G[56] = in1[69] & in2[69];
    assign P[56] = in1[69] ^ in2[69];
    assign G[57] = in1[68] & in2[68];
    assign P[57] = in1[68] ^ in2[68];
    assign G[58] = in1[67] & in2[67];
    assign P[58] = in1[67] ^ in2[67];
    assign G[59] = in1[66] & in2[66];
    assign P[59] = in1[66] ^ in2[66];
    assign G[60] = in1[65] & in2[65];
    assign P[60] = in1[65] ^ in2[65];
    assign G[61] = in1[64] & in2[64];
    assign P[61] = in1[64] ^ in2[64];
    assign G[62] = in1[63] & in2[63];
    assign P[62] = in1[63] ^ in2[63];
    assign G[63] = in1[62] & in2[62];
    assign P[63] = in1[62] ^ in2[62];
    assign G[64] = in1[61] & in2[61];
    assign P[64] = in1[61] ^ in2[61];
    assign G[65] = in1[60] & in2[60];
    assign P[65] = in1[60] ^ in2[60];
    assign G[66] = in1[59] & in2[59];
    assign P[66] = in1[59] ^ in2[59];
    assign G[67] = in1[58] & in2[58];
    assign P[67] = in1[58] ^ in2[58];
    assign G[68] = in1[57] & in2[57];
    assign P[68] = in1[57] ^ in2[57];
    assign G[69] = in1[56] & in2[56];
    assign P[69] = in1[56] ^ in2[56];
    assign G[70] = in1[55] & in2[55];
    assign P[70] = in1[55] ^ in2[55];
    assign G[71] = in1[54] & in2[54];
    assign P[71] = in1[54] ^ in2[54];
    assign G[72] = in1[53] & in2[53];
    assign P[72] = in1[53] ^ in2[53];
    assign G[73] = in1[52] & in2[52];
    assign P[73] = in1[52] ^ in2[52];
    assign G[74] = in1[51] & in2[51];
    assign P[74] = in1[51] ^ in2[51];
    assign G[75] = in1[50] & in2[50];
    assign P[75] = in1[50] ^ in2[50];
    assign G[76] = in1[49] & in2[49];
    assign P[76] = in1[49] ^ in2[49];
    assign G[77] = in1[48] & in2[48];
    assign P[77] = in1[48] ^ in2[48];
    assign G[78] = in1[47] & in2[47];
    assign P[78] = in1[47] ^ in2[47];
    assign G[79] = in1[46] & in2[46];
    assign P[79] = in1[46] ^ in2[46];
    assign G[80] = in1[45] & in2[45];
    assign P[80] = in1[45] ^ in2[45];
    assign G[81] = in1[44] & in2[44];
    assign P[81] = in1[44] ^ in2[44];
    assign G[82] = in1[43] & in2[43];
    assign P[82] = in1[43] ^ in2[43];
    assign G[83] = in1[42] & in2[42];
    assign P[83] = in1[42] ^ in2[42];
    assign G[84] = in1[41] & in2[41];
    assign P[84] = in1[41] ^ in2[41];
    assign G[85] = in1[40] & in2[40];
    assign P[85] = in1[40] ^ in2[40];
    assign G[86] = in1[39] & in2[39];
    assign P[86] = in1[39] ^ in2[39];
    assign G[87] = in1[38] & in2[38];
    assign P[87] = in1[38] ^ in2[38];
    assign G[88] = in1[37] & in2[37];
    assign P[88] = in1[37] ^ in2[37];
    assign G[89] = in1[36] & in2[36];
    assign P[89] = in1[36] ^ in2[36];
    assign G[90] = in1[35] & in2[35];
    assign P[90] = in1[35] ^ in2[35];
    assign G[91] = in1[34] & in2[34];
    assign P[91] = in1[34] ^ in2[34];
    assign G[92] = in1[33] & in2[33];
    assign P[92] = in1[33] ^ in2[33];
    assign G[93] = in1[32] & in2[32];
    assign P[93] = in1[32] ^ in2[32];
    assign G[94] = in1[31] & in2[31];
    assign P[94] = in1[31] ^ in2[31];
    assign G[95] = in1[30] & in2[30];
    assign P[95] = in1[30] ^ in2[30];
    assign G[96] = in1[29] & in2[29];
    assign P[96] = in1[29] ^ in2[29];
    assign G[97] = in1[28] & in2[28];
    assign P[97] = in1[28] ^ in2[28];
    assign G[98] = in1[27] & in2[27];
    assign P[98] = in1[27] ^ in2[27];
    assign G[99] = in1[26] & in2[26];
    assign P[99] = in1[26] ^ in2[26];
    assign G[100] = in1[25] & in2[25];
    assign P[100] = in1[25] ^ in2[25];
    assign G[101] = in1[24] & in2[24];
    assign P[101] = in1[24] ^ in2[24];
    assign G[102] = in1[23] & in2[23];
    assign P[102] = in1[23] ^ in2[23];
    assign G[103] = in1[22] & in2[22];
    assign P[103] = in1[22] ^ in2[22];
    assign G[104] = in1[21] & in2[21];
    assign P[104] = in1[21] ^ in2[21];
    assign G[105] = in1[20] & in2[20];
    assign P[105] = in1[20] ^ in2[20];
    assign G[106] = in1[19] & in2[19];
    assign P[106] = in1[19] ^ in2[19];
    assign G[107] = in1[18] & in2[18];
    assign P[107] = in1[18] ^ in2[18];
    assign G[108] = in1[17] & in2[17];
    assign P[108] = in1[17] ^ in2[17];
    assign G[109] = in1[16] & in2[16];
    assign P[109] = in1[16] ^ in2[16];
    assign G[110] = in1[15] & in2[15];
    assign P[110] = in1[15] ^ in2[15];
    assign G[111] = in1[14] & in2[14];
    assign P[111] = in1[14] ^ in2[14];
    assign G[112] = in1[13] & in2[13];
    assign P[112] = in1[13] ^ in2[13];
    assign G[113] = in1[12] & in2[12];
    assign P[113] = in1[12] ^ in2[12];
    assign G[114] = in1[11] & in2[11];
    assign P[114] = in1[11] ^ in2[11];
    assign G[115] = in1[10] & in2[10];
    assign P[115] = in1[10] ^ in2[10];
    assign G[116] = in1[9] & in2[9];
    assign P[116] = in1[9] ^ in2[9];
    assign G[117] = in1[8] & in2[8];
    assign P[117] = in1[8] ^ in2[8];
    assign G[118] = in1[7] & in2[7];
    assign P[118] = in1[7] ^ in2[7];
    assign G[119] = in1[6] & in2[6];
    assign P[119] = in1[6] ^ in2[6];
    assign G[120] = in1[5] & in2[5];
    assign P[120] = in1[5] ^ in2[5];
    assign G[121] = in1[4] & in2[4];
    assign P[121] = in1[4] ^ in2[4];
    assign G[122] = in1[3] & in2[3];
    assign P[122] = in1[3] ^ in2[3];
    assign G[123] = in1[2] & in2[2];
    assign P[123] = in1[2] ^ in2[2];
    assign G[124] = in1[1] & in2[1];
    assign P[124] = in1[1] ^ in2[1];
    assign G[125] = in1[0] & in2[0];
    assign P[125] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign cout = G[125] | (P[125] & C[125]);
    assign sum = P ^ C;
endmodule

