module multiplier_32bits_version14(product, A, B);

    output [63:0] product;
    input [31:0] A, B;

    /*
     * Area: 19245.053832
     * Power: 15.7174mW
     * Timing: 4.19ns
     */

    wire [31:0] pp0;
    wire [31:0] pp1;
    wire [31:0] pp2;
    wire [31:0] pp3;
    wire [31:0] pp4;
    wire [31:0] pp5;
    wire [31:0] pp6;
    wire [31:0] pp7;
    wire [31:0] pp8;
    wire [31:0] pp9;
    wire [31:0] pp10;
    wire [31:0] pp11;
    wire [31:0] pp12;
    wire [31:0] pp13;
    wire [31:0] pp14;
    wire [31:0] pp15;
    wire [31:0] pp16;
    wire [31:0] pp17;
    wire [31:0] pp18;
    wire [31:0] pp19;
    wire [31:0] pp20;
    wire [31:0] pp21;
    wire [31:0] pp22;
    wire [31:0] pp23;
    wire [31:0] pp24;
    wire [31:0] pp25;
    wire [31:0] pp26;
    wire [31:0] pp27;
    wire [31:0] pp28;
    wire [31:0] pp29;
    wire [31:0] pp30;
    wire [31:0] pp31;


    assign pp0 = A[0] ? B: 32'b00000000000000000000000000000000;
    assign pp1 = A[1] ? B: 32'b00000000000000000000000000000000;
    assign pp2 = A[2] ? B: 32'b00000000000000000000000000000000;
    assign pp3 = A[3] ? B: 32'b00000000000000000000000000000000;
    assign pp4 = A[4] ? B: 32'b00000000000000000000000000000000;
    assign pp5 = A[5] ? B: 32'b00000000000000000000000000000000;
    assign pp6 = A[6] ? B: 32'b00000000000000000000000000000000;
    assign pp7 = A[7] ? B: 32'b00000000000000000000000000000000;
    assign pp8 = A[8] ? B: 32'b00000000000000000000000000000000;
    assign pp9 = A[9] ? B: 32'b00000000000000000000000000000000;
    assign pp10 = A[10] ? B: 32'b00000000000000000000000000000000;
    assign pp11 = A[11] ? B: 32'b00000000000000000000000000000000;
    assign pp12 = A[12] ? B: 32'b00000000000000000000000000000000;
    assign pp13 = A[13] ? B: 32'b00000000000000000000000000000000;
    assign pp14 = A[14] ? B: 32'b00000000000000000000000000000000;
    assign pp15 = A[15] ? B: 32'b00000000000000000000000000000000;
    assign pp16 = A[16] ? B: 32'b00000000000000000000000000000000;
    assign pp17 = A[17] ? B: 32'b00000000000000000000000000000000;
    assign pp18 = A[18] ? B: 32'b00000000000000000000000000000000;
    assign pp19 = A[19] ? B: 32'b00000000000000000000000000000000;
    assign pp20 = A[20] ? B: 32'b00000000000000000000000000000000;
    assign pp21 = A[21] ? B: 32'b00000000000000000000000000000000;
    assign pp22 = A[22] ? B: 32'b00000000000000000000000000000000;
    assign pp23 = A[23] ? B: 32'b00000000000000000000000000000000;
    assign pp24 = A[24] ? B: 32'b00000000000000000000000000000000;
    assign pp25 = A[25] ? B: 32'b00000000000000000000000000000000;
    assign pp26 = A[26] ? B: 32'b00000000000000000000000000000000;
    assign pp27 = A[27] ? B: 32'b00000000000000000000000000000000;
    assign pp28 = A[28] ? B: 32'b00000000000000000000000000000000;
    assign pp29 = A[29] ? B: 32'b00000000000000000000000000000000;
    assign pp30 = A[30] ? B: 32'b00000000000000000000000000000000;
    assign pp31 = A[31] ? B: 32'b00000000000000000000000000000000;


    /*Stage 1*/
    wire[0:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[22]};
    assign in1_2 = {pp1[21]};
    Half_Adder HA_1(s1, c1, in1_1, in1_2);
    wire[0:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp1[22]};
    assign in2_2 = {pp2[21]};
    Full_Adder FA_2(s2, c2, in2_1, in2_2, pp0[23]);
    wire[0:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp3[20]};
    assign in3_2 = {pp4[19]};
    Half_Adder HA_3(s3, c3, in3_1, in3_2);
    wire[0:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp1[23]};
    assign in4_2 = {pp2[22]};
    Full_Adder FA_4(s4, c4, in4_1, in4_2, pp0[24]);
    wire[0:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp4[20]};
    assign in5_2 = {pp5[19]};
    Full_Adder FA_5(s5, c5, in5_1, in5_2, pp3[21]);
    wire[0:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp6[18]};
    assign in6_2 = {pp7[17]};
    Half_Adder HA_6(s6, c6, in6_1, in6_2);
    wire[0:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp1[24]};
    assign in7_2 = {pp2[23]};
    Full_Adder FA_7(s7, c7, in7_1, in7_2, pp0[25]);
    wire[0:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp4[21]};
    assign in8_2 = {pp5[20]};
    Full_Adder FA_8(s8, c8, in8_1, in8_2, pp3[22]);
    wire[0:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp7[18]};
    assign in9_2 = {pp8[17]};
    Full_Adder FA_9(s9, c9, in9_1, in9_2, pp6[19]);
    wire[0:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp9[16]};
    assign in10_2 = {pp10[15]};
    Half_Adder HA_10(s10, c10, in10_1, in10_2);
    wire[0:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp1[25]};
    assign in11_2 = {pp2[24]};
    Full_Adder FA_11(s11, c11, in11_1, in11_2, pp0[26]);
    wire[0:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp4[22]};
    assign in12_2 = {pp5[21]};
    Full_Adder FA_12(s12, c12, in12_1, in12_2, pp3[23]);
    wire[0:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp7[19]};
    assign in13_2 = {pp8[18]};
    Full_Adder FA_13(s13, c13, in13_1, in13_2, pp6[20]);
    wire[0:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp10[16]};
    assign in14_2 = {pp11[15]};
    Full_Adder FA_14(s14, c14, in14_1, in14_2, pp9[17]);
    wire[0:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp12[14]};
    assign in15_2 = {pp13[13]};
    Half_Adder HA_15(s15, c15, in15_1, in15_2);
    wire[0:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp1[26]};
    assign in16_2 = {pp2[25]};
    Full_Adder FA_16(s16, c16, in16_1, in16_2, pp0[27]);
    wire[0:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp4[23]};
    assign in17_2 = {pp5[22]};
    Full_Adder FA_17(s17, c17, in17_1, in17_2, pp3[24]);
    wire[0:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp7[20]};
    assign in18_2 = {pp8[19]};
    Full_Adder FA_18(s18, c18, in18_1, in18_2, pp6[21]);
    wire[0:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp10[17]};
    assign in19_2 = {pp11[16]};
    Full_Adder FA_19(s19, c19, in19_1, in19_2, pp9[18]);
    wire[0:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp13[14]};
    assign in20_2 = {pp14[13]};
    Full_Adder FA_20(s20, c20, in20_1, in20_2, pp12[15]);
    wire[0:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp15[12]};
    assign in21_2 = {pp16[11]};
    Half_Adder HA_21(s21, c21, in21_1, in21_2);
    wire[0:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp1[27]};
    assign in22_2 = {pp2[26]};
    Full_Adder FA_22(s22, c22, in22_1, in22_2, pp0[28]);
    wire[0:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp4[24]};
    assign in23_2 = {pp5[23]};
    Full_Adder FA_23(s23, c23, in23_1, in23_2, pp3[25]);
    wire[0:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp7[21]};
    assign in24_2 = {pp8[20]};
    Full_Adder FA_24(s24, c24, in24_1, in24_2, pp6[22]);
    wire[0:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp10[18]};
    assign in25_2 = {pp11[17]};
    Full_Adder FA_25(s25, c25, in25_1, in25_2, pp9[19]);
    wire[0:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp13[15]};
    assign in26_2 = {pp14[14]};
    Full_Adder FA_26(s26, c26, in26_1, in26_2, pp12[16]);
    wire[0:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp16[12]};
    assign in27_2 = {pp17[11]};
    Full_Adder FA_27(s27, c27, in27_1, in27_2, pp15[13]);
    wire[0:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp18[10]};
    assign in28_2 = {pp19[9]};
    Half_Adder HA_28(s28, c28, in28_1, in28_2);
    wire[0:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp1[28]};
    assign in29_2 = {pp2[27]};
    Full_Adder FA_29(s29, c29, in29_1, in29_2, pp0[29]);
    wire[0:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp4[25]};
    assign in30_2 = {pp5[24]};
    Full_Adder FA_30(s30, c30, in30_1, in30_2, pp3[26]);
    wire[0:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp7[22]};
    assign in31_2 = {pp8[21]};
    Full_Adder FA_31(s31, c31, in31_1, in31_2, pp6[23]);
    wire[0:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp10[19]};
    assign in32_2 = {pp11[18]};
    Full_Adder FA_32(s32, c32, in32_1, in32_2, pp9[20]);
    wire[0:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp13[16]};
    assign in33_2 = {pp14[15]};
    Full_Adder FA_33(s33, c33, in33_1, in33_2, pp12[17]);
    wire[0:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp16[13]};
    assign in34_2 = {pp17[12]};
    Full_Adder FA_34(s34, c34, in34_1, in34_2, pp15[14]);
    wire[0:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp19[10]};
    assign in35_2 = {pp20[9]};
    Full_Adder FA_35(s35, c35, in35_1, in35_2, pp18[11]);
    wire[0:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp21[8]};
    assign in36_2 = {pp22[7]};
    Half_Adder HA_36(s36, c36, in36_1, in36_2);
    wire[0:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp1[29]};
    assign in37_2 = {pp2[28]};
    Full_Adder FA_37(s37, c37, in37_1, in37_2, pp0[30]);
    wire[0:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp4[26]};
    assign in38_2 = {pp5[25]};
    Full_Adder FA_38(s38, c38, in38_1, in38_2, pp3[27]);
    wire[0:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp7[23]};
    assign in39_2 = {pp8[22]};
    Full_Adder FA_39(s39, c39, in39_1, in39_2, pp6[24]);
    wire[0:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp10[20]};
    assign in40_2 = {pp11[19]};
    Full_Adder FA_40(s40, c40, in40_1, in40_2, pp9[21]);
    wire[0:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp13[17]};
    assign in41_2 = {pp14[16]};
    Full_Adder FA_41(s41, c41, in41_1, in41_2, pp12[18]);
    wire[0:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp16[14]};
    assign in42_2 = {pp17[13]};
    Full_Adder FA_42(s42, c42, in42_1, in42_2, pp15[15]);
    wire[0:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp19[11]};
    assign in43_2 = {pp20[10]};
    Full_Adder FA_43(s43, c43, in43_1, in43_2, pp18[12]);
    wire[0:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[8]};
    assign in44_2 = {pp23[7]};
    Full_Adder FA_44(s44, c44, in44_1, in44_2, pp21[9]);
    wire[0:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[6]};
    assign in45_2 = {pp25[5]};
    Half_Adder HA_45(s45, c45, in45_1, in45_2);
    wire[0:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp1[30]};
    assign in46_2 = {pp2[29]};
    Full_Adder FA_46(s46, c46, in46_1, in46_2, pp0[31]);
    wire[0:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp4[27]};
    assign in47_2 = {pp5[26]};
    Full_Adder FA_47(s47, c47, in47_1, in47_2, pp3[28]);
    wire[0:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp7[24]};
    assign in48_2 = {pp8[23]};
    Full_Adder FA_48(s48, c48, in48_1, in48_2, pp6[25]);
    wire[0:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp10[21]};
    assign in49_2 = {pp11[20]};
    Full_Adder FA_49(s49, c49, in49_1, in49_2, pp9[22]);
    wire[0:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp13[18]};
    assign in50_2 = {pp14[17]};
    Full_Adder FA_50(s50, c50, in50_1, in50_2, pp12[19]);
    wire[0:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp16[15]};
    assign in51_2 = {pp17[14]};
    Full_Adder FA_51(s51, c51, in51_1, in51_2, pp15[16]);
    wire[0:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp19[12]};
    assign in52_2 = {pp20[11]};
    Full_Adder FA_52(s52, c52, in52_1, in52_2, pp18[13]);
    wire[0:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp22[9]};
    assign in53_2 = {pp23[8]};
    Full_Adder FA_53(s53, c53, in53_1, in53_2, pp21[10]);
    wire[0:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp25[6]};
    assign in54_2 = {pp26[5]};
    Full_Adder FA_54(s54, c54, in54_1, in54_2, pp24[7]);
    wire[0:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp27[4]};
    assign in55_2 = {pp28[3]};
    Half_Adder HA_55(s55, c55, in55_1, in55_2);
    wire[0:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp2[30]};
    assign in56_2 = {pp3[29]};
    Full_Adder FA_56(s56, c56, in56_1, in56_2, pp1[31]);
    wire[0:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp5[27]};
    assign in57_2 = {pp6[26]};
    Full_Adder FA_57(s57, c57, in57_1, in57_2, pp4[28]);
    wire[0:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp8[24]};
    assign in58_2 = {pp9[23]};
    Full_Adder FA_58(s58, c58, in58_1, in58_2, pp7[25]);
    wire[0:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp11[21]};
    assign in59_2 = {pp12[20]};
    Full_Adder FA_59(s59, c59, in59_1, in59_2, pp10[22]);
    wire[0:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp14[18]};
    assign in60_2 = {pp15[17]};
    Full_Adder FA_60(s60, c60, in60_1, in60_2, pp13[19]);
    wire[0:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp17[15]};
    assign in61_2 = {pp18[14]};
    Full_Adder FA_61(s61, c61, in61_1, in61_2, pp16[16]);
    wire[0:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp20[12]};
    assign in62_2 = {pp21[11]};
    Full_Adder FA_62(s62, c62, in62_1, in62_2, pp19[13]);
    wire[0:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp23[9]};
    assign in63_2 = {pp24[8]};
    Full_Adder FA_63(s63, c63, in63_1, in63_2, pp22[10]);
    wire[0:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp26[6]};
    assign in64_2 = {pp27[5]};
    Full_Adder FA_64(s64, c64, in64_1, in64_2, pp25[7]);
    wire[0:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp28[4]};
    assign in65_2 = {pp29[3]};
    Half_Adder HA_65(s65, c65, in65_1, in65_2);
    wire[0:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp3[30]};
    assign in66_2 = {pp4[29]};
    Full_Adder FA_66(s66, c66, in66_1, in66_2, pp2[31]);
    wire[0:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp6[27]};
    assign in67_2 = {pp7[26]};
    Full_Adder FA_67(s67, c67, in67_1, in67_2, pp5[28]);
    wire[0:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp9[24]};
    assign in68_2 = {pp10[23]};
    Full_Adder FA_68(s68, c68, in68_1, in68_2, pp8[25]);
    wire[0:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp12[21]};
    assign in69_2 = {pp13[20]};
    Full_Adder FA_69(s69, c69, in69_1, in69_2, pp11[22]);
    wire[0:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp15[18]};
    assign in70_2 = {pp16[17]};
    Full_Adder FA_70(s70, c70, in70_1, in70_2, pp14[19]);
    wire[0:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp18[15]};
    assign in71_2 = {pp19[14]};
    Full_Adder FA_71(s71, c71, in71_1, in71_2, pp17[16]);
    wire[0:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp21[12]};
    assign in72_2 = {pp22[11]};
    Full_Adder FA_72(s72, c72, in72_1, in72_2, pp20[13]);
    wire[0:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp24[9]};
    assign in73_2 = {pp25[8]};
    Full_Adder FA_73(s73, c73, in73_1, in73_2, pp23[10]);
    wire[0:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp27[6]};
    assign in74_2 = {pp28[5]};
    Full_Adder FA_74(s74, c74, in74_1, in74_2, pp26[7]);
    wire[0:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp4[30]};
    assign in75_2 = {pp5[29]};
    Full_Adder FA_75(s75, c75, in75_1, in75_2, pp3[31]);
    wire[0:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp7[27]};
    assign in76_2 = {pp8[26]};
    Full_Adder FA_76(s76, c76, in76_1, in76_2, pp6[28]);
    wire[0:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp10[24]};
    assign in77_2 = {pp11[23]};
    Full_Adder FA_77(s77, c77, in77_1, in77_2, pp9[25]);
    wire[0:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp13[21]};
    assign in78_2 = {pp14[20]};
    Full_Adder FA_78(s78, c78, in78_1, in78_2, pp12[22]);
    wire[0:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp16[18]};
    assign in79_2 = {pp17[17]};
    Full_Adder FA_79(s79, c79, in79_1, in79_2, pp15[19]);
    wire[0:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp19[15]};
    assign in80_2 = {pp20[14]};
    Full_Adder FA_80(s80, c80, in80_1, in80_2, pp18[16]);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp22[12]};
    assign in81_2 = {pp23[11]};
    Full_Adder FA_81(s81, c81, in81_1, in81_2, pp21[13]);
    wire[0:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp25[9]};
    assign in82_2 = {pp26[8]};
    Full_Adder FA_82(s82, c82, in82_1, in82_2, pp24[10]);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp5[30]};
    assign in83_2 = {pp6[29]};
    Full_Adder FA_83(s83, c83, in83_1, in83_2, pp4[31]);
    wire[0:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp8[27]};
    assign in84_2 = {pp9[26]};
    Full_Adder FA_84(s84, c84, in84_1, in84_2, pp7[28]);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp11[24]};
    assign in85_2 = {pp12[23]};
    Full_Adder FA_85(s85, c85, in85_1, in85_2, pp10[25]);
    wire[0:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp14[21]};
    assign in86_2 = {pp15[20]};
    Full_Adder FA_86(s86, c86, in86_1, in86_2, pp13[22]);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp17[18]};
    assign in87_2 = {pp18[17]};
    Full_Adder FA_87(s87, c87, in87_1, in87_2, pp16[19]);
    wire[0:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp20[15]};
    assign in88_2 = {pp21[14]};
    Full_Adder FA_88(s88, c88, in88_1, in88_2, pp19[16]);
    wire[0:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp23[12]};
    assign in89_2 = {pp24[11]};
    Full_Adder FA_89(s89, c89, in89_1, in89_2, pp22[13]);
    wire[0:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp6[30]};
    assign in90_2 = {pp7[29]};
    Full_Adder FA_90(s90, c90, in90_1, in90_2, pp5[31]);
    wire[0:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp9[27]};
    assign in91_2 = {pp10[26]};
    Full_Adder FA_91(s91, c91, in91_1, in91_2, pp8[28]);
    wire[0:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp12[24]};
    assign in92_2 = {pp13[23]};
    Full_Adder FA_92(s92, c92, in92_1, in92_2, pp11[25]);
    wire[0:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp15[21]};
    assign in93_2 = {pp16[20]};
    Full_Adder FA_93(s93, c93, in93_1, in93_2, pp14[22]);
    wire[0:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp18[18]};
    assign in94_2 = {pp19[17]};
    Full_Adder FA_94(s94, c94, in94_1, in94_2, pp17[19]);
    wire[0:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp21[15]};
    assign in95_2 = {pp22[14]};
    Full_Adder FA_95(s95, c95, in95_1, in95_2, pp20[16]);
    wire[0:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp7[30]};
    assign in96_2 = {pp8[29]};
    Full_Adder FA_96(s96, c96, in96_1, in96_2, pp6[31]);
    wire[0:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp10[27]};
    assign in97_2 = {pp11[26]};
    Full_Adder FA_97(s97, c97, in97_1, in97_2, pp9[28]);
    wire[0:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp13[24]};
    assign in98_2 = {pp14[23]};
    Full_Adder FA_98(s98, c98, in98_1, in98_2, pp12[25]);
    wire[0:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp16[21]};
    assign in99_2 = {pp17[20]};
    Full_Adder FA_99(s99, c99, in99_1, in99_2, pp15[22]);
    wire[0:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp19[18]};
    assign in100_2 = {pp20[17]};
    Full_Adder FA_100(s100, c100, in100_1, in100_2, pp18[19]);
    wire[0:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp8[30]};
    assign in101_2 = {pp9[29]};
    Full_Adder FA_101(s101, c101, in101_1, in101_2, pp7[31]);
    wire[0:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp11[27]};
    assign in102_2 = {pp12[26]};
    Full_Adder FA_102(s102, c102, in102_1, in102_2, pp10[28]);
    wire[0:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp14[24]};
    assign in103_2 = {pp15[23]};
    Full_Adder FA_103(s103, c103, in103_1, in103_2, pp13[25]);
    wire[0:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp17[21]};
    assign in104_2 = {pp18[20]};
    Full_Adder FA_104(s104, c104, in104_1, in104_2, pp16[22]);
    wire[0:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp9[30]};
    assign in105_2 = {pp10[29]};
    Full_Adder FA_105(s105, c105, in105_1, in105_2, pp8[31]);
    wire[0:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp12[27]};
    assign in106_2 = {pp13[26]};
    Full_Adder FA_106(s106, c106, in106_1, in106_2, pp11[28]);
    wire[0:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp15[24]};
    assign in107_2 = {pp16[23]};
    Full_Adder FA_107(s107, c107, in107_1, in107_2, pp14[25]);
    wire[0:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp10[30]};
    assign in108_2 = {pp11[29]};
    Full_Adder FA_108(s108, c108, in108_1, in108_2, pp9[31]);
    wire[0:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp13[27]};
    assign in109_2 = {pp14[26]};
    Full_Adder FA_109(s109, c109, in109_1, in109_2, pp12[28]);
    wire[0:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp11[30]};
    assign in110_2 = {pp12[29]};
    Full_Adder FA_110(s110, c110, in110_1, in110_2, pp10[31]);

    /*Stage 2*/
    wire[0:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp0[15]};
    assign in111_2 = {pp1[14]};
    Half_Adder HA_111(s111, c111, in111_1, in111_2);
    wire[0:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp1[15]};
    assign in112_2 = {pp2[14]};
    Full_Adder FA_112(s112, c112, in112_1, in112_2, pp0[16]);
    wire[0:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp3[13]};
    assign in113_2 = {pp4[12]};
    Half_Adder HA_113(s113, c113, in113_1, in113_2);
    wire[0:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp1[16]};
    assign in114_2 = {pp2[15]};
    Full_Adder FA_114(s114, c114, in114_1, in114_2, pp0[17]);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp4[13]};
    assign in115_2 = {pp5[12]};
    Full_Adder FA_115(s115, c115, in115_1, in115_2, pp3[14]);
    wire[0:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp6[11]};
    assign in116_2 = {pp7[10]};
    Half_Adder HA_116(s116, c116, in116_1, in116_2);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp1[17]};
    assign in117_2 = {pp2[16]};
    Full_Adder FA_117(s117, c117, in117_1, in117_2, pp0[18]);
    wire[0:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp4[14]};
    assign in118_2 = {pp5[13]};
    Full_Adder FA_118(s118, c118, in118_1, in118_2, pp3[15]);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp7[11]};
    assign in119_2 = {pp8[10]};
    Full_Adder FA_119(s119, c119, in119_1, in119_2, pp6[12]);
    wire[0:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {pp9[9]};
    assign in120_2 = {pp10[8]};
    Half_Adder HA_120(s120, c120, in120_1, in120_2);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp1[18]};
    assign in121_2 = {pp2[17]};
    Full_Adder FA_121(s121, c121, in121_1, in121_2, pp0[19]);
    wire[0:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp4[15]};
    assign in122_2 = {pp5[14]};
    Full_Adder FA_122(s122, c122, in122_1, in122_2, pp3[16]);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp7[12]};
    assign in123_2 = {pp8[11]};
    Full_Adder FA_123(s123, c123, in123_1, in123_2, pp6[13]);
    wire[0:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp10[9]};
    assign in124_2 = {pp11[8]};
    Full_Adder FA_124(s124, c124, in124_1, in124_2, pp9[10]);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp12[7]};
    assign in125_2 = {pp13[6]};
    Half_Adder HA_125(s125, c125, in125_1, in125_2);
    wire[0:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp1[19]};
    assign in126_2 = {pp2[18]};
    Full_Adder FA_126(s126, c126, in126_1, in126_2, pp0[20]);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {pp4[16]};
    assign in127_2 = {pp5[15]};
    Full_Adder FA_127(s127, c127, in127_1, in127_2, pp3[17]);
    wire[0:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {pp7[13]};
    assign in128_2 = {pp8[12]};
    Full_Adder FA_128(s128, c128, in128_1, in128_2, pp6[14]);
    wire[0:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp10[10]};
    assign in129_2 = {pp11[9]};
    Full_Adder FA_129(s129, c129, in129_1, in129_2, pp9[11]);
    wire[0:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp13[7]};
    assign in130_2 = {pp14[6]};
    Full_Adder FA_130(s130, c130, in130_1, in130_2, pp12[8]);
    wire[0:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp15[5]};
    assign in131_2 = {pp16[4]};
    Half_Adder HA_131(s131, c131, in131_1, in131_2);
    wire[0:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp1[20]};
    assign in132_2 = {pp2[19]};
    Full_Adder FA_132(s132, c132, in132_1, in132_2, pp0[21]);
    wire[0:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp4[17]};
    assign in133_2 = {pp5[16]};
    Full_Adder FA_133(s133, c133, in133_1, in133_2, pp3[18]);
    wire[0:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp7[14]};
    assign in134_2 = {pp8[13]};
    Full_Adder FA_134(s134, c134, in134_1, in134_2, pp6[15]);
    wire[0:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp10[11]};
    assign in135_2 = {pp11[10]};
    Full_Adder FA_135(s135, c135, in135_1, in135_2, pp9[12]);
    wire[0:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp13[8]};
    assign in136_2 = {pp14[7]};
    Full_Adder FA_136(s136, c136, in136_1, in136_2, pp12[9]);
    wire[0:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp16[5]};
    assign in137_2 = {pp17[4]};
    Full_Adder FA_137(s137, c137, in137_1, in137_2, pp15[6]);
    wire[0:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp18[3]};
    assign in138_2 = {pp19[2]};
    Half_Adder HA_138(s138, c138, in138_1, in138_2);
    wire[0:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp3[19]};
    assign in139_2 = {pp4[18]};
    Full_Adder FA_139(s139, c139, in139_1, in139_2, pp2[20]);
    wire[0:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp6[16]};
    assign in140_2 = {pp7[15]};
    Full_Adder FA_140(s140, c140, in140_1, in140_2, pp5[17]);
    wire[0:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp9[13]};
    assign in141_2 = {pp10[12]};
    Full_Adder FA_141(s141, c141, in141_1, in141_2, pp8[14]);
    wire[0:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp12[10]};
    assign in142_2 = {pp13[9]};
    Full_Adder FA_142(s142, c142, in142_1, in142_2, pp11[11]);
    wire[0:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp15[7]};
    assign in143_2 = {pp16[6]};
    Full_Adder FA_143(s143, c143, in143_1, in143_2, pp14[8]);
    wire[0:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp18[4]};
    assign in144_2 = {pp19[3]};
    Full_Adder FA_144(s144, c144, in144_1, in144_2, pp17[5]);
    wire[0:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp21[1]};
    assign in145_2 = {pp22[0]};
    Full_Adder FA_145(s145, c145, in145_1, in145_2, pp20[2]);
    wire[0:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp6[17]};
    assign in146_2 = {pp7[16]};
    Full_Adder FA_146(s146, c146, in146_1, in146_2, pp5[18]);
    wire[0:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp9[14]};
    assign in147_2 = {pp10[13]};
    Full_Adder FA_147(s147, c147, in147_1, in147_2, pp8[15]);
    wire[0:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp12[11]};
    assign in148_2 = {pp13[10]};
    Full_Adder FA_148(s148, c148, in148_1, in148_2, pp11[12]);
    wire[0:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp15[8]};
    assign in149_2 = {pp16[7]};
    Full_Adder FA_149(s149, c149, in149_1, in149_2, pp14[9]);
    wire[0:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp18[5]};
    assign in150_2 = {pp19[4]};
    Full_Adder FA_150(s150, c150, in150_1, in150_2, pp17[6]);
    wire[0:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp21[2]};
    assign in151_2 = {pp22[1]};
    Full_Adder FA_151(s151, c151, in151_1, in151_2, pp20[3]);
    wire[0:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {c1};
    assign in152_2 = {s2[0]};
    Full_Adder FA_152(s152, c152, in152_1, in152_2, pp23[0]);
    wire[0:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp9[15]};
    assign in153_2 = {pp10[14]};
    Full_Adder FA_153(s153, c153, in153_1, in153_2, pp8[16]);
    wire[0:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp12[12]};
    assign in154_2 = {pp13[11]};
    Full_Adder FA_154(s154, c154, in154_1, in154_2, pp11[13]);
    wire[0:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp15[9]};
    assign in155_2 = {pp16[8]};
    Full_Adder FA_155(s155, c155, in155_1, in155_2, pp14[10]);
    wire[0:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp18[6]};
    assign in156_2 = {pp19[5]};
    Full_Adder FA_156(s156, c156, in156_1, in156_2, pp17[7]);
    wire[0:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp21[3]};
    assign in157_2 = {pp22[2]};
    Full_Adder FA_157(s157, c157, in157_1, in157_2, pp20[4]);
    wire[0:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp24[0]};
    assign in158_2 = {c2};
    Full_Adder FA_158(s158, c158, in158_1, in158_2, pp23[1]);
    wire[0:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {s4[0]};
    assign in159_2 = {s5[0]};
    Full_Adder FA_159(s159, c159, in159_1, in159_2, c3);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp12[13]};
    assign in160_2 = {pp13[12]};
    Full_Adder FA_160(s160, c160, in160_1, in160_2, pp11[14]);
    wire[0:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp15[10]};
    assign in161_2 = {pp16[9]};
    Full_Adder FA_161(s161, c161, in161_1, in161_2, pp14[11]);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp18[7]};
    assign in162_2 = {pp19[6]};
    Full_Adder FA_162(s162, c162, in162_1, in162_2, pp17[8]);
    wire[0:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp21[4]};
    assign in163_2 = {pp22[3]};
    Full_Adder FA_163(s163, c163, in163_1, in163_2, pp20[5]);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp24[1]};
    assign in164_2 = {pp25[0]};
    Full_Adder FA_164(s164, c164, in164_1, in164_2, pp23[2]);
    wire[0:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {c5};
    assign in165_2 = {c6};
    Full_Adder FA_165(s165, c165, in165_1, in165_2, c4);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {s8[0]};
    assign in166_2 = {s9[0]};
    Full_Adder FA_166(s166, c166, in166_1, in166_2, s7[0]);
    wire[0:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {pp15[11]};
    assign in167_2 = {pp16[10]};
    Full_Adder FA_167(s167, c167, in167_1, in167_2, pp14[12]);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {pp18[8]};
    assign in168_2 = {pp19[7]};
    Full_Adder FA_168(s168, c168, in168_1, in168_2, pp17[9]);
    wire[0:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {pp21[5]};
    assign in169_2 = {pp22[4]};
    Full_Adder FA_169(s169, c169, in169_1, in169_2, pp20[6]);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {pp24[2]};
    assign in170_2 = {pp25[1]};
    Full_Adder FA_170(s170, c170, in170_1, in170_2, pp23[3]);
    wire[0:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {c7};
    assign in171_2 = {c8};
    Full_Adder FA_171(s171, c171, in171_1, in171_2, pp26[0]);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {c10};
    assign in172_2 = {s11[0]};
    Full_Adder FA_172(s172, c172, in172_1, in172_2, c9);
    wire[0:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {s13[0]};
    assign in173_2 = {s14[0]};
    Full_Adder FA_173(s173, c173, in173_1, in173_2, s12[0]);
    wire[0:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp18[9]};
    assign in174_2 = {pp19[8]};
    Full_Adder FA_174(s174, c174, in174_1, in174_2, pp17[10]);
    wire[0:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp21[6]};
    assign in175_2 = {pp22[5]};
    Full_Adder FA_175(s175, c175, in175_1, in175_2, pp20[7]);
    wire[0:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp24[3]};
    assign in176_2 = {pp25[2]};
    Full_Adder FA_176(s176, c176, in176_1, in176_2, pp23[4]);
    wire[0:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp27[0]};
    assign in177_2 = {c11};
    Full_Adder FA_177(s177, c177, in177_1, in177_2, pp26[1]);
    wire[0:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {c13};
    assign in178_2 = {c14};
    Full_Adder FA_178(s178, c178, in178_1, in178_2, c12);
    wire[0:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {s16[0]};
    assign in179_2 = {s17[0]};
    Full_Adder FA_179(s179, c179, in179_1, in179_2, c15);
    wire[0:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {s19[0]};
    assign in180_2 = {s20[0]};
    Full_Adder FA_180(s180, c180, in180_1, in180_2, s18[0]);
    wire[0:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp21[7]};
    assign in181_2 = {pp22[6]};
    Full_Adder FA_181(s181, c181, in181_1, in181_2, pp20[8]);
    wire[0:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp24[4]};
    assign in182_2 = {pp25[3]};
    Full_Adder FA_182(s182, c182, in182_1, in182_2, pp23[5]);
    wire[0:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp27[1]};
    assign in183_2 = {pp28[0]};
    Full_Adder FA_183(s183, c183, in183_1, in183_2, pp26[2]);
    wire[0:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {c17};
    assign in184_2 = {c18};
    Full_Adder FA_184(s184, c184, in184_1, in184_2, c16);
    wire[0:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {c20};
    assign in185_2 = {c21};
    Full_Adder FA_185(s185, c185, in185_1, in185_2, c19);
    wire[0:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {s23[0]};
    assign in186_2 = {s24[0]};
    Full_Adder FA_186(s186, c186, in186_1, in186_2, s22[0]);
    wire[0:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {s26[0]};
    assign in187_2 = {s27[0]};
    Full_Adder FA_187(s187, c187, in187_1, in187_2, s25[0]);
    wire[0:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp24[5]};
    assign in188_2 = {pp25[4]};
    Full_Adder FA_188(s188, c188, in188_1, in188_2, pp23[6]);
    wire[0:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp27[2]};
    assign in189_2 = {pp28[1]};
    Full_Adder FA_189(s189, c189, in189_1, in189_2, pp26[3]);
    wire[0:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {c22};
    assign in190_2 = {c23};
    Full_Adder FA_190(s190, c190, in190_1, in190_2, pp29[0]);
    wire[0:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {c25};
    assign in191_2 = {c26};
    Full_Adder FA_191(s191, c191, in191_1, in191_2, c24);
    wire[0:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {c28};
    assign in192_2 = {s29[0]};
    Full_Adder FA_192(s192, c192, in192_1, in192_2, c27);
    wire[0:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {s31[0]};
    assign in193_2 = {s32[0]};
    Full_Adder FA_193(s193, c193, in193_1, in193_2, s30[0]);
    wire[0:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {s34[0]};
    assign in194_2 = {s35[0]};
    Full_Adder FA_194(s194, c194, in194_1, in194_2, s33[0]);
    wire[0:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp27[3]};
    assign in195_2 = {pp28[2]};
    Full_Adder FA_195(s195, c195, in195_1, in195_2, pp26[4]);
    wire[0:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp30[0]};
    assign in196_2 = {c29};
    Full_Adder FA_196(s196, c196, in196_1, in196_2, pp29[1]);
    wire[0:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {c31};
    assign in197_2 = {c32};
    Full_Adder FA_197(s197, c197, in197_1, in197_2, c30);
    wire[0:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {c34};
    assign in198_2 = {c35};
    Full_Adder FA_198(s198, c198, in198_1, in198_2, c33);
    wire[0:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {s37[0]};
    assign in199_2 = {s38[0]};
    Full_Adder FA_199(s199, c199, in199_1, in199_2, c36);
    wire[0:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {s40[0]};
    assign in200_2 = {s41[0]};
    Full_Adder FA_200(s200, c200, in200_1, in200_2, s39[0]);
    wire[0:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {s43[0]};
    assign in201_2 = {s44[0]};
    Full_Adder FA_201(s201, c201, in201_1, in201_2, s42[0]);
    wire[0:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp30[1]};
    assign in202_2 = {pp31[0]};
    Full_Adder FA_202(s202, c202, in202_1, in202_2, pp29[2]);
    wire[0:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {c38};
    assign in203_2 = {c39};
    Full_Adder FA_203(s203, c203, in203_1, in203_2, c37);
    wire[0:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {c41};
    assign in204_2 = {c42};
    Full_Adder FA_204(s204, c204, in204_1, in204_2, c40);
    wire[0:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {c44};
    assign in205_2 = {c45};
    Full_Adder FA_205(s205, c205, in205_1, in205_2, c43);
    wire[0:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {s47[0]};
    assign in206_2 = {s48[0]};
    Full_Adder FA_206(s206, c206, in206_1, in206_2, s46[0]);
    wire[0:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {s50[0]};
    assign in207_2 = {s51[0]};
    Full_Adder FA_207(s207, c207, in207_1, in207_2, s49[0]);
    wire[0:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {s53[0]};
    assign in208_2 = {s54[0]};
    Full_Adder FA_208(s208, c208, in208_1, in208_2, s52[0]);
    wire[0:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {pp31[1]};
    assign in209_2 = {c46};
    Full_Adder FA_209(s209, c209, in209_1, in209_2, pp30[2]);
    wire[0:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {c48};
    assign in210_2 = {c49};
    Full_Adder FA_210(s210, c210, in210_1, in210_2, c47);
    wire[0:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {c51};
    assign in211_2 = {c52};
    Full_Adder FA_211(s211, c211, in211_1, in211_2, c50);
    wire[0:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {c54};
    assign in212_2 = {c55};
    Full_Adder FA_212(s212, c212, in212_1, in212_2, c53);
    wire[0:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {s57[0]};
    assign in213_2 = {s58[0]};
    Full_Adder FA_213(s213, c213, in213_1, in213_2, s56[0]);
    wire[0:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {s60[0]};
    assign in214_2 = {s61[0]};
    Full_Adder FA_214(s214, c214, in214_1, in214_2, s59[0]);
    wire[0:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {s63[0]};
    assign in215_2 = {s64[0]};
    Full_Adder FA_215(s215, c215, in215_1, in215_2, s62[0]);
    wire[0:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {pp30[3]};
    assign in216_2 = {pp31[2]};
    Full_Adder FA_216(s216, c216, in216_1, in216_2, pp29[4]);
    wire[0:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {c57};
    assign in217_2 = {c58};
    Full_Adder FA_217(s217, c217, in217_1, in217_2, c56);
    wire[0:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {c60};
    assign in218_2 = {c61};
    Full_Adder FA_218(s218, c218, in218_1, in218_2, c59);
    wire[0:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {c63};
    assign in219_2 = {c64};
    Full_Adder FA_219(s219, c219, in219_1, in219_2, c62);
    wire[0:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {s66[0]};
    assign in220_2 = {s67[0]};
    Full_Adder FA_220(s220, c220, in220_1, in220_2, c65);
    wire[0:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {s69[0]};
    assign in221_2 = {s70[0]};
    Full_Adder FA_221(s221, c221, in221_1, in221_2, s68[0]);
    wire[0:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {s72[0]};
    assign in222_2 = {s73[0]};
    Full_Adder FA_222(s222, c222, in222_1, in222_2, s71[0]);
    wire[0:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {pp28[6]};
    assign in223_2 = {pp29[5]};
    Full_Adder FA_223(s223, c223, in223_1, in223_2, pp27[7]);
    wire[0:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {pp31[3]};
    assign in224_2 = {c66};
    Full_Adder FA_224(s224, c224, in224_1, in224_2, pp30[4]);
    wire[0:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {c68};
    assign in225_2 = {c69};
    Full_Adder FA_225(s225, c225, in225_1, in225_2, c67);
    wire[0:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {c71};
    assign in226_2 = {c72};
    Full_Adder FA_226(s226, c226, in226_1, in226_2, c70);
    wire[0:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {c74};
    assign in227_2 = {s75[0]};
    Full_Adder FA_227(s227, c227, in227_1, in227_2, c73);
    wire[0:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {s77[0]};
    assign in228_2 = {s78[0]};
    Full_Adder FA_228(s228, c228, in228_1, in228_2, s76[0]);
    wire[0:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {s80[0]};
    assign in229_2 = {s81[0]};
    Full_Adder FA_229(s229, c229, in229_1, in229_2, s79[0]);
    wire[0:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp26[9]};
    assign in230_2 = {pp27[8]};
    Full_Adder FA_230(s230, c230, in230_1, in230_2, pp25[10]);
    wire[0:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp29[6]};
    assign in231_2 = {pp30[5]};
    Full_Adder FA_231(s231, c231, in231_1, in231_2, pp28[7]);
    wire[0:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {c75};
    assign in232_2 = {c76};
    Full_Adder FA_232(s232, c232, in232_1, in232_2, pp31[4]);
    wire[0:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {c78};
    assign in233_2 = {c79};
    Full_Adder FA_233(s233, c233, in233_1, in233_2, c77);
    wire[0:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {c81};
    assign in234_2 = {c82};
    Full_Adder FA_234(s234, c234, in234_1, in234_2, c80);
    wire[0:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {s84[0]};
    assign in235_2 = {s85[0]};
    Full_Adder FA_235(s235, c235, in235_1, in235_2, s83[0]);
    wire[0:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {s87[0]};
    assign in236_2 = {s88[0]};
    Full_Adder FA_236(s236, c236, in236_1, in236_2, s86[0]);
    wire[0:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {pp24[12]};
    assign in237_2 = {pp25[11]};
    Full_Adder FA_237(s237, c237, in237_1, in237_2, pp23[13]);
    wire[0:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {pp27[9]};
    assign in238_2 = {pp28[8]};
    Full_Adder FA_238(s238, c238, in238_1, in238_2, pp26[10]);
    wire[0:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {pp30[6]};
    assign in239_2 = {pp31[5]};
    Full_Adder FA_239(s239, c239, in239_1, in239_2, pp29[7]);
    wire[0:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {c84};
    assign in240_2 = {c85};
    Full_Adder FA_240(s240, c240, in240_1, in240_2, c83);
    wire[0:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {c87};
    assign in241_2 = {c88};
    Full_Adder FA_241(s241, c241, in241_1, in241_2, c86);
    wire[0:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {s90[0]};
    assign in242_2 = {s91[0]};
    Full_Adder FA_242(s242, c242, in242_1, in242_2, c89);
    wire[0:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {s93[0]};
    assign in243_2 = {s94[0]};
    Full_Adder FA_243(s243, c243, in243_1, in243_2, s92[0]);
    wire[0:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp22[15]};
    assign in244_2 = {pp23[14]};
    Full_Adder FA_244(s244, c244, in244_1, in244_2, pp21[16]);
    wire[0:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {pp25[12]};
    assign in245_2 = {pp26[11]};
    Full_Adder FA_245(s245, c245, in245_1, in245_2, pp24[13]);
    wire[0:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {pp28[9]};
    assign in246_2 = {pp29[8]};
    Full_Adder FA_246(s246, c246, in246_1, in246_2, pp27[10]);
    wire[0:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {pp31[6]};
    assign in247_2 = {c90};
    Full_Adder FA_247(s247, c247, in247_1, in247_2, pp30[7]);
    wire[0:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {c92};
    assign in248_2 = {c93};
    Full_Adder FA_248(s248, c248, in248_1, in248_2, c91);
    wire[0:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {c95};
    assign in249_2 = {s96[0]};
    Full_Adder FA_249(s249, c249, in249_1, in249_2, c94);
    wire[0:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {s98[0]};
    assign in250_2 = {s99[0]};
    Full_Adder FA_250(s250, c250, in250_1, in250_2, s97[0]);
    wire[0:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp20[18]};
    assign in251_2 = {pp21[17]};
    Full_Adder FA_251(s251, c251, in251_1, in251_2, pp19[19]);
    wire[0:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp23[15]};
    assign in252_2 = {pp24[14]};
    Full_Adder FA_252(s252, c252, in252_1, in252_2, pp22[16]);
    wire[0:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp26[12]};
    assign in253_2 = {pp27[11]};
    Full_Adder FA_253(s253, c253, in253_1, in253_2, pp25[13]);
    wire[0:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp29[9]};
    assign in254_2 = {pp30[8]};
    Full_Adder FA_254(s254, c254, in254_1, in254_2, pp28[10]);
    wire[0:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {c96};
    assign in255_2 = {c97};
    Full_Adder FA_255(s255, c255, in255_1, in255_2, pp31[7]);
    wire[0:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {c99};
    assign in256_2 = {c100};
    Full_Adder FA_256(s256, c256, in256_1, in256_2, c98);
    wire[0:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {s102[0]};
    assign in257_2 = {s103[0]};
    Full_Adder FA_257(s257, c257, in257_1, in257_2, s101[0]);
    wire[0:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {pp18[21]};
    assign in258_2 = {pp19[20]};
    Full_Adder FA_258(s258, c258, in258_1, in258_2, pp17[22]);
    wire[0:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {pp21[18]};
    assign in259_2 = {pp22[17]};
    Full_Adder FA_259(s259, c259, in259_1, in259_2, pp20[19]);
    wire[0:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {pp24[15]};
    assign in260_2 = {pp25[14]};
    Full_Adder FA_260(s260, c260, in260_1, in260_2, pp23[16]);
    wire[0:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {pp27[12]};
    assign in261_2 = {pp28[11]};
    Full_Adder FA_261(s261, c261, in261_1, in261_2, pp26[13]);
    wire[0:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {pp30[9]};
    assign in262_2 = {pp31[8]};
    Full_Adder FA_262(s262, c262, in262_1, in262_2, pp29[10]);
    wire[0:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {c102};
    assign in263_2 = {c103};
    Full_Adder FA_263(s263, c263, in263_1, in263_2, c101);
    wire[0:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {s105[0]};
    assign in264_2 = {s106[0]};
    Full_Adder FA_264(s264, c264, in264_1, in264_2, c104);
    wire[0:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {pp16[24]};
    assign in265_2 = {pp17[23]};
    Full_Adder FA_265(s265, c265, in265_1, in265_2, pp15[25]);
    wire[0:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {pp19[21]};
    assign in266_2 = {pp20[20]};
    Full_Adder FA_266(s266, c266, in266_1, in266_2, pp18[22]);
    wire[0:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {pp22[18]};
    assign in267_2 = {pp23[17]};
    Full_Adder FA_267(s267, c267, in267_1, in267_2, pp21[19]);
    wire[0:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {pp25[15]};
    assign in268_2 = {pp26[14]};
    Full_Adder FA_268(s268, c268, in268_1, in268_2, pp24[16]);
    wire[0:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {pp28[12]};
    assign in269_2 = {pp29[11]};
    Full_Adder FA_269(s269, c269, in269_1, in269_2, pp27[13]);
    wire[0:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {pp31[9]};
    assign in270_2 = {c105};
    Full_Adder FA_270(s270, c270, in270_1, in270_2, pp30[10]);
    wire[0:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {c107};
    assign in271_2 = {s108[0]};
    Full_Adder FA_271(s271, c271, in271_1, in271_2, c106);
    wire[0:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {pp14[27]};
    assign in272_2 = {pp15[26]};
    Full_Adder FA_272(s272, c272, in272_1, in272_2, pp13[28]);
    wire[0:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {pp17[24]};
    assign in273_2 = {pp18[23]};
    Full_Adder FA_273(s273, c273, in273_1, in273_2, pp16[25]);
    wire[0:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {pp20[21]};
    assign in274_2 = {pp21[20]};
    Full_Adder FA_274(s274, c274, in274_1, in274_2, pp19[22]);
    wire[0:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp23[18]};
    assign in275_2 = {pp24[17]};
    Full_Adder FA_275(s275, c275, in275_1, in275_2, pp22[19]);
    wire[0:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {pp26[15]};
    assign in276_2 = {pp27[14]};
    Full_Adder FA_276(s276, c276, in276_1, in276_2, pp25[16]);
    wire[0:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {pp29[12]};
    assign in277_2 = {pp30[11]};
    Full_Adder FA_277(s277, c277, in277_1, in277_2, pp28[13]);
    wire[0:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {c108};
    assign in278_2 = {c109};
    Full_Adder FA_278(s278, c278, in278_1, in278_2, pp31[10]);
    wire[0:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {pp12[30]};
    assign in279_2 = {pp13[29]};
    Full_Adder FA_279(s279, c279, in279_1, in279_2, pp11[31]);
    wire[0:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {pp15[27]};
    assign in280_2 = {pp16[26]};
    Full_Adder FA_280(s280, c280, in280_1, in280_2, pp14[28]);
    wire[0:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {pp18[24]};
    assign in281_2 = {pp19[23]};
    Full_Adder FA_281(s281, c281, in281_1, in281_2, pp17[25]);
    wire[0:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {pp21[21]};
    assign in282_2 = {pp22[20]};
    Full_Adder FA_282(s282, c282, in282_1, in282_2, pp20[22]);
    wire[0:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {pp24[18]};
    assign in283_2 = {pp25[17]};
    Full_Adder FA_283(s283, c283, in283_1, in283_2, pp23[19]);
    wire[0:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {pp27[15]};
    assign in284_2 = {pp28[14]};
    Full_Adder FA_284(s284, c284, in284_1, in284_2, pp26[16]);
    wire[0:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {pp30[12]};
    assign in285_2 = {pp31[11]};
    Full_Adder FA_285(s285, c285, in285_1, in285_2, pp29[13]);
    wire[0:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {pp13[30]};
    assign in286_2 = {pp14[29]};
    Full_Adder FA_286(s286, c286, in286_1, in286_2, pp12[31]);
    wire[0:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {pp16[27]};
    assign in287_2 = {pp17[26]};
    Full_Adder FA_287(s287, c287, in287_1, in287_2, pp15[28]);
    wire[0:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {pp19[24]};
    assign in288_2 = {pp20[23]};
    Full_Adder FA_288(s288, c288, in288_1, in288_2, pp18[25]);
    wire[0:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {pp22[21]};
    assign in289_2 = {pp23[20]};
    Full_Adder FA_289(s289, c289, in289_1, in289_2, pp21[22]);
    wire[0:0] s290, in290_1, in290_2;
    wire c290;
    assign in290_1 = {pp25[18]};
    assign in290_2 = {pp26[17]};
    Full_Adder FA_290(s290, c290, in290_1, in290_2, pp24[19]);
    wire[0:0] s291, in291_1, in291_2;
    wire c291;
    assign in291_1 = {pp28[15]};
    assign in291_2 = {pp29[14]};
    Full_Adder FA_291(s291, c291, in291_1, in291_2, pp27[16]);
    wire[0:0] s292, in292_1, in292_2;
    wire c292;
    assign in292_1 = {pp14[30]};
    assign in292_2 = {pp15[29]};
    Full_Adder FA_292(s292, c292, in292_1, in292_2, pp13[31]);
    wire[0:0] s293, in293_1, in293_2;
    wire c293;
    assign in293_1 = {pp17[27]};
    assign in293_2 = {pp18[26]};
    Full_Adder FA_293(s293, c293, in293_1, in293_2, pp16[28]);
    wire[0:0] s294, in294_1, in294_2;
    wire c294;
    assign in294_1 = {pp20[24]};
    assign in294_2 = {pp21[23]};
    Full_Adder FA_294(s294, c294, in294_1, in294_2, pp19[25]);
    wire[0:0] s295, in295_1, in295_2;
    wire c295;
    assign in295_1 = {pp23[21]};
    assign in295_2 = {pp24[20]};
    Full_Adder FA_295(s295, c295, in295_1, in295_2, pp22[22]);
    wire[0:0] s296, in296_1, in296_2;
    wire c296;
    assign in296_1 = {pp26[18]};
    assign in296_2 = {pp27[17]};
    Full_Adder FA_296(s296, c296, in296_1, in296_2, pp25[19]);
    wire[0:0] s297, in297_1, in297_2;
    wire c297;
    assign in297_1 = {pp15[30]};
    assign in297_2 = {pp16[29]};
    Full_Adder FA_297(s297, c297, in297_1, in297_2, pp14[31]);
    wire[0:0] s298, in298_1, in298_2;
    wire c298;
    assign in298_1 = {pp18[27]};
    assign in298_2 = {pp19[26]};
    Full_Adder FA_298(s298, c298, in298_1, in298_2, pp17[28]);
    wire[0:0] s299, in299_1, in299_2;
    wire c299;
    assign in299_1 = {pp21[24]};
    assign in299_2 = {pp22[23]};
    Full_Adder FA_299(s299, c299, in299_1, in299_2, pp20[25]);
    wire[0:0] s300, in300_1, in300_2;
    wire c300;
    assign in300_1 = {pp24[21]};
    assign in300_2 = {pp25[20]};
    Full_Adder FA_300(s300, c300, in300_1, in300_2, pp23[22]);
    wire[0:0] s301, in301_1, in301_2;
    wire c301;
    assign in301_1 = {pp16[30]};
    assign in301_2 = {pp17[29]};
    Full_Adder FA_301(s301, c301, in301_1, in301_2, pp15[31]);
    wire[0:0] s302, in302_1, in302_2;
    wire c302;
    assign in302_1 = {pp19[27]};
    assign in302_2 = {pp20[26]};
    Full_Adder FA_302(s302, c302, in302_1, in302_2, pp18[28]);
    wire[0:0] s303, in303_1, in303_2;
    wire c303;
    assign in303_1 = {pp22[24]};
    assign in303_2 = {pp23[23]};
    Full_Adder FA_303(s303, c303, in303_1, in303_2, pp21[25]);
    wire[0:0] s304, in304_1, in304_2;
    wire c304;
    assign in304_1 = {pp17[30]};
    assign in304_2 = {pp18[29]};
    Full_Adder FA_304(s304, c304, in304_1, in304_2, pp16[31]);
    wire[0:0] s305, in305_1, in305_2;
    wire c305;
    assign in305_1 = {pp20[27]};
    assign in305_2 = {pp21[26]};
    Full_Adder FA_305(s305, c305, in305_1, in305_2, pp19[28]);
    wire[0:0] s306, in306_1, in306_2;
    wire c306;
    assign in306_1 = {pp18[30]};
    assign in306_2 = {pp19[29]};
    Full_Adder FA_306(s306, c306, in306_1, in306_2, pp17[31]);

    /*Stage 3*/
    wire[0:0] s307, in307_1, in307_2;
    wire c307;
    assign in307_1 = {pp0[10]};
    assign in307_2 = {pp1[9]};
    Half_Adder HA_307(s307, c307, in307_1, in307_2);
    wire[0:0] s308, in308_1, in308_2;
    wire c308;
    assign in308_1 = {pp1[10]};
    assign in308_2 = {pp2[9]};
    Full_Adder FA_308(s308, c308, in308_1, in308_2, pp0[11]);
    wire[0:0] s309, in309_1, in309_2;
    wire c309;
    assign in309_1 = {pp3[8]};
    assign in309_2 = {pp4[7]};
    Half_Adder HA_309(s309, c309, in309_1, in309_2);
    wire[0:0] s310, in310_1, in310_2;
    wire c310;
    assign in310_1 = {pp1[11]};
    assign in310_2 = {pp2[10]};
    Full_Adder FA_310(s310, c310, in310_1, in310_2, pp0[12]);
    wire[0:0] s311, in311_1, in311_2;
    wire c311;
    assign in311_1 = {pp4[8]};
    assign in311_2 = {pp5[7]};
    Full_Adder FA_311(s311, c311, in311_1, in311_2, pp3[9]);
    wire[0:0] s312, in312_1, in312_2;
    wire c312;
    assign in312_1 = {pp6[6]};
    assign in312_2 = {pp7[5]};
    Half_Adder HA_312(s312, c312, in312_1, in312_2);
    wire[0:0] s313, in313_1, in313_2;
    wire c313;
    assign in313_1 = {pp1[12]};
    assign in313_2 = {pp2[11]};
    Full_Adder FA_313(s313, c313, in313_1, in313_2, pp0[13]);
    wire[0:0] s314, in314_1, in314_2;
    wire c314;
    assign in314_1 = {pp4[9]};
    assign in314_2 = {pp5[8]};
    Full_Adder FA_314(s314, c314, in314_1, in314_2, pp3[10]);
    wire[0:0] s315, in315_1, in315_2;
    wire c315;
    assign in315_1 = {pp7[6]};
    assign in315_2 = {pp8[5]};
    Full_Adder FA_315(s315, c315, in315_1, in315_2, pp6[7]);
    wire[0:0] s316, in316_1, in316_2;
    wire c316;
    assign in316_1 = {pp9[4]};
    assign in316_2 = {pp10[3]};
    Half_Adder HA_316(s316, c316, in316_1, in316_2);
    wire[0:0] s317, in317_1, in317_2;
    wire c317;
    assign in317_1 = {pp1[13]};
    assign in317_2 = {pp2[12]};
    Full_Adder FA_317(s317, c317, in317_1, in317_2, pp0[14]);
    wire[0:0] s318, in318_1, in318_2;
    wire c318;
    assign in318_1 = {pp4[10]};
    assign in318_2 = {pp5[9]};
    Full_Adder FA_318(s318, c318, in318_1, in318_2, pp3[11]);
    wire[0:0] s319, in319_1, in319_2;
    wire c319;
    assign in319_1 = {pp7[7]};
    assign in319_2 = {pp8[6]};
    Full_Adder FA_319(s319, c319, in319_1, in319_2, pp6[8]);
    wire[0:0] s320, in320_1, in320_2;
    wire c320;
    assign in320_1 = {pp10[4]};
    assign in320_2 = {pp11[3]};
    Full_Adder FA_320(s320, c320, in320_1, in320_2, pp9[5]);
    wire[0:0] s321, in321_1, in321_2;
    wire c321;
    assign in321_1 = {pp12[2]};
    assign in321_2 = {pp13[1]};
    Half_Adder HA_321(s321, c321, in321_1, in321_2);
    wire[0:0] s322, in322_1, in322_2;
    wire c322;
    assign in322_1 = {pp3[12]};
    assign in322_2 = {pp4[11]};
    Full_Adder FA_322(s322, c322, in322_1, in322_2, pp2[13]);
    wire[0:0] s323, in323_1, in323_2;
    wire c323;
    assign in323_1 = {pp6[9]};
    assign in323_2 = {pp7[8]};
    Full_Adder FA_323(s323, c323, in323_1, in323_2, pp5[10]);
    wire[0:0] s324, in324_1, in324_2;
    wire c324;
    assign in324_1 = {pp9[6]};
    assign in324_2 = {pp10[5]};
    Full_Adder FA_324(s324, c324, in324_1, in324_2, pp8[7]);
    wire[0:0] s325, in325_1, in325_2;
    wire c325;
    assign in325_1 = {pp12[3]};
    assign in325_2 = {pp13[2]};
    Full_Adder FA_325(s325, c325, in325_1, in325_2, pp11[4]);
    wire[0:0] s326, in326_1, in326_2;
    wire c326;
    assign in326_1 = {pp15[0]};
    assign in326_2 = {s111[0]};
    Full_Adder FA_326(s326, c326, in326_1, in326_2, pp14[1]);
    wire[0:0] s327, in327_1, in327_2;
    wire c327;
    assign in327_1 = {pp6[10]};
    assign in327_2 = {pp7[9]};
    Full_Adder FA_327(s327, c327, in327_1, in327_2, pp5[11]);
    wire[0:0] s328, in328_1, in328_2;
    wire c328;
    assign in328_1 = {pp9[7]};
    assign in328_2 = {pp10[6]};
    Full_Adder FA_328(s328, c328, in328_1, in328_2, pp8[8]);
    wire[0:0] s329, in329_1, in329_2;
    wire c329;
    assign in329_1 = {pp12[4]};
    assign in329_2 = {pp13[3]};
    Full_Adder FA_329(s329, c329, in329_1, in329_2, pp11[5]);
    wire[0:0] s330, in330_1, in330_2;
    wire c330;
    assign in330_1 = {pp15[1]};
    assign in330_2 = {pp16[0]};
    Full_Adder FA_330(s330, c330, in330_1, in330_2, pp14[2]);
    wire[0:0] s331, in331_1, in331_2;
    wire c331;
    assign in331_1 = {s112[0]};
    assign in331_2 = {s113[0]};
    Full_Adder FA_331(s331, c331, in331_1, in331_2, c111);
    wire[0:0] s332, in332_1, in332_2;
    wire c332;
    assign in332_1 = {pp9[8]};
    assign in332_2 = {pp10[7]};
    Full_Adder FA_332(s332, c332, in332_1, in332_2, pp8[9]);
    wire[0:0] s333, in333_1, in333_2;
    wire c333;
    assign in333_1 = {pp12[5]};
    assign in333_2 = {pp13[4]};
    Full_Adder FA_333(s333, c333, in333_1, in333_2, pp11[6]);
    wire[0:0] s334, in334_1, in334_2;
    wire c334;
    assign in334_1 = {pp15[2]};
    assign in334_2 = {pp16[1]};
    Full_Adder FA_334(s334, c334, in334_1, in334_2, pp14[3]);
    wire[0:0] s335, in335_1, in335_2;
    wire c335;
    assign in335_1 = {c112};
    assign in335_2 = {c113};
    Full_Adder FA_335(s335, c335, in335_1, in335_2, pp17[0]);
    wire[0:0] s336, in336_1, in336_2;
    wire c336;
    assign in336_1 = {s115[0]};
    assign in336_2 = {s116[0]};
    Full_Adder FA_336(s336, c336, in336_1, in336_2, s114[0]);
    wire[0:0] s337, in337_1, in337_2;
    wire c337;
    assign in337_1 = {pp12[6]};
    assign in337_2 = {pp13[5]};
    Full_Adder FA_337(s337, c337, in337_1, in337_2, pp11[7]);
    wire[0:0] s338, in338_1, in338_2;
    wire c338;
    assign in338_1 = {pp15[3]};
    assign in338_2 = {pp16[2]};
    Full_Adder FA_338(s338, c338, in338_1, in338_2, pp14[4]);
    wire[0:0] s339, in339_1, in339_2;
    wire c339;
    assign in339_1 = {pp18[0]};
    assign in339_2 = {c114};
    Full_Adder FA_339(s339, c339, in339_1, in339_2, pp17[1]);
    wire[0:0] s340, in340_1, in340_2;
    wire c340;
    assign in340_1 = {c116};
    assign in340_2 = {s117[0]};
    Full_Adder FA_340(s340, c340, in340_1, in340_2, c115);
    wire[0:0] s341, in341_1, in341_2;
    wire c341;
    assign in341_1 = {s119[0]};
    assign in341_2 = {s120[0]};
    Full_Adder FA_341(s341, c341, in341_1, in341_2, s118[0]);
    wire[0:0] s342, in342_1, in342_2;
    wire c342;
    assign in342_1 = {pp15[4]};
    assign in342_2 = {pp16[3]};
    Full_Adder FA_342(s342, c342, in342_1, in342_2, pp14[5]);
    wire[0:0] s343, in343_1, in343_2;
    wire c343;
    assign in343_1 = {pp18[1]};
    assign in343_2 = {pp19[0]};
    Full_Adder FA_343(s343, c343, in343_1, in343_2, pp17[2]);
    wire[0:0] s344, in344_1, in344_2;
    wire c344;
    assign in344_1 = {c118};
    assign in344_2 = {c119};
    Full_Adder FA_344(s344, c344, in344_1, in344_2, c117);
    wire[0:0] s345, in345_1, in345_2;
    wire c345;
    assign in345_1 = {s121[0]};
    assign in345_2 = {s122[0]};
    Full_Adder FA_345(s345, c345, in345_1, in345_2, c120);
    wire[0:0] s346, in346_1, in346_2;
    wire c346;
    assign in346_1 = {s124[0]};
    assign in346_2 = {s125[0]};
    Full_Adder FA_346(s346, c346, in346_1, in346_2, s123[0]);
    wire[0:0] s347, in347_1, in347_2;
    wire c347;
    assign in347_1 = {pp18[2]};
    assign in347_2 = {pp19[1]};
    Full_Adder FA_347(s347, c347, in347_1, in347_2, pp17[3]);
    wire[0:0] s348, in348_1, in348_2;
    wire c348;
    assign in348_1 = {c121};
    assign in348_2 = {c122};
    Full_Adder FA_348(s348, c348, in348_1, in348_2, pp20[0]);
    wire[0:0] s349, in349_1, in349_2;
    wire c349;
    assign in349_1 = {c124};
    assign in349_2 = {c125};
    Full_Adder FA_349(s349, c349, in349_1, in349_2, c123);
    wire[0:0] s350, in350_1, in350_2;
    wire c350;
    assign in350_1 = {s127[0]};
    assign in350_2 = {s128[0]};
    Full_Adder FA_350(s350, c350, in350_1, in350_2, s126[0]);
    wire[0:0] s351, in351_1, in351_2;
    wire c351;
    assign in351_1 = {s130[0]};
    assign in351_2 = {s131[0]};
    Full_Adder FA_351(s351, c351, in351_1, in351_2, s129[0]);
    wire[0:0] s352, in352_1, in352_2;
    wire c352;
    assign in352_1 = {pp21[0]};
    assign in352_2 = {c126};
    Full_Adder FA_352(s352, c352, in352_1, in352_2, pp20[1]);
    wire[0:0] s353, in353_1, in353_2;
    wire c353;
    assign in353_1 = {c128};
    assign in353_2 = {c129};
    Full_Adder FA_353(s353, c353, in353_1, in353_2, c127);
    wire[0:0] s354, in354_1, in354_2;
    wire c354;
    assign in354_1 = {c131};
    assign in354_2 = {s132[0]};
    Full_Adder FA_354(s354, c354, in354_1, in354_2, c130);
    wire[0:0] s355, in355_1, in355_2;
    wire c355;
    assign in355_1 = {s134[0]};
    assign in355_2 = {s135[0]};
    Full_Adder FA_355(s355, c355, in355_1, in355_2, s133[0]);
    wire[0:0] s356, in356_1, in356_2;
    wire c356;
    assign in356_1 = {s137[0]};
    assign in356_2 = {s138[0]};
    Full_Adder FA_356(s356, c356, in356_1, in356_2, s136[0]);
    wire[0:0] s357, in357_1, in357_2;
    wire c357;
    assign in357_1 = {c132};
    assign in357_2 = {c133};
    Full_Adder FA_357(s357, c357, in357_1, in357_2, s1[0]);
    wire[0:0] s358, in358_1, in358_2;
    wire c358;
    assign in358_1 = {c135};
    assign in358_2 = {c136};
    Full_Adder FA_358(s358, c358, in358_1, in358_2, c134);
    wire[0:0] s359, in359_1, in359_2;
    wire c359;
    assign in359_1 = {c138};
    assign in359_2 = {s139[0]};
    Full_Adder FA_359(s359, c359, in359_1, in359_2, c137);
    wire[0:0] s360, in360_1, in360_2;
    wire c360;
    assign in360_1 = {s141[0]};
    assign in360_2 = {s142[0]};
    Full_Adder FA_360(s360, c360, in360_1, in360_2, s140[0]);
    wire[0:0] s361, in361_1, in361_2;
    wire c361;
    assign in361_1 = {s144[0]};
    assign in361_2 = {s145[0]};
    Full_Adder FA_361(s361, c361, in361_1, in361_2, s143[0]);
    wire[0:0] s362, in362_1, in362_2;
    wire c362;
    assign in362_1 = {c139};
    assign in362_2 = {c140};
    Full_Adder FA_362(s362, c362, in362_1, in362_2, s3[0]);
    wire[0:0] s363, in363_1, in363_2;
    wire c363;
    assign in363_1 = {c142};
    assign in363_2 = {c143};
    Full_Adder FA_363(s363, c363, in363_1, in363_2, c141);
    wire[0:0] s364, in364_1, in364_2;
    wire c364;
    assign in364_1 = {c145};
    assign in364_2 = {s146[0]};
    Full_Adder FA_364(s364, c364, in364_1, in364_2, c144);
    wire[0:0] s365, in365_1, in365_2;
    wire c365;
    assign in365_1 = {s148[0]};
    assign in365_2 = {s149[0]};
    Full_Adder FA_365(s365, c365, in365_1, in365_2, s147[0]);
    wire[0:0] s366, in366_1, in366_2;
    wire c366;
    assign in366_1 = {s151[0]};
    assign in366_2 = {s152[0]};
    Full_Adder FA_366(s366, c366, in366_1, in366_2, s150[0]);
    wire[0:0] s367, in367_1, in367_2;
    wire c367;
    assign in367_1 = {c146};
    assign in367_2 = {c147};
    Full_Adder FA_367(s367, c367, in367_1, in367_2, s6[0]);
    wire[0:0] s368, in368_1, in368_2;
    wire c368;
    assign in368_1 = {c149};
    assign in368_2 = {c150};
    Full_Adder FA_368(s368, c368, in368_1, in368_2, c148);
    wire[0:0] s369, in369_1, in369_2;
    wire c369;
    assign in369_1 = {c152};
    assign in369_2 = {s153[0]};
    Full_Adder FA_369(s369, c369, in369_1, in369_2, c151);
    wire[0:0] s370, in370_1, in370_2;
    wire c370;
    assign in370_1 = {s155[0]};
    assign in370_2 = {s156[0]};
    Full_Adder FA_370(s370, c370, in370_1, in370_2, s154[0]);
    wire[0:0] s371, in371_1, in371_2;
    wire c371;
    assign in371_1 = {s158[0]};
    assign in371_2 = {s159[0]};
    Full_Adder FA_371(s371, c371, in371_1, in371_2, s157[0]);
    wire[0:0] s372, in372_1, in372_2;
    wire c372;
    assign in372_1 = {c153};
    assign in372_2 = {c154};
    Full_Adder FA_372(s372, c372, in372_1, in372_2, s10[0]);
    wire[0:0] s373, in373_1, in373_2;
    wire c373;
    assign in373_1 = {c156};
    assign in373_2 = {c157};
    Full_Adder FA_373(s373, c373, in373_1, in373_2, c155);
    wire[0:0] s374, in374_1, in374_2;
    wire c374;
    assign in374_1 = {c159};
    assign in374_2 = {s160[0]};
    Full_Adder FA_374(s374, c374, in374_1, in374_2, c158);
    wire[0:0] s375, in375_1, in375_2;
    wire c375;
    assign in375_1 = {s162[0]};
    assign in375_2 = {s163[0]};
    Full_Adder FA_375(s375, c375, in375_1, in375_2, s161[0]);
    wire[0:0] s376, in376_1, in376_2;
    wire c376;
    assign in376_1 = {s165[0]};
    assign in376_2 = {s166[0]};
    Full_Adder FA_376(s376, c376, in376_1, in376_2, s164[0]);
    wire[0:0] s377, in377_1, in377_2;
    wire c377;
    assign in377_1 = {c160};
    assign in377_2 = {c161};
    Full_Adder FA_377(s377, c377, in377_1, in377_2, s15[0]);
    wire[0:0] s378, in378_1, in378_2;
    wire c378;
    assign in378_1 = {c163};
    assign in378_2 = {c164};
    Full_Adder FA_378(s378, c378, in378_1, in378_2, c162);
    wire[0:0] s379, in379_1, in379_2;
    wire c379;
    assign in379_1 = {c166};
    assign in379_2 = {s167[0]};
    Full_Adder FA_379(s379, c379, in379_1, in379_2, c165);
    wire[0:0] s380, in380_1, in380_2;
    wire c380;
    assign in380_1 = {s169[0]};
    assign in380_2 = {s170[0]};
    Full_Adder FA_380(s380, c380, in380_1, in380_2, s168[0]);
    wire[0:0] s381, in381_1, in381_2;
    wire c381;
    assign in381_1 = {s172[0]};
    assign in381_2 = {s173[0]};
    Full_Adder FA_381(s381, c381, in381_1, in381_2, s171[0]);
    wire[0:0] s382, in382_1, in382_2;
    wire c382;
    assign in382_1 = {c167};
    assign in382_2 = {c168};
    Full_Adder FA_382(s382, c382, in382_1, in382_2, s21[0]);
    wire[0:0] s383, in383_1, in383_2;
    wire c383;
    assign in383_1 = {c170};
    assign in383_2 = {c171};
    Full_Adder FA_383(s383, c383, in383_1, in383_2, c169);
    wire[0:0] s384, in384_1, in384_2;
    wire c384;
    assign in384_1 = {c173};
    assign in384_2 = {s174[0]};
    Full_Adder FA_384(s384, c384, in384_1, in384_2, c172);
    wire[0:0] s385, in385_1, in385_2;
    wire c385;
    assign in385_1 = {s176[0]};
    assign in385_2 = {s177[0]};
    Full_Adder FA_385(s385, c385, in385_1, in385_2, s175[0]);
    wire[0:0] s386, in386_1, in386_2;
    wire c386;
    assign in386_1 = {s179[0]};
    assign in386_2 = {s180[0]};
    Full_Adder FA_386(s386, c386, in386_1, in386_2, s178[0]);
    wire[0:0] s387, in387_1, in387_2;
    wire c387;
    assign in387_1 = {c174};
    assign in387_2 = {c175};
    Full_Adder FA_387(s387, c387, in387_1, in387_2, s28[0]);
    wire[0:0] s388, in388_1, in388_2;
    wire c388;
    assign in388_1 = {c177};
    assign in388_2 = {c178};
    Full_Adder FA_388(s388, c388, in388_1, in388_2, c176);
    wire[0:0] s389, in389_1, in389_2;
    wire c389;
    assign in389_1 = {c180};
    assign in389_2 = {s181[0]};
    Full_Adder FA_389(s389, c389, in389_1, in389_2, c179);
    wire[0:0] s390, in390_1, in390_2;
    wire c390;
    assign in390_1 = {s183[0]};
    assign in390_2 = {s184[0]};
    Full_Adder FA_390(s390, c390, in390_1, in390_2, s182[0]);
    wire[0:0] s391, in391_1, in391_2;
    wire c391;
    assign in391_1 = {s186[0]};
    assign in391_2 = {s187[0]};
    Full_Adder FA_391(s391, c391, in391_1, in391_2, s185[0]);
    wire[0:0] s392, in392_1, in392_2;
    wire c392;
    assign in392_1 = {c181};
    assign in392_2 = {c182};
    Full_Adder FA_392(s392, c392, in392_1, in392_2, s36[0]);
    wire[0:0] s393, in393_1, in393_2;
    wire c393;
    assign in393_1 = {c184};
    assign in393_2 = {c185};
    Full_Adder FA_393(s393, c393, in393_1, in393_2, c183);
    wire[0:0] s394, in394_1, in394_2;
    wire c394;
    assign in394_1 = {c187};
    assign in394_2 = {s188[0]};
    Full_Adder FA_394(s394, c394, in394_1, in394_2, c186);
    wire[0:0] s395, in395_1, in395_2;
    wire c395;
    assign in395_1 = {s190[0]};
    assign in395_2 = {s191[0]};
    Full_Adder FA_395(s395, c395, in395_1, in395_2, s189[0]);
    wire[0:0] s396, in396_1, in396_2;
    wire c396;
    assign in396_1 = {s193[0]};
    assign in396_2 = {s194[0]};
    Full_Adder FA_396(s396, c396, in396_1, in396_2, s192[0]);
    wire[0:0] s397, in397_1, in397_2;
    wire c397;
    assign in397_1 = {c188};
    assign in397_2 = {c189};
    Full_Adder FA_397(s397, c397, in397_1, in397_2, s45[0]);
    wire[0:0] s398, in398_1, in398_2;
    wire c398;
    assign in398_1 = {c191};
    assign in398_2 = {c192};
    Full_Adder FA_398(s398, c398, in398_1, in398_2, c190);
    wire[0:0] s399, in399_1, in399_2;
    wire c399;
    assign in399_1 = {c194};
    assign in399_2 = {s195[0]};
    Full_Adder FA_399(s399, c399, in399_1, in399_2, c193);
    wire[0:0] s400, in400_1, in400_2;
    wire c400;
    assign in400_1 = {s197[0]};
    assign in400_2 = {s198[0]};
    Full_Adder FA_400(s400, c400, in400_1, in400_2, s196[0]);
    wire[0:0] s401, in401_1, in401_2;
    wire c401;
    assign in401_1 = {s200[0]};
    assign in401_2 = {s201[0]};
    Full_Adder FA_401(s401, c401, in401_1, in401_2, s199[0]);
    wire[0:0] s402, in402_1, in402_2;
    wire c402;
    assign in402_1 = {c195};
    assign in402_2 = {c196};
    Full_Adder FA_402(s402, c402, in402_1, in402_2, s55[0]);
    wire[0:0] s403, in403_1, in403_2;
    wire c403;
    assign in403_1 = {c198};
    assign in403_2 = {c199};
    Full_Adder FA_403(s403, c403, in403_1, in403_2, c197);
    wire[0:0] s404, in404_1, in404_2;
    wire c404;
    assign in404_1 = {c201};
    assign in404_2 = {s202[0]};
    Full_Adder FA_404(s404, c404, in404_1, in404_2, c200);
    wire[0:0] s405, in405_1, in405_2;
    wire c405;
    assign in405_1 = {s204[0]};
    assign in405_2 = {s205[0]};
    Full_Adder FA_405(s405, c405, in405_1, in405_2, s203[0]);
    wire[0:0] s406, in406_1, in406_2;
    wire c406;
    assign in406_1 = {s207[0]};
    assign in406_2 = {s208[0]};
    Full_Adder FA_406(s406, c406, in406_1, in406_2, s206[0]);
    wire[0:0] s407, in407_1, in407_2;
    wire c407;
    assign in407_1 = {c202};
    assign in407_2 = {c203};
    Full_Adder FA_407(s407, c407, in407_1, in407_2, s65[0]);
    wire[0:0] s408, in408_1, in408_2;
    wire c408;
    assign in408_1 = {c205};
    assign in408_2 = {c206};
    Full_Adder FA_408(s408, c408, in408_1, in408_2, c204);
    wire[0:0] s409, in409_1, in409_2;
    wire c409;
    assign in409_1 = {c208};
    assign in409_2 = {s209[0]};
    Full_Adder FA_409(s409, c409, in409_1, in409_2, c207);
    wire[0:0] s410, in410_1, in410_2;
    wire c410;
    assign in410_1 = {s211[0]};
    assign in410_2 = {s212[0]};
    Full_Adder FA_410(s410, c410, in410_1, in410_2, s210[0]);
    wire[0:0] s411, in411_1, in411_2;
    wire c411;
    assign in411_1 = {s214[0]};
    assign in411_2 = {s215[0]};
    Full_Adder FA_411(s411, c411, in411_1, in411_2, s213[0]);
    wire[0:0] s412, in412_1, in412_2;
    wire c412;
    assign in412_1 = {c209};
    assign in412_2 = {c210};
    Full_Adder FA_412(s412, c412, in412_1, in412_2, s74[0]);
    wire[0:0] s413, in413_1, in413_2;
    wire c413;
    assign in413_1 = {c212};
    assign in413_2 = {c213};
    Full_Adder FA_413(s413, c413, in413_1, in413_2, c211);
    wire[0:0] s414, in414_1, in414_2;
    wire c414;
    assign in414_1 = {c215};
    assign in414_2 = {s216[0]};
    Full_Adder FA_414(s414, c414, in414_1, in414_2, c214);
    wire[0:0] s415, in415_1, in415_2;
    wire c415;
    assign in415_1 = {s218[0]};
    assign in415_2 = {s219[0]};
    Full_Adder FA_415(s415, c415, in415_1, in415_2, s217[0]);
    wire[0:0] s416, in416_1, in416_2;
    wire c416;
    assign in416_1 = {s221[0]};
    assign in416_2 = {s222[0]};
    Full_Adder FA_416(s416, c416, in416_1, in416_2, s220[0]);
    wire[0:0] s417, in417_1, in417_2;
    wire c417;
    assign in417_1 = {c216};
    assign in417_2 = {c217};
    Full_Adder FA_417(s417, c417, in417_1, in417_2, s82[0]);
    wire[0:0] s418, in418_1, in418_2;
    wire c418;
    assign in418_1 = {c219};
    assign in418_2 = {c220};
    Full_Adder FA_418(s418, c418, in418_1, in418_2, c218);
    wire[0:0] s419, in419_1, in419_2;
    wire c419;
    assign in419_1 = {c222};
    assign in419_2 = {s223[0]};
    Full_Adder FA_419(s419, c419, in419_1, in419_2, c221);
    wire[0:0] s420, in420_1, in420_2;
    wire c420;
    assign in420_1 = {s225[0]};
    assign in420_2 = {s226[0]};
    Full_Adder FA_420(s420, c420, in420_1, in420_2, s224[0]);
    wire[0:0] s421, in421_1, in421_2;
    wire c421;
    assign in421_1 = {s228[0]};
    assign in421_2 = {s229[0]};
    Full_Adder FA_421(s421, c421, in421_1, in421_2, s227[0]);
    wire[0:0] s422, in422_1, in422_2;
    wire c422;
    assign in422_1 = {c223};
    assign in422_2 = {c224};
    Full_Adder FA_422(s422, c422, in422_1, in422_2, s89[0]);
    wire[0:0] s423, in423_1, in423_2;
    wire c423;
    assign in423_1 = {c226};
    assign in423_2 = {c227};
    Full_Adder FA_423(s423, c423, in423_1, in423_2, c225);
    wire[0:0] s424, in424_1, in424_2;
    wire c424;
    assign in424_1 = {c229};
    assign in424_2 = {s230[0]};
    Full_Adder FA_424(s424, c424, in424_1, in424_2, c228);
    wire[0:0] s425, in425_1, in425_2;
    wire c425;
    assign in425_1 = {s232[0]};
    assign in425_2 = {s233[0]};
    Full_Adder FA_425(s425, c425, in425_1, in425_2, s231[0]);
    wire[0:0] s426, in426_1, in426_2;
    wire c426;
    assign in426_1 = {s235[0]};
    assign in426_2 = {s236[0]};
    Full_Adder FA_426(s426, c426, in426_1, in426_2, s234[0]);
    wire[0:0] s427, in427_1, in427_2;
    wire c427;
    assign in427_1 = {c230};
    assign in427_2 = {c231};
    Full_Adder FA_427(s427, c427, in427_1, in427_2, s95[0]);
    wire[0:0] s428, in428_1, in428_2;
    wire c428;
    assign in428_1 = {c233};
    assign in428_2 = {c234};
    Full_Adder FA_428(s428, c428, in428_1, in428_2, c232);
    wire[0:0] s429, in429_1, in429_2;
    wire c429;
    assign in429_1 = {c236};
    assign in429_2 = {s237[0]};
    Full_Adder FA_429(s429, c429, in429_1, in429_2, c235);
    wire[0:0] s430, in430_1, in430_2;
    wire c430;
    assign in430_1 = {s239[0]};
    assign in430_2 = {s240[0]};
    Full_Adder FA_430(s430, c430, in430_1, in430_2, s238[0]);
    wire[0:0] s431, in431_1, in431_2;
    wire c431;
    assign in431_1 = {s242[0]};
    assign in431_2 = {s243[0]};
    Full_Adder FA_431(s431, c431, in431_1, in431_2, s241[0]);
    wire[0:0] s432, in432_1, in432_2;
    wire c432;
    assign in432_1 = {c237};
    assign in432_2 = {c238};
    Full_Adder FA_432(s432, c432, in432_1, in432_2, s100[0]);
    wire[0:0] s433, in433_1, in433_2;
    wire c433;
    assign in433_1 = {c240};
    assign in433_2 = {c241};
    Full_Adder FA_433(s433, c433, in433_1, in433_2, c239);
    wire[0:0] s434, in434_1, in434_2;
    wire c434;
    assign in434_1 = {c243};
    assign in434_2 = {s244[0]};
    Full_Adder FA_434(s434, c434, in434_1, in434_2, c242);
    wire[0:0] s435, in435_1, in435_2;
    wire c435;
    assign in435_1 = {s246[0]};
    assign in435_2 = {s247[0]};
    Full_Adder FA_435(s435, c435, in435_1, in435_2, s245[0]);
    wire[0:0] s436, in436_1, in436_2;
    wire c436;
    assign in436_1 = {s249[0]};
    assign in436_2 = {s250[0]};
    Full_Adder FA_436(s436, c436, in436_1, in436_2, s248[0]);
    wire[0:0] s437, in437_1, in437_2;
    wire c437;
    assign in437_1 = {c244};
    assign in437_2 = {c245};
    Full_Adder FA_437(s437, c437, in437_1, in437_2, s104[0]);
    wire[0:0] s438, in438_1, in438_2;
    wire c438;
    assign in438_1 = {c247};
    assign in438_2 = {c248};
    Full_Adder FA_438(s438, c438, in438_1, in438_2, c246);
    wire[0:0] s439, in439_1, in439_2;
    wire c439;
    assign in439_1 = {c250};
    assign in439_2 = {s251[0]};
    Full_Adder FA_439(s439, c439, in439_1, in439_2, c249);
    wire[0:0] s440, in440_1, in440_2;
    wire c440;
    assign in440_1 = {s253[0]};
    assign in440_2 = {s254[0]};
    Full_Adder FA_440(s440, c440, in440_1, in440_2, s252[0]);
    wire[0:0] s441, in441_1, in441_2;
    wire c441;
    assign in441_1 = {s256[0]};
    assign in441_2 = {s257[0]};
    Full_Adder FA_441(s441, c441, in441_1, in441_2, s255[0]);
    wire[0:0] s442, in442_1, in442_2;
    wire c442;
    assign in442_1 = {c251};
    assign in442_2 = {c252};
    Full_Adder FA_442(s442, c442, in442_1, in442_2, s107[0]);
    wire[0:0] s443, in443_1, in443_2;
    wire c443;
    assign in443_1 = {c254};
    assign in443_2 = {c255};
    Full_Adder FA_443(s443, c443, in443_1, in443_2, c253);
    wire[0:0] s444, in444_1, in444_2;
    wire c444;
    assign in444_1 = {c257};
    assign in444_2 = {s258[0]};
    Full_Adder FA_444(s444, c444, in444_1, in444_2, c256);
    wire[0:0] s445, in445_1, in445_2;
    wire c445;
    assign in445_1 = {s260[0]};
    assign in445_2 = {s261[0]};
    Full_Adder FA_445(s445, c445, in445_1, in445_2, s259[0]);
    wire[0:0] s446, in446_1, in446_2;
    wire c446;
    assign in446_1 = {s263[0]};
    assign in446_2 = {s264[0]};
    Full_Adder FA_446(s446, c446, in446_1, in446_2, s262[0]);
    wire[0:0] s447, in447_1, in447_2;
    wire c447;
    assign in447_1 = {c258};
    assign in447_2 = {c259};
    Full_Adder FA_447(s447, c447, in447_1, in447_2, s109[0]);
    wire[0:0] s448, in448_1, in448_2;
    wire c448;
    assign in448_1 = {c261};
    assign in448_2 = {c262};
    Full_Adder FA_448(s448, c448, in448_1, in448_2, c260);
    wire[0:0] s449, in449_1, in449_2;
    wire c449;
    assign in449_1 = {c264};
    assign in449_2 = {s265[0]};
    Full_Adder FA_449(s449, c449, in449_1, in449_2, c263);
    wire[0:0] s450, in450_1, in450_2;
    wire c450;
    assign in450_1 = {s267[0]};
    assign in450_2 = {s268[0]};
    Full_Adder FA_450(s450, c450, in450_1, in450_2, s266[0]);
    wire[0:0] s451, in451_1, in451_2;
    wire c451;
    assign in451_1 = {s270[0]};
    assign in451_2 = {s271[0]};
    Full_Adder FA_451(s451, c451, in451_1, in451_2, s269[0]);
    wire[0:0] s452, in452_1, in452_2;
    wire c452;
    assign in452_1 = {c265};
    assign in452_2 = {c266};
    Full_Adder FA_452(s452, c452, in452_1, in452_2, s110[0]);
    wire[0:0] s453, in453_1, in453_2;
    wire c453;
    assign in453_1 = {c268};
    assign in453_2 = {c269};
    Full_Adder FA_453(s453, c453, in453_1, in453_2, c267);
    wire[0:0] s454, in454_1, in454_2;
    wire c454;
    assign in454_1 = {c271};
    assign in454_2 = {s272[0]};
    Full_Adder FA_454(s454, c454, in454_1, in454_2, c270);
    wire[0:0] s455, in455_1, in455_2;
    wire c455;
    assign in455_1 = {s274[0]};
    assign in455_2 = {s275[0]};
    Full_Adder FA_455(s455, c455, in455_1, in455_2, s273[0]);
    wire[0:0] s456, in456_1, in456_2;
    wire c456;
    assign in456_1 = {s277[0]};
    assign in456_2 = {s278[0]};
    Full_Adder FA_456(s456, c456, in456_1, in456_2, s276[0]);
    wire[0:0] s457, in457_1, in457_2;
    wire c457;
    assign in457_1 = {c272};
    assign in457_2 = {c273};
    Full_Adder FA_457(s457, c457, in457_1, in457_2, c110);
    wire[0:0] s458, in458_1, in458_2;
    wire c458;
    assign in458_1 = {c275};
    assign in458_2 = {c276};
    Full_Adder FA_458(s458, c458, in458_1, in458_2, c274);
    wire[0:0] s459, in459_1, in459_2;
    wire c459;
    assign in459_1 = {c278};
    assign in459_2 = {s279[0]};
    Full_Adder FA_459(s459, c459, in459_1, in459_2, c277);
    wire[0:0] s460, in460_1, in460_2;
    wire c460;
    assign in460_1 = {s281[0]};
    assign in460_2 = {s282[0]};
    Full_Adder FA_460(s460, c460, in460_1, in460_2, s280[0]);
    wire[0:0] s461, in461_1, in461_2;
    wire c461;
    assign in461_1 = {s284[0]};
    assign in461_2 = {s285[0]};
    Full_Adder FA_461(s461, c461, in461_1, in461_2, s283[0]);
    wire[0:0] s462, in462_1, in462_2;
    wire c462;
    assign in462_1 = {pp31[12]};
    assign in462_2 = {c279};
    Full_Adder FA_462(s462, c462, in462_1, in462_2, pp30[13]);
    wire[0:0] s463, in463_1, in463_2;
    wire c463;
    assign in463_1 = {c281};
    assign in463_2 = {c282};
    Full_Adder FA_463(s463, c463, in463_1, in463_2, c280);
    wire[0:0] s464, in464_1, in464_2;
    wire c464;
    assign in464_1 = {c284};
    assign in464_2 = {c285};
    Full_Adder FA_464(s464, c464, in464_1, in464_2, c283);
    wire[0:0] s465, in465_1, in465_2;
    wire c465;
    assign in465_1 = {s287[0]};
    assign in465_2 = {s288[0]};
    Full_Adder FA_465(s465, c465, in465_1, in465_2, s286[0]);
    wire[0:0] s466, in466_1, in466_2;
    wire c466;
    assign in466_1 = {s290[0]};
    assign in466_2 = {s291[0]};
    Full_Adder FA_466(s466, c466, in466_1, in466_2, s289[0]);
    wire[0:0] s467, in467_1, in467_2;
    wire c467;
    assign in467_1 = {pp29[15]};
    assign in467_2 = {pp30[14]};
    Full_Adder FA_467(s467, c467, in467_1, in467_2, pp28[16]);
    wire[0:0] s468, in468_1, in468_2;
    wire c468;
    assign in468_1 = {c286};
    assign in468_2 = {c287};
    Full_Adder FA_468(s468, c468, in468_1, in468_2, pp31[13]);
    wire[0:0] s469, in469_1, in469_2;
    wire c469;
    assign in469_1 = {c289};
    assign in469_2 = {c290};
    Full_Adder FA_469(s469, c469, in469_1, in469_2, c288);
    wire[0:0] s470, in470_1, in470_2;
    wire c470;
    assign in470_1 = {s292[0]};
    assign in470_2 = {s293[0]};
    Full_Adder FA_470(s470, c470, in470_1, in470_2, c291);
    wire[0:0] s471, in471_1, in471_2;
    wire c471;
    assign in471_1 = {s295[0]};
    assign in471_2 = {s296[0]};
    Full_Adder FA_471(s471, c471, in471_1, in471_2, s294[0]);
    wire[0:0] s472, in472_1, in472_2;
    wire c472;
    assign in472_1 = {pp27[18]};
    assign in472_2 = {pp28[17]};
    Full_Adder FA_472(s472, c472, in472_1, in472_2, pp26[19]);
    wire[0:0] s473, in473_1, in473_2;
    wire c473;
    assign in473_1 = {pp30[15]};
    assign in473_2 = {pp31[14]};
    Full_Adder FA_473(s473, c473, in473_1, in473_2, pp29[16]);
    wire[0:0] s474, in474_1, in474_2;
    wire c474;
    assign in474_1 = {c293};
    assign in474_2 = {c294};
    Full_Adder FA_474(s474, c474, in474_1, in474_2, c292);
    wire[0:0] s475, in475_1, in475_2;
    wire c475;
    assign in475_1 = {c296};
    assign in475_2 = {s297[0]};
    Full_Adder FA_475(s475, c475, in475_1, in475_2, c295);
    wire[0:0] s476, in476_1, in476_2;
    wire c476;
    assign in476_1 = {s299[0]};
    assign in476_2 = {s300[0]};
    Full_Adder FA_476(s476, c476, in476_1, in476_2, s298[0]);
    wire[0:0] s477, in477_1, in477_2;
    wire c477;
    assign in477_1 = {pp25[21]};
    assign in477_2 = {pp26[20]};
    Full_Adder FA_477(s477, c477, in477_1, in477_2, pp24[22]);
    wire[0:0] s478, in478_1, in478_2;
    wire c478;
    assign in478_1 = {pp28[18]};
    assign in478_2 = {pp29[17]};
    Full_Adder FA_478(s478, c478, in478_1, in478_2, pp27[19]);
    wire[0:0] s479, in479_1, in479_2;
    wire c479;
    assign in479_1 = {pp31[15]};
    assign in479_2 = {c297};
    Full_Adder FA_479(s479, c479, in479_1, in479_2, pp30[16]);
    wire[0:0] s480, in480_1, in480_2;
    wire c480;
    assign in480_1 = {c299};
    assign in480_2 = {c300};
    Full_Adder FA_480(s480, c480, in480_1, in480_2, c298);
    wire[0:0] s481, in481_1, in481_2;
    wire c481;
    assign in481_1 = {s302[0]};
    assign in481_2 = {s303[0]};
    Full_Adder FA_481(s481, c481, in481_1, in481_2, s301[0]);
    wire[0:0] s482, in482_1, in482_2;
    wire c482;
    assign in482_1 = {pp23[24]};
    assign in482_2 = {pp24[23]};
    Full_Adder FA_482(s482, c482, in482_1, in482_2, pp22[25]);
    wire[0:0] s483, in483_1, in483_2;
    wire c483;
    assign in483_1 = {pp26[21]};
    assign in483_2 = {pp27[20]};
    Full_Adder FA_483(s483, c483, in483_1, in483_2, pp25[22]);
    wire[0:0] s484, in484_1, in484_2;
    wire c484;
    assign in484_1 = {pp29[18]};
    assign in484_2 = {pp30[17]};
    Full_Adder FA_484(s484, c484, in484_1, in484_2, pp28[19]);
    wire[0:0] s485, in485_1, in485_2;
    wire c485;
    assign in485_1 = {c301};
    assign in485_2 = {c302};
    Full_Adder FA_485(s485, c485, in485_1, in485_2, pp31[16]);
    wire[0:0] s486, in486_1, in486_2;
    wire c486;
    assign in486_1 = {s304[0]};
    assign in486_2 = {s305[0]};
    Full_Adder FA_486(s486, c486, in486_1, in486_2, c303);
    wire[0:0] s487, in487_1, in487_2;
    wire c487;
    assign in487_1 = {pp21[27]};
    assign in487_2 = {pp22[26]};
    Full_Adder FA_487(s487, c487, in487_1, in487_2, pp20[28]);
    wire[0:0] s488, in488_1, in488_2;
    wire c488;
    assign in488_1 = {pp24[24]};
    assign in488_2 = {pp25[23]};
    Full_Adder FA_488(s488, c488, in488_1, in488_2, pp23[25]);
    wire[0:0] s489, in489_1, in489_2;
    wire c489;
    assign in489_1 = {pp27[21]};
    assign in489_2 = {pp28[20]};
    Full_Adder FA_489(s489, c489, in489_1, in489_2, pp26[22]);
    wire[0:0] s490, in490_1, in490_2;
    wire c490;
    assign in490_1 = {pp30[18]};
    assign in490_2 = {pp31[17]};
    Full_Adder FA_490(s490, c490, in490_1, in490_2, pp29[19]);
    wire[0:0] s491, in491_1, in491_2;
    wire c491;
    assign in491_1 = {c305};
    assign in491_2 = {s306[0]};
    Full_Adder FA_491(s491, c491, in491_1, in491_2, c304);
    wire[0:0] s492, in492_1, in492_2;
    wire c492;
    assign in492_1 = {pp19[30]};
    assign in492_2 = {pp20[29]};
    Full_Adder FA_492(s492, c492, in492_1, in492_2, pp18[31]);
    wire[0:0] s493, in493_1, in493_2;
    wire c493;
    assign in493_1 = {pp22[27]};
    assign in493_2 = {pp23[26]};
    Full_Adder FA_493(s493, c493, in493_1, in493_2, pp21[28]);
    wire[0:0] s494, in494_1, in494_2;
    wire c494;
    assign in494_1 = {pp25[24]};
    assign in494_2 = {pp26[23]};
    Full_Adder FA_494(s494, c494, in494_1, in494_2, pp24[25]);
    wire[0:0] s495, in495_1, in495_2;
    wire c495;
    assign in495_1 = {pp28[21]};
    assign in495_2 = {pp29[20]};
    Full_Adder FA_495(s495, c495, in495_1, in495_2, pp27[22]);
    wire[0:0] s496, in496_1, in496_2;
    wire c496;
    assign in496_1 = {pp31[18]};
    assign in496_2 = {c306};
    Full_Adder FA_496(s496, c496, in496_1, in496_2, pp30[19]);
    wire[0:0] s497, in497_1, in497_2;
    wire c497;
    assign in497_1 = {pp20[30]};
    assign in497_2 = {pp21[29]};
    Full_Adder FA_497(s497, c497, in497_1, in497_2, pp19[31]);
    wire[0:0] s498, in498_1, in498_2;
    wire c498;
    assign in498_1 = {pp23[27]};
    assign in498_2 = {pp24[26]};
    Full_Adder FA_498(s498, c498, in498_1, in498_2, pp22[28]);
    wire[0:0] s499, in499_1, in499_2;
    wire c499;
    assign in499_1 = {pp26[24]};
    assign in499_2 = {pp27[23]};
    Full_Adder FA_499(s499, c499, in499_1, in499_2, pp25[25]);
    wire[0:0] s500, in500_1, in500_2;
    wire c500;
    assign in500_1 = {pp29[21]};
    assign in500_2 = {pp30[20]};
    Full_Adder FA_500(s500, c500, in500_1, in500_2, pp28[22]);
    wire[0:0] s501, in501_1, in501_2;
    wire c501;
    assign in501_1 = {pp21[30]};
    assign in501_2 = {pp22[29]};
    Full_Adder FA_501(s501, c501, in501_1, in501_2, pp20[31]);
    wire[0:0] s502, in502_1, in502_2;
    wire c502;
    assign in502_1 = {pp24[27]};
    assign in502_2 = {pp25[26]};
    Full_Adder FA_502(s502, c502, in502_1, in502_2, pp23[28]);
    wire[0:0] s503, in503_1, in503_2;
    wire c503;
    assign in503_1 = {pp27[24]};
    assign in503_2 = {pp28[23]};
    Full_Adder FA_503(s503, c503, in503_1, in503_2, pp26[25]);
    wire[0:0] s504, in504_1, in504_2;
    wire c504;
    assign in504_1 = {pp22[30]};
    assign in504_2 = {pp23[29]};
    Full_Adder FA_504(s504, c504, in504_1, in504_2, pp21[31]);
    wire[0:0] s505, in505_1, in505_2;
    wire c505;
    assign in505_1 = {pp25[27]};
    assign in505_2 = {pp26[26]};
    Full_Adder FA_505(s505, c505, in505_1, in505_2, pp24[28]);
    wire[0:0] s506, in506_1, in506_2;
    wire c506;
    assign in506_1 = {pp23[30]};
    assign in506_2 = {pp24[29]};
    Full_Adder FA_506(s506, c506, in506_1, in506_2, pp22[31]);

    /*Stage 4*/
    wire[0:0] s507, in507_1, in507_2;
    wire c507;
    assign in507_1 = {pp0[7]};
    assign in507_2 = {pp1[6]};
    Half_Adder HA_507(s507, c507, in507_1, in507_2);
    wire[0:0] s508, in508_1, in508_2;
    wire c508;
    assign in508_1 = {pp1[7]};
    assign in508_2 = {pp2[6]};
    Full_Adder FA_508(s508, c508, in508_1, in508_2, pp0[8]);
    wire[0:0] s509, in509_1, in509_2;
    wire c509;
    assign in509_1 = {pp3[5]};
    assign in509_2 = {pp4[4]};
    Half_Adder HA_509(s509, c509, in509_1, in509_2);
    wire[0:0] s510, in510_1, in510_2;
    wire c510;
    assign in510_1 = {pp1[8]};
    assign in510_2 = {pp2[7]};
    Full_Adder FA_510(s510, c510, in510_1, in510_2, pp0[9]);
    wire[0:0] s511, in511_1, in511_2;
    wire c511;
    assign in511_1 = {pp4[5]};
    assign in511_2 = {pp5[4]};
    Full_Adder FA_511(s511, c511, in511_1, in511_2, pp3[6]);
    wire[0:0] s512, in512_1, in512_2;
    wire c512;
    assign in512_1 = {pp6[3]};
    assign in512_2 = {pp7[2]};
    Half_Adder HA_512(s512, c512, in512_1, in512_2);
    wire[0:0] s513, in513_1, in513_2;
    wire c513;
    assign in513_1 = {pp3[7]};
    assign in513_2 = {pp4[6]};
    Full_Adder FA_513(s513, c513, in513_1, in513_2, pp2[8]);
    wire[0:0] s514, in514_1, in514_2;
    wire c514;
    assign in514_1 = {pp6[4]};
    assign in514_2 = {pp7[3]};
    Full_Adder FA_514(s514, c514, in514_1, in514_2, pp5[5]);
    wire[0:0] s515, in515_1, in515_2;
    wire c515;
    assign in515_1 = {pp9[1]};
    assign in515_2 = {pp10[0]};
    Full_Adder FA_515(s515, c515, in515_1, in515_2, pp8[2]);
    wire[0:0] s516, in516_1, in516_2;
    wire c516;
    assign in516_1 = {pp6[5]};
    assign in516_2 = {pp7[4]};
    Full_Adder FA_516(s516, c516, in516_1, in516_2, pp5[6]);
    wire[0:0] s517, in517_1, in517_2;
    wire c517;
    assign in517_1 = {pp9[2]};
    assign in517_2 = {pp10[1]};
    Full_Adder FA_517(s517, c517, in517_1, in517_2, pp8[3]);
    wire[0:0] s518, in518_1, in518_2;
    wire c518;
    assign in518_1 = {c307};
    assign in518_2 = {s308[0]};
    Full_Adder FA_518(s518, c518, in518_1, in518_2, pp11[0]);
    wire[0:0] s519, in519_1, in519_2;
    wire c519;
    assign in519_1 = {pp9[3]};
    assign in519_2 = {pp10[2]};
    Full_Adder FA_519(s519, c519, in519_1, in519_2, pp8[4]);
    wire[0:0] s520, in520_1, in520_2;
    wire c520;
    assign in520_1 = {pp12[0]};
    assign in520_2 = {c308};
    Full_Adder FA_520(s520, c520, in520_1, in520_2, pp11[1]);
    wire[0:0] s521, in521_1, in521_2;
    wire c521;
    assign in521_1 = {s310[0]};
    assign in521_2 = {s311[0]};
    Full_Adder FA_521(s521, c521, in521_1, in521_2, c309);
    wire[0:0] s522, in522_1, in522_2;
    wire c522;
    assign in522_1 = {pp12[1]};
    assign in522_2 = {pp13[0]};
    Full_Adder FA_522(s522, c522, in522_1, in522_2, pp11[2]);
    wire[0:0] s523, in523_1, in523_2;
    wire c523;
    assign in523_1 = {c311};
    assign in523_2 = {c312};
    Full_Adder FA_523(s523, c523, in523_1, in523_2, c310);
    wire[0:0] s524, in524_1, in524_2;
    wire c524;
    assign in524_1 = {s314[0]};
    assign in524_2 = {s315[0]};
    Full_Adder FA_524(s524, c524, in524_1, in524_2, s313[0]);
    wire[0:0] s525, in525_1, in525_2;
    wire c525;
    assign in525_1 = {c313};
    assign in525_2 = {c314};
    Full_Adder FA_525(s525, c525, in525_1, in525_2, pp14[0]);
    wire[0:0] s526, in526_1, in526_2;
    wire c526;
    assign in526_1 = {c316};
    assign in526_2 = {s317[0]};
    Full_Adder FA_526(s526, c526, in526_1, in526_2, c315);
    wire[0:0] s527, in527_1, in527_2;
    wire c527;
    assign in527_1 = {s319[0]};
    assign in527_2 = {s320[0]};
    Full_Adder FA_527(s527, c527, in527_1, in527_2, s318[0]);
    wire[0:0] s528, in528_1, in528_2;
    wire c528;
    assign in528_1 = {c318};
    assign in528_2 = {c319};
    Full_Adder FA_528(s528, c528, in528_1, in528_2, c317);
    wire[0:0] s529, in529_1, in529_2;
    wire c529;
    assign in529_1 = {c321};
    assign in529_2 = {s322[0]};
    Full_Adder FA_529(s529, c529, in529_1, in529_2, c320);
    wire[0:0] s530, in530_1, in530_2;
    wire c530;
    assign in530_1 = {s324[0]};
    assign in530_2 = {s325[0]};
    Full_Adder FA_530(s530, c530, in530_1, in530_2, s323[0]);
    wire[0:0] s531, in531_1, in531_2;
    wire c531;
    assign in531_1 = {c323};
    assign in531_2 = {c324};
    Full_Adder FA_531(s531, c531, in531_1, in531_2, c322);
    wire[0:0] s532, in532_1, in532_2;
    wire c532;
    assign in532_1 = {c326};
    assign in532_2 = {s327[0]};
    Full_Adder FA_532(s532, c532, in532_1, in532_2, c325);
    wire[0:0] s533, in533_1, in533_2;
    wire c533;
    assign in533_1 = {s329[0]};
    assign in533_2 = {s330[0]};
    Full_Adder FA_533(s533, c533, in533_1, in533_2, s328[0]);
    wire[0:0] s534, in534_1, in534_2;
    wire c534;
    assign in534_1 = {c328};
    assign in534_2 = {c329};
    Full_Adder FA_534(s534, c534, in534_1, in534_2, c327);
    wire[0:0] s535, in535_1, in535_2;
    wire c535;
    assign in535_1 = {c331};
    assign in535_2 = {s332[0]};
    Full_Adder FA_535(s535, c535, in535_1, in535_2, c330);
    wire[0:0] s536, in536_1, in536_2;
    wire c536;
    assign in536_1 = {s334[0]};
    assign in536_2 = {s335[0]};
    Full_Adder FA_536(s536, c536, in536_1, in536_2, s333[0]);
    wire[0:0] s537, in537_1, in537_2;
    wire c537;
    assign in537_1 = {c333};
    assign in537_2 = {c334};
    Full_Adder FA_537(s537, c537, in537_1, in537_2, c332);
    wire[0:0] s538, in538_1, in538_2;
    wire c538;
    assign in538_1 = {c336};
    assign in538_2 = {s337[0]};
    Full_Adder FA_538(s538, c538, in538_1, in538_2, c335);
    wire[0:0] s539, in539_1, in539_2;
    wire c539;
    assign in539_1 = {s339[0]};
    assign in539_2 = {s340[0]};
    Full_Adder FA_539(s539, c539, in539_1, in539_2, s338[0]);
    wire[0:0] s540, in540_1, in540_2;
    wire c540;
    assign in540_1 = {c338};
    assign in540_2 = {c339};
    Full_Adder FA_540(s540, c540, in540_1, in540_2, c337);
    wire[0:0] s541, in541_1, in541_2;
    wire c541;
    assign in541_1 = {c341};
    assign in541_2 = {s342[0]};
    Full_Adder FA_541(s541, c541, in541_1, in541_2, c340);
    wire[0:0] s542, in542_1, in542_2;
    wire c542;
    assign in542_1 = {s344[0]};
    assign in542_2 = {s345[0]};
    Full_Adder FA_542(s542, c542, in542_1, in542_2, s343[0]);
    wire[0:0] s543, in543_1, in543_2;
    wire c543;
    assign in543_1 = {c343};
    assign in543_2 = {c344};
    Full_Adder FA_543(s543, c543, in543_1, in543_2, c342);
    wire[0:0] s544, in544_1, in544_2;
    wire c544;
    assign in544_1 = {c346};
    assign in544_2 = {s347[0]};
    Full_Adder FA_544(s544, c544, in544_1, in544_2, c345);
    wire[0:0] s545, in545_1, in545_2;
    wire c545;
    assign in545_1 = {s349[0]};
    assign in545_2 = {s350[0]};
    Full_Adder FA_545(s545, c545, in545_1, in545_2, s348[0]);
    wire[0:0] s546, in546_1, in546_2;
    wire c546;
    assign in546_1 = {c348};
    assign in546_2 = {c349};
    Full_Adder FA_546(s546, c546, in546_1, in546_2, c347);
    wire[0:0] s547, in547_1, in547_2;
    wire c547;
    assign in547_1 = {c351};
    assign in547_2 = {s352[0]};
    Full_Adder FA_547(s547, c547, in547_1, in547_2, c350);
    wire[0:0] s548, in548_1, in548_2;
    wire c548;
    assign in548_1 = {s354[0]};
    assign in548_2 = {s355[0]};
    Full_Adder FA_548(s548, c548, in548_1, in548_2, s353[0]);
    wire[0:0] s549, in549_1, in549_2;
    wire c549;
    assign in549_1 = {c353};
    assign in549_2 = {c354};
    Full_Adder FA_549(s549, c549, in549_1, in549_2, c352);
    wire[0:0] s550, in550_1, in550_2;
    wire c550;
    assign in550_1 = {c356};
    assign in550_2 = {s357[0]};
    Full_Adder FA_550(s550, c550, in550_1, in550_2, c355);
    wire[0:0] s551, in551_1, in551_2;
    wire c551;
    assign in551_1 = {s359[0]};
    assign in551_2 = {s360[0]};
    Full_Adder FA_551(s551, c551, in551_1, in551_2, s358[0]);
    wire[0:0] s552, in552_1, in552_2;
    wire c552;
    assign in552_1 = {c358};
    assign in552_2 = {c359};
    Full_Adder FA_552(s552, c552, in552_1, in552_2, c357);
    wire[0:0] s553, in553_1, in553_2;
    wire c553;
    assign in553_1 = {c361};
    assign in553_2 = {s362[0]};
    Full_Adder FA_553(s553, c553, in553_1, in553_2, c360);
    wire[0:0] s554, in554_1, in554_2;
    wire c554;
    assign in554_1 = {s364[0]};
    assign in554_2 = {s365[0]};
    Full_Adder FA_554(s554, c554, in554_1, in554_2, s363[0]);
    wire[0:0] s555, in555_1, in555_2;
    wire c555;
    assign in555_1 = {c363};
    assign in555_2 = {c364};
    Full_Adder FA_555(s555, c555, in555_1, in555_2, c362);
    wire[0:0] s556, in556_1, in556_2;
    wire c556;
    assign in556_1 = {c366};
    assign in556_2 = {s367[0]};
    Full_Adder FA_556(s556, c556, in556_1, in556_2, c365);
    wire[0:0] s557, in557_1, in557_2;
    wire c557;
    assign in557_1 = {s369[0]};
    assign in557_2 = {s370[0]};
    Full_Adder FA_557(s557, c557, in557_1, in557_2, s368[0]);
    wire[0:0] s558, in558_1, in558_2;
    wire c558;
    assign in558_1 = {c368};
    assign in558_2 = {c369};
    Full_Adder FA_558(s558, c558, in558_1, in558_2, c367);
    wire[0:0] s559, in559_1, in559_2;
    wire c559;
    assign in559_1 = {c371};
    assign in559_2 = {s372[0]};
    Full_Adder FA_559(s559, c559, in559_1, in559_2, c370);
    wire[0:0] s560, in560_1, in560_2;
    wire c560;
    assign in560_1 = {s374[0]};
    assign in560_2 = {s375[0]};
    Full_Adder FA_560(s560, c560, in560_1, in560_2, s373[0]);
    wire[0:0] s561, in561_1, in561_2;
    wire c561;
    assign in561_1 = {c373};
    assign in561_2 = {c374};
    Full_Adder FA_561(s561, c561, in561_1, in561_2, c372);
    wire[0:0] s562, in562_1, in562_2;
    wire c562;
    assign in562_1 = {c376};
    assign in562_2 = {s377[0]};
    Full_Adder FA_562(s562, c562, in562_1, in562_2, c375);
    wire[0:0] s563, in563_1, in563_2;
    wire c563;
    assign in563_1 = {s379[0]};
    assign in563_2 = {s380[0]};
    Full_Adder FA_563(s563, c563, in563_1, in563_2, s378[0]);
    wire[0:0] s564, in564_1, in564_2;
    wire c564;
    assign in564_1 = {c378};
    assign in564_2 = {c379};
    Full_Adder FA_564(s564, c564, in564_1, in564_2, c377);
    wire[0:0] s565, in565_1, in565_2;
    wire c565;
    assign in565_1 = {c381};
    assign in565_2 = {s382[0]};
    Full_Adder FA_565(s565, c565, in565_1, in565_2, c380);
    wire[0:0] s566, in566_1, in566_2;
    wire c566;
    assign in566_1 = {s384[0]};
    assign in566_2 = {s385[0]};
    Full_Adder FA_566(s566, c566, in566_1, in566_2, s383[0]);
    wire[0:0] s567, in567_1, in567_2;
    wire c567;
    assign in567_1 = {c383};
    assign in567_2 = {c384};
    Full_Adder FA_567(s567, c567, in567_1, in567_2, c382);
    wire[0:0] s568, in568_1, in568_2;
    wire c568;
    assign in568_1 = {c386};
    assign in568_2 = {s387[0]};
    Full_Adder FA_568(s568, c568, in568_1, in568_2, c385);
    wire[0:0] s569, in569_1, in569_2;
    wire c569;
    assign in569_1 = {s389[0]};
    assign in569_2 = {s390[0]};
    Full_Adder FA_569(s569, c569, in569_1, in569_2, s388[0]);
    wire[0:0] s570, in570_1, in570_2;
    wire c570;
    assign in570_1 = {c388};
    assign in570_2 = {c389};
    Full_Adder FA_570(s570, c570, in570_1, in570_2, c387);
    wire[0:0] s571, in571_1, in571_2;
    wire c571;
    assign in571_1 = {c391};
    assign in571_2 = {s392[0]};
    Full_Adder FA_571(s571, c571, in571_1, in571_2, c390);
    wire[0:0] s572, in572_1, in572_2;
    wire c572;
    assign in572_1 = {s394[0]};
    assign in572_2 = {s395[0]};
    Full_Adder FA_572(s572, c572, in572_1, in572_2, s393[0]);
    wire[0:0] s573, in573_1, in573_2;
    wire c573;
    assign in573_1 = {c393};
    assign in573_2 = {c394};
    Full_Adder FA_573(s573, c573, in573_1, in573_2, c392);
    wire[0:0] s574, in574_1, in574_2;
    wire c574;
    assign in574_1 = {c396};
    assign in574_2 = {s397[0]};
    Full_Adder FA_574(s574, c574, in574_1, in574_2, c395);
    wire[0:0] s575, in575_1, in575_2;
    wire c575;
    assign in575_1 = {s399[0]};
    assign in575_2 = {s400[0]};
    Full_Adder FA_575(s575, c575, in575_1, in575_2, s398[0]);
    wire[0:0] s576, in576_1, in576_2;
    wire c576;
    assign in576_1 = {c398};
    assign in576_2 = {c399};
    Full_Adder FA_576(s576, c576, in576_1, in576_2, c397);
    wire[0:0] s577, in577_1, in577_2;
    wire c577;
    assign in577_1 = {c401};
    assign in577_2 = {s402[0]};
    Full_Adder FA_577(s577, c577, in577_1, in577_2, c400);
    wire[0:0] s578, in578_1, in578_2;
    wire c578;
    assign in578_1 = {s404[0]};
    assign in578_2 = {s405[0]};
    Full_Adder FA_578(s578, c578, in578_1, in578_2, s403[0]);
    wire[0:0] s579, in579_1, in579_2;
    wire c579;
    assign in579_1 = {c403};
    assign in579_2 = {c404};
    Full_Adder FA_579(s579, c579, in579_1, in579_2, c402);
    wire[0:0] s580, in580_1, in580_2;
    wire c580;
    assign in580_1 = {c406};
    assign in580_2 = {s407[0]};
    Full_Adder FA_580(s580, c580, in580_1, in580_2, c405);
    wire[0:0] s581, in581_1, in581_2;
    wire c581;
    assign in581_1 = {s409[0]};
    assign in581_2 = {s410[0]};
    Full_Adder FA_581(s581, c581, in581_1, in581_2, s408[0]);
    wire[0:0] s582, in582_1, in582_2;
    wire c582;
    assign in582_1 = {c408};
    assign in582_2 = {c409};
    Full_Adder FA_582(s582, c582, in582_1, in582_2, c407);
    wire[0:0] s583, in583_1, in583_2;
    wire c583;
    assign in583_1 = {c411};
    assign in583_2 = {s412[0]};
    Full_Adder FA_583(s583, c583, in583_1, in583_2, c410);
    wire[0:0] s584, in584_1, in584_2;
    wire c584;
    assign in584_1 = {s414[0]};
    assign in584_2 = {s415[0]};
    Full_Adder FA_584(s584, c584, in584_1, in584_2, s413[0]);
    wire[0:0] s585, in585_1, in585_2;
    wire c585;
    assign in585_1 = {c413};
    assign in585_2 = {c414};
    Full_Adder FA_585(s585, c585, in585_1, in585_2, c412);
    wire[0:0] s586, in586_1, in586_2;
    wire c586;
    assign in586_1 = {c416};
    assign in586_2 = {s417[0]};
    Full_Adder FA_586(s586, c586, in586_1, in586_2, c415);
    wire[0:0] s587, in587_1, in587_2;
    wire c587;
    assign in587_1 = {s419[0]};
    assign in587_2 = {s420[0]};
    Full_Adder FA_587(s587, c587, in587_1, in587_2, s418[0]);
    wire[0:0] s588, in588_1, in588_2;
    wire c588;
    assign in588_1 = {c418};
    assign in588_2 = {c419};
    Full_Adder FA_588(s588, c588, in588_1, in588_2, c417);
    wire[0:0] s589, in589_1, in589_2;
    wire c589;
    assign in589_1 = {c421};
    assign in589_2 = {s422[0]};
    Full_Adder FA_589(s589, c589, in589_1, in589_2, c420);
    wire[0:0] s590, in590_1, in590_2;
    wire c590;
    assign in590_1 = {s424[0]};
    assign in590_2 = {s425[0]};
    Full_Adder FA_590(s590, c590, in590_1, in590_2, s423[0]);
    wire[0:0] s591, in591_1, in591_2;
    wire c591;
    assign in591_1 = {c423};
    assign in591_2 = {c424};
    Full_Adder FA_591(s591, c591, in591_1, in591_2, c422);
    wire[0:0] s592, in592_1, in592_2;
    wire c592;
    assign in592_1 = {c426};
    assign in592_2 = {s427[0]};
    Full_Adder FA_592(s592, c592, in592_1, in592_2, c425);
    wire[0:0] s593, in593_1, in593_2;
    wire c593;
    assign in593_1 = {s429[0]};
    assign in593_2 = {s430[0]};
    Full_Adder FA_593(s593, c593, in593_1, in593_2, s428[0]);
    wire[0:0] s594, in594_1, in594_2;
    wire c594;
    assign in594_1 = {c428};
    assign in594_2 = {c429};
    Full_Adder FA_594(s594, c594, in594_1, in594_2, c427);
    wire[0:0] s595, in595_1, in595_2;
    wire c595;
    assign in595_1 = {c431};
    assign in595_2 = {s432[0]};
    Full_Adder FA_595(s595, c595, in595_1, in595_2, c430);
    wire[0:0] s596, in596_1, in596_2;
    wire c596;
    assign in596_1 = {s434[0]};
    assign in596_2 = {s435[0]};
    Full_Adder FA_596(s596, c596, in596_1, in596_2, s433[0]);
    wire[0:0] s597, in597_1, in597_2;
    wire c597;
    assign in597_1 = {c433};
    assign in597_2 = {c434};
    Full_Adder FA_597(s597, c597, in597_1, in597_2, c432);
    wire[0:0] s598, in598_1, in598_2;
    wire c598;
    assign in598_1 = {c436};
    assign in598_2 = {s437[0]};
    Full_Adder FA_598(s598, c598, in598_1, in598_2, c435);
    wire[0:0] s599, in599_1, in599_2;
    wire c599;
    assign in599_1 = {s439[0]};
    assign in599_2 = {s440[0]};
    Full_Adder FA_599(s599, c599, in599_1, in599_2, s438[0]);
    wire[0:0] s600, in600_1, in600_2;
    wire c600;
    assign in600_1 = {c438};
    assign in600_2 = {c439};
    Full_Adder FA_600(s600, c600, in600_1, in600_2, c437);
    wire[0:0] s601, in601_1, in601_2;
    wire c601;
    assign in601_1 = {c441};
    assign in601_2 = {s442[0]};
    Full_Adder FA_601(s601, c601, in601_1, in601_2, c440);
    wire[0:0] s602, in602_1, in602_2;
    wire c602;
    assign in602_1 = {s444[0]};
    assign in602_2 = {s445[0]};
    Full_Adder FA_602(s602, c602, in602_1, in602_2, s443[0]);
    wire[0:0] s603, in603_1, in603_2;
    wire c603;
    assign in603_1 = {c443};
    assign in603_2 = {c444};
    Full_Adder FA_603(s603, c603, in603_1, in603_2, c442);
    wire[0:0] s604, in604_1, in604_2;
    wire c604;
    assign in604_1 = {c446};
    assign in604_2 = {s447[0]};
    Full_Adder FA_604(s604, c604, in604_1, in604_2, c445);
    wire[0:0] s605, in605_1, in605_2;
    wire c605;
    assign in605_1 = {s449[0]};
    assign in605_2 = {s450[0]};
    Full_Adder FA_605(s605, c605, in605_1, in605_2, s448[0]);
    wire[0:0] s606, in606_1, in606_2;
    wire c606;
    assign in606_1 = {c448};
    assign in606_2 = {c449};
    Full_Adder FA_606(s606, c606, in606_1, in606_2, c447);
    wire[0:0] s607, in607_1, in607_2;
    wire c607;
    assign in607_1 = {c451};
    assign in607_2 = {s452[0]};
    Full_Adder FA_607(s607, c607, in607_1, in607_2, c450);
    wire[0:0] s608, in608_1, in608_2;
    wire c608;
    assign in608_1 = {s454[0]};
    assign in608_2 = {s455[0]};
    Full_Adder FA_608(s608, c608, in608_1, in608_2, s453[0]);
    wire[0:0] s609, in609_1, in609_2;
    wire c609;
    assign in609_1 = {c453};
    assign in609_2 = {c454};
    Full_Adder FA_609(s609, c609, in609_1, in609_2, c452);
    wire[0:0] s610, in610_1, in610_2;
    wire c610;
    assign in610_1 = {c456};
    assign in610_2 = {s457[0]};
    Full_Adder FA_610(s610, c610, in610_1, in610_2, c455);
    wire[0:0] s611, in611_1, in611_2;
    wire c611;
    assign in611_1 = {s459[0]};
    assign in611_2 = {s460[0]};
    Full_Adder FA_611(s611, c611, in611_1, in611_2, s458[0]);
    wire[0:0] s612, in612_1, in612_2;
    wire c612;
    assign in612_1 = {c458};
    assign in612_2 = {c459};
    Full_Adder FA_612(s612, c612, in612_1, in612_2, c457);
    wire[0:0] s613, in613_1, in613_2;
    wire c613;
    assign in613_1 = {c461};
    assign in613_2 = {s462[0]};
    Full_Adder FA_613(s613, c613, in613_1, in613_2, c460);
    wire[0:0] s614, in614_1, in614_2;
    wire c614;
    assign in614_1 = {s464[0]};
    assign in614_2 = {s465[0]};
    Full_Adder FA_614(s614, c614, in614_1, in614_2, s463[0]);
    wire[0:0] s615, in615_1, in615_2;
    wire c615;
    assign in615_1 = {c463};
    assign in615_2 = {c464};
    Full_Adder FA_615(s615, c615, in615_1, in615_2, c462);
    wire[0:0] s616, in616_1, in616_2;
    wire c616;
    assign in616_1 = {c466};
    assign in616_2 = {s467[0]};
    Full_Adder FA_616(s616, c616, in616_1, in616_2, c465);
    wire[0:0] s617, in617_1, in617_2;
    wire c617;
    assign in617_1 = {s469[0]};
    assign in617_2 = {s470[0]};
    Full_Adder FA_617(s617, c617, in617_1, in617_2, s468[0]);
    wire[0:0] s618, in618_1, in618_2;
    wire c618;
    assign in618_1 = {c468};
    assign in618_2 = {c469};
    Full_Adder FA_618(s618, c618, in618_1, in618_2, c467);
    wire[0:0] s619, in619_1, in619_2;
    wire c619;
    assign in619_1 = {c471};
    assign in619_2 = {s472[0]};
    Full_Adder FA_619(s619, c619, in619_1, in619_2, c470);
    wire[0:0] s620, in620_1, in620_2;
    wire c620;
    assign in620_1 = {s474[0]};
    assign in620_2 = {s475[0]};
    Full_Adder FA_620(s620, c620, in620_1, in620_2, s473[0]);
    wire[0:0] s621, in621_1, in621_2;
    wire c621;
    assign in621_1 = {c473};
    assign in621_2 = {c474};
    Full_Adder FA_621(s621, c621, in621_1, in621_2, c472);
    wire[0:0] s622, in622_1, in622_2;
    wire c622;
    assign in622_1 = {c476};
    assign in622_2 = {s477[0]};
    Full_Adder FA_622(s622, c622, in622_1, in622_2, c475);
    wire[0:0] s623, in623_1, in623_2;
    wire c623;
    assign in623_1 = {s479[0]};
    assign in623_2 = {s480[0]};
    Full_Adder FA_623(s623, c623, in623_1, in623_2, s478[0]);
    wire[0:0] s624, in624_1, in624_2;
    wire c624;
    assign in624_1 = {c478};
    assign in624_2 = {c479};
    Full_Adder FA_624(s624, c624, in624_1, in624_2, c477);
    wire[0:0] s625, in625_1, in625_2;
    wire c625;
    assign in625_1 = {c481};
    assign in625_2 = {s482[0]};
    Full_Adder FA_625(s625, c625, in625_1, in625_2, c480);
    wire[0:0] s626, in626_1, in626_2;
    wire c626;
    assign in626_1 = {s484[0]};
    assign in626_2 = {s485[0]};
    Full_Adder FA_626(s626, c626, in626_1, in626_2, s483[0]);
    wire[0:0] s627, in627_1, in627_2;
    wire c627;
    assign in627_1 = {c483};
    assign in627_2 = {c484};
    Full_Adder FA_627(s627, c627, in627_1, in627_2, c482);
    wire[0:0] s628, in628_1, in628_2;
    wire c628;
    assign in628_1 = {c486};
    assign in628_2 = {s487[0]};
    Full_Adder FA_628(s628, c628, in628_1, in628_2, c485);
    wire[0:0] s629, in629_1, in629_2;
    wire c629;
    assign in629_1 = {s489[0]};
    assign in629_2 = {s490[0]};
    Full_Adder FA_629(s629, c629, in629_1, in629_2, s488[0]);
    wire[0:0] s630, in630_1, in630_2;
    wire c630;
    assign in630_1 = {c488};
    assign in630_2 = {c489};
    Full_Adder FA_630(s630, c630, in630_1, in630_2, c487);
    wire[0:0] s631, in631_1, in631_2;
    wire c631;
    assign in631_1 = {c491};
    assign in631_2 = {s492[0]};
    Full_Adder FA_631(s631, c631, in631_1, in631_2, c490);
    wire[0:0] s632, in632_1, in632_2;
    wire c632;
    assign in632_1 = {s494[0]};
    assign in632_2 = {s495[0]};
    Full_Adder FA_632(s632, c632, in632_1, in632_2, s493[0]);
    wire[0:0] s633, in633_1, in633_2;
    wire c633;
    assign in633_1 = {c492};
    assign in633_2 = {c493};
    Full_Adder FA_633(s633, c633, in633_1, in633_2, pp31[19]);
    wire[0:0] s634, in634_1, in634_2;
    wire c634;
    assign in634_1 = {c495};
    assign in634_2 = {c496};
    Full_Adder FA_634(s634, c634, in634_1, in634_2, c494);
    wire[0:0] s635, in635_1, in635_2;
    wire c635;
    assign in635_1 = {s498[0]};
    assign in635_2 = {s499[0]};
    Full_Adder FA_635(s635, c635, in635_1, in635_2, s497[0]);
    wire[0:0] s636, in636_1, in636_2;
    wire c636;
    assign in636_1 = {pp30[21]};
    assign in636_2 = {pp31[20]};
    Full_Adder FA_636(s636, c636, in636_1, in636_2, pp29[22]);
    wire[0:0] s637, in637_1, in637_2;
    wire c637;
    assign in637_1 = {c498};
    assign in637_2 = {c499};
    Full_Adder FA_637(s637, c637, in637_1, in637_2, c497);
    wire[0:0] s638, in638_1, in638_2;
    wire c638;
    assign in638_1 = {s501[0]};
    assign in638_2 = {s502[0]};
    Full_Adder FA_638(s638, c638, in638_1, in638_2, c500);
    wire[0:0] s639, in639_1, in639_2;
    wire c639;
    assign in639_1 = {pp28[24]};
    assign in639_2 = {pp29[23]};
    Full_Adder FA_639(s639, c639, in639_1, in639_2, pp27[25]);
    wire[0:0] s640, in640_1, in640_2;
    wire c640;
    assign in640_1 = {pp31[21]};
    assign in640_2 = {c501};
    Full_Adder FA_640(s640, c640, in640_1, in640_2, pp30[22]);
    wire[0:0] s641, in641_1, in641_2;
    wire c641;
    assign in641_1 = {c503};
    assign in641_2 = {s504[0]};
    Full_Adder FA_641(s641, c641, in641_1, in641_2, c502);
    wire[0:0] s642, in642_1, in642_2;
    wire c642;
    assign in642_1 = {pp26[27]};
    assign in642_2 = {pp27[26]};
    Full_Adder FA_642(s642, c642, in642_1, in642_2, pp25[28]);
    wire[0:0] s643, in643_1, in643_2;
    wire c643;
    assign in643_1 = {pp29[24]};
    assign in643_2 = {pp30[23]};
    Full_Adder FA_643(s643, c643, in643_1, in643_2, pp28[25]);
    wire[0:0] s644, in644_1, in644_2;
    wire c644;
    assign in644_1 = {c504};
    assign in644_2 = {c505};
    Full_Adder FA_644(s644, c644, in644_1, in644_2, pp31[22]);
    wire[0:0] s645, in645_1, in645_2;
    wire c645;
    assign in645_1 = {pp24[30]};
    assign in645_2 = {pp25[29]};
    Full_Adder FA_645(s645, c645, in645_1, in645_2, pp23[31]);
    wire[0:0] s646, in646_1, in646_2;
    wire c646;
    assign in646_1 = {pp27[27]};
    assign in646_2 = {pp28[26]};
    Full_Adder FA_646(s646, c646, in646_1, in646_2, pp26[28]);
    wire[0:0] s647, in647_1, in647_2;
    wire c647;
    assign in647_1 = {pp30[24]};
    assign in647_2 = {pp31[23]};
    Full_Adder FA_647(s647, c647, in647_1, in647_2, pp29[25]);
    wire[0:0] s648, in648_1, in648_2;
    wire c648;
    assign in648_1 = {pp25[30]};
    assign in648_2 = {pp26[29]};
    Full_Adder FA_648(s648, c648, in648_1, in648_2, pp24[31]);
    wire[0:0] s649, in649_1, in649_2;
    wire c649;
    assign in649_1 = {pp28[27]};
    assign in649_2 = {pp29[26]};
    Full_Adder FA_649(s649, c649, in649_1, in649_2, pp27[28]);
    wire[0:0] s650, in650_1, in650_2;
    wire c650;
    assign in650_1 = {pp26[30]};
    assign in650_2 = {pp27[29]};
    Full_Adder FA_650(s650, c650, in650_1, in650_2, pp25[31]);

    /*Stage 5*/
    wire[0:0] s651, in651_1, in651_2;
    wire c651;
    assign in651_1 = {pp0[5]};
    assign in651_2 = {pp1[4]};
    Half_Adder HA_651(s651, c651, in651_1, in651_2);
    wire[0:0] s652, in652_1, in652_2;
    wire c652;
    assign in652_1 = {pp1[5]};
    assign in652_2 = {pp2[4]};
    Full_Adder FA_652(s652, c652, in652_1, in652_2, pp0[6]);
    wire[0:0] s653, in653_1, in653_2;
    wire c653;
    assign in653_1 = {pp3[3]};
    assign in653_2 = {pp4[2]};
    Half_Adder HA_653(s653, c653, in653_1, in653_2);
    wire[0:0] s654, in654_1, in654_2;
    wire c654;
    assign in654_1 = {pp3[4]};
    assign in654_2 = {pp4[3]};
    Full_Adder FA_654(s654, c654, in654_1, in654_2, pp2[5]);
    wire[0:0] s655, in655_1, in655_2;
    wire c655;
    assign in655_1 = {pp6[1]};
    assign in655_2 = {pp7[0]};
    Full_Adder FA_655(s655, c655, in655_1, in655_2, pp5[2]);
    wire[0:0] s656, in656_1, in656_2;
    wire c656;
    assign in656_1 = {pp6[2]};
    assign in656_2 = {pp7[1]};
    Full_Adder FA_656(s656, c656, in656_1, in656_2, pp5[3]);
    wire[0:0] s657, in657_1, in657_2;
    wire c657;
    assign in657_1 = {c507};
    assign in657_2 = {s508[0]};
    Full_Adder FA_657(s657, c657, in657_1, in657_2, pp8[0]);
    wire[0:0] s658, in658_1, in658_2;
    wire c658;
    assign in658_1 = {pp9[0]};
    assign in658_2 = {c508};
    Full_Adder FA_658(s658, c658, in658_1, in658_2, pp8[1]);
    wire[0:0] s659, in659_1, in659_2;
    wire c659;
    assign in659_1 = {s510[0]};
    assign in659_2 = {s511[0]};
    Full_Adder FA_659(s659, c659, in659_1, in659_2, c509);
    wire[0:0] s660, in660_1, in660_2;
    wire c660;
    assign in660_1 = {c510};
    assign in660_2 = {c511};
    Full_Adder FA_660(s660, c660, in660_1, in660_2, s307[0]);
    wire[0:0] s661, in661_1, in661_2;
    wire c661;
    assign in661_1 = {s513[0]};
    assign in661_2 = {s514[0]};
    Full_Adder FA_661(s661, c661, in661_1, in661_2, c512);
    wire[0:0] s662, in662_1, in662_2;
    wire c662;
    assign in662_1 = {c513};
    assign in662_2 = {c514};
    Full_Adder FA_662(s662, c662, in662_1, in662_2, s309[0]);
    wire[0:0] s663, in663_1, in663_2;
    wire c663;
    assign in663_1 = {s516[0]};
    assign in663_2 = {s517[0]};
    Full_Adder FA_663(s663, c663, in663_1, in663_2, c515);
    wire[0:0] s664, in664_1, in664_2;
    wire c664;
    assign in664_1 = {c516};
    assign in664_2 = {c517};
    Full_Adder FA_664(s664, c664, in664_1, in664_2, s312[0]);
    wire[0:0] s665, in665_1, in665_2;
    wire c665;
    assign in665_1 = {s519[0]};
    assign in665_2 = {s520[0]};
    Full_Adder FA_665(s665, c665, in665_1, in665_2, c518);
    wire[0:0] s666, in666_1, in666_2;
    wire c666;
    assign in666_1 = {c519};
    assign in666_2 = {c520};
    Full_Adder FA_666(s666, c666, in666_1, in666_2, s316[0]);
    wire[0:0] s667, in667_1, in667_2;
    wire c667;
    assign in667_1 = {s522[0]};
    assign in667_2 = {s523[0]};
    Full_Adder FA_667(s667, c667, in667_1, in667_2, c521);
    wire[0:0] s668, in668_1, in668_2;
    wire c668;
    assign in668_1 = {c522};
    assign in668_2 = {c523};
    Full_Adder FA_668(s668, c668, in668_1, in668_2, s321[0]);
    wire[0:0] s669, in669_1, in669_2;
    wire c669;
    assign in669_1 = {s525[0]};
    assign in669_2 = {s526[0]};
    Full_Adder FA_669(s669, c669, in669_1, in669_2, c524);
    wire[0:0] s670, in670_1, in670_2;
    wire c670;
    assign in670_1 = {c525};
    assign in670_2 = {c526};
    Full_Adder FA_670(s670, c670, in670_1, in670_2, s326[0]);
    wire[0:0] s671, in671_1, in671_2;
    wire c671;
    assign in671_1 = {s528[0]};
    assign in671_2 = {s529[0]};
    Full_Adder FA_671(s671, c671, in671_1, in671_2, c527);
    wire[0:0] s672, in672_1, in672_2;
    wire c672;
    assign in672_1 = {c528};
    assign in672_2 = {c529};
    Full_Adder FA_672(s672, c672, in672_1, in672_2, s331[0]);
    wire[0:0] s673, in673_1, in673_2;
    wire c673;
    assign in673_1 = {s531[0]};
    assign in673_2 = {s532[0]};
    Full_Adder FA_673(s673, c673, in673_1, in673_2, c530);
    wire[0:0] s674, in674_1, in674_2;
    wire c674;
    assign in674_1 = {c531};
    assign in674_2 = {c532};
    Full_Adder FA_674(s674, c674, in674_1, in674_2, s336[0]);
    wire[0:0] s675, in675_1, in675_2;
    wire c675;
    assign in675_1 = {s534[0]};
    assign in675_2 = {s535[0]};
    Full_Adder FA_675(s675, c675, in675_1, in675_2, c533);
    wire[0:0] s676, in676_1, in676_2;
    wire c676;
    assign in676_1 = {c534};
    assign in676_2 = {c535};
    Full_Adder FA_676(s676, c676, in676_1, in676_2, s341[0]);
    wire[0:0] s677, in677_1, in677_2;
    wire c677;
    assign in677_1 = {s537[0]};
    assign in677_2 = {s538[0]};
    Full_Adder FA_677(s677, c677, in677_1, in677_2, c536);
    wire[0:0] s678, in678_1, in678_2;
    wire c678;
    assign in678_1 = {c537};
    assign in678_2 = {c538};
    Full_Adder FA_678(s678, c678, in678_1, in678_2, s346[0]);
    wire[0:0] s679, in679_1, in679_2;
    wire c679;
    assign in679_1 = {s540[0]};
    assign in679_2 = {s541[0]};
    Full_Adder FA_679(s679, c679, in679_1, in679_2, c539);
    wire[0:0] s680, in680_1, in680_2;
    wire c680;
    assign in680_1 = {c540};
    assign in680_2 = {c541};
    Full_Adder FA_680(s680, c680, in680_1, in680_2, s351[0]);
    wire[0:0] s681, in681_1, in681_2;
    wire c681;
    assign in681_1 = {s543[0]};
    assign in681_2 = {s544[0]};
    Full_Adder FA_681(s681, c681, in681_1, in681_2, c542);
    wire[0:0] s682, in682_1, in682_2;
    wire c682;
    assign in682_1 = {c543};
    assign in682_2 = {c544};
    Full_Adder FA_682(s682, c682, in682_1, in682_2, s356[0]);
    wire[0:0] s683, in683_1, in683_2;
    wire c683;
    assign in683_1 = {s546[0]};
    assign in683_2 = {s547[0]};
    Full_Adder FA_683(s683, c683, in683_1, in683_2, c545);
    wire[0:0] s684, in684_1, in684_2;
    wire c684;
    assign in684_1 = {c546};
    assign in684_2 = {c547};
    Full_Adder FA_684(s684, c684, in684_1, in684_2, s361[0]);
    wire[0:0] s685, in685_1, in685_2;
    wire c685;
    assign in685_1 = {s549[0]};
    assign in685_2 = {s550[0]};
    Full_Adder FA_685(s685, c685, in685_1, in685_2, c548);
    wire[0:0] s686, in686_1, in686_2;
    wire c686;
    assign in686_1 = {c549};
    assign in686_2 = {c550};
    Full_Adder FA_686(s686, c686, in686_1, in686_2, s366[0]);
    wire[0:0] s687, in687_1, in687_2;
    wire c687;
    assign in687_1 = {s552[0]};
    assign in687_2 = {s553[0]};
    Full_Adder FA_687(s687, c687, in687_1, in687_2, c551);
    wire[0:0] s688, in688_1, in688_2;
    wire c688;
    assign in688_1 = {c552};
    assign in688_2 = {c553};
    Full_Adder FA_688(s688, c688, in688_1, in688_2, s371[0]);
    wire[0:0] s689, in689_1, in689_2;
    wire c689;
    assign in689_1 = {s555[0]};
    assign in689_2 = {s556[0]};
    Full_Adder FA_689(s689, c689, in689_1, in689_2, c554);
    wire[0:0] s690, in690_1, in690_2;
    wire c690;
    assign in690_1 = {c555};
    assign in690_2 = {c556};
    Full_Adder FA_690(s690, c690, in690_1, in690_2, s376[0]);
    wire[0:0] s691, in691_1, in691_2;
    wire c691;
    assign in691_1 = {s558[0]};
    assign in691_2 = {s559[0]};
    Full_Adder FA_691(s691, c691, in691_1, in691_2, c557);
    wire[0:0] s692, in692_1, in692_2;
    wire c692;
    assign in692_1 = {c558};
    assign in692_2 = {c559};
    Full_Adder FA_692(s692, c692, in692_1, in692_2, s381[0]);
    wire[0:0] s693, in693_1, in693_2;
    wire c693;
    assign in693_1 = {s561[0]};
    assign in693_2 = {s562[0]};
    Full_Adder FA_693(s693, c693, in693_1, in693_2, c560);
    wire[0:0] s694, in694_1, in694_2;
    wire c694;
    assign in694_1 = {c561};
    assign in694_2 = {c562};
    Full_Adder FA_694(s694, c694, in694_1, in694_2, s386[0]);
    wire[0:0] s695, in695_1, in695_2;
    wire c695;
    assign in695_1 = {s564[0]};
    assign in695_2 = {s565[0]};
    Full_Adder FA_695(s695, c695, in695_1, in695_2, c563);
    wire[0:0] s696, in696_1, in696_2;
    wire c696;
    assign in696_1 = {c564};
    assign in696_2 = {c565};
    Full_Adder FA_696(s696, c696, in696_1, in696_2, s391[0]);
    wire[0:0] s697, in697_1, in697_2;
    wire c697;
    assign in697_1 = {s567[0]};
    assign in697_2 = {s568[0]};
    Full_Adder FA_697(s697, c697, in697_1, in697_2, c566);
    wire[0:0] s698, in698_1, in698_2;
    wire c698;
    assign in698_1 = {c567};
    assign in698_2 = {c568};
    Full_Adder FA_698(s698, c698, in698_1, in698_2, s396[0]);
    wire[0:0] s699, in699_1, in699_2;
    wire c699;
    assign in699_1 = {s570[0]};
    assign in699_2 = {s571[0]};
    Full_Adder FA_699(s699, c699, in699_1, in699_2, c569);
    wire[0:0] s700, in700_1, in700_2;
    wire c700;
    assign in700_1 = {c570};
    assign in700_2 = {c571};
    Full_Adder FA_700(s700, c700, in700_1, in700_2, s401[0]);
    wire[0:0] s701, in701_1, in701_2;
    wire c701;
    assign in701_1 = {s573[0]};
    assign in701_2 = {s574[0]};
    Full_Adder FA_701(s701, c701, in701_1, in701_2, c572);
    wire[0:0] s702, in702_1, in702_2;
    wire c702;
    assign in702_1 = {c573};
    assign in702_2 = {c574};
    Full_Adder FA_702(s702, c702, in702_1, in702_2, s406[0]);
    wire[0:0] s703, in703_1, in703_2;
    wire c703;
    assign in703_1 = {s576[0]};
    assign in703_2 = {s577[0]};
    Full_Adder FA_703(s703, c703, in703_1, in703_2, c575);
    wire[0:0] s704, in704_1, in704_2;
    wire c704;
    assign in704_1 = {c576};
    assign in704_2 = {c577};
    Full_Adder FA_704(s704, c704, in704_1, in704_2, s411[0]);
    wire[0:0] s705, in705_1, in705_2;
    wire c705;
    assign in705_1 = {s579[0]};
    assign in705_2 = {s580[0]};
    Full_Adder FA_705(s705, c705, in705_1, in705_2, c578);
    wire[0:0] s706, in706_1, in706_2;
    wire c706;
    assign in706_1 = {c579};
    assign in706_2 = {c580};
    Full_Adder FA_706(s706, c706, in706_1, in706_2, s416[0]);
    wire[0:0] s707, in707_1, in707_2;
    wire c707;
    assign in707_1 = {s582[0]};
    assign in707_2 = {s583[0]};
    Full_Adder FA_707(s707, c707, in707_1, in707_2, c581);
    wire[0:0] s708, in708_1, in708_2;
    wire c708;
    assign in708_1 = {c582};
    assign in708_2 = {c583};
    Full_Adder FA_708(s708, c708, in708_1, in708_2, s421[0]);
    wire[0:0] s709, in709_1, in709_2;
    wire c709;
    assign in709_1 = {s585[0]};
    assign in709_2 = {s586[0]};
    Full_Adder FA_709(s709, c709, in709_1, in709_2, c584);
    wire[0:0] s710, in710_1, in710_2;
    wire c710;
    assign in710_1 = {c585};
    assign in710_2 = {c586};
    Full_Adder FA_710(s710, c710, in710_1, in710_2, s426[0]);
    wire[0:0] s711, in711_1, in711_2;
    wire c711;
    assign in711_1 = {s588[0]};
    assign in711_2 = {s589[0]};
    Full_Adder FA_711(s711, c711, in711_1, in711_2, c587);
    wire[0:0] s712, in712_1, in712_2;
    wire c712;
    assign in712_1 = {c588};
    assign in712_2 = {c589};
    Full_Adder FA_712(s712, c712, in712_1, in712_2, s431[0]);
    wire[0:0] s713, in713_1, in713_2;
    wire c713;
    assign in713_1 = {s591[0]};
    assign in713_2 = {s592[0]};
    Full_Adder FA_713(s713, c713, in713_1, in713_2, c590);
    wire[0:0] s714, in714_1, in714_2;
    wire c714;
    assign in714_1 = {c591};
    assign in714_2 = {c592};
    Full_Adder FA_714(s714, c714, in714_1, in714_2, s436[0]);
    wire[0:0] s715, in715_1, in715_2;
    wire c715;
    assign in715_1 = {s594[0]};
    assign in715_2 = {s595[0]};
    Full_Adder FA_715(s715, c715, in715_1, in715_2, c593);
    wire[0:0] s716, in716_1, in716_2;
    wire c716;
    assign in716_1 = {c594};
    assign in716_2 = {c595};
    Full_Adder FA_716(s716, c716, in716_1, in716_2, s441[0]);
    wire[0:0] s717, in717_1, in717_2;
    wire c717;
    assign in717_1 = {s597[0]};
    assign in717_2 = {s598[0]};
    Full_Adder FA_717(s717, c717, in717_1, in717_2, c596);
    wire[0:0] s718, in718_1, in718_2;
    wire c718;
    assign in718_1 = {c597};
    assign in718_2 = {c598};
    Full_Adder FA_718(s718, c718, in718_1, in718_2, s446[0]);
    wire[0:0] s719, in719_1, in719_2;
    wire c719;
    assign in719_1 = {s600[0]};
    assign in719_2 = {s601[0]};
    Full_Adder FA_719(s719, c719, in719_1, in719_2, c599);
    wire[0:0] s720, in720_1, in720_2;
    wire c720;
    assign in720_1 = {c600};
    assign in720_2 = {c601};
    Full_Adder FA_720(s720, c720, in720_1, in720_2, s451[0]);
    wire[0:0] s721, in721_1, in721_2;
    wire c721;
    assign in721_1 = {s603[0]};
    assign in721_2 = {s604[0]};
    Full_Adder FA_721(s721, c721, in721_1, in721_2, c602);
    wire[0:0] s722, in722_1, in722_2;
    wire c722;
    assign in722_1 = {c603};
    assign in722_2 = {c604};
    Full_Adder FA_722(s722, c722, in722_1, in722_2, s456[0]);
    wire[0:0] s723, in723_1, in723_2;
    wire c723;
    assign in723_1 = {s606[0]};
    assign in723_2 = {s607[0]};
    Full_Adder FA_723(s723, c723, in723_1, in723_2, c605);
    wire[0:0] s724, in724_1, in724_2;
    wire c724;
    assign in724_1 = {c606};
    assign in724_2 = {c607};
    Full_Adder FA_724(s724, c724, in724_1, in724_2, s461[0]);
    wire[0:0] s725, in725_1, in725_2;
    wire c725;
    assign in725_1 = {s609[0]};
    assign in725_2 = {s610[0]};
    Full_Adder FA_725(s725, c725, in725_1, in725_2, c608);
    wire[0:0] s726, in726_1, in726_2;
    wire c726;
    assign in726_1 = {c609};
    assign in726_2 = {c610};
    Full_Adder FA_726(s726, c726, in726_1, in726_2, s466[0]);
    wire[0:0] s727, in727_1, in727_2;
    wire c727;
    assign in727_1 = {s612[0]};
    assign in727_2 = {s613[0]};
    Full_Adder FA_727(s727, c727, in727_1, in727_2, c611);
    wire[0:0] s728, in728_1, in728_2;
    wire c728;
    assign in728_1 = {c612};
    assign in728_2 = {c613};
    Full_Adder FA_728(s728, c728, in728_1, in728_2, s471[0]);
    wire[0:0] s729, in729_1, in729_2;
    wire c729;
    assign in729_1 = {s615[0]};
    assign in729_2 = {s616[0]};
    Full_Adder FA_729(s729, c729, in729_1, in729_2, c614);
    wire[0:0] s730, in730_1, in730_2;
    wire c730;
    assign in730_1 = {c615};
    assign in730_2 = {c616};
    Full_Adder FA_730(s730, c730, in730_1, in730_2, s476[0]);
    wire[0:0] s731, in731_1, in731_2;
    wire c731;
    assign in731_1 = {s618[0]};
    assign in731_2 = {s619[0]};
    Full_Adder FA_731(s731, c731, in731_1, in731_2, c617);
    wire[0:0] s732, in732_1, in732_2;
    wire c732;
    assign in732_1 = {c618};
    assign in732_2 = {c619};
    Full_Adder FA_732(s732, c732, in732_1, in732_2, s481[0]);
    wire[0:0] s733, in733_1, in733_2;
    wire c733;
    assign in733_1 = {s621[0]};
    assign in733_2 = {s622[0]};
    Full_Adder FA_733(s733, c733, in733_1, in733_2, c620);
    wire[0:0] s734, in734_1, in734_2;
    wire c734;
    assign in734_1 = {c621};
    assign in734_2 = {c622};
    Full_Adder FA_734(s734, c734, in734_1, in734_2, s486[0]);
    wire[0:0] s735, in735_1, in735_2;
    wire c735;
    assign in735_1 = {s624[0]};
    assign in735_2 = {s625[0]};
    Full_Adder FA_735(s735, c735, in735_1, in735_2, c623);
    wire[0:0] s736, in736_1, in736_2;
    wire c736;
    assign in736_1 = {c624};
    assign in736_2 = {c625};
    Full_Adder FA_736(s736, c736, in736_1, in736_2, s491[0]);
    wire[0:0] s737, in737_1, in737_2;
    wire c737;
    assign in737_1 = {s627[0]};
    assign in737_2 = {s628[0]};
    Full_Adder FA_737(s737, c737, in737_1, in737_2, c626);
    wire[0:0] s738, in738_1, in738_2;
    wire c738;
    assign in738_1 = {c627};
    assign in738_2 = {c628};
    Full_Adder FA_738(s738, c738, in738_1, in738_2, s496[0]);
    wire[0:0] s739, in739_1, in739_2;
    wire c739;
    assign in739_1 = {s630[0]};
    assign in739_2 = {s631[0]};
    Full_Adder FA_739(s739, c739, in739_1, in739_2, c629);
    wire[0:0] s740, in740_1, in740_2;
    wire c740;
    assign in740_1 = {c630};
    assign in740_2 = {c631};
    Full_Adder FA_740(s740, c740, in740_1, in740_2, s500[0]);
    wire[0:0] s741, in741_1, in741_2;
    wire c741;
    assign in741_1 = {s633[0]};
    assign in741_2 = {s634[0]};
    Full_Adder FA_741(s741, c741, in741_1, in741_2, c632);
    wire[0:0] s742, in742_1, in742_2;
    wire c742;
    assign in742_1 = {c633};
    assign in742_2 = {c634};
    Full_Adder FA_742(s742, c742, in742_1, in742_2, s503[0]);
    wire[0:0] s743, in743_1, in743_2;
    wire c743;
    assign in743_1 = {s636[0]};
    assign in743_2 = {s637[0]};
    Full_Adder FA_743(s743, c743, in743_1, in743_2, c635);
    wire[0:0] s744, in744_1, in744_2;
    wire c744;
    assign in744_1 = {c636};
    assign in744_2 = {c637};
    Full_Adder FA_744(s744, c744, in744_1, in744_2, s505[0]);
    wire[0:0] s745, in745_1, in745_2;
    wire c745;
    assign in745_1 = {s639[0]};
    assign in745_2 = {s640[0]};
    Full_Adder FA_745(s745, c745, in745_1, in745_2, c638);
    wire[0:0] s746, in746_1, in746_2;
    wire c746;
    assign in746_1 = {c639};
    assign in746_2 = {c640};
    Full_Adder FA_746(s746, c746, in746_1, in746_2, s506[0]);
    wire[0:0] s747, in747_1, in747_2;
    wire c747;
    assign in747_1 = {s642[0]};
    assign in747_2 = {s643[0]};
    Full_Adder FA_747(s747, c747, in747_1, in747_2, c641);
    wire[0:0] s748, in748_1, in748_2;
    wire c748;
    assign in748_1 = {c642};
    assign in748_2 = {c643};
    Full_Adder FA_748(s748, c748, in748_1, in748_2, c506);
    wire[0:0] s749, in749_1, in749_2;
    wire c749;
    assign in749_1 = {s645[0]};
    assign in749_2 = {s646[0]};
    Full_Adder FA_749(s749, c749, in749_1, in749_2, c644);
    wire[0:0] s750, in750_1, in750_2;
    wire c750;
    assign in750_1 = {pp31[24]};
    assign in750_2 = {c645};
    Full_Adder FA_750(s750, c750, in750_1, in750_2, pp30[25]);
    wire[0:0] s751, in751_1, in751_2;
    wire c751;
    assign in751_1 = {c647};
    assign in751_2 = {s648[0]};
    Full_Adder FA_751(s751, c751, in751_1, in751_2, c646);
    wire[0:0] s752, in752_1, in752_2;
    wire c752;
    assign in752_1 = {pp29[27]};
    assign in752_2 = {pp30[26]};
    Full_Adder FA_752(s752, c752, in752_1, in752_2, pp28[28]);
    wire[0:0] s753, in753_1, in753_2;
    wire c753;
    assign in753_1 = {c648};
    assign in753_2 = {c649};
    Full_Adder FA_753(s753, c753, in753_1, in753_2, pp31[25]);
    wire[0:0] s754, in754_1, in754_2;
    wire c754;
    assign in754_1 = {pp27[30]};
    assign in754_2 = {pp28[29]};
    Full_Adder FA_754(s754, c754, in754_1, in754_2, pp26[31]);
    wire[0:0] s755, in755_1, in755_2;
    wire c755;
    assign in755_1 = {pp30[27]};
    assign in755_2 = {pp31[26]};
    Full_Adder FA_755(s755, c755, in755_1, in755_2, pp29[28]);
    wire[0:0] s756, in756_1, in756_2;
    wire c756;
    assign in756_1 = {pp28[30]};
    assign in756_2 = {pp29[29]};
    Full_Adder FA_756(s756, c756, in756_1, in756_2, pp27[31]);

    /*Stage 6*/
    wire[0:0] s757, in757_1, in757_2;
    wire c757;
    assign in757_1 = {pp0[4]};
    assign in757_2 = {pp1[3]};
    Half_Adder HA_757(s757, c757, in757_1, in757_2);
    wire[0:0] s758, in758_1, in758_2;
    wire c758;
    assign in758_1 = {pp3[2]};
    assign in758_2 = {pp4[1]};
    Full_Adder FA_758(s758, c758, in758_1, in758_2, pp2[3]);
    wire[0:0] s759, in759_1, in759_2;
    wire c759;
    assign in759_1 = {pp6[0]};
    assign in759_2 = {c651};
    Full_Adder FA_759(s759, c759, in759_1, in759_2, pp5[1]);
    wire[0:0] s760, in760_1, in760_2;
    wire c760;
    assign in760_1 = {c652};
    assign in760_2 = {c653};
    Full_Adder FA_760(s760, c760, in760_1, in760_2, s507[0]);
    wire[0:0] s761, in761_1, in761_2;
    wire c761;
    assign in761_1 = {c654};
    assign in761_2 = {c655};
    Full_Adder FA_761(s761, c761, in761_1, in761_2, s509[0]);
    wire[0:0] s762, in762_1, in762_2;
    wire c762;
    assign in762_1 = {c656};
    assign in762_2 = {c657};
    Full_Adder FA_762(s762, c762, in762_1, in762_2, s512[0]);
    wire[0:0] s763, in763_1, in763_2;
    wire c763;
    assign in763_1 = {c658};
    assign in763_2 = {c659};
    Full_Adder FA_763(s763, c763, in763_1, in763_2, s515[0]);
    wire[0:0] s764, in764_1, in764_2;
    wire c764;
    assign in764_1 = {c660};
    assign in764_2 = {c661};
    Full_Adder FA_764(s764, c764, in764_1, in764_2, s518[0]);
    wire[0:0] s765, in765_1, in765_2;
    wire c765;
    assign in765_1 = {c662};
    assign in765_2 = {c663};
    Full_Adder FA_765(s765, c765, in765_1, in765_2, s521[0]);
    wire[0:0] s766, in766_1, in766_2;
    wire c766;
    assign in766_1 = {c664};
    assign in766_2 = {c665};
    Full_Adder FA_766(s766, c766, in766_1, in766_2, s524[0]);
    wire[0:0] s767, in767_1, in767_2;
    wire c767;
    assign in767_1 = {c666};
    assign in767_2 = {c667};
    Full_Adder FA_767(s767, c767, in767_1, in767_2, s527[0]);
    wire[0:0] s768, in768_1, in768_2;
    wire c768;
    assign in768_1 = {c668};
    assign in768_2 = {c669};
    Full_Adder FA_768(s768, c768, in768_1, in768_2, s530[0]);
    wire[0:0] s769, in769_1, in769_2;
    wire c769;
    assign in769_1 = {c670};
    assign in769_2 = {c671};
    Full_Adder FA_769(s769, c769, in769_1, in769_2, s533[0]);
    wire[0:0] s770, in770_1, in770_2;
    wire c770;
    assign in770_1 = {c672};
    assign in770_2 = {c673};
    Full_Adder FA_770(s770, c770, in770_1, in770_2, s536[0]);
    wire[0:0] s771, in771_1, in771_2;
    wire c771;
    assign in771_1 = {c674};
    assign in771_2 = {c675};
    Full_Adder FA_771(s771, c771, in771_1, in771_2, s539[0]);
    wire[0:0] s772, in772_1, in772_2;
    wire c772;
    assign in772_1 = {c676};
    assign in772_2 = {c677};
    Full_Adder FA_772(s772, c772, in772_1, in772_2, s542[0]);
    wire[0:0] s773, in773_1, in773_2;
    wire c773;
    assign in773_1 = {c678};
    assign in773_2 = {c679};
    Full_Adder FA_773(s773, c773, in773_1, in773_2, s545[0]);
    wire[0:0] s774, in774_1, in774_2;
    wire c774;
    assign in774_1 = {c680};
    assign in774_2 = {c681};
    Full_Adder FA_774(s774, c774, in774_1, in774_2, s548[0]);
    wire[0:0] s775, in775_1, in775_2;
    wire c775;
    assign in775_1 = {c682};
    assign in775_2 = {c683};
    Full_Adder FA_775(s775, c775, in775_1, in775_2, s551[0]);
    wire[0:0] s776, in776_1, in776_2;
    wire c776;
    assign in776_1 = {c684};
    assign in776_2 = {c685};
    Full_Adder FA_776(s776, c776, in776_1, in776_2, s554[0]);
    wire[0:0] s777, in777_1, in777_2;
    wire c777;
    assign in777_1 = {c686};
    assign in777_2 = {c687};
    Full_Adder FA_777(s777, c777, in777_1, in777_2, s557[0]);
    wire[0:0] s778, in778_1, in778_2;
    wire c778;
    assign in778_1 = {c688};
    assign in778_2 = {c689};
    Full_Adder FA_778(s778, c778, in778_1, in778_2, s560[0]);
    wire[0:0] s779, in779_1, in779_2;
    wire c779;
    assign in779_1 = {c690};
    assign in779_2 = {c691};
    Full_Adder FA_779(s779, c779, in779_1, in779_2, s563[0]);
    wire[0:0] s780, in780_1, in780_2;
    wire c780;
    assign in780_1 = {c692};
    assign in780_2 = {c693};
    Full_Adder FA_780(s780, c780, in780_1, in780_2, s566[0]);
    wire[0:0] s781, in781_1, in781_2;
    wire c781;
    assign in781_1 = {c694};
    assign in781_2 = {c695};
    Full_Adder FA_781(s781, c781, in781_1, in781_2, s569[0]);
    wire[0:0] s782, in782_1, in782_2;
    wire c782;
    assign in782_1 = {c696};
    assign in782_2 = {c697};
    Full_Adder FA_782(s782, c782, in782_1, in782_2, s572[0]);
    wire[0:0] s783, in783_1, in783_2;
    wire c783;
    assign in783_1 = {c698};
    assign in783_2 = {c699};
    Full_Adder FA_783(s783, c783, in783_1, in783_2, s575[0]);
    wire[0:0] s784, in784_1, in784_2;
    wire c784;
    assign in784_1 = {c700};
    assign in784_2 = {c701};
    Full_Adder FA_784(s784, c784, in784_1, in784_2, s578[0]);
    wire[0:0] s785, in785_1, in785_2;
    wire c785;
    assign in785_1 = {c702};
    assign in785_2 = {c703};
    Full_Adder FA_785(s785, c785, in785_1, in785_2, s581[0]);
    wire[0:0] s786, in786_1, in786_2;
    wire c786;
    assign in786_1 = {c704};
    assign in786_2 = {c705};
    Full_Adder FA_786(s786, c786, in786_1, in786_2, s584[0]);
    wire[0:0] s787, in787_1, in787_2;
    wire c787;
    assign in787_1 = {c706};
    assign in787_2 = {c707};
    Full_Adder FA_787(s787, c787, in787_1, in787_2, s587[0]);
    wire[0:0] s788, in788_1, in788_2;
    wire c788;
    assign in788_1 = {c708};
    assign in788_2 = {c709};
    Full_Adder FA_788(s788, c788, in788_1, in788_2, s590[0]);
    wire[0:0] s789, in789_1, in789_2;
    wire c789;
    assign in789_1 = {c710};
    assign in789_2 = {c711};
    Full_Adder FA_789(s789, c789, in789_1, in789_2, s593[0]);
    wire[0:0] s790, in790_1, in790_2;
    wire c790;
    assign in790_1 = {c712};
    assign in790_2 = {c713};
    Full_Adder FA_790(s790, c790, in790_1, in790_2, s596[0]);
    wire[0:0] s791, in791_1, in791_2;
    wire c791;
    assign in791_1 = {c714};
    assign in791_2 = {c715};
    Full_Adder FA_791(s791, c791, in791_1, in791_2, s599[0]);
    wire[0:0] s792, in792_1, in792_2;
    wire c792;
    assign in792_1 = {c716};
    assign in792_2 = {c717};
    Full_Adder FA_792(s792, c792, in792_1, in792_2, s602[0]);
    wire[0:0] s793, in793_1, in793_2;
    wire c793;
    assign in793_1 = {c718};
    assign in793_2 = {c719};
    Full_Adder FA_793(s793, c793, in793_1, in793_2, s605[0]);
    wire[0:0] s794, in794_1, in794_2;
    wire c794;
    assign in794_1 = {c720};
    assign in794_2 = {c721};
    Full_Adder FA_794(s794, c794, in794_1, in794_2, s608[0]);
    wire[0:0] s795, in795_1, in795_2;
    wire c795;
    assign in795_1 = {c722};
    assign in795_2 = {c723};
    Full_Adder FA_795(s795, c795, in795_1, in795_2, s611[0]);
    wire[0:0] s796, in796_1, in796_2;
    wire c796;
    assign in796_1 = {c724};
    assign in796_2 = {c725};
    Full_Adder FA_796(s796, c796, in796_1, in796_2, s614[0]);
    wire[0:0] s797, in797_1, in797_2;
    wire c797;
    assign in797_1 = {c726};
    assign in797_2 = {c727};
    Full_Adder FA_797(s797, c797, in797_1, in797_2, s617[0]);
    wire[0:0] s798, in798_1, in798_2;
    wire c798;
    assign in798_1 = {c728};
    assign in798_2 = {c729};
    Full_Adder FA_798(s798, c798, in798_1, in798_2, s620[0]);
    wire[0:0] s799, in799_1, in799_2;
    wire c799;
    assign in799_1 = {c730};
    assign in799_2 = {c731};
    Full_Adder FA_799(s799, c799, in799_1, in799_2, s623[0]);
    wire[0:0] s800, in800_1, in800_2;
    wire c800;
    assign in800_1 = {c732};
    assign in800_2 = {c733};
    Full_Adder FA_800(s800, c800, in800_1, in800_2, s626[0]);
    wire[0:0] s801, in801_1, in801_2;
    wire c801;
    assign in801_1 = {c734};
    assign in801_2 = {c735};
    Full_Adder FA_801(s801, c801, in801_1, in801_2, s629[0]);
    wire[0:0] s802, in802_1, in802_2;
    wire c802;
    assign in802_1 = {c736};
    assign in802_2 = {c737};
    Full_Adder FA_802(s802, c802, in802_1, in802_2, s632[0]);
    wire[0:0] s803, in803_1, in803_2;
    wire c803;
    assign in803_1 = {c738};
    assign in803_2 = {c739};
    Full_Adder FA_803(s803, c803, in803_1, in803_2, s635[0]);
    wire[0:0] s804, in804_1, in804_2;
    wire c804;
    assign in804_1 = {c740};
    assign in804_2 = {c741};
    Full_Adder FA_804(s804, c804, in804_1, in804_2, s638[0]);
    wire[0:0] s805, in805_1, in805_2;
    wire c805;
    assign in805_1 = {c742};
    assign in805_2 = {c743};
    Full_Adder FA_805(s805, c805, in805_1, in805_2, s641[0]);
    wire[0:0] s806, in806_1, in806_2;
    wire c806;
    assign in806_1 = {c744};
    assign in806_2 = {c745};
    Full_Adder FA_806(s806, c806, in806_1, in806_2, s644[0]);
    wire[0:0] s807, in807_1, in807_2;
    wire c807;
    assign in807_1 = {c746};
    assign in807_2 = {c747};
    Full_Adder FA_807(s807, c807, in807_1, in807_2, s647[0]);
    wire[0:0] s808, in808_1, in808_2;
    wire c808;
    assign in808_1 = {c748};
    assign in808_2 = {c749};
    Full_Adder FA_808(s808, c808, in808_1, in808_2, s649[0]);
    wire[0:0] s809, in809_1, in809_2;
    wire c809;
    assign in809_1 = {c750};
    assign in809_2 = {c751};
    Full_Adder FA_809(s809, c809, in809_1, in809_2, s650[0]);
    wire[0:0] s810, in810_1, in810_2;
    wire c810;
    assign in810_1 = {c752};
    assign in810_2 = {c753};
    Full_Adder FA_810(s810, c810, in810_1, in810_2, c650);
    wire[0:0] s811, in811_1, in811_2;
    wire c811;
    assign in811_1 = {pp31[27]};
    assign in811_2 = {c754};
    Full_Adder FA_811(s811, c811, in811_1, in811_2, pp30[28]);
    wire[0:0] s812, in812_1, in812_2;
    wire c812;
    assign in812_1 = {pp29[30]};
    assign in812_2 = {pp30[29]};
    Full_Adder FA_812(s812, c812, in812_1, in812_2, pp28[31]);

    /*Stage 7*/
    wire[0:0] s813, in813_1, in813_2;
    wire c813;
    assign in813_1 = {pp0[3]};
    assign in813_2 = {pp1[2]};
    Half_Adder HA_813(s813, c813, in813_1, in813_2);
    wire[0:0] s814, in814_1, in814_2;
    wire c814;
    assign in814_1 = {pp3[1]};
    assign in814_2 = {pp4[0]};
    Full_Adder FA_814(s814, c814, in814_1, in814_2, pp2[2]);
    wire[0:0] s815, in815_1, in815_2;
    wire c815;
    assign in815_1 = {s651[0]};
    assign in815_2 = {c757};
    Full_Adder FA_815(s815, c815, in815_1, in815_2, pp5[0]);
    wire[0:0] s816, in816_1, in816_2;
    wire c816;
    assign in816_1 = {s653[0]};
    assign in816_2 = {c758};
    Full_Adder FA_816(s816, c816, in816_1, in816_2, s652[0]);
    wire[0:0] s817, in817_1, in817_2;
    wire c817;
    assign in817_1 = {s655[0]};
    assign in817_2 = {c759};
    Full_Adder FA_817(s817, c817, in817_1, in817_2, s654[0]);
    wire[0:0] s818, in818_1, in818_2;
    wire c818;
    assign in818_1 = {s657[0]};
    assign in818_2 = {c760};
    Full_Adder FA_818(s818, c818, in818_1, in818_2, s656[0]);
    wire[0:0] s819, in819_1, in819_2;
    wire c819;
    assign in819_1 = {s659[0]};
    assign in819_2 = {c761};
    Full_Adder FA_819(s819, c819, in819_1, in819_2, s658[0]);
    wire[0:0] s820, in820_1, in820_2;
    wire c820;
    assign in820_1 = {s661[0]};
    assign in820_2 = {c762};
    Full_Adder FA_820(s820, c820, in820_1, in820_2, s660[0]);
    wire[0:0] s821, in821_1, in821_2;
    wire c821;
    assign in821_1 = {s663[0]};
    assign in821_2 = {c763};
    Full_Adder FA_821(s821, c821, in821_1, in821_2, s662[0]);
    wire[0:0] s822, in822_1, in822_2;
    wire c822;
    assign in822_1 = {s665[0]};
    assign in822_2 = {c764};
    Full_Adder FA_822(s822, c822, in822_1, in822_2, s664[0]);
    wire[0:0] s823, in823_1, in823_2;
    wire c823;
    assign in823_1 = {s667[0]};
    assign in823_2 = {c765};
    Full_Adder FA_823(s823, c823, in823_1, in823_2, s666[0]);
    wire[0:0] s824, in824_1, in824_2;
    wire c824;
    assign in824_1 = {s669[0]};
    assign in824_2 = {c766};
    Full_Adder FA_824(s824, c824, in824_1, in824_2, s668[0]);
    wire[0:0] s825, in825_1, in825_2;
    wire c825;
    assign in825_1 = {s671[0]};
    assign in825_2 = {c767};
    Full_Adder FA_825(s825, c825, in825_1, in825_2, s670[0]);
    wire[0:0] s826, in826_1, in826_2;
    wire c826;
    assign in826_1 = {s673[0]};
    assign in826_2 = {c768};
    Full_Adder FA_826(s826, c826, in826_1, in826_2, s672[0]);
    wire[0:0] s827, in827_1, in827_2;
    wire c827;
    assign in827_1 = {s675[0]};
    assign in827_2 = {c769};
    Full_Adder FA_827(s827, c827, in827_1, in827_2, s674[0]);
    wire[0:0] s828, in828_1, in828_2;
    wire c828;
    assign in828_1 = {s677[0]};
    assign in828_2 = {c770};
    Full_Adder FA_828(s828, c828, in828_1, in828_2, s676[0]);
    wire[0:0] s829, in829_1, in829_2;
    wire c829;
    assign in829_1 = {s679[0]};
    assign in829_2 = {c771};
    Full_Adder FA_829(s829, c829, in829_1, in829_2, s678[0]);
    wire[0:0] s830, in830_1, in830_2;
    wire c830;
    assign in830_1 = {s681[0]};
    assign in830_2 = {c772};
    Full_Adder FA_830(s830, c830, in830_1, in830_2, s680[0]);
    wire[0:0] s831, in831_1, in831_2;
    wire c831;
    assign in831_1 = {s683[0]};
    assign in831_2 = {c773};
    Full_Adder FA_831(s831, c831, in831_1, in831_2, s682[0]);
    wire[0:0] s832, in832_1, in832_2;
    wire c832;
    assign in832_1 = {s685[0]};
    assign in832_2 = {c774};
    Full_Adder FA_832(s832, c832, in832_1, in832_2, s684[0]);
    wire[0:0] s833, in833_1, in833_2;
    wire c833;
    assign in833_1 = {s687[0]};
    assign in833_2 = {c775};
    Full_Adder FA_833(s833, c833, in833_1, in833_2, s686[0]);
    wire[0:0] s834, in834_1, in834_2;
    wire c834;
    assign in834_1 = {s689[0]};
    assign in834_2 = {c776};
    Full_Adder FA_834(s834, c834, in834_1, in834_2, s688[0]);
    wire[0:0] s835, in835_1, in835_2;
    wire c835;
    assign in835_1 = {s691[0]};
    assign in835_2 = {c777};
    Full_Adder FA_835(s835, c835, in835_1, in835_2, s690[0]);
    wire[0:0] s836, in836_1, in836_2;
    wire c836;
    assign in836_1 = {s693[0]};
    assign in836_2 = {c778};
    Full_Adder FA_836(s836, c836, in836_1, in836_2, s692[0]);
    wire[0:0] s837, in837_1, in837_2;
    wire c837;
    assign in837_1 = {s695[0]};
    assign in837_2 = {c779};
    Full_Adder FA_837(s837, c837, in837_1, in837_2, s694[0]);
    wire[0:0] s838, in838_1, in838_2;
    wire c838;
    assign in838_1 = {s697[0]};
    assign in838_2 = {c780};
    Full_Adder FA_838(s838, c838, in838_1, in838_2, s696[0]);
    wire[0:0] s839, in839_1, in839_2;
    wire c839;
    assign in839_1 = {s699[0]};
    assign in839_2 = {c781};
    Full_Adder FA_839(s839, c839, in839_1, in839_2, s698[0]);
    wire[0:0] s840, in840_1, in840_2;
    wire c840;
    assign in840_1 = {s701[0]};
    assign in840_2 = {c782};
    Full_Adder FA_840(s840, c840, in840_1, in840_2, s700[0]);
    wire[0:0] s841, in841_1, in841_2;
    wire c841;
    assign in841_1 = {s703[0]};
    assign in841_2 = {c783};
    Full_Adder FA_841(s841, c841, in841_1, in841_2, s702[0]);
    wire[0:0] s842, in842_1, in842_2;
    wire c842;
    assign in842_1 = {s705[0]};
    assign in842_2 = {c784};
    Full_Adder FA_842(s842, c842, in842_1, in842_2, s704[0]);
    wire[0:0] s843, in843_1, in843_2;
    wire c843;
    assign in843_1 = {s707[0]};
    assign in843_2 = {c785};
    Full_Adder FA_843(s843, c843, in843_1, in843_2, s706[0]);
    wire[0:0] s844, in844_1, in844_2;
    wire c844;
    assign in844_1 = {s709[0]};
    assign in844_2 = {c786};
    Full_Adder FA_844(s844, c844, in844_1, in844_2, s708[0]);
    wire[0:0] s845, in845_1, in845_2;
    wire c845;
    assign in845_1 = {s711[0]};
    assign in845_2 = {c787};
    Full_Adder FA_845(s845, c845, in845_1, in845_2, s710[0]);
    wire[0:0] s846, in846_1, in846_2;
    wire c846;
    assign in846_1 = {s713[0]};
    assign in846_2 = {c788};
    Full_Adder FA_846(s846, c846, in846_1, in846_2, s712[0]);
    wire[0:0] s847, in847_1, in847_2;
    wire c847;
    assign in847_1 = {s715[0]};
    assign in847_2 = {c789};
    Full_Adder FA_847(s847, c847, in847_1, in847_2, s714[0]);
    wire[0:0] s848, in848_1, in848_2;
    wire c848;
    assign in848_1 = {s717[0]};
    assign in848_2 = {c790};
    Full_Adder FA_848(s848, c848, in848_1, in848_2, s716[0]);
    wire[0:0] s849, in849_1, in849_2;
    wire c849;
    assign in849_1 = {s719[0]};
    assign in849_2 = {c791};
    Full_Adder FA_849(s849, c849, in849_1, in849_2, s718[0]);
    wire[0:0] s850, in850_1, in850_2;
    wire c850;
    assign in850_1 = {s721[0]};
    assign in850_2 = {c792};
    Full_Adder FA_850(s850, c850, in850_1, in850_2, s720[0]);
    wire[0:0] s851, in851_1, in851_2;
    wire c851;
    assign in851_1 = {s723[0]};
    assign in851_2 = {c793};
    Full_Adder FA_851(s851, c851, in851_1, in851_2, s722[0]);
    wire[0:0] s852, in852_1, in852_2;
    wire c852;
    assign in852_1 = {s725[0]};
    assign in852_2 = {c794};
    Full_Adder FA_852(s852, c852, in852_1, in852_2, s724[0]);
    wire[0:0] s853, in853_1, in853_2;
    wire c853;
    assign in853_1 = {s727[0]};
    assign in853_2 = {c795};
    Full_Adder FA_853(s853, c853, in853_1, in853_2, s726[0]);
    wire[0:0] s854, in854_1, in854_2;
    wire c854;
    assign in854_1 = {s729[0]};
    assign in854_2 = {c796};
    Full_Adder FA_854(s854, c854, in854_1, in854_2, s728[0]);
    wire[0:0] s855, in855_1, in855_2;
    wire c855;
    assign in855_1 = {s731[0]};
    assign in855_2 = {c797};
    Full_Adder FA_855(s855, c855, in855_1, in855_2, s730[0]);
    wire[0:0] s856, in856_1, in856_2;
    wire c856;
    assign in856_1 = {s733[0]};
    assign in856_2 = {c798};
    Full_Adder FA_856(s856, c856, in856_1, in856_2, s732[0]);
    wire[0:0] s857, in857_1, in857_2;
    wire c857;
    assign in857_1 = {s735[0]};
    assign in857_2 = {c799};
    Full_Adder FA_857(s857, c857, in857_1, in857_2, s734[0]);
    wire[0:0] s858, in858_1, in858_2;
    wire c858;
    assign in858_1 = {s737[0]};
    assign in858_2 = {c800};
    Full_Adder FA_858(s858, c858, in858_1, in858_2, s736[0]);
    wire[0:0] s859, in859_1, in859_2;
    wire c859;
    assign in859_1 = {s739[0]};
    assign in859_2 = {c801};
    Full_Adder FA_859(s859, c859, in859_1, in859_2, s738[0]);
    wire[0:0] s860, in860_1, in860_2;
    wire c860;
    assign in860_1 = {s741[0]};
    assign in860_2 = {c802};
    Full_Adder FA_860(s860, c860, in860_1, in860_2, s740[0]);
    wire[0:0] s861, in861_1, in861_2;
    wire c861;
    assign in861_1 = {s743[0]};
    assign in861_2 = {c803};
    Full_Adder FA_861(s861, c861, in861_1, in861_2, s742[0]);
    wire[0:0] s862, in862_1, in862_2;
    wire c862;
    assign in862_1 = {s745[0]};
    assign in862_2 = {c804};
    Full_Adder FA_862(s862, c862, in862_1, in862_2, s744[0]);
    wire[0:0] s863, in863_1, in863_2;
    wire c863;
    assign in863_1 = {s747[0]};
    assign in863_2 = {c805};
    Full_Adder FA_863(s863, c863, in863_1, in863_2, s746[0]);
    wire[0:0] s864, in864_1, in864_2;
    wire c864;
    assign in864_1 = {s749[0]};
    assign in864_2 = {c806};
    Full_Adder FA_864(s864, c864, in864_1, in864_2, s748[0]);
    wire[0:0] s865, in865_1, in865_2;
    wire c865;
    assign in865_1 = {s751[0]};
    assign in865_2 = {c807};
    Full_Adder FA_865(s865, c865, in865_1, in865_2, s750[0]);
    wire[0:0] s866, in866_1, in866_2;
    wire c866;
    assign in866_1 = {s753[0]};
    assign in866_2 = {c808};
    Full_Adder FA_866(s866, c866, in866_1, in866_2, s752[0]);
    wire[0:0] s867, in867_1, in867_2;
    wire c867;
    assign in867_1 = {s755[0]};
    assign in867_2 = {c809};
    Full_Adder FA_867(s867, c867, in867_1, in867_2, s754[0]);
    wire[0:0] s868, in868_1, in868_2;
    wire c868;
    assign in868_1 = {s756[0]};
    assign in868_2 = {c810};
    Full_Adder FA_868(s868, c868, in868_1, in868_2, c755);
    wire[0:0] s869, in869_1, in869_2;
    wire c869;
    assign in869_1 = {c756};
    assign in869_2 = {c811};
    Full_Adder FA_869(s869, c869, in869_1, in869_2, pp31[28]);
    wire[0:0] s870, in870_1, in870_2;
    wire c870;
    assign in870_1 = {pp30[30]};
    assign in870_2 = {pp31[29]};
    Full_Adder FA_870(s870, c870, in870_1, in870_2, pp29[31]);

    /*Stage 8*/
    wire[0:0] s871, in871_1, in871_2;
    wire c871;
    assign in871_1 = {pp0[2]};
    assign in871_2 = {pp1[1]};
    Half_Adder HA_871(s871, c871, in871_1, in871_2);
    wire[0:0] s872, in872_1, in872_2;
    wire c872;
    assign in872_1 = {pp3[0]};
    assign in872_2 = {s813[0]};
    Full_Adder FA_872(s872, c872, in872_1, in872_2, pp2[1]);
    wire[0:0] s873, in873_1, in873_2;
    wire c873;
    assign in873_1 = {c813};
    assign in873_2 = {s814[0]};
    Full_Adder FA_873(s873, c873, in873_1, in873_2, s757[0]);
    wire[0:0] s874, in874_1, in874_2;
    wire c874;
    assign in874_1 = {c814};
    assign in874_2 = {s815[0]};
    Full_Adder FA_874(s874, c874, in874_1, in874_2, s758[0]);
    wire[0:0] s875, in875_1, in875_2;
    wire c875;
    assign in875_1 = {c815};
    assign in875_2 = {s816[0]};
    Full_Adder FA_875(s875, c875, in875_1, in875_2, s759[0]);
    wire[0:0] s876, in876_1, in876_2;
    wire c876;
    assign in876_1 = {c816};
    assign in876_2 = {s817[0]};
    Full_Adder FA_876(s876, c876, in876_1, in876_2, s760[0]);
    wire[0:0] s877, in877_1, in877_2;
    wire c877;
    assign in877_1 = {c817};
    assign in877_2 = {s818[0]};
    Full_Adder FA_877(s877, c877, in877_1, in877_2, s761[0]);
    wire[0:0] s878, in878_1, in878_2;
    wire c878;
    assign in878_1 = {c818};
    assign in878_2 = {s819[0]};
    Full_Adder FA_878(s878, c878, in878_1, in878_2, s762[0]);
    wire[0:0] s879, in879_1, in879_2;
    wire c879;
    assign in879_1 = {c819};
    assign in879_2 = {s820[0]};
    Full_Adder FA_879(s879, c879, in879_1, in879_2, s763[0]);
    wire[0:0] s880, in880_1, in880_2;
    wire c880;
    assign in880_1 = {c820};
    assign in880_2 = {s821[0]};
    Full_Adder FA_880(s880, c880, in880_1, in880_2, s764[0]);
    wire[0:0] s881, in881_1, in881_2;
    wire c881;
    assign in881_1 = {c821};
    assign in881_2 = {s822[0]};
    Full_Adder FA_881(s881, c881, in881_1, in881_2, s765[0]);
    wire[0:0] s882, in882_1, in882_2;
    wire c882;
    assign in882_1 = {c822};
    assign in882_2 = {s823[0]};
    Full_Adder FA_882(s882, c882, in882_1, in882_2, s766[0]);
    wire[0:0] s883, in883_1, in883_2;
    wire c883;
    assign in883_1 = {c823};
    assign in883_2 = {s824[0]};
    Full_Adder FA_883(s883, c883, in883_1, in883_2, s767[0]);
    wire[0:0] s884, in884_1, in884_2;
    wire c884;
    assign in884_1 = {c824};
    assign in884_2 = {s825[0]};
    Full_Adder FA_884(s884, c884, in884_1, in884_2, s768[0]);
    wire[0:0] s885, in885_1, in885_2;
    wire c885;
    assign in885_1 = {c825};
    assign in885_2 = {s826[0]};
    Full_Adder FA_885(s885, c885, in885_1, in885_2, s769[0]);
    wire[0:0] s886, in886_1, in886_2;
    wire c886;
    assign in886_1 = {c826};
    assign in886_2 = {s827[0]};
    Full_Adder FA_886(s886, c886, in886_1, in886_2, s770[0]);
    wire[0:0] s887, in887_1, in887_2;
    wire c887;
    assign in887_1 = {c827};
    assign in887_2 = {s828[0]};
    Full_Adder FA_887(s887, c887, in887_1, in887_2, s771[0]);
    wire[0:0] s888, in888_1, in888_2;
    wire c888;
    assign in888_1 = {c828};
    assign in888_2 = {s829[0]};
    Full_Adder FA_888(s888, c888, in888_1, in888_2, s772[0]);
    wire[0:0] s889, in889_1, in889_2;
    wire c889;
    assign in889_1 = {c829};
    assign in889_2 = {s830[0]};
    Full_Adder FA_889(s889, c889, in889_1, in889_2, s773[0]);
    wire[0:0] s890, in890_1, in890_2;
    wire c890;
    assign in890_1 = {c830};
    assign in890_2 = {s831[0]};
    Full_Adder FA_890(s890, c890, in890_1, in890_2, s774[0]);
    wire[0:0] s891, in891_1, in891_2;
    wire c891;
    assign in891_1 = {c831};
    assign in891_2 = {s832[0]};
    Full_Adder FA_891(s891, c891, in891_1, in891_2, s775[0]);
    wire[0:0] s892, in892_1, in892_2;
    wire c892;
    assign in892_1 = {c832};
    assign in892_2 = {s833[0]};
    Full_Adder FA_892(s892, c892, in892_1, in892_2, s776[0]);
    wire[0:0] s893, in893_1, in893_2;
    wire c893;
    assign in893_1 = {c833};
    assign in893_2 = {s834[0]};
    Full_Adder FA_893(s893, c893, in893_1, in893_2, s777[0]);
    wire[0:0] s894, in894_1, in894_2;
    wire c894;
    assign in894_1 = {c834};
    assign in894_2 = {s835[0]};
    Full_Adder FA_894(s894, c894, in894_1, in894_2, s778[0]);
    wire[0:0] s895, in895_1, in895_2;
    wire c895;
    assign in895_1 = {c835};
    assign in895_2 = {s836[0]};
    Full_Adder FA_895(s895, c895, in895_1, in895_2, s779[0]);
    wire[0:0] s896, in896_1, in896_2;
    wire c896;
    assign in896_1 = {c836};
    assign in896_2 = {s837[0]};
    Full_Adder FA_896(s896, c896, in896_1, in896_2, s780[0]);
    wire[0:0] s897, in897_1, in897_2;
    wire c897;
    assign in897_1 = {c837};
    assign in897_2 = {s838[0]};
    Full_Adder FA_897(s897, c897, in897_1, in897_2, s781[0]);
    wire[0:0] s898, in898_1, in898_2;
    wire c898;
    assign in898_1 = {c838};
    assign in898_2 = {s839[0]};
    Full_Adder FA_898(s898, c898, in898_1, in898_2, s782[0]);
    wire[0:0] s899, in899_1, in899_2;
    wire c899;
    assign in899_1 = {c839};
    assign in899_2 = {s840[0]};
    Full_Adder FA_899(s899, c899, in899_1, in899_2, s783[0]);
    wire[0:0] s900, in900_1, in900_2;
    wire c900;
    assign in900_1 = {c840};
    assign in900_2 = {s841[0]};
    Full_Adder FA_900(s900, c900, in900_1, in900_2, s784[0]);
    wire[0:0] s901, in901_1, in901_2;
    wire c901;
    assign in901_1 = {c841};
    assign in901_2 = {s842[0]};
    Full_Adder FA_901(s901, c901, in901_1, in901_2, s785[0]);
    wire[0:0] s902, in902_1, in902_2;
    wire c902;
    assign in902_1 = {c842};
    assign in902_2 = {s843[0]};
    Full_Adder FA_902(s902, c902, in902_1, in902_2, s786[0]);
    wire[0:0] s903, in903_1, in903_2;
    wire c903;
    assign in903_1 = {c843};
    assign in903_2 = {s844[0]};
    Full_Adder FA_903(s903, c903, in903_1, in903_2, s787[0]);
    wire[0:0] s904, in904_1, in904_2;
    wire c904;
    assign in904_1 = {c844};
    assign in904_2 = {s845[0]};
    Full_Adder FA_904(s904, c904, in904_1, in904_2, s788[0]);
    wire[0:0] s905, in905_1, in905_2;
    wire c905;
    assign in905_1 = {c845};
    assign in905_2 = {s846[0]};
    Full_Adder FA_905(s905, c905, in905_1, in905_2, s789[0]);
    wire[0:0] s906, in906_1, in906_2;
    wire c906;
    assign in906_1 = {c846};
    assign in906_2 = {s847[0]};
    Full_Adder FA_906(s906, c906, in906_1, in906_2, s790[0]);
    wire[0:0] s907, in907_1, in907_2;
    wire c907;
    assign in907_1 = {c847};
    assign in907_2 = {s848[0]};
    Full_Adder FA_907(s907, c907, in907_1, in907_2, s791[0]);
    wire[0:0] s908, in908_1, in908_2;
    wire c908;
    assign in908_1 = {c848};
    assign in908_2 = {s849[0]};
    Full_Adder FA_908(s908, c908, in908_1, in908_2, s792[0]);
    wire[0:0] s909, in909_1, in909_2;
    wire c909;
    assign in909_1 = {c849};
    assign in909_2 = {s850[0]};
    Full_Adder FA_909(s909, c909, in909_1, in909_2, s793[0]);
    wire[0:0] s910, in910_1, in910_2;
    wire c910;
    assign in910_1 = {c850};
    assign in910_2 = {s851[0]};
    Full_Adder FA_910(s910, c910, in910_1, in910_2, s794[0]);
    wire[0:0] s911, in911_1, in911_2;
    wire c911;
    assign in911_1 = {c851};
    assign in911_2 = {s852[0]};
    Full_Adder FA_911(s911, c911, in911_1, in911_2, s795[0]);
    wire[0:0] s912, in912_1, in912_2;
    wire c912;
    assign in912_1 = {c852};
    assign in912_2 = {s853[0]};
    Full_Adder FA_912(s912, c912, in912_1, in912_2, s796[0]);
    wire[0:0] s913, in913_1, in913_2;
    wire c913;
    assign in913_1 = {c853};
    assign in913_2 = {s854[0]};
    Full_Adder FA_913(s913, c913, in913_1, in913_2, s797[0]);
    wire[0:0] s914, in914_1, in914_2;
    wire c914;
    assign in914_1 = {c854};
    assign in914_2 = {s855[0]};
    Full_Adder FA_914(s914, c914, in914_1, in914_2, s798[0]);
    wire[0:0] s915, in915_1, in915_2;
    wire c915;
    assign in915_1 = {c855};
    assign in915_2 = {s856[0]};
    Full_Adder FA_915(s915, c915, in915_1, in915_2, s799[0]);
    wire[0:0] s916, in916_1, in916_2;
    wire c916;
    assign in916_1 = {c856};
    assign in916_2 = {s857[0]};
    Full_Adder FA_916(s916, c916, in916_1, in916_2, s800[0]);
    wire[0:0] s917, in917_1, in917_2;
    wire c917;
    assign in917_1 = {c857};
    assign in917_2 = {s858[0]};
    Full_Adder FA_917(s917, c917, in917_1, in917_2, s801[0]);
    wire[0:0] s918, in918_1, in918_2;
    wire c918;
    assign in918_1 = {c858};
    assign in918_2 = {s859[0]};
    Full_Adder FA_918(s918, c918, in918_1, in918_2, s802[0]);
    wire[0:0] s919, in919_1, in919_2;
    wire c919;
    assign in919_1 = {c859};
    assign in919_2 = {s860[0]};
    Full_Adder FA_919(s919, c919, in919_1, in919_2, s803[0]);
    wire[0:0] s920, in920_1, in920_2;
    wire c920;
    assign in920_1 = {c860};
    assign in920_2 = {s861[0]};
    Full_Adder FA_920(s920, c920, in920_1, in920_2, s804[0]);
    wire[0:0] s921, in921_1, in921_2;
    wire c921;
    assign in921_1 = {c861};
    assign in921_2 = {s862[0]};
    Full_Adder FA_921(s921, c921, in921_1, in921_2, s805[0]);
    wire[0:0] s922, in922_1, in922_2;
    wire c922;
    assign in922_1 = {c862};
    assign in922_2 = {s863[0]};
    Full_Adder FA_922(s922, c922, in922_1, in922_2, s806[0]);
    wire[0:0] s923, in923_1, in923_2;
    wire c923;
    assign in923_1 = {c863};
    assign in923_2 = {s864[0]};
    Full_Adder FA_923(s923, c923, in923_1, in923_2, s807[0]);
    wire[0:0] s924, in924_1, in924_2;
    wire c924;
    assign in924_1 = {c864};
    assign in924_2 = {s865[0]};
    Full_Adder FA_924(s924, c924, in924_1, in924_2, s808[0]);
    wire[0:0] s925, in925_1, in925_2;
    wire c925;
    assign in925_1 = {c865};
    assign in925_2 = {s866[0]};
    Full_Adder FA_925(s925, c925, in925_1, in925_2, s809[0]);
    wire[0:0] s926, in926_1, in926_2;
    wire c926;
    assign in926_1 = {c866};
    assign in926_2 = {s867[0]};
    Full_Adder FA_926(s926, c926, in926_1, in926_2, s810[0]);
    wire[0:0] s927, in927_1, in927_2;
    wire c927;
    assign in927_1 = {c867};
    assign in927_2 = {s868[0]};
    Full_Adder FA_927(s927, c927, in927_1, in927_2, s811[0]);
    wire[0:0] s928, in928_1, in928_2;
    wire c928;
    assign in928_1 = {c868};
    assign in928_2 = {s869[0]};
    Full_Adder FA_928(s928, c928, in928_1, in928_2, s812[0]);
    wire[0:0] s929, in929_1, in929_2;
    wire c929;
    assign in929_1 = {c869};
    assign in929_2 = {s870[0]};
    Full_Adder FA_929(s929, c929, in929_1, in929_2, c812);
    wire[0:0] s930, in930_1, in930_2;
    wire c930;
    assign in930_1 = {pp31[30]};
    assign in930_2 = {c870};
    Full_Adder FA_930(s930, c930, in930_1, in930_2, pp30[31]);


    /*Final Stage 8*/
    wire[61:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],c871,c872,c873,c874,c875,c876,c877,c878,c879,c880,c881,c882,c883,c884,c885,c886,c887,c888,c889,c890,c891,c892,c893,c894,c895,c896,c897,c898,c899,c900,c901,c902,c903,c904,c905,c906,c907,c908,c909,c910,c911,c912,c913,c914,c915,c916,c917,c918,c919,c920,c921,c922,c923,c924,c925,c926,c927,c928,c929,pp31[31]};
    assign in_2 = {pp1[0],s871[0],s872[0],s873[0],s874[0],s875[0],s876[0],s877[0],s878[0],s879[0],s880[0],s881[0],s882[0],s883[0],s884[0],s885[0],s886[0],s887[0],s888[0],s889[0],s890[0],s891[0],s892[0],s893[0],s894[0],s895[0],s896[0],s897[0],s898[0],s899[0],s900[0],s901[0],s902[0],s903[0],s904[0],s905[0],s906[0],s907[0],s908[0],s909[0],s910[0],s911[0],s912[0],s913[0],s914[0],s915[0],s916[0],s917[0],s918[0],s919[0],s920[0],s921[0],s922[0],s923[0],s924[0],s925[0],s926[0],s927[0],s928[0],s929[0],s930[0],c930};
    CLA_62(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = c;
endmodule


module CLA_62(output [61:0] sum, output cout, input [61:0] in1, input [61:0] in2);

    wire[61:0] G;
    wire[61:0] C;
    wire[61:0] P;

    assign G[0] = in1[61] & in2[61];
    assign P[0] = in1[61] ^ in2[61];
    assign G[1] = in1[60] & in2[60];
    assign P[1] = in1[60] ^ in2[60];
    assign G[2] = in1[59] & in2[59];
    assign P[2] = in1[59] ^ in2[59];
    assign G[3] = in1[58] & in2[58];
    assign P[3] = in1[58] ^ in2[58];
    assign G[4] = in1[57] & in2[57];
    assign P[4] = in1[57] ^ in2[57];
    assign G[5] = in1[56] & in2[56];
    assign P[5] = in1[56] ^ in2[56];
    assign G[6] = in1[55] & in2[55];
    assign P[6] = in1[55] ^ in2[55];
    assign G[7] = in1[54] & in2[54];
    assign P[7] = in1[54] ^ in2[54];
    assign G[8] = in1[53] & in2[53];
    assign P[8] = in1[53] ^ in2[53];
    assign G[9] = in1[52] & in2[52];
    assign P[9] = in1[52] ^ in2[52];
    assign G[10] = in1[51] & in2[51];
    assign P[10] = in1[51] ^ in2[51];
    assign G[11] = in1[50] & in2[50];
    assign P[11] = in1[50] ^ in2[50];
    assign G[12] = in1[49] & in2[49];
    assign P[12] = in1[49] ^ in2[49];
    assign G[13] = in1[48] & in2[48];
    assign P[13] = in1[48] ^ in2[48];
    assign G[14] = in1[47] & in2[47];
    assign P[14] = in1[47] ^ in2[47];
    assign G[15] = in1[46] & in2[46];
    assign P[15] = in1[46] ^ in2[46];
    assign G[16] = in1[45] & in2[45];
    assign P[16] = in1[45] ^ in2[45];
    assign G[17] = in1[44] & in2[44];
    assign P[17] = in1[44] ^ in2[44];
    assign G[18] = in1[43] & in2[43];
    assign P[18] = in1[43] ^ in2[43];
    assign G[19] = in1[42] & in2[42];
    assign P[19] = in1[42] ^ in2[42];
    assign G[20] = in1[41] & in2[41];
    assign P[20] = in1[41] ^ in2[41];
    assign G[21] = in1[40] & in2[40];
    assign P[21] = in1[40] ^ in2[40];
    assign G[22] = in1[39] & in2[39];
    assign P[22] = in1[39] ^ in2[39];
    assign G[23] = in1[38] & in2[38];
    assign P[23] = in1[38] ^ in2[38];
    assign G[24] = in1[37] & in2[37];
    assign P[24] = in1[37] ^ in2[37];
    assign G[25] = in1[36] & in2[36];
    assign P[25] = in1[36] ^ in2[36];
    assign G[26] = in1[35] & in2[35];
    assign P[26] = in1[35] ^ in2[35];
    assign G[27] = in1[34] & in2[34];
    assign P[27] = in1[34] ^ in2[34];
    assign G[28] = in1[33] & in2[33];
    assign P[28] = in1[33] ^ in2[33];
    assign G[29] = in1[32] & in2[32];
    assign P[29] = in1[32] ^ in2[32];
    assign G[30] = in1[31] & in2[31];
    assign P[30] = in1[31] ^ in2[31];
    assign G[31] = in1[30] & in2[30];
    assign P[31] = in1[30] ^ in2[30];
    assign G[32] = in1[29] & in2[29];
    assign P[32] = in1[29] ^ in2[29];
    assign G[33] = in1[28] & in2[28];
    assign P[33] = in1[28] ^ in2[28];
    assign G[34] = in1[27] & in2[27];
    assign P[34] = in1[27] ^ in2[27];
    assign G[35] = in1[26] & in2[26];
    assign P[35] = in1[26] ^ in2[26];
    assign G[36] = in1[25] & in2[25];
    assign P[36] = in1[25] ^ in2[25];
    assign G[37] = in1[24] & in2[24];
    assign P[37] = in1[24] ^ in2[24];
    assign G[38] = in1[23] & in2[23];
    assign P[38] = in1[23] ^ in2[23];
    assign G[39] = in1[22] & in2[22];
    assign P[39] = in1[22] ^ in2[22];
    assign G[40] = in1[21] & in2[21];
    assign P[40] = in1[21] ^ in2[21];
    assign G[41] = in1[20] & in2[20];
    assign P[41] = in1[20] ^ in2[20];
    assign G[42] = in1[19] & in2[19];
    assign P[42] = in1[19] ^ in2[19];
    assign G[43] = in1[18] & in2[18];
    assign P[43] = in1[18] ^ in2[18];
    assign G[44] = in1[17] & in2[17];
    assign P[44] = in1[17] ^ in2[17];
    assign G[45] = in1[16] & in2[16];
    assign P[45] = in1[16] ^ in2[16];
    assign G[46] = in1[15] & in2[15];
    assign P[46] = in1[15] ^ in2[15];
    assign G[47] = in1[14] & in2[14];
    assign P[47] = in1[14] ^ in2[14];
    assign G[48] = in1[13] & in2[13];
    assign P[48] = in1[13] ^ in2[13];
    assign G[49] = in1[12] & in2[12];
    assign P[49] = in1[12] ^ in2[12];
    assign G[50] = in1[11] & in2[11];
    assign P[50] = in1[11] ^ in2[11];
    assign G[51] = in1[10] & in2[10];
    assign P[51] = in1[10] ^ in2[10];
    assign G[52] = in1[9] & in2[9];
    assign P[52] = in1[9] ^ in2[9];
    assign G[53] = in1[8] & in2[8];
    assign P[53] = in1[8] ^ in2[8];
    assign G[54] = in1[7] & in2[7];
    assign P[54] = in1[7] ^ in2[7];
    assign G[55] = in1[6] & in2[6];
    assign P[55] = in1[6] ^ in2[6];
    assign G[56] = in1[5] & in2[5];
    assign P[56] = in1[5] ^ in2[5];
    assign G[57] = in1[4] & in2[4];
    assign P[57] = in1[4] ^ in2[4];
    assign G[58] = in1[3] & in2[3];
    assign P[58] = in1[3] ^ in2[3];
    assign G[59] = in1[2] & in2[2];
    assign P[59] = in1[2] ^ in2[2];
    assign G[60] = in1[1] & in2[1];
    assign P[60] = in1[1] ^ in2[1];
    assign G[61] = in1[0] & in2[0];
    assign P[61] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign cout = G[61] | (P[61] & C[61]);
    assign sum = P ^ C;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule

