module multiplier_128bits_version12(product, A, B);

    output [255:0] product;
    input [127:0] A, B;

    wire [127:0] pp0;
    wire [127:0] pp1;
    wire [127:0] pp2;
    wire [127:0] pp3;
    wire [127:0] pp4;
    wire [127:0] pp5;
    wire [127:0] pp6;
    wire [127:0] pp7;
    wire [127:0] pp8;
    wire [127:0] pp9;
    wire [127:0] pp10;
    wire [127:0] pp11;
    wire [127:0] pp12;
    wire [127:0] pp13;
    wire [127:0] pp14;
    wire [127:0] pp15;
    wire [127:0] pp16;
    wire [127:0] pp17;
    wire [127:0] pp18;
    wire [127:0] pp19;
    wire [127:0] pp20;
    wire [127:0] pp21;
    wire [127:0] pp22;
    wire [127:0] pp23;
    wire [127:0] pp24;
    wire [127:0] pp25;
    wire [127:0] pp26;
    wire [127:0] pp27;
    wire [127:0] pp28;
    wire [127:0] pp29;
    wire [127:0] pp30;
    wire [127:0] pp31;
    wire [127:0] pp32;
    wire [127:0] pp33;
    wire [127:0] pp34;
    wire [127:0] pp35;
    wire [127:0] pp36;
    wire [127:0] pp37;
    wire [127:0] pp38;
    wire [127:0] pp39;
    wire [127:0] pp40;
    wire [127:0] pp41;
    wire [127:0] pp42;
    wire [127:0] pp43;
    wire [127:0] pp44;
    wire [127:0] pp45;
    wire [127:0] pp46;
    wire [127:0] pp47;
    wire [127:0] pp48;
    wire [127:0] pp49;
    wire [127:0] pp50;
    wire [127:0] pp51;
    wire [127:0] pp52;
    wire [127:0] pp53;
    wire [127:0] pp54;
    wire [127:0] pp55;
    wire [127:0] pp56;
    wire [127:0] pp57;
    wire [127:0] pp58;
    wire [127:0] pp59;
    wire [127:0] pp60;
    wire [127:0] pp61;
    wire [127:0] pp62;
    wire [127:0] pp63;
    wire [127:0] pp64;
    wire [127:0] pp65;
    wire [127:0] pp66;
    wire [127:0] pp67;
    wire [127:0] pp68;
    wire [127:0] pp69;
    wire [127:0] pp70;
    wire [127:0] pp71;
    wire [127:0] pp72;
    wire [127:0] pp73;
    wire [127:0] pp74;
    wire [127:0] pp75;
    wire [127:0] pp76;
    wire [127:0] pp77;
    wire [127:0] pp78;
    wire [127:0] pp79;
    wire [127:0] pp80;
    wire [127:0] pp81;
    wire [127:0] pp82;
    wire [127:0] pp83;
    wire [127:0] pp84;
    wire [127:0] pp85;
    wire [127:0] pp86;
    wire [127:0] pp87;
    wire [127:0] pp88;
    wire [127:0] pp89;
    wire [127:0] pp90;
    wire [127:0] pp91;
    wire [127:0] pp92;
    wire [127:0] pp93;
    wire [127:0] pp94;
    wire [127:0] pp95;
    wire [127:0] pp96;
    wire [127:0] pp97;
    wire [127:0] pp98;
    wire [127:0] pp99;
    wire [127:0] pp100;
    wire [127:0] pp101;
    wire [127:0] pp102;
    wire [127:0] pp103;
    wire [127:0] pp104;
    wire [127:0] pp105;
    wire [127:0] pp106;
    wire [127:0] pp107;
    wire [127:0] pp108;
    wire [127:0] pp109;
    wire [127:0] pp110;
    wire [127:0] pp111;
    wire [127:0] pp112;
    wire [127:0] pp113;
    wire [127:0] pp114;
    wire [127:0] pp115;
    wire [127:0] pp116;
    wire [127:0] pp117;
    wire [127:0] pp118;
    wire [127:0] pp119;
    wire [127:0] pp120;
    wire [127:0] pp121;
    wire [127:0] pp122;
    wire [127:0] pp123;
    wire [127:0] pp124;
    wire [127:0] pp125;
    wire [127:0] pp126;
    wire [127:0] pp127;


    assign pp0 = A[0] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp64 = A[64] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp65 = A[65] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp66 = A[66] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp67 = A[67] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp68 = A[68] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp69 = A[69] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp70 = A[70] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp71 = A[71] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp72 = A[72] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp73 = A[73] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp74 = A[74] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp75 = A[75] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp76 = A[76] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp77 = A[77] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp78 = A[78] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp79 = A[79] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp80 = A[80] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp81 = A[81] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp82 = A[82] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp83 = A[83] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp84 = A[84] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp85 = A[85] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp86 = A[86] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp87 = A[87] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp88 = A[88] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp89 = A[89] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp90 = A[90] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp91 = A[91] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp92 = A[92] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp93 = A[93] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp94 = A[94] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp95 = A[95] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp96 = A[96] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp97 = A[97] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp98 = A[98] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp99 = A[99] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp100 = A[100] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp101 = A[101] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp102 = A[102] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp103 = A[103] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp104 = A[104] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp105 = A[105] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp106 = A[106] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp107 = A[107] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp108 = A[108] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp109 = A[109] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp110 = A[110] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp111 = A[111] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp112 = A[112] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp113 = A[113] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp114 = A[114] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp115 = A[115] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp116 = A[116] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp117 = A[117] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp118 = A[118] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp119 = A[119] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp120 = A[120] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp121 = A[121] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp122 = A[122] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp123 = A[123] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp124 = A[124] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp125 = A[125] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp126 = A[126] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp127 = A[127] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[3:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[76],pp0[77],pp0[78],pp0[79]};
    assign in1_2 = {pp1[75],pp1[76],pp1[77],pp1[78]};
    CLA_4 KS_1(s1, c1, in1_1, in1_2);
    wire[3:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp2[75],pp2[76],pp2[77],pp0[80]};
    assign in2_2 = {pp3[74],pp3[75],pp3[76],pp1[79]};
    CLA_4 KS_2(s2, c2, in2_1, in2_2);
    wire[3:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp4[74],pp4[75],pp2[78],pp0[81]};
    assign in3_2 = {pp5[73],pp5[74],pp3[77],pp1[80]};
    CLA_4 KS_3(s3, c3, in3_1, in3_2);
    wire[3:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp6[73],pp4[76],pp2[79],pp0[82]};
    assign in4_2 = {pp7[72],pp5[75],pp3[78],pp1[81]};
    CLA_4 KS_4(s4, c4, in4_1, in4_2);
    wire[3:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp6[74],pp4[77],pp2[80],pp0[83]};
    assign in5_2 = {pp7[73],pp5[76],pp3[79],pp1[82]};
    CLA_4 KS_5(s5, c5, in5_1, in5_2);
    wire[3:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp9[71],pp6[75],pp4[78],pp2[81]};
    assign in6_2 = {pp10[70],pp7[74],pp5[77],pp3[80]};
    CLA_4_c KS_6(s6, c6, in6_1, in6_2, pp8[72]);
    wire[3:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp8[73],pp6[76],pp4[79],pp0[84]};
    assign in7_2 = {pp9[72],pp7[75],pp5[78],pp1[83]};
    CLA_4 KS_7(s7, c7, in7_1, in7_2);
    wire[3:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp11[70],pp8[74],pp6[77],pp2[82]};
    assign in8_2 = {pp12[69],pp9[73],pp7[76],pp3[81]};
    CLA_4_c KS_8(s8, c8, in8_1, in8_2, pp10[71]);
    wire[3:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp10[72],pp8[75],pp4[80],pp0[85]};
    assign in9_2 = {pp11[71],pp9[74],pp5[79],pp1[84]};
    CLA_4 KS_9(s9, c9, in9_1, in9_2);
    wire[3:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp13[69],pp10[73],pp6[78],pp2[83]};
    assign in10_2 = {pp14[68],pp11[72],pp7[77],pp3[82]};
    CLA_4_c KS_10(s10, c10, in10_1, in10_2, pp12[70]);
    wire[3:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp12[71],pp8[76],pp4[81],pp0[86]};
    assign in11_2 = {pp13[70],pp9[75],pp5[80],pp1[85]};
    CLA_4 KS_11(s11, c11, in11_1, in11_2);
    wire[3:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp15[68],pp10[74],pp6[79],pp2[84]};
    assign in12_2 = {pp16[67],pp11[73],pp7[78],pp3[83]};
    CLA_4_c KS_12(s12, c12, in12_1, in12_2, pp14[69]);
    wire[3:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp12[72],pp8[77],pp4[82],pp0[87]};
    assign in13_2 = {pp13[71],pp9[76],pp5[81],pp1[86]};
    CLA_4 KS_13(s13, c13, in13_1, in13_2);
    wire[3:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp14[70],pp10[75],pp6[80],pp2[85]};
    assign in14_2 = {pp15[69],pp11[74],pp7[79],pp3[84]};
    CLA_4 KS_14(s14, c14, in14_1, in14_2);
    wire[3:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp16[68],pp12[73],pp8[78],pp4[83]};
    assign in15_2 = {pp17[67],pp13[72],pp9[77],pp5[82]};
    CLA_4 KS_15(s15, c15, in15_1, in15_2);
    wire[3:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp19[65],pp14[71],pp10[76],pp6[81]};
    assign in16_2 = {pp20[64],pp15[70],pp11[75],pp7[80]};
    CLA_4_c KS_16(s16, c16, in16_1, in16_2, pp18[66]);
    wire[3:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp16[69],pp12[74],pp8[79],pp0[88]};
    assign in17_2 = {pp17[68],pp13[73],pp9[78],pp1[87]};
    CLA_4 KS_17(s17, c17, in17_1, in17_2);
    wire[3:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp18[67],pp14[72],pp10[77],pp2[86]};
    assign in18_2 = {pp19[66],pp15[71],pp11[76],pp3[85]};
    CLA_4 KS_18(s18, c18, in18_1, in18_2);
    wire[3:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp21[64],pp16[70],pp12[75],pp4[84]};
    assign in19_2 = {pp22[63],pp17[69],pp13[74],pp5[83]};
    CLA_4_c KS_19(s19, c19, in19_1, in19_2, pp20[65]);
    wire[3:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp18[68],pp14[73],pp6[82],pp0[89]};
    assign in20_2 = {pp19[67],pp15[72],pp7[81],pp1[88]};
    CLA_4 KS_20(s20, c20, in20_1, in20_2);
    wire[3:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp20[66],pp16[71],pp8[80],pp2[87]};
    assign in21_2 = {pp21[65],pp17[70],pp9[79],pp3[86]};
    CLA_4 KS_21(s21, c21, in21_1, in21_2);
    wire[3:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp23[63],pp18[69],pp10[78],pp4[85]};
    assign in22_2 = {pp24[62],pp19[68],pp11[77],pp5[84]};
    CLA_4_c KS_22(s22, c22, in22_1, in22_2, pp22[64]);
    wire[3:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp20[67],pp12[76],pp6[83],pp0[90]};
    assign in23_2 = {pp21[66],pp13[75],pp7[82],pp1[89]};
    CLA_4 KS_23(s23, c23, in23_1, in23_2);
    wire[3:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp22[65],pp14[74],pp8[81],pp2[88]};
    assign in24_2 = {pp23[64],pp15[73],pp9[80],pp3[87]};
    CLA_4 KS_24(s24, c24, in24_1, in24_2);
    wire[3:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp25[62],pp16[72],pp10[79],pp4[86]};
    assign in25_2 = {pp26[61],pp17[71],pp11[78],pp5[85]};
    CLA_4_c KS_25(s25, c25, in25_1, in25_2, pp24[63]);
    wire[3:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp18[70],pp12[77],pp6[84],pp0[91]};
    assign in26_2 = {pp19[69],pp13[76],pp7[83],pp1[90]};
    CLA_4 KS_26(s26, c26, in26_1, in26_2);
    wire[3:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp20[68],pp14[75],pp8[82],pp2[89]};
    assign in27_2 = {pp21[67],pp15[74],pp9[81],pp3[88]};
    CLA_4 KS_27(s27, c27, in27_1, in27_2);
    wire[3:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp22[66],pp16[73],pp10[80],pp4[87]};
    assign in28_2 = {pp23[65],pp17[72],pp11[79],pp5[86]};
    CLA_4 KS_28(s28, c28, in28_1, in28_2);
    wire[3:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp24[64],pp18[71],pp12[78],pp6[85]};
    assign in29_2 = {pp25[63],pp19[70],pp13[77],pp7[84]};
    CLA_4 KS_29(s29, c29, in29_1, in29_2);
    wire[3:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp26[62],pp20[69],pp14[76],pp8[83]};
    assign in30_2 = {pp27[61],pp21[68],pp15[75],pp9[82]};
    CLA_4 KS_30(s30, c30, in30_1, in30_2);
    wire[3:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp28[60],pp22[67],pp16[74],pp10[81]};
    assign in31_2 = {pp29[59],pp23[66],pp17[73],pp11[80]};
    CLA_4 KS_31(s31, c31, in31_1, in31_2);
    wire[3:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp31[57],pp24[65],pp18[72],pp12[79]};
    assign in32_2 = {pp32[56],pp25[64],pp19[71],pp13[78]};
    CLA_4_c KS_32(s32, c32, in32_1, in32_2, pp30[58]);
    wire[3:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp26[63],pp20[70],pp14[77],pp0[92]};
    assign in33_2 = {pp27[62],pp21[69],pp15[76],pp1[91]};
    CLA_4 KS_33(s33, c33, in33_1, in33_2);
    wire[3:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp28[61],pp22[68],pp16[75],pp2[90]};
    assign in34_2 = {pp29[60],pp23[67],pp17[74],pp3[89]};
    CLA_4 KS_34(s34, c34, in34_1, in34_2);
    wire[3:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp31[58],pp24[66],pp18[73],pp4[88]};
    assign in35_2 = {pp32[57],pp25[65],pp19[72],pp5[87]};
    CLA_4_c KS_35(s35, c35, in35_1, in35_2, pp30[59]);
    wire[3:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp26[64],pp20[71],pp6[86],pp0[93]};
    assign in36_2 = {pp27[63],pp21[70],pp7[85],pp1[92]};
    CLA_4 KS_36(s36, c36, in36_1, in36_2);
    wire[3:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp28[62],pp22[69],pp8[84],pp2[91]};
    assign in37_2 = {pp29[61],pp23[68],pp9[83],pp3[90]};
    CLA_4 KS_37(s37, c37, in37_1, in37_2);
    wire[3:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp30[60],pp24[67],pp10[82],pp4[89]};
    assign in38_2 = {pp31[59],pp25[66],pp11[81],pp5[88]};
    CLA_4 KS_38(s38, c38, in38_1, in38_2);
    wire[3:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp33[57],pp26[65],pp12[80],pp6[87]};
    assign in39_2 = {pp34[56],pp27[64],pp13[79],pp7[86]};
    CLA_4_c KS_39(s39, c39, in39_1, in39_2, pp32[58]);
    wire[3:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp28[63],pp14[78],pp8[85],pp0[94]};
    assign in40_2 = {pp29[62],pp15[77],pp9[84],pp1[93]};
    CLA_4 KS_40(s40, c40, in40_1, in40_2);
    wire[3:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp30[61],pp16[76],pp10[83],pp2[92]};
    assign in41_2 = {pp31[60],pp17[75],pp11[82],pp3[91]};
    CLA_4 KS_41(s41, c41, in41_1, in41_2);
    wire[3:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp32[59],pp18[74],pp12[81],pp4[90]};
    assign in42_2 = {pp33[58],pp19[73],pp13[80],pp5[89]};
    CLA_4 KS_42(s42, c42, in42_1, in42_2);
    wire[3:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp35[56],pp20[72],pp14[79],pp6[88]};
    assign in43_2 = {pp36[55],pp21[71],pp15[78],pp7[87]};
    CLA_4_c KS_43(s43, c43, in43_1, in43_2, pp34[57]);
    wire[3:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[70],pp16[77],pp8[86],pp0[95]};
    assign in44_2 = {pp23[69],pp17[76],pp9[85],pp1[94]};
    CLA_4 KS_44(s44, c44, in44_1, in44_2);
    wire[3:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[68],pp18[75],pp10[84],pp2[93]};
    assign in45_2 = {pp25[67],pp19[74],pp11[83],pp3[92]};
    CLA_4 KS_45(s45, c45, in45_1, in45_2);
    wire[3:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp26[66],pp20[73],pp12[82],pp4[91]};
    assign in46_2 = {pp27[65],pp21[72],pp13[81],pp5[90]};
    CLA_4 KS_46(s46, c46, in46_1, in46_2);
    wire[3:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp28[64],pp22[71],pp14[80],pp6[89]};
    assign in47_2 = {pp29[63],pp23[70],pp15[79],pp7[88]};
    CLA_4 KS_47(s47, c47, in47_1, in47_2);
    wire[3:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp30[62],pp24[69],pp16[78],pp8[87]};
    assign in48_2 = {pp31[61],pp25[68],pp17[77],pp9[86]};
    CLA_4 KS_48(s48, c48, in48_1, in48_2);
    wire[3:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp32[60],pp26[67],pp18[76],pp10[85]};
    assign in49_2 = {pp33[59],pp27[66],pp19[75],pp11[84]};
    CLA_4 KS_49(s49, c49, in49_1, in49_2);
    wire[3:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp34[58],pp28[65],pp20[74],pp12[83]};
    assign in50_2 = {pp35[57],pp29[64],pp21[73],pp13[82]};
    CLA_4 KS_50(s50, c50, in50_1, in50_2);
    wire[3:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp36[56],pp30[63],pp22[72],pp14[81]};
    assign in51_2 = {pp37[55],pp31[62],pp23[71],pp15[80]};
    CLA_4 KS_51(s51, c51, in51_1, in51_2);
    wire[3:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp38[54],pp32[61],pp24[70],pp16[79]};
    assign in52_2 = {pp39[53],pp33[60],pp25[69],pp17[78]};
    CLA_4 KS_52(s52, c52, in52_1, in52_2);
    wire[3:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp40[52],pp34[59],pp26[68],pp18[77]};
    assign in53_2 = {pp41[51],pp35[58],pp27[67],pp19[76]};
    CLA_4 KS_53(s53, c53, in53_1, in53_2);
    wire[3:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp42[50],pp36[57],pp28[66],pp20[75]};
    assign in54_2 = {pp43[49],pp37[56],pp29[65],pp21[74]};
    CLA_4 KS_54(s54, c54, in54_1, in54_2);
    wire[3:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp45[47],pp38[55],pp30[64],pp22[73]};
    assign in55_2 = {pp46[46],pp39[54],pp31[63],pp23[72]};
    CLA_4_c KS_55(s55, c55, in55_1, in55_2, pp44[48]);
    wire[3:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp40[53],pp32[62],pp24[71],pp0[96]};
    assign in56_2 = {pp41[52],pp33[61],pp25[70],pp1[95]};
    CLA_4 KS_56(s56, c56, in56_1, in56_2);
    wire[3:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp34[60],pp26[69],pp2[94],pp0[97]};
    assign in57_2 = {pp35[59],pp27[68],pp3[93],pp1[96]};
    CLA_4 KS_57(s57, c57, in57_1, in57_2);
    wire[3:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp36[58],pp28[67],pp4[92],pp2[95]};
    assign in58_2 = {pp37[57],pp29[66],pp5[91],pp3[94]};
    CLA_4 KS_58(s58, c58, in58_1, in58_2);
    wire[3:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp38[56],pp30[65],pp6[90],pp4[93]};
    assign in59_2 = {pp39[55],pp31[64],pp7[89],pp5[92]};
    CLA_4 KS_59(s59, c59, in59_1, in59_2);
    wire[3:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp40[54],pp32[63],pp8[88],pp6[91]};
    assign in60_2 = {pp41[53],pp33[62],pp9[87],pp7[90]};
    CLA_4 KS_60(s60, c60, in60_1, in60_2);
    wire[3:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp43[51],pp34[61],pp10[86],pp8[89]};
    assign in61_2 = {pp44[50],pp35[60],pp11[85],pp9[88]};
    CLA_4_c KS_61(s61, c61, in61_1, in61_2, pp42[52]);
    wire[3:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp36[59],pp12[84],pp10[87],pp0[98]};
    assign in62_2 = {pp37[58],pp13[83],pp11[86],pp1[97]};
    CLA_4 KS_62(s62, c62, in62_1, in62_2);
    wire[3:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp38[57],pp14[82],pp12[85],pp2[96]};
    assign in63_2 = {pp39[56],pp15[81],pp13[84],pp3[95]};
    CLA_4 KS_63(s63, c63, in63_1, in63_2);
    wire[3:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp40[55],pp16[80],pp14[83],pp4[94]};
    assign in64_2 = {pp41[54],pp17[79],pp15[82],pp5[93]};
    CLA_4 KS_64(s64, c64, in64_1, in64_2);
    wire[3:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp42[53],pp18[78],pp16[81],pp6[92]};
    assign in65_2 = {pp43[52],pp19[77],pp17[80],pp7[91]};
    CLA_4 KS_65(s65, c65, in65_1, in65_2);
    wire[3:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp45[50],pp20[76],pp18[79],pp8[90]};
    assign in66_2 = {pp46[49],pp21[75],pp19[78],pp9[89]};
    CLA_4_c KS_66(s66, c66, in66_1, in66_2, pp44[51]);
    wire[3:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp22[74],pp20[77],pp10[88],pp0[99]};
    assign in67_2 = {pp23[73],pp21[76],pp11[87],pp1[98]};
    CLA_4 KS_67(s67, c67, in67_1, in67_2);
    wire[3:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp24[72],pp22[75],pp12[86],pp2[97]};
    assign in68_2 = {pp25[71],pp23[74],pp13[85],pp3[96]};
    CLA_4 KS_68(s68, c68, in68_1, in68_2);
    wire[3:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp26[70],pp24[73],pp14[84],pp4[95]};
    assign in69_2 = {pp27[69],pp25[72],pp15[83],pp5[94]};
    CLA_4 KS_69(s69, c69, in69_1, in69_2);
    wire[3:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp28[68],pp26[71],pp16[82],pp6[93]};
    assign in70_2 = {pp29[67],pp27[70],pp17[81],pp7[92]};
    CLA_4 KS_70(s70, c70, in70_1, in70_2);
    wire[3:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp30[66],pp28[69],pp18[80],pp8[91]};
    assign in71_2 = {pp31[65],pp29[68],pp19[79],pp9[90]};
    CLA_4 KS_71(s71, c71, in71_1, in71_2);
    wire[3:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp32[64],pp30[67],pp20[78],pp10[89]};
    assign in72_2 = {pp33[63],pp31[66],pp21[77],pp11[88]};
    CLA_4 KS_72(s72, c72, in72_1, in72_2);
    wire[3:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp34[62],pp32[65],pp22[76],pp12[87]};
    assign in73_2 = {pp35[61],pp33[64],pp23[75],pp13[86]};
    CLA_4 KS_73(s73, c73, in73_1, in73_2);
    wire[3:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp36[60],pp34[63],pp24[74],pp14[85]};
    assign in74_2 = {pp37[59],pp35[62],pp25[73],pp15[84]};
    CLA_4 KS_74(s74, c74, in74_1, in74_2);
    wire[3:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp38[58],pp36[61],pp26[72],pp16[83]};
    assign in75_2 = {pp39[57],pp37[60],pp27[71],pp17[82]};
    CLA_4 KS_75(s75, c75, in75_1, in75_2);
    wire[3:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp40[56],pp38[59],pp28[70],pp18[81]};
    assign in76_2 = {pp41[55],pp39[58],pp29[69],pp19[80]};
    CLA_4 KS_76(s76, c76, in76_1, in76_2);
    wire[3:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp42[54],pp40[57],pp30[68],pp20[79]};
    assign in77_2 = {pp43[53],pp41[56],pp31[67],pp21[78]};
    CLA_4 KS_77(s77, c77, in77_1, in77_2);
    wire[3:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp44[52],pp42[55],pp32[66],pp22[77]};
    assign in78_2 = {pp45[51],pp43[54],pp33[65],pp23[76]};
    CLA_4 KS_78(s78, c78, in78_1, in78_2);
    wire[3:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp46[50],pp44[53],pp34[64],pp24[75]};
    assign in79_2 = {pp47[49],pp45[52],pp35[63],pp25[74]};
    CLA_4 KS_79(s79, c79, in79_1, in79_2);
    wire[3:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp48[48],pp46[51],pp36[62],pp26[73]};
    assign in80_2 = {pp49[47],pp47[50],pp37[61],pp27[72]};
    CLA_4 KS_80(s80, c80, in80_1, in80_2);
    wire[0:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp50[46]};
    assign in81_2 = {pp51[45]};
    Half_Adder KS_81(s81, c81, in81_1, in81_2);
    wire[3:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp52[44],pp48[49],pp38[60],pp28[71]};
    assign in82_2 = {pp53[43],pp49[48],pp39[59],pp29[70]};
    CLA_4 KS_82(s82, c82, in82_1, in82_2);
    wire[0:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp54[42]};
    assign in83_2 = {pp55[41]};
    Half_Adder KS_83(s83, c83, in83_1, in83_2);
    wire[3:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp56[40],pp50[47],pp40[58],pp30[69]};
    assign in84_2 = {pp57[39],pp51[46],pp41[57],pp31[68]};
    CLA_4 KS_84(s84, c84, in84_1, in84_2);
    wire[0:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp58[38]};
    assign in85_2 = {pp59[37]};
    Half_Adder KS_85(s85, c85, in85_1, in85_2);
    wire[3:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp60[36],pp52[45],pp42[56],pp32[67]};
    assign in86_2 = {pp61[35],pp53[44],pp43[55],pp33[66]};
    CLA_4 KS_86(s86, c86, in86_1, in86_2);
    wire[0:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp63[33]};
    assign in87_2 = {pp64[32]};
    Full_Adder KS_87(s87, c87, in87_1, in87_2, pp62[34]);
    wire[3:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp44[54],pp34[65],pp0[100],pp0[101]};
    assign in88_2 = {pp45[53],pp35[64],pp1[99],pp1[100]};
    CLA_4 KS_88(s88, c88, in88_1, in88_2);
    wire[3:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp46[52],pp36[63],pp2[98],pp2[99]};
    assign in89_2 = {pp47[51],pp37[62],pp3[97],pp3[98]};
    CLA_4 KS_89(s89, c89, in89_1, in89_2);
    wire[3:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp48[50],pp38[61],pp4[96],pp4[97]};
    assign in90_2 = {pp49[49],pp39[60],pp5[95],pp5[96]};
    CLA_4 KS_90(s90, c90, in90_1, in90_2);
    wire[3:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp50[48],pp40[59],pp6[94],pp6[95]};
    assign in91_2 = {pp51[47],pp41[58],pp7[93],pp7[94]};
    CLA_4 KS_91(s91, c91, in91_1, in91_2);
    wire[3:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp53[45],pp42[57],pp8[92],pp8[93]};
    assign in92_2 = {pp54[44],pp43[56],pp9[91],pp9[92]};
    CLA_4_c KS_92(s92, c92, in92_1, in92_2, pp52[46]);
    wire[3:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp44[55],pp10[90],pp10[91],pp0[102]};
    assign in93_2 = {pp45[54],pp11[89],pp11[90],pp1[101]};
    CLA_4 KS_93(s93, c93, in93_1, in93_2);
    wire[3:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp46[53],pp12[88],pp12[89],pp2[100]};
    assign in94_2 = {pp47[52],pp13[87],pp13[88],pp3[99]};
    CLA_4 KS_94(s94, c94, in94_1, in94_2);
    wire[3:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp48[51],pp14[86],pp14[87],pp4[98]};
    assign in95_2 = {pp49[50],pp15[85],pp15[86],pp5[97]};
    CLA_4 KS_95(s95, c95, in95_1, in95_2);
    wire[3:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp50[49],pp16[84],pp16[85],pp6[96]};
    assign in96_2 = {pp51[48],pp17[83],pp17[84],pp7[95]};
    CLA_4 KS_96(s96, c96, in96_1, in96_2);
    wire[3:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp52[47],pp18[82],pp18[83],pp8[94]};
    assign in97_2 = {pp53[46],pp19[81],pp19[82],pp9[93]};
    CLA_4 KS_97(s97, c97, in97_1, in97_2);
    wire[3:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp55[44],pp20[80],pp20[81],pp10[92]};
    assign in98_2 = {pp56[43],pp21[79],pp21[80],pp11[91]};
    CLA_4_c KS_98(s98, c98, in98_1, in98_2, pp54[45]);
    wire[3:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp22[78],pp22[79],pp12[90],pp0[103]};
    assign in99_2 = {pp23[77],pp23[78],pp13[89],pp1[102]};
    CLA_4 KS_99(s99, c99, in99_1, in99_2);
    wire[3:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp24[76],pp24[77],pp14[88],pp2[101]};
    assign in100_2 = {pp25[75],pp25[76],pp15[87],pp3[100]};
    CLA_4 KS_100(s100, c100, in100_1, in100_2);
    wire[3:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp26[74],pp26[75],pp16[86],pp4[99]};
    assign in101_2 = {pp27[73],pp27[74],pp17[85],pp5[98]};
    CLA_4 KS_101(s101, c101, in101_1, in101_2);
    wire[3:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp28[72],pp28[73],pp18[84],pp6[97]};
    assign in102_2 = {pp29[71],pp29[72],pp19[83],pp7[96]};
    CLA_4 KS_102(s102, c102, in102_1, in102_2);
    wire[3:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp30[70],pp30[71],pp20[82],pp8[95]};
    assign in103_2 = {pp31[69],pp31[70],pp21[81],pp9[94]};
    CLA_4 KS_103(s103, c103, in103_1, in103_2);
    wire[3:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp32[68],pp32[69],pp22[80],pp10[93]};
    assign in104_2 = {pp33[67],pp33[68],pp23[79],pp11[92]};
    CLA_4 KS_104(s104, c104, in104_1, in104_2);
    wire[3:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp34[66],pp34[67],pp24[78],pp12[91]};
    assign in105_2 = {pp35[65],pp35[66],pp25[77],pp13[90]};
    CLA_4 KS_105(s105, c105, in105_1, in105_2);
    wire[3:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp36[64],pp36[65],pp26[76],pp14[89]};
    assign in106_2 = {pp37[63],pp37[64],pp27[75],pp15[88]};
    CLA_4 KS_106(s106, c106, in106_1, in106_2);
    wire[3:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp38[62],pp38[63],pp28[74],pp16[87]};
    assign in107_2 = {pp39[61],pp39[62],pp29[73],pp17[86]};
    CLA_4 KS_107(s107, c107, in107_1, in107_2);
    wire[3:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp40[60],pp40[61],pp30[72],pp18[85]};
    assign in108_2 = {pp41[59],pp41[60],pp31[71],pp19[84]};
    CLA_4 KS_108(s108, c108, in108_1, in108_2);
    wire[3:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp42[58],pp42[59],pp32[70],pp20[83]};
    assign in109_2 = {pp43[57],pp43[58],pp33[69],pp21[82]};
    CLA_4 KS_109(s109, c109, in109_1, in109_2);
    wire[3:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp44[56],pp44[57],pp34[68],pp22[81]};
    assign in110_2 = {pp45[55],pp45[56],pp35[67],pp23[80]};
    CLA_4 KS_110(s110, c110, in110_1, in110_2);
    wire[3:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp46[54],pp46[55],pp36[66],pp24[79]};
    assign in111_2 = {pp47[53],pp47[54],pp37[65],pp25[78]};
    CLA_4 KS_111(s111, c111, in111_1, in111_2);
    wire[3:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp48[52],pp48[53],pp38[64],pp26[77]};
    assign in112_2 = {pp49[51],pp49[52],pp39[63],pp27[76]};
    CLA_4 KS_112(s112, c112, in112_1, in112_2);
    wire[3:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp50[50],pp50[51],pp40[62],pp28[75]};
    assign in113_2 = {pp51[49],pp51[50],pp41[61],pp29[74]};
    CLA_4 KS_113(s113, c113, in113_1, in113_2);
    wire[3:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp52[48],pp52[49],pp42[60],pp30[73]};
    assign in114_2 = {pp53[47],pp53[48],pp43[59],pp31[72]};
    CLA_4 KS_114(s114, c114, in114_1, in114_2);
    wire[0:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp54[46]};
    assign in115_2 = {pp55[45]};
    Half_Adder KS_115(s115, c115, in115_1, in115_2);
    wire[3:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp56[44],pp54[47],pp44[58],pp32[71]};
    assign in116_2 = {pp57[43],pp55[46],pp45[57],pp33[70]};
    CLA_4 KS_116(s116, c116, in116_1, in116_2);
    wire[0:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {pp58[42]};
    assign in117_2 = {pp59[41]};
    Half_Adder KS_117(s117, c117, in117_1, in117_2);
    wire[3:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {pp60[40],pp56[45],pp46[56],pp34[69]};
    assign in118_2 = {pp61[39],pp57[44],pp47[55],pp35[68]};
    CLA_4 KS_118(s118, c118, in118_1, in118_2);
    wire[0:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {pp62[38]};
    assign in119_2 = {pp63[37]};
    Half_Adder KS_119(s119, c119, in119_1, in119_2);
    wire[3:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {pp64[36],pp58[43],pp48[54],pp36[67]};
    assign in120_2 = {pp65[35],pp59[42],pp49[53],pp37[66]};
    CLA_4 KS_120(s120, c120, in120_1, in120_2);
    wire[0:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp66[34]};
    assign in121_2 = {pp67[33]};
    Half_Adder KS_121(s121, c121, in121_1, in121_2);
    wire[3:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp68[32],pp60[41],pp50[52],pp38[65]};
    assign in122_2 = {pp69[31],pp61[40],pp51[51],pp39[64]};
    CLA_4 KS_122(s122, c122, in122_1, in122_2);
    wire[0:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp70[30]};
    assign in123_2 = {pp71[29]};
    Half_Adder KS_123(s123, c123, in123_1, in123_2);
    wire[3:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp72[28],pp62[39],pp52[50],pp40[63]};
    assign in124_2 = {pp73[27],pp63[38],pp53[49],pp41[62]};
    CLA_4 KS_124(s124, c124, in124_1, in124_2);
    wire[0:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp74[26]};
    assign in125_2 = {pp75[25]};
    Half_Adder KS_125(s125, c125, in125_1, in125_2);
    wire[3:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp76[24],pp64[37],pp54[48],pp42[61]};
    assign in126_2 = {pp77[23],pp65[36],pp55[47],pp43[60]};
    CLA_4 KS_126(s126, c126, in126_1, in126_2);
    wire[0:0] s127, in127_1, in127_2;
    wire c127;
    assign in127_1 = {pp78[22]};
    assign in127_2 = {pp79[21]};
    Half_Adder KS_127(s127, c127, in127_1, in127_2);
    wire[3:0] s128, in128_1, in128_2;
    wire c128;
    assign in128_1 = {pp81[19],pp66[35],pp56[46],pp44[59]};
    assign in128_2 = {pp82[18],pp67[34],pp57[45],pp45[58]};
    CLA_4_c KS_128(s128, c128, in128_1, in128_2, pp80[20]);
    wire[3:0] s129, in129_1, in129_2;
    wire c129;
    assign in129_1 = {pp58[44],pp46[57],pp0[104],pp0[105]};
    assign in129_2 = {pp59[43],pp47[56],pp1[103],pp1[104]};
    CLA_4 KS_129(s129, c129, in129_1, in129_2);
    wire[3:0] s130, in130_1, in130_2;
    wire c130;
    assign in130_1 = {pp61[41],pp48[55],pp2[102],pp2[103]};
    assign in130_2 = {pp62[40],pp49[54],pp3[101],pp3[102]};
    CLA_4_c KS_130(s130, c130, in130_1, in130_2, pp60[42]);
    wire[3:0] s131, in131_1, in131_2;
    wire c131;
    assign in131_1 = {pp50[53],pp4[100],pp4[101],pp0[106]};
    assign in131_2 = {pp51[52],pp5[99],pp5[100],pp1[105]};
    CLA_4 KS_131(s131, c131, in131_1, in131_2);
    wire[3:0] s132, in132_1, in132_2;
    wire c132;
    assign in132_1 = {pp52[51],pp6[98],pp6[99],pp2[104]};
    assign in132_2 = {pp53[50],pp7[97],pp7[98],pp3[103]};
    CLA_4 KS_132(s132, c132, in132_1, in132_2);
    wire[3:0] s133, in133_1, in133_2;
    wire c133;
    assign in133_1 = {pp54[49],pp8[96],pp8[97],pp4[102]};
    assign in133_2 = {pp55[48],pp9[95],pp9[96],pp5[101]};
    CLA_4 KS_133(s133, c133, in133_1, in133_2);
    wire[3:0] s134, in134_1, in134_2;
    wire c134;
    assign in134_1 = {pp56[47],pp10[94],pp10[95],pp6[100]};
    assign in134_2 = {pp57[46],pp11[93],pp11[94],pp7[99]};
    CLA_4 KS_134(s134, c134, in134_1, in134_2);
    wire[3:0] s135, in135_1, in135_2;
    wire c135;
    assign in135_1 = {pp58[45],pp12[92],pp12[93],pp8[98]};
    assign in135_2 = {pp59[44],pp13[91],pp13[92],pp9[97]};
    CLA_4 KS_135(s135, c135, in135_1, in135_2);
    wire[3:0] s136, in136_1, in136_2;
    wire c136;
    assign in136_1 = {pp60[43],pp14[90],pp14[91],pp10[96]};
    assign in136_2 = {pp61[42],pp15[89],pp15[90],pp11[95]};
    CLA_4 KS_136(s136, c136, in136_1, in136_2);
    wire[3:0] s137, in137_1, in137_2;
    wire c137;
    assign in137_1 = {pp62[41],pp16[88],pp16[89],pp12[94]};
    assign in137_2 = {pp63[40],pp17[87],pp17[88],pp13[93]};
    CLA_4 KS_137(s137, c137, in137_1, in137_2);
    wire[3:0] s138, in138_1, in138_2;
    wire c138;
    assign in138_1 = {pp65[38],pp18[86],pp18[87],pp14[92]};
    assign in138_2 = {pp66[37],pp19[85],pp19[86],pp15[91]};
    CLA_4_c KS_138(s138, c138, in138_1, in138_2, pp64[39]);
    wire[3:0] s139, in139_1, in139_2;
    wire c139;
    assign in139_1 = {pp20[84],pp20[85],pp16[90],pp0[107]};
    assign in139_2 = {pp21[83],pp21[84],pp17[89],pp1[106]};
    CLA_4 KS_139(s139, c139, in139_1, in139_2);
    wire[3:0] s140, in140_1, in140_2;
    wire c140;
    assign in140_1 = {pp22[82],pp22[83],pp18[88],pp2[105]};
    assign in140_2 = {pp23[81],pp23[82],pp19[87],pp3[104]};
    CLA_4 KS_140(s140, c140, in140_1, in140_2);
    wire[3:0] s141, in141_1, in141_2;
    wire c141;
    assign in141_1 = {pp24[80],pp24[81],pp20[86],pp4[103]};
    assign in141_2 = {pp25[79],pp25[80],pp21[85],pp5[102]};
    CLA_4 KS_141(s141, c141, in141_1, in141_2);
    wire[3:0] s142, in142_1, in142_2;
    wire c142;
    assign in142_1 = {pp26[78],pp26[79],pp22[84],pp6[101]};
    assign in142_2 = {pp27[77],pp27[78],pp23[83],pp7[100]};
    CLA_4 KS_142(s142, c142, in142_1, in142_2);
    wire[3:0] s143, in143_1, in143_2;
    wire c143;
    assign in143_1 = {pp28[76],pp28[77],pp24[82],pp8[99]};
    assign in143_2 = {pp29[75],pp29[76],pp25[81],pp9[98]};
    CLA_4 KS_143(s143, c143, in143_1, in143_2);
    wire[3:0] s144, in144_1, in144_2;
    wire c144;
    assign in144_1 = {pp30[74],pp30[75],pp26[80],pp10[97]};
    assign in144_2 = {pp31[73],pp31[74],pp27[79],pp11[96]};
    CLA_4 KS_144(s144, c144, in144_1, in144_2);
    wire[3:0] s145, in145_1, in145_2;
    wire c145;
    assign in145_1 = {pp32[72],pp32[73],pp28[78],pp12[95]};
    assign in145_2 = {pp33[71],pp33[72],pp29[77],pp13[94]};
    CLA_4 KS_145(s145, c145, in145_1, in145_2);
    wire[3:0] s146, in146_1, in146_2;
    wire c146;
    assign in146_1 = {pp34[70],pp34[71],pp30[76],pp14[93]};
    assign in146_2 = {pp35[69],pp35[70],pp31[75],pp15[92]};
    CLA_4 KS_146(s146, c146, in146_1, in146_2);
    wire[3:0] s147, in147_1, in147_2;
    wire c147;
    assign in147_1 = {pp36[68],pp36[69],pp32[74],pp16[91]};
    assign in147_2 = {pp37[67],pp37[68],pp33[73],pp17[90]};
    CLA_4 KS_147(s147, c147, in147_1, in147_2);
    wire[3:0] s148, in148_1, in148_2;
    wire c148;
    assign in148_1 = {pp38[66],pp38[67],pp34[72],pp18[89]};
    assign in148_2 = {pp39[65],pp39[66],pp35[71],pp19[88]};
    CLA_4 KS_148(s148, c148, in148_1, in148_2);
    wire[3:0] s149, in149_1, in149_2;
    wire c149;
    assign in149_1 = {pp40[64],pp40[65],pp36[70],pp20[87]};
    assign in149_2 = {pp41[63],pp41[64],pp37[69],pp21[86]};
    CLA_4 KS_149(s149, c149, in149_1, in149_2);
    wire[3:0] s150, in150_1, in150_2;
    wire c150;
    assign in150_1 = {pp42[62],pp42[63],pp38[68],pp22[85]};
    assign in150_2 = {pp43[61],pp43[62],pp39[67],pp23[84]};
    CLA_4 KS_150(s150, c150, in150_1, in150_2);
    wire[3:0] s151, in151_1, in151_2;
    wire c151;
    assign in151_1 = {pp44[60],pp44[61],pp40[66],pp24[83]};
    assign in151_2 = {pp45[59],pp45[60],pp41[65],pp25[82]};
    CLA_4 KS_151(s151, c151, in151_1, in151_2);
    wire[3:0] s152, in152_1, in152_2;
    wire c152;
    assign in152_1 = {pp46[58],pp46[59],pp42[64],pp26[81]};
    assign in152_2 = {pp47[57],pp47[58],pp43[63],pp27[80]};
    CLA_4 KS_152(s152, c152, in152_1, in152_2);
    wire[3:0] s153, in153_1, in153_2;
    wire c153;
    assign in153_1 = {pp48[56],pp48[57],pp44[62],pp28[79]};
    assign in153_2 = {pp49[55],pp49[56],pp45[61],pp29[78]};
    CLA_4 KS_153(s153, c153, in153_1, in153_2);
    wire[3:0] s154, in154_1, in154_2;
    wire c154;
    assign in154_1 = {pp50[54],pp50[55],pp46[60],pp30[77]};
    assign in154_2 = {pp51[53],pp51[54],pp47[59],pp31[76]};
    CLA_4 KS_154(s154, c154, in154_1, in154_2);
    wire[3:0] s155, in155_1, in155_2;
    wire c155;
    assign in155_1 = {pp52[52],pp52[53],pp48[58],pp32[75]};
    assign in155_2 = {pp53[51],pp53[52],pp49[57],pp33[74]};
    CLA_4 KS_155(s155, c155, in155_1, in155_2);
    wire[3:0] s156, in156_1, in156_2;
    wire c156;
    assign in156_1 = {pp54[50],pp54[51],pp50[56],pp34[73]};
    assign in156_2 = {pp55[49],pp55[50],pp51[55],pp35[72]};
    CLA_4 KS_156(s156, c156, in156_1, in156_2);
    wire[3:0] s157, in157_1, in157_2;
    wire c157;
    assign in157_1 = {pp56[48],pp56[49],pp52[54],pp36[71]};
    assign in157_2 = {pp57[47],pp57[48],pp53[53],pp37[70]};
    CLA_4 KS_157(s157, c157, in157_1, in157_2);
    wire[3:0] s158, in158_1, in158_2;
    wire c158;
    assign in158_1 = {pp58[46],pp58[47],pp54[52],pp38[69]};
    assign in158_2 = {pp59[45],pp59[46],pp55[51],pp39[68]};
    CLA_4 KS_158(s158, c158, in158_1, in158_2);
    wire[3:0] s159, in159_1, in159_2;
    wire c159;
    assign in159_1 = {pp60[44],pp60[45],pp56[50],pp40[67]};
    assign in159_2 = {pp61[43],pp61[44],pp57[49],pp41[66]};
    CLA_4 KS_159(s159, c159, in159_1, in159_2);
    wire[0:0] s160, in160_1, in160_2;
    wire c160;
    assign in160_1 = {pp62[42]};
    assign in160_2 = {pp63[41]};
    Half_Adder KS_160(s160, c160, in160_1, in160_2);
    wire[3:0] s161, in161_1, in161_2;
    wire c161;
    assign in161_1 = {pp64[40],pp62[43],pp58[48],pp42[65]};
    assign in161_2 = {pp65[39],pp63[42],pp59[47],pp43[64]};
    CLA_4 KS_161(s161, c161, in161_1, in161_2);
    wire[0:0] s162, in162_1, in162_2;
    wire c162;
    assign in162_1 = {pp66[38]};
    assign in162_2 = {pp67[37]};
    Half_Adder KS_162(s162, c162, in162_1, in162_2);
    wire[3:0] s163, in163_1, in163_2;
    wire c163;
    assign in163_1 = {pp68[36],pp64[41],pp60[46],pp44[63]};
    assign in163_2 = {pp69[35],pp65[40],pp61[45],pp45[62]};
    CLA_4 KS_163(s163, c163, in163_1, in163_2);
    wire[0:0] s164, in164_1, in164_2;
    wire c164;
    assign in164_1 = {pp70[34]};
    assign in164_2 = {pp71[33]};
    Half_Adder KS_164(s164, c164, in164_1, in164_2);
    wire[3:0] s165, in165_1, in165_2;
    wire c165;
    assign in165_1 = {pp72[32],pp66[39],pp62[44],pp46[61]};
    assign in165_2 = {pp73[31],pp67[38],pp63[43],pp47[60]};
    CLA_4 KS_165(s165, c165, in165_1, in165_2);
    wire[0:0] s166, in166_1, in166_2;
    wire c166;
    assign in166_1 = {pp74[30]};
    assign in166_2 = {pp75[29]};
    Half_Adder KS_166(s166, c166, in166_1, in166_2);
    wire[3:0] s167, in167_1, in167_2;
    wire c167;
    assign in167_1 = {pp76[28],pp68[37],pp64[42],pp48[59]};
    assign in167_2 = {pp77[27],pp69[36],pp65[41],pp49[58]};
    CLA_4 KS_167(s167, c167, in167_1, in167_2);
    wire[0:0] s168, in168_1, in168_2;
    wire c168;
    assign in168_1 = {pp78[26]};
    assign in168_2 = {pp79[25]};
    Half_Adder KS_168(s168, c168, in168_1, in168_2);
    wire[3:0] s169, in169_1, in169_2;
    wire c169;
    assign in169_1 = {pp80[24],pp70[35],pp66[40],pp50[57]};
    assign in169_2 = {pp81[23],pp71[34],pp67[39],pp51[56]};
    CLA_4 KS_169(s169, c169, in169_1, in169_2);
    wire[0:0] s170, in170_1, in170_2;
    wire c170;
    assign in170_1 = {pp82[22]};
    assign in170_2 = {pp83[21]};
    Half_Adder KS_170(s170, c170, in170_1, in170_2);
    wire[1:0] s171, in171_1, in171_2;
    wire c171;
    assign in171_1 = {pp84[20],pp72[33]};
    assign in171_2 = {pp85[19],pp73[32]};
    CLA_2 KS_171(s171, c171, in171_1, in171_2);
    wire[0:0] s172, in172_1, in172_2;
    wire c172;
    assign in172_1 = {pp86[18]};
    assign in172_2 = {pp87[17]};
    Half_Adder KS_172(s172, c172, in172_1, in172_2);
    wire[3:0] s173, in173_1, in173_2;
    wire c173;
    assign in173_1 = {pp88[16],pp74[31],pp68[38],pp52[55]};
    assign in173_2 = {pp89[15],pp75[30],pp69[37],pp53[54]};
    CLA_4 KS_173(s173, c173, in173_1, in173_2);
    wire[0:0] s174, in174_1, in174_2;
    wire c174;
    assign in174_1 = {pp90[14]};
    assign in174_2 = {pp91[13]};
    Half_Adder KS_174(s174, c174, in174_1, in174_2);
    wire[1:0] s175, in175_1, in175_2;
    wire c175;
    assign in175_1 = {pp92[12],pp76[29]};
    assign in175_2 = {pp93[11],pp77[28]};
    CLA_2 KS_175(s175, c175, in175_1, in175_2);
    wire[0:0] s176, in176_1, in176_2;
    wire c176;
    assign in176_1 = {pp94[10]};
    assign in176_2 = {pp95[9]};
    Half_Adder KS_176(s176, c176, in176_1, in176_2);
    wire[3:0] s177, in177_1, in177_2;
    wire c177;
    assign in177_1 = {pp96[8],pp78[27],pp70[36],pp54[53]};
    assign in177_2 = {pp97[7],pp79[26],pp71[35],pp55[52]};
    CLA_4 KS_177(s177, c177, in177_1, in177_2);
    wire[0:0] s178, in178_1, in178_2;
    wire c178;
    assign in178_1 = {pp98[6]};
    assign in178_2 = {pp99[5]};
    Half_Adder KS_178(s178, c178, in178_1, in178_2);
    wire[1:0] s179, in179_1, in179_2;
    wire c179;
    assign in179_1 = {pp101[3],pp80[25]};
    assign in179_2 = {pp102[2],pp81[24]};
    CLA_2_c KS_179(s179, c179, in179_1, in179_2, pp100[4]);
    wire[3:0] s180, in180_1, in180_2;
    wire c180;
    assign in180_1 = {pp56[51],pp0[108],pp0[109],pp0[110]};
    assign in180_2 = {pp57[50],pp1[107],pp1[108],pp1[109]};
    CLA_4 KS_180(s180, c180, in180_1, in180_2);
    wire[3:0] s181, in181_1, in181_2;
    wire c181;
    assign in181_1 = {pp58[49],pp2[106],pp2[107],pp2[108]};
    assign in181_2 = {pp59[48],pp3[105],pp3[106],pp3[107]};
    CLA_4 KS_181(s181, c181, in181_1, in181_2);
    wire[3:0] s182, in182_1, in182_2;
    wire c182;
    assign in182_1 = {pp60[47],pp4[104],pp4[105],pp4[106]};
    assign in182_2 = {pp61[46],pp5[103],pp5[104],pp5[105]};
    CLA_4 KS_182(s182, c182, in182_1, in182_2);
    wire[3:0] s183, in183_1, in183_2;
    wire c183;
    assign in183_1 = {pp62[45],pp6[102],pp6[103],pp6[104]};
    assign in183_2 = {pp63[44],pp7[101],pp7[102],pp7[103]};
    CLA_4 KS_183(s183, c183, in183_1, in183_2);
    wire[3:0] s184, in184_1, in184_2;
    wire c184;
    assign in184_1 = {pp64[43],pp8[100],pp8[101],pp8[102]};
    assign in184_2 = {pp65[42],pp9[99],pp9[100],pp9[101]};
    CLA_4 KS_184(s184, c184, in184_1, in184_2);
    wire[3:0] s185, in185_1, in185_2;
    wire c185;
    assign in185_1 = {pp66[41],pp10[98],pp10[99],pp10[100]};
    assign in185_2 = {pp67[40],pp11[97],pp11[98],pp11[99]};
    CLA_4 KS_185(s185, c185, in185_1, in185_2);
    wire[3:0] s186, in186_1, in186_2;
    wire c186;
    assign in186_1 = {pp68[39],pp12[96],pp12[97],pp12[98]};
    assign in186_2 = {pp69[38],pp13[95],pp13[96],pp13[97]};
    CLA_4 KS_186(s186, c186, in186_1, in186_2);
    wire[3:0] s187, in187_1, in187_2;
    wire c187;
    assign in187_1 = {pp70[37],pp14[94],pp14[95],pp14[96]};
    assign in187_2 = {pp71[36],pp15[93],pp15[94],pp15[95]};
    CLA_4 KS_187(s187, c187, in187_1, in187_2);
    wire[3:0] s188, in188_1, in188_2;
    wire c188;
    assign in188_1 = {pp72[35],pp16[92],pp16[93],pp16[94]};
    assign in188_2 = {pp73[34],pp17[91],pp17[92],pp17[93]};
    CLA_4 KS_188(s188, c188, in188_1, in188_2);
    wire[3:0] s189, in189_1, in189_2;
    wire c189;
    assign in189_1 = {pp74[33],pp18[90],pp18[91],pp18[92]};
    assign in189_2 = {pp75[32],pp19[89],pp19[90],pp19[91]};
    CLA_4 KS_189(s189, c189, in189_1, in189_2);
    wire[3:0] s190, in190_1, in190_2;
    wire c190;
    assign in190_1 = {pp77[30],pp20[88],pp20[89],pp20[90]};
    assign in190_2 = {pp78[29],pp21[87],pp21[88],pp21[89]};
    CLA_4_c KS_190(s190, c190, in190_1, in190_2, pp76[31]);
    wire[3:0] s191, in191_1, in191_2;
    wire c191;
    assign in191_1 = {pp22[86],pp22[87],pp22[88],pp0[111]};
    assign in191_2 = {pp23[85],pp23[86],pp23[87],pp1[110]};
    CLA_4 KS_191(s191, c191, in191_1, in191_2);
    wire[3:0] s192, in192_1, in192_2;
    wire c192;
    assign in192_1 = {pp24[84],pp24[85],pp24[86],pp2[109]};
    assign in192_2 = {pp25[83],pp25[84],pp25[85],pp3[108]};
    CLA_4 KS_192(s192, c192, in192_1, in192_2);
    wire[3:0] s193, in193_1, in193_2;
    wire c193;
    assign in193_1 = {pp26[82],pp26[83],pp26[84],pp4[107]};
    assign in193_2 = {pp27[81],pp27[82],pp27[83],pp5[106]};
    CLA_4 KS_193(s193, c193, in193_1, in193_2);
    wire[3:0] s194, in194_1, in194_2;
    wire c194;
    assign in194_1 = {pp28[80],pp28[81],pp28[82],pp6[105]};
    assign in194_2 = {pp29[79],pp29[80],pp29[81],pp7[104]};
    CLA_4 KS_194(s194, c194, in194_1, in194_2);
    wire[3:0] s195, in195_1, in195_2;
    wire c195;
    assign in195_1 = {pp30[78],pp30[79],pp30[80],pp8[103]};
    assign in195_2 = {pp31[77],pp31[78],pp31[79],pp9[102]};
    CLA_4 KS_195(s195, c195, in195_1, in195_2);
    wire[3:0] s196, in196_1, in196_2;
    wire c196;
    assign in196_1 = {pp32[76],pp32[77],pp32[78],pp10[101]};
    assign in196_2 = {pp33[75],pp33[76],pp33[77],pp11[100]};
    CLA_4 KS_196(s196, c196, in196_1, in196_2);
    wire[3:0] s197, in197_1, in197_2;
    wire c197;
    assign in197_1 = {pp34[74],pp34[75],pp34[76],pp12[99]};
    assign in197_2 = {pp35[73],pp35[74],pp35[75],pp13[98]};
    CLA_4 KS_197(s197, c197, in197_1, in197_2);
    wire[3:0] s198, in198_1, in198_2;
    wire c198;
    assign in198_1 = {pp36[72],pp36[73],pp36[74],pp14[97]};
    assign in198_2 = {pp37[71],pp37[72],pp37[73],pp15[96]};
    CLA_4 KS_198(s198, c198, in198_1, in198_2);
    wire[3:0] s199, in199_1, in199_2;
    wire c199;
    assign in199_1 = {pp38[70],pp38[71],pp38[72],pp16[95]};
    assign in199_2 = {pp39[69],pp39[70],pp39[71],pp17[94]};
    CLA_4 KS_199(s199, c199, in199_1, in199_2);
    wire[3:0] s200, in200_1, in200_2;
    wire c200;
    assign in200_1 = {pp40[68],pp40[69],pp40[70],pp18[93]};
    assign in200_2 = {pp41[67],pp41[68],pp41[69],pp19[92]};
    CLA_4 KS_200(s200, c200, in200_1, in200_2);
    wire[3:0] s201, in201_1, in201_2;
    wire c201;
    assign in201_1 = {pp42[66],pp42[67],pp42[68],pp20[91]};
    assign in201_2 = {pp43[65],pp43[66],pp43[67],pp21[90]};
    CLA_4 KS_201(s201, c201, in201_1, in201_2);
    wire[3:0] s202, in202_1, in202_2;
    wire c202;
    assign in202_1 = {pp44[64],pp44[65],pp44[66],pp22[89]};
    assign in202_2 = {pp45[63],pp45[64],pp45[65],pp23[88]};
    CLA_4 KS_202(s202, c202, in202_1, in202_2);
    wire[3:0] s203, in203_1, in203_2;
    wire c203;
    assign in203_1 = {pp46[62],pp46[63],pp46[64],pp24[87]};
    assign in203_2 = {pp47[61],pp47[62],pp47[63],pp25[86]};
    CLA_4 KS_203(s203, c203, in203_1, in203_2);
    wire[3:0] s204, in204_1, in204_2;
    wire c204;
    assign in204_1 = {pp48[60],pp48[61],pp48[62],pp26[85]};
    assign in204_2 = {pp49[59],pp49[60],pp49[61],pp27[84]};
    CLA_4 KS_204(s204, c204, in204_1, in204_2);
    wire[3:0] s205, in205_1, in205_2;
    wire c205;
    assign in205_1 = {pp50[58],pp50[59],pp50[60],pp28[83]};
    assign in205_2 = {pp51[57],pp51[58],pp51[59],pp29[82]};
    CLA_4 KS_205(s205, c205, in205_1, in205_2);
    wire[3:0] s206, in206_1, in206_2;
    wire c206;
    assign in206_1 = {pp52[56],pp52[57],pp52[58],pp30[81]};
    assign in206_2 = {pp53[55],pp53[56],pp53[57],pp31[80]};
    CLA_4 KS_206(s206, c206, in206_1, in206_2);
    wire[3:0] s207, in207_1, in207_2;
    wire c207;
    assign in207_1 = {pp54[54],pp54[55],pp54[56],pp32[79]};
    assign in207_2 = {pp55[53],pp55[54],pp55[55],pp33[78]};
    CLA_4 KS_207(s207, c207, in207_1, in207_2);
    wire[3:0] s208, in208_1, in208_2;
    wire c208;
    assign in208_1 = {pp56[52],pp56[53],pp56[54],pp34[77]};
    assign in208_2 = {pp57[51],pp57[52],pp57[53],pp35[76]};
    CLA_4 KS_208(s208, c208, in208_1, in208_2);
    wire[3:0] s209, in209_1, in209_2;
    wire c209;
    assign in209_1 = {pp58[50],pp58[51],pp58[52],pp36[75]};
    assign in209_2 = {pp59[49],pp59[50],pp59[51],pp37[74]};
    CLA_4 KS_209(s209, c209, in209_1, in209_2);
    wire[3:0] s210, in210_1, in210_2;
    wire c210;
    assign in210_1 = {pp60[48],pp60[49],pp60[50],pp38[73]};
    assign in210_2 = {pp61[47],pp61[48],pp61[49],pp39[72]};
    CLA_4 KS_210(s210, c210, in210_1, in210_2);
    wire[3:0] s211, in211_1, in211_2;
    wire c211;
    assign in211_1 = {pp62[46],pp62[47],pp62[48],pp40[71]};
    assign in211_2 = {pp63[45],pp63[46],pp63[47],pp41[70]};
    CLA_4 KS_211(s211, c211, in211_1, in211_2);
    wire[3:0] s212, in212_1, in212_2;
    wire c212;
    assign in212_1 = {pp64[44],pp64[45],pp64[46],pp42[69]};
    assign in212_2 = {pp65[43],pp65[44],pp65[45],pp43[68]};
    CLA_4 KS_212(s212, c212, in212_1, in212_2);
    wire[3:0] s213, in213_1, in213_2;
    wire c213;
    assign in213_1 = {pp66[42],pp66[43],pp66[44],pp44[67]};
    assign in213_2 = {pp67[41],pp67[42],pp67[43],pp45[66]};
    CLA_4 KS_213(s213, c213, in213_1, in213_2);
    wire[3:0] s214, in214_1, in214_2;
    wire c214;
    assign in214_1 = {pp68[40],pp68[41],pp68[42],pp46[65]};
    assign in214_2 = {pp69[39],pp69[40],pp69[41],pp47[64]};
    CLA_4 KS_214(s214, c214, in214_1, in214_2);
    wire[0:0] s215, in215_1, in215_2;
    wire c215;
    assign in215_1 = {pp70[38]};
    assign in215_2 = {pp71[37]};
    Half_Adder KS_215(s215, c215, in215_1, in215_2);
    wire[3:0] s216, in216_1, in216_2;
    wire c216;
    assign in216_1 = {pp72[36],pp70[39],pp70[40],pp48[63]};
    assign in216_2 = {pp73[35],pp71[38],pp71[39],pp49[62]};
    CLA_4 KS_216(s216, c216, in216_1, in216_2);
    wire[0:0] s217, in217_1, in217_2;
    wire c217;
    assign in217_1 = {pp74[34]};
    assign in217_2 = {pp75[33]};
    Half_Adder KS_217(s217, c217, in217_1, in217_2);
    wire[1:0] s218, in218_1, in218_2;
    wire c218;
    assign in218_1 = {pp76[32],pp72[37]};
    assign in218_2 = {pp77[31],pp73[36]};
    CLA_2 KS_218(s218, c218, in218_1, in218_2);
    wire[0:0] s219, in219_1, in219_2;
    wire c219;
    assign in219_1 = {pp78[30]};
    assign in219_2 = {pp79[29]};
    Half_Adder KS_219(s219, c219, in219_1, in219_2);
    wire[3:0] s220, in220_1, in220_2;
    wire c220;
    assign in220_1 = {pp80[28],pp74[35],pp72[38],pp50[61]};
    assign in220_2 = {pp81[27],pp75[34],pp73[37],pp51[60]};
    CLA_4 KS_220(s220, c220, in220_1, in220_2);
    wire[0:0] s221, in221_1, in221_2;
    wire c221;
    assign in221_1 = {pp82[26]};
    assign in221_2 = {pp83[25]};
    Half_Adder KS_221(s221, c221, in221_1, in221_2);
    wire[1:0] s222, in222_1, in222_2;
    wire c222;
    assign in222_1 = {pp84[24],pp76[33]};
    assign in222_2 = {pp85[23],pp77[32]};
    CLA_2 KS_222(s222, c222, in222_1, in222_2);
    wire[0:0] s223, in223_1, in223_2;
    wire c223;
    assign in223_1 = {pp86[22]};
    assign in223_2 = {pp87[21]};
    Half_Adder KS_223(s223, c223, in223_1, in223_2);
    wire[3:0] s224, in224_1, in224_2;
    wire c224;
    assign in224_1 = {pp88[20],pp78[31],pp74[36],pp52[59]};
    assign in224_2 = {pp89[19],pp79[30],pp75[35],pp53[58]};
    CLA_4 KS_224(s224, c224, in224_1, in224_2);
    wire[0:0] s225, in225_1, in225_2;
    wire c225;
    assign in225_1 = {pp90[18]};
    assign in225_2 = {pp91[17]};
    Half_Adder KS_225(s225, c225, in225_1, in225_2);
    wire[1:0] s226, in226_1, in226_2;
    wire c226;
    assign in226_1 = {pp92[16],pp80[29]};
    assign in226_2 = {pp93[15],pp81[28]};
    CLA_2 KS_226(s226, c226, in226_1, in226_2);
    wire[0:0] s227, in227_1, in227_2;
    wire c227;
    assign in227_1 = {pp94[14]};
    assign in227_2 = {pp95[13]};
    Half_Adder KS_227(s227, c227, in227_1, in227_2);
    wire[3:0] s228, in228_1, in228_2;
    wire c228;
    assign in228_1 = {pp96[12],pp82[27],pp76[34],pp54[57]};
    assign in228_2 = {pp97[11],pp83[26],pp77[33],pp55[56]};
    CLA_4 KS_228(s228, c228, in228_1, in228_2);
    wire[0:0] s229, in229_1, in229_2;
    wire c229;
    assign in229_1 = {pp98[10]};
    assign in229_2 = {pp99[9]};
    Half_Adder KS_229(s229, c229, in229_1, in229_2);
    wire[1:0] s230, in230_1, in230_2;
    wire c230;
    assign in230_1 = {pp100[8],pp84[25]};
    assign in230_2 = {pp101[7],pp85[24]};
    CLA_2 KS_230(s230, c230, in230_1, in230_2);
    wire[0:0] s231, in231_1, in231_2;
    wire c231;
    assign in231_1 = {pp102[6]};
    assign in231_2 = {pp103[5]};
    Half_Adder KS_231(s231, c231, in231_1, in231_2);
    wire[3:0] s232, in232_1, in232_2;
    wire c232;
    assign in232_1 = {pp104[4],pp86[23],pp78[32],pp56[55]};
    assign in232_2 = {pp105[3],pp87[22],pp79[31],pp57[54]};
    CLA_4 KS_232(s232, c232, in232_1, in232_2);
    wire[0:0] s233, in233_1, in233_2;
    wire c233;
    assign in233_1 = {pp106[2]};
    assign in233_2 = {pp107[1]};
    Half_Adder KS_233(s233, c233, in233_1, in233_2);
    wire[1:0] s234, in234_1, in234_2;
    wire c234;
    assign in234_1 = {pp108[0],pp88[21]};
    assign in234_2 = {c139,pp89[20]};
    CLA_2 KS_234(s234, c234, in234_1, in234_2);
    wire[0:0] s235, in235_1, in235_2;
    wire c235;
    assign in235_1 = {c140};
    assign in235_2 = {c141};
    Half_Adder KS_235(s235, c235, in235_1, in235_2);
    wire[3:0] s236, in236_1, in236_2;
    wire c236;
    assign in236_1 = {c142,pp90[19],pp80[30],pp58[53]};
    assign in236_2 = {c143,pp91[18],pp81[29],pp59[52]};
    CLA_4 KS_236(s236, c236, in236_1, in236_2);
    wire[0:0] s237, in237_1, in237_2;
    wire c237;
    assign in237_1 = {c144};
    assign in237_2 = {c145};
    Half_Adder KS_237(s237, c237, in237_1, in237_2);
    wire[1:0] s238, in238_1, in238_2;
    wire c238;
    assign in238_1 = {c146,pp92[17]};
    assign in238_2 = {c147,pp93[16]};
    CLA_2 KS_238(s238, c238, in238_1, in238_2);
    wire[0:0] s239, in239_1, in239_2;
    wire c239;
    assign in239_1 = {c149};
    assign in239_2 = {c150};
    Full_Adder KS_239(s239, c239, in239_1, in239_2, c148);
    wire[3:0] s240, in240_1, in240_2;
    wire c240;
    assign in240_1 = {pp60[51],pp0[112],pp0[113],pp0[114]};
    assign in240_2 = {pp61[50],pp1[111],pp1[112],pp1[113]};
    CLA_4 KS_240(s240, c240, in240_1, in240_2);
    wire[3:0] s241, in241_1, in241_2;
    wire c241;
    assign in241_1 = {pp62[49],pp2[110],pp2[111],pp2[112]};
    assign in241_2 = {pp63[48],pp3[109],pp3[110],pp3[111]};
    CLA_4 KS_241(s241, c241, in241_1, in241_2);
    wire[3:0] s242, in242_1, in242_2;
    wire c242;
    assign in242_1 = {pp64[47],pp4[108],pp4[109],pp4[110]};
    assign in242_2 = {pp65[46],pp5[107],pp5[108],pp5[109]};
    CLA_4 KS_242(s242, c242, in242_1, in242_2);
    wire[3:0] s243, in243_1, in243_2;
    wire c243;
    assign in243_1 = {pp66[45],pp6[106],pp6[107],pp6[108]};
    assign in243_2 = {pp67[44],pp7[105],pp7[106],pp7[107]};
    CLA_4 KS_243(s243, c243, in243_1, in243_2);
    wire[3:0] s244, in244_1, in244_2;
    wire c244;
    assign in244_1 = {pp68[43],pp8[104],pp8[105],pp8[106]};
    assign in244_2 = {pp69[42],pp9[103],pp9[104],pp9[105]};
    CLA_4 KS_244(s244, c244, in244_1, in244_2);
    wire[3:0] s245, in245_1, in245_2;
    wire c245;
    assign in245_1 = {pp70[41],pp10[102],pp10[103],pp10[104]};
    assign in245_2 = {pp71[40],pp11[101],pp11[102],pp11[103]};
    CLA_4 KS_245(s245, c245, in245_1, in245_2);
    wire[3:0] s246, in246_1, in246_2;
    wire c246;
    assign in246_1 = {pp72[39],pp12[100],pp12[101],pp12[102]};
    assign in246_2 = {pp73[38],pp13[99],pp13[100],pp13[101]};
    CLA_4 KS_246(s246, c246, in246_1, in246_2);
    wire[3:0] s247, in247_1, in247_2;
    wire c247;
    assign in247_1 = {pp74[37],pp14[98],pp14[99],pp14[100]};
    assign in247_2 = {pp75[36],pp15[97],pp15[98],pp15[99]};
    CLA_4 KS_247(s247, c247, in247_1, in247_2);
    wire[3:0] s248, in248_1, in248_2;
    wire c248;
    assign in248_1 = {pp76[35],pp16[96],pp16[97],pp16[98]};
    assign in248_2 = {pp77[34],pp17[95],pp17[96],pp17[97]};
    CLA_4 KS_248(s248, c248, in248_1, in248_2);
    wire[3:0] s249, in249_1, in249_2;
    wire c249;
    assign in249_1 = {pp78[33],pp18[94],pp18[95],pp18[96]};
    assign in249_2 = {pp79[32],pp19[93],pp19[94],pp19[95]};
    CLA_4 KS_249(s249, c249, in249_1, in249_2);
    wire[3:0] s250, in250_1, in250_2;
    wire c250;
    assign in250_1 = {pp80[31],pp20[92],pp20[93],pp20[94]};
    assign in250_2 = {pp81[30],pp21[91],pp21[92],pp21[93]};
    CLA_4 KS_250(s250, c250, in250_1, in250_2);
    wire[3:0] s251, in251_1, in251_2;
    wire c251;
    assign in251_1 = {pp82[29],pp22[90],pp22[91],pp22[92]};
    assign in251_2 = {pp83[28],pp23[89],pp23[90],pp23[91]};
    CLA_4 KS_251(s251, c251, in251_1, in251_2);
    wire[3:0] s252, in252_1, in252_2;
    wire c252;
    assign in252_1 = {pp84[27],pp24[88],pp24[89],pp24[90]};
    assign in252_2 = {pp85[26],pp25[87],pp25[88],pp25[89]};
    CLA_4 KS_252(s252, c252, in252_1, in252_2);
    wire[3:0] s253, in253_1, in253_2;
    wire c253;
    assign in253_1 = {pp86[25],pp26[86],pp26[87],pp26[88]};
    assign in253_2 = {pp87[24],pp27[85],pp27[86],pp27[87]};
    CLA_4 KS_253(s253, c253, in253_1, in253_2);
    wire[3:0] s254, in254_1, in254_2;
    wire c254;
    assign in254_1 = {pp88[23],pp28[84],pp28[85],pp28[86]};
    assign in254_2 = {pp89[22],pp29[83],pp29[84],pp29[85]};
    CLA_4 KS_254(s254, c254, in254_1, in254_2);
    wire[3:0] s255, in255_1, in255_2;
    wire c255;
    assign in255_1 = {pp91[20],pp30[82],pp30[83],pp30[84]};
    assign in255_2 = {pp92[19],pp31[81],pp31[82],pp31[83]};
    CLA_4_c KS_255(s255, c255, in255_1, in255_2, pp90[21]);
    wire[3:0] s256, in256_1, in256_2;
    wire c256;
    assign in256_1 = {pp32[80],pp32[81],pp32[82],pp0[115]};
    assign in256_2 = {pp33[79],pp33[80],pp33[81],pp1[114]};
    CLA_4 KS_256(s256, c256, in256_1, in256_2);
    wire[3:0] s257, in257_1, in257_2;
    wire c257;
    assign in257_1 = {pp34[78],pp34[79],pp34[80],pp2[113]};
    assign in257_2 = {pp35[77],pp35[78],pp35[79],pp3[112]};
    CLA_4 KS_257(s257, c257, in257_1, in257_2);
    wire[3:0] s258, in258_1, in258_2;
    wire c258;
    assign in258_1 = {pp36[76],pp36[77],pp36[78],pp4[111]};
    assign in258_2 = {pp37[75],pp37[76],pp37[77],pp5[110]};
    CLA_4 KS_258(s258, c258, in258_1, in258_2);
    wire[3:0] s259, in259_1, in259_2;
    wire c259;
    assign in259_1 = {pp38[74],pp38[75],pp38[76],pp6[109]};
    assign in259_2 = {pp39[73],pp39[74],pp39[75],pp7[108]};
    CLA_4 KS_259(s259, c259, in259_1, in259_2);
    wire[3:0] s260, in260_1, in260_2;
    wire c260;
    assign in260_1 = {pp40[72],pp40[73],pp40[74],pp8[107]};
    assign in260_2 = {pp41[71],pp41[72],pp41[73],pp9[106]};
    CLA_4 KS_260(s260, c260, in260_1, in260_2);
    wire[3:0] s261, in261_1, in261_2;
    wire c261;
    assign in261_1 = {pp42[70],pp42[71],pp42[72],pp10[105]};
    assign in261_2 = {pp43[69],pp43[70],pp43[71],pp11[104]};
    CLA_4 KS_261(s261, c261, in261_1, in261_2);
    wire[3:0] s262, in262_1, in262_2;
    wire c262;
    assign in262_1 = {pp44[68],pp44[69],pp44[70],pp12[103]};
    assign in262_2 = {pp45[67],pp45[68],pp45[69],pp13[102]};
    CLA_4 KS_262(s262, c262, in262_1, in262_2);
    wire[3:0] s263, in263_1, in263_2;
    wire c263;
    assign in263_1 = {pp46[66],pp46[67],pp46[68],pp14[101]};
    assign in263_2 = {pp47[65],pp47[66],pp47[67],pp15[100]};
    CLA_4 KS_263(s263, c263, in263_1, in263_2);
    wire[3:0] s264, in264_1, in264_2;
    wire c264;
    assign in264_1 = {pp48[64],pp48[65],pp48[66],pp16[99]};
    assign in264_2 = {pp49[63],pp49[64],pp49[65],pp17[98]};
    CLA_4 KS_264(s264, c264, in264_1, in264_2);
    wire[3:0] s265, in265_1, in265_2;
    wire c265;
    assign in265_1 = {pp50[62],pp50[63],pp50[64],pp18[97]};
    assign in265_2 = {pp51[61],pp51[62],pp51[63],pp19[96]};
    CLA_4 KS_265(s265, c265, in265_1, in265_2);
    wire[3:0] s266, in266_1, in266_2;
    wire c266;
    assign in266_1 = {pp52[60],pp52[61],pp52[62],pp20[95]};
    assign in266_2 = {pp53[59],pp53[60],pp53[61],pp21[94]};
    CLA_4 KS_266(s266, c266, in266_1, in266_2);
    wire[3:0] s267, in267_1, in267_2;
    wire c267;
    assign in267_1 = {pp54[58],pp54[59],pp54[60],pp22[93]};
    assign in267_2 = {pp55[57],pp55[58],pp55[59],pp23[92]};
    CLA_4 KS_267(s267, c267, in267_1, in267_2);
    wire[3:0] s268, in268_1, in268_2;
    wire c268;
    assign in268_1 = {pp56[56],pp56[57],pp56[58],pp24[91]};
    assign in268_2 = {pp57[55],pp57[56],pp57[57],pp25[90]};
    CLA_4 KS_268(s268, c268, in268_1, in268_2);
    wire[3:0] s269, in269_1, in269_2;
    wire c269;
    assign in269_1 = {pp58[54],pp58[55],pp58[56],pp26[89]};
    assign in269_2 = {pp59[53],pp59[54],pp59[55],pp27[88]};
    CLA_4 KS_269(s269, c269, in269_1, in269_2);
    wire[3:0] s270, in270_1, in270_2;
    wire c270;
    assign in270_1 = {pp60[52],pp60[53],pp60[54],pp28[87]};
    assign in270_2 = {pp61[51],pp61[52],pp61[53],pp29[86]};
    CLA_4 KS_270(s270, c270, in270_1, in270_2);
    wire[3:0] s271, in271_1, in271_2;
    wire c271;
    assign in271_1 = {pp62[50],pp62[51],pp62[52],pp30[85]};
    assign in271_2 = {pp63[49],pp63[50],pp63[51],pp31[84]};
    CLA_4 KS_271(s271, c271, in271_1, in271_2);
    wire[3:0] s272, in272_1, in272_2;
    wire c272;
    assign in272_1 = {pp64[48],pp64[49],pp64[50],pp32[83]};
    assign in272_2 = {pp65[47],pp65[48],pp65[49],pp33[82]};
    CLA_4 KS_272(s272, c272, in272_1, in272_2);
    wire[3:0] s273, in273_1, in273_2;
    wire c273;
    assign in273_1 = {pp66[46],pp66[47],pp66[48],pp34[81]};
    assign in273_2 = {pp67[45],pp67[46],pp67[47],pp35[80]};
    CLA_4 KS_273(s273, c273, in273_1, in273_2);
    wire[3:0] s274, in274_1, in274_2;
    wire c274;
    assign in274_1 = {pp68[44],pp68[45],pp68[46],pp36[79]};
    assign in274_2 = {pp69[43],pp69[44],pp69[45],pp37[78]};
    CLA_4 KS_274(s274, c274, in274_1, in274_2);
    wire[3:0] s275, in275_1, in275_2;
    wire c275;
    assign in275_1 = {pp70[42],pp70[43],pp70[44],pp38[77]};
    assign in275_2 = {pp71[41],pp71[42],pp71[43],pp39[76]};
    CLA_4 KS_275(s275, c275, in275_1, in275_2);
    wire[3:0] s276, in276_1, in276_2;
    wire c276;
    assign in276_1 = {pp72[40],pp72[41],pp72[42],pp40[75]};
    assign in276_2 = {pp73[39],pp73[40],pp73[41],pp41[74]};
    CLA_4 KS_276(s276, c276, in276_1, in276_2);
    wire[3:0] s277, in277_1, in277_2;
    wire c277;
    assign in277_1 = {pp74[38],pp74[39],pp74[40],pp42[73]};
    assign in277_2 = {pp75[37],pp75[38],pp75[39],pp43[72]};
    CLA_4 KS_277(s277, c277, in277_1, in277_2);
    wire[3:0] s278, in278_1, in278_2;
    wire c278;
    assign in278_1 = {pp76[36],pp76[37],pp76[38],pp44[71]};
    assign in278_2 = {pp77[35],pp77[36],pp77[37],pp45[70]};
    CLA_4 KS_278(s278, c278, in278_1, in278_2);
    wire[0:0] s279, in279_1, in279_2;
    wire c279;
    assign in279_1 = {pp78[34]};
    assign in279_2 = {pp79[33]};
    Half_Adder KS_279(s279, c279, in279_1, in279_2);
    wire[3:0] s280, in280_1, in280_2;
    wire c280;
    assign in280_1 = {pp80[32],pp78[35],pp78[36],pp46[69]};
    assign in280_2 = {pp81[31],pp79[34],pp79[35],pp47[68]};
    CLA_4 KS_280(s280, c280, in280_1, in280_2);
    wire[0:0] s281, in281_1, in281_2;
    wire c281;
    assign in281_1 = {pp82[30]};
    assign in281_2 = {pp83[29]};
    Half_Adder KS_281(s281, c281, in281_1, in281_2);
    wire[1:0] s282, in282_1, in282_2;
    wire c282;
    assign in282_1 = {pp84[28],pp80[33]};
    assign in282_2 = {pp85[27],pp81[32]};
    CLA_2 KS_282(s282, c282, in282_1, in282_2);
    wire[0:0] s283, in283_1, in283_2;
    wire c283;
    assign in283_1 = {pp86[26]};
    assign in283_2 = {pp87[25]};
    Half_Adder KS_283(s283, c283, in283_1, in283_2);
    wire[3:0] s284, in284_1, in284_2;
    wire c284;
    assign in284_1 = {pp88[24],pp82[31],pp80[34],pp48[67]};
    assign in284_2 = {pp89[23],pp83[30],pp81[33],pp49[66]};
    CLA_4 KS_284(s284, c284, in284_1, in284_2);
    wire[0:0] s285, in285_1, in285_2;
    wire c285;
    assign in285_1 = {pp90[22]};
    assign in285_2 = {pp91[21]};
    Half_Adder KS_285(s285, c285, in285_1, in285_2);
    wire[1:0] s286, in286_1, in286_2;
    wire c286;
    assign in286_1 = {pp92[20],pp84[29]};
    assign in286_2 = {pp93[19],pp85[28]};
    CLA_2 KS_286(s286, c286, in286_1, in286_2);
    wire[0:0] s287, in287_1, in287_2;
    wire c287;
    assign in287_1 = {pp94[18]};
    assign in287_2 = {pp95[17]};
    Half_Adder KS_287(s287, c287, in287_1, in287_2);
    wire[3:0] s288, in288_1, in288_2;
    wire c288;
    assign in288_1 = {pp96[16],pp86[27],pp82[32],pp50[65]};
    assign in288_2 = {pp97[15],pp87[26],pp83[31],pp51[64]};
    CLA_4 KS_288(s288, c288, in288_1, in288_2);
    wire[0:0] s289, in289_1, in289_2;
    wire c289;
    assign in289_1 = {pp98[14]};
    assign in289_2 = {pp99[13]};
    Half_Adder KS_289(s289, c289, in289_1, in289_2);
    wire[1:0] s290, in290_1, in290_2;
    wire c290;
    assign in290_1 = {pp100[12],pp88[25]};
    assign in290_2 = {pp101[11],pp89[24]};
    CLA_2 KS_290(s290, c290, in290_1, in290_2);
    wire[0:0] s291, in291_1, in291_2;
    wire c291;
    assign in291_1 = {pp102[10]};
    assign in291_2 = {pp103[9]};
    Half_Adder KS_291(s291, c291, in291_1, in291_2);
    wire[3:0] s292, in292_1, in292_2;
    wire c292;
    assign in292_1 = {pp104[8],pp90[23],pp84[30],pp52[63]};
    assign in292_2 = {pp105[7],pp91[22],pp85[29],pp53[62]};
    CLA_4 KS_292(s292, c292, in292_1, in292_2);
    wire[0:0] s293, in293_1, in293_2;
    wire c293;
    assign in293_1 = {pp106[6]};
    assign in293_2 = {pp107[5]};
    Half_Adder KS_293(s293, c293, in293_1, in293_2);
    wire[1:0] s294, in294_1, in294_2;
    wire c294;
    assign in294_1 = {pp108[4],pp92[21]};
    assign in294_2 = {pp109[3],pp93[20]};
    CLA_2 KS_294(s294, c294, in294_1, in294_2);
    wire[0:0] s295, in295_1, in295_2;
    wire c295;
    assign in295_1 = {pp110[2]};
    assign in295_2 = {pp111[1]};
    Half_Adder KS_295(s295, c295, in295_1, in295_2);
    wire[3:0] s296, in296_1, in296_2;
    wire c296;
    assign in296_1 = {pp112[0],pp94[19],pp86[28],pp54[61]};
    assign in296_2 = {c191,pp95[18],pp87[27],pp55[60]};
    CLA_4 KS_296(s296, c296, in296_1, in296_2);
    wire[0:0] s297, in297_1, in297_2;
    wire c297;
    assign in297_1 = {c192};
    assign in297_2 = {c193};
    Half_Adder KS_297(s297, c297, in297_1, in297_2);
    wire[1:0] s298, in298_1, in298_2;
    wire c298;
    assign in298_1 = {c194,pp96[17]};
    assign in298_2 = {c195,pp97[16]};
    CLA_2 KS_298(s298, c298, in298_1, in298_2);
    wire[0:0] s299, in299_1, in299_2;
    wire c299;
    assign in299_1 = {c196};
    assign in299_2 = {c197};
    Half_Adder KS_299(s299, c299, in299_1, in299_2);
    wire[3:0] s300, in300_1, in300_2;
    wire c300;
    assign in300_1 = {c198,pp98[15],pp88[26],pp56[59]};
    assign in300_2 = {c199,pp99[14],pp89[25],pp57[58]};
    CLA_4 KS_300(s300, c300, in300_1, in300_2);
    wire[0:0] s301, in301_1, in301_2;
    wire c301;
    assign in301_1 = {c200};
    assign in301_2 = {c201};
    Half_Adder KS_301(s301, c301, in301_1, in301_2);
    wire[1:0] s302, in302_1, in302_2;
    wire c302;
    assign in302_1 = {c202,pp100[13]};
    assign in302_2 = {c203,pp101[12]};
    CLA_2 KS_302(s302, c302, in302_1, in302_2);
    wire[0:0] s303, in303_1, in303_2;
    wire c303;
    assign in303_1 = {c204};
    assign in303_2 = {c205};
    Half_Adder KS_303(s303, c303, in303_1, in303_2);
    wire[3:0] s304, in304_1, in304_2;
    wire c304;
    assign in304_1 = {c206,pp102[11],pp90[24],pp58[57]};
    assign in304_2 = {c207,pp103[10],pp91[23],pp59[56]};
    CLA_4 KS_304(s304, c304, in304_1, in304_2);
    wire[0:0] s305, in305_1, in305_2;
    wire c305;
    assign in305_1 = {c209};
    assign in305_2 = {c210};
    Full_Adder KS_305(s305, c305, in305_1, in305_2, c208);
    wire[3:0] s306, in306_1, in306_2;
    wire c306;
    assign in306_1 = {pp60[55],pp0[116],pp0[117],pp0[118]};
    assign in306_2 = {pp61[54],pp1[115],pp1[116],pp1[117]};
    CLA_4 KS_306(s306, c306, in306_1, in306_2);
    wire[3:0] s307, in307_1, in307_2;
    wire c307;
    assign in307_1 = {pp62[53],pp2[114],pp2[115],pp2[116]};
    assign in307_2 = {pp63[52],pp3[113],pp3[114],pp3[115]};
    CLA_4 KS_307(s307, c307, in307_1, in307_2);
    wire[3:0] s308, in308_1, in308_2;
    wire c308;
    assign in308_1 = {pp64[51],pp4[112],pp4[113],pp4[114]};
    assign in308_2 = {pp65[50],pp5[111],pp5[112],pp5[113]};
    CLA_4 KS_308(s308, c308, in308_1, in308_2);
    wire[3:0] s309, in309_1, in309_2;
    wire c309;
    assign in309_1 = {pp66[49],pp6[110],pp6[111],pp6[112]};
    assign in309_2 = {pp67[48],pp7[109],pp7[110],pp7[111]};
    CLA_4 KS_309(s309, c309, in309_1, in309_2);
    wire[3:0] s310, in310_1, in310_2;
    wire c310;
    assign in310_1 = {pp68[47],pp8[108],pp8[109],pp8[110]};
    assign in310_2 = {pp69[46],pp9[107],pp9[108],pp9[109]};
    CLA_4 KS_310(s310, c310, in310_1, in310_2);
    wire[3:0] s311, in311_1, in311_2;
    wire c311;
    assign in311_1 = {pp70[45],pp10[106],pp10[107],pp10[108]};
    assign in311_2 = {pp71[44],pp11[105],pp11[106],pp11[107]};
    CLA_4 KS_311(s311, c311, in311_1, in311_2);
    wire[3:0] s312, in312_1, in312_2;
    wire c312;
    assign in312_1 = {pp72[43],pp12[104],pp12[105],pp12[106]};
    assign in312_2 = {pp73[42],pp13[103],pp13[104],pp13[105]};
    CLA_4 KS_312(s312, c312, in312_1, in312_2);
    wire[3:0] s313, in313_1, in313_2;
    wire c313;
    assign in313_1 = {pp74[41],pp14[102],pp14[103],pp14[104]};
    assign in313_2 = {pp75[40],pp15[101],pp15[102],pp15[103]};
    CLA_4 KS_313(s313, c313, in313_1, in313_2);
    wire[3:0] s314, in314_1, in314_2;
    wire c314;
    assign in314_1 = {pp76[39],pp16[100],pp16[101],pp16[102]};
    assign in314_2 = {pp77[38],pp17[99],pp17[100],pp17[101]};
    CLA_4 KS_314(s314, c314, in314_1, in314_2);
    wire[3:0] s315, in315_1, in315_2;
    wire c315;
    assign in315_1 = {pp78[37],pp18[98],pp18[99],pp18[100]};
    assign in315_2 = {pp79[36],pp19[97],pp19[98],pp19[99]};
    CLA_4 KS_315(s315, c315, in315_1, in315_2);
    wire[3:0] s316, in316_1, in316_2;
    wire c316;
    assign in316_1 = {pp80[35],pp20[96],pp20[97],pp20[98]};
    assign in316_2 = {pp81[34],pp21[95],pp21[96],pp21[97]};
    CLA_4 KS_316(s316, c316, in316_1, in316_2);
    wire[3:0] s317, in317_1, in317_2;
    wire c317;
    assign in317_1 = {pp82[33],pp22[94],pp22[95],pp22[96]};
    assign in317_2 = {pp83[32],pp23[93],pp23[94],pp23[95]};
    CLA_4 KS_317(s317, c317, in317_1, in317_2);
    wire[3:0] s318, in318_1, in318_2;
    wire c318;
    assign in318_1 = {pp84[31],pp24[92],pp24[93],pp24[94]};
    assign in318_2 = {pp85[30],pp25[91],pp25[92],pp25[93]};
    CLA_4 KS_318(s318, c318, in318_1, in318_2);
    wire[3:0] s319, in319_1, in319_2;
    wire c319;
    assign in319_1 = {pp86[29],pp26[90],pp26[91],pp26[92]};
    assign in319_2 = {pp87[28],pp27[89],pp27[90],pp27[91]};
    CLA_4 KS_319(s319, c319, in319_1, in319_2);
    wire[3:0] s320, in320_1, in320_2;
    wire c320;
    assign in320_1 = {pp88[27],pp28[88],pp28[89],pp28[90]};
    assign in320_2 = {pp89[26],pp29[87],pp29[88],pp29[89]};
    CLA_4 KS_320(s320, c320, in320_1, in320_2);
    wire[3:0] s321, in321_1, in321_2;
    wire c321;
    assign in321_1 = {pp90[25],pp30[86],pp30[87],pp30[88]};
    assign in321_2 = {pp91[24],pp31[85],pp31[86],pp31[87]};
    CLA_4 KS_321(s321, c321, in321_1, in321_2);
    wire[3:0] s322, in322_1, in322_2;
    wire c322;
    assign in322_1 = {pp92[23],pp32[84],pp32[85],pp32[86]};
    assign in322_2 = {pp93[22],pp33[83],pp33[84],pp33[85]};
    CLA_4 KS_322(s322, c322, in322_1, in322_2);
    wire[3:0] s323, in323_1, in323_2;
    wire c323;
    assign in323_1 = {pp94[21],pp34[82],pp34[83],pp34[84]};
    assign in323_2 = {pp95[20],pp35[81],pp35[82],pp35[83]};
    CLA_4 KS_323(s323, c323, in323_1, in323_2);
    wire[3:0] s324, in324_1, in324_2;
    wire c324;
    assign in324_1 = {pp96[19],pp36[80],pp36[81],pp36[82]};
    assign in324_2 = {pp97[18],pp37[79],pp37[80],pp37[81]};
    CLA_4 KS_324(s324, c324, in324_1, in324_2);
    wire[3:0] s325, in325_1, in325_2;
    wire c325;
    assign in325_1 = {pp98[17],pp38[78],pp38[79],pp38[80]};
    assign in325_2 = {pp99[16],pp39[77],pp39[78],pp39[79]};
    CLA_4 KS_325(s325, c325, in325_1, in325_2);
    wire[3:0] s326, in326_1, in326_2;
    wire c326;
    assign in326_1 = {pp100[15],pp40[76],pp40[77],pp40[78]};
    assign in326_2 = {pp101[14],pp41[75],pp41[76],pp41[77]};
    CLA_4 KS_326(s326, c326, in326_1, in326_2);
    wire[3:0] s327, in327_1, in327_2;
    wire c327;
    assign in327_1 = {pp102[13],pp42[74],pp42[75],pp42[76]};
    assign in327_2 = {pp103[12],pp43[73],pp43[74],pp43[75]};
    CLA_4 KS_327(s327, c327, in327_1, in327_2);
    wire[3:0] s328, in328_1, in328_2;
    wire c328;
    assign in328_1 = {pp104[11],pp44[72],pp44[73],pp44[74]};
    assign in328_2 = {pp105[10],pp45[71],pp45[72],pp45[73]};
    CLA_4 KS_328(s328, c328, in328_1, in328_2);
    wire[3:0] s329, in329_1, in329_2;
    wire c329;
    assign in329_1 = {pp106[9],pp46[70],pp46[71],pp46[72]};
    assign in329_2 = {pp107[8],pp47[69],pp47[70],pp47[71]};
    CLA_4 KS_329(s329, c329, in329_1, in329_2);
    wire[3:0] s330, in330_1, in330_2;
    wire c330;
    assign in330_1 = {pp109[6],pp48[68],pp48[69],pp48[70]};
    assign in330_2 = {pp110[5],pp49[67],pp49[68],pp49[69]};
    CLA_4_c KS_330(s330, c330, in330_1, in330_2, pp108[7]);
    wire[3:0] s331, in331_1, in331_2;
    wire c331;
    assign in331_1 = {pp50[66],pp50[67],pp50[68],pp0[119]};
    assign in331_2 = {pp51[65],pp51[66],pp51[67],pp1[118]};
    CLA_4 KS_331(s331, c331, in331_1, in331_2);
    wire[3:0] s332, in332_1, in332_2;
    wire c332;
    assign in332_1 = {pp52[64],pp52[65],pp52[66],pp2[117]};
    assign in332_2 = {pp53[63],pp53[64],pp53[65],pp3[116]};
    CLA_4 KS_332(s332, c332, in332_1, in332_2);
    wire[3:0] s333, in333_1, in333_2;
    wire c333;
    assign in333_1 = {pp54[62],pp54[63],pp54[64],pp4[115]};
    assign in333_2 = {pp55[61],pp55[62],pp55[63],pp5[114]};
    CLA_4 KS_333(s333, c333, in333_1, in333_2);
    wire[3:0] s334, in334_1, in334_2;
    wire c334;
    assign in334_1 = {pp56[60],pp56[61],pp56[62],pp6[113]};
    assign in334_2 = {pp57[59],pp57[60],pp57[61],pp7[112]};
    CLA_4 KS_334(s334, c334, in334_1, in334_2);
    wire[3:0] s335, in335_1, in335_2;
    wire c335;
    assign in335_1 = {pp58[58],pp58[59],pp58[60],pp8[111]};
    assign in335_2 = {pp59[57],pp59[58],pp59[59],pp9[110]};
    CLA_4 KS_335(s335, c335, in335_1, in335_2);
    wire[3:0] s336, in336_1, in336_2;
    wire c336;
    assign in336_1 = {pp60[56],pp60[57],pp60[58],pp10[109]};
    assign in336_2 = {pp61[55],pp61[56],pp61[57],pp11[108]};
    CLA_4 KS_336(s336, c336, in336_1, in336_2);
    wire[3:0] s337, in337_1, in337_2;
    wire c337;
    assign in337_1 = {pp62[54],pp62[55],pp62[56],pp12[107]};
    assign in337_2 = {pp63[53],pp63[54],pp63[55],pp13[106]};
    CLA_4 KS_337(s337, c337, in337_1, in337_2);
    wire[3:0] s338, in338_1, in338_2;
    wire c338;
    assign in338_1 = {pp64[52],pp64[53],pp64[54],pp14[105]};
    assign in338_2 = {pp65[51],pp65[52],pp65[53],pp15[104]};
    CLA_4 KS_338(s338, c338, in338_1, in338_2);
    wire[3:0] s339, in339_1, in339_2;
    wire c339;
    assign in339_1 = {pp66[50],pp66[51],pp66[52],pp16[103]};
    assign in339_2 = {pp67[49],pp67[50],pp67[51],pp17[102]};
    CLA_4 KS_339(s339, c339, in339_1, in339_2);
    wire[3:0] s340, in340_1, in340_2;
    wire c340;
    assign in340_1 = {pp68[48],pp68[49],pp68[50],pp18[101]};
    assign in340_2 = {pp69[47],pp69[48],pp69[49],pp19[100]};
    CLA_4 KS_340(s340, c340, in340_1, in340_2);
    wire[3:0] s341, in341_1, in341_2;
    wire c341;
    assign in341_1 = {pp70[46],pp70[47],pp70[48],pp20[99]};
    assign in341_2 = {pp71[45],pp71[46],pp71[47],pp21[98]};
    CLA_4 KS_341(s341, c341, in341_1, in341_2);
    wire[3:0] s342, in342_1, in342_2;
    wire c342;
    assign in342_1 = {pp72[44],pp72[45],pp72[46],pp22[97]};
    assign in342_2 = {pp73[43],pp73[44],pp73[45],pp23[96]};
    CLA_4 KS_342(s342, c342, in342_1, in342_2);
    wire[3:0] s343, in343_1, in343_2;
    wire c343;
    assign in343_1 = {pp74[42],pp74[43],pp74[44],pp24[95]};
    assign in343_2 = {pp75[41],pp75[42],pp75[43],pp25[94]};
    CLA_4 KS_343(s343, c343, in343_1, in343_2);
    wire[3:0] s344, in344_1, in344_2;
    wire c344;
    assign in344_1 = {pp76[40],pp76[41],pp76[42],pp26[93]};
    assign in344_2 = {pp77[39],pp77[40],pp77[41],pp27[92]};
    CLA_4 KS_344(s344, c344, in344_1, in344_2);
    wire[3:0] s345, in345_1, in345_2;
    wire c345;
    assign in345_1 = {pp78[38],pp78[39],pp78[40],pp28[91]};
    assign in345_2 = {pp79[37],pp79[38],pp79[39],pp29[90]};
    CLA_4 KS_345(s345, c345, in345_1, in345_2);
    wire[3:0] s346, in346_1, in346_2;
    wire c346;
    assign in346_1 = {pp80[36],pp80[37],pp80[38],pp30[89]};
    assign in346_2 = {pp81[35],pp81[36],pp81[37],pp31[88]};
    CLA_4 KS_346(s346, c346, in346_1, in346_2);
    wire[3:0] s347, in347_1, in347_2;
    wire c347;
    assign in347_1 = {pp82[34],pp82[35],pp82[36],pp32[87]};
    assign in347_2 = {pp83[33],pp83[34],pp83[35],pp33[86]};
    CLA_4 KS_347(s347, c347, in347_1, in347_2);
    wire[3:0] s348, in348_1, in348_2;
    wire c348;
    assign in348_1 = {pp84[32],pp84[33],pp84[34],pp34[85]};
    assign in348_2 = {pp85[31],pp85[32],pp85[33],pp35[84]};
    CLA_4 KS_348(s348, c348, in348_1, in348_2);
    wire[0:0] s349, in349_1, in349_2;
    wire c349;
    assign in349_1 = {pp86[30]};
    assign in349_2 = {pp87[29]};
    Half_Adder KS_349(s349, c349, in349_1, in349_2);
    wire[3:0] s350, in350_1, in350_2;
    wire c350;
    assign in350_1 = {pp88[28],pp86[31],pp86[32],pp36[83]};
    assign in350_2 = {pp89[27],pp87[30],pp87[31],pp37[82]};
    CLA_4 KS_350(s350, c350, in350_1, in350_2);
    wire[0:0] s351, in351_1, in351_2;
    wire c351;
    assign in351_1 = {pp90[26]};
    assign in351_2 = {pp91[25]};
    Half_Adder KS_351(s351, c351, in351_1, in351_2);
    wire[1:0] s352, in352_1, in352_2;
    wire c352;
    assign in352_1 = {pp92[24],pp88[29]};
    assign in352_2 = {pp93[23],pp89[28]};
    CLA_2 KS_352(s352, c352, in352_1, in352_2);
    wire[0:0] s353, in353_1, in353_2;
    wire c353;
    assign in353_1 = {pp94[22]};
    assign in353_2 = {pp95[21]};
    Half_Adder KS_353(s353, c353, in353_1, in353_2);
    wire[3:0] s354, in354_1, in354_2;
    wire c354;
    assign in354_1 = {pp96[20],pp90[27],pp88[30],pp38[81]};
    assign in354_2 = {pp97[19],pp91[26],pp89[29],pp39[80]};
    CLA_4 KS_354(s354, c354, in354_1, in354_2);
    wire[0:0] s355, in355_1, in355_2;
    wire c355;
    assign in355_1 = {pp98[18]};
    assign in355_2 = {pp99[17]};
    Half_Adder KS_355(s355, c355, in355_1, in355_2);
    wire[1:0] s356, in356_1, in356_2;
    wire c356;
    assign in356_1 = {pp100[16],pp92[25]};
    assign in356_2 = {pp101[15],pp93[24]};
    CLA_2 KS_356(s356, c356, in356_1, in356_2);
    wire[0:0] s357, in357_1, in357_2;
    wire c357;
    assign in357_1 = {pp102[14]};
    assign in357_2 = {pp103[13]};
    Half_Adder KS_357(s357, c357, in357_1, in357_2);
    wire[3:0] s358, in358_1, in358_2;
    wire c358;
    assign in358_1 = {pp104[12],pp94[23],pp90[28],pp40[79]};
    assign in358_2 = {pp105[11],pp95[22],pp91[27],pp41[78]};
    CLA_4 KS_358(s358, c358, in358_1, in358_2);
    wire[0:0] s359, in359_1, in359_2;
    wire c359;
    assign in359_1 = {pp106[10]};
    assign in359_2 = {pp107[9]};
    Half_Adder KS_359(s359, c359, in359_1, in359_2);
    wire[1:0] s360, in360_1, in360_2;
    wire c360;
    assign in360_1 = {pp108[8],pp96[21]};
    assign in360_2 = {pp109[7],pp97[20]};
    CLA_2 KS_360(s360, c360, in360_1, in360_2);
    wire[0:0] s361, in361_1, in361_2;
    wire c361;
    assign in361_1 = {pp110[6]};
    assign in361_2 = {pp111[5]};
    Half_Adder KS_361(s361, c361, in361_1, in361_2);
    wire[3:0] s362, in362_1, in362_2;
    wire c362;
    assign in362_1 = {pp112[4],pp98[19],pp92[26],pp42[77]};
    assign in362_2 = {pp113[3],pp99[18],pp93[25],pp43[76]};
    CLA_4 KS_362(s362, c362, in362_1, in362_2);
    wire[0:0] s363, in363_1, in363_2;
    wire c363;
    assign in363_1 = {pp114[2]};
    assign in363_2 = {pp115[1]};
    Half_Adder KS_363(s363, c363, in363_1, in363_2);
    wire[1:0] s364, in364_1, in364_2;
    wire c364;
    assign in364_1 = {pp116[0],pp100[17]};
    assign in364_2 = {c256,pp101[16]};
    CLA_2 KS_364(s364, c364, in364_1, in364_2);
    wire[0:0] s365, in365_1, in365_2;
    wire c365;
    assign in365_1 = {c257};
    assign in365_2 = {c258};
    Half_Adder KS_365(s365, c365, in365_1, in365_2);
    wire[3:0] s366, in366_1, in366_2;
    wire c366;
    assign in366_1 = {c259,pp102[15],pp94[24],pp44[75]};
    assign in366_2 = {c260,pp103[14],pp95[23],pp45[74]};
    CLA_4 KS_366(s366, c366, in366_1, in366_2);
    wire[0:0] s367, in367_1, in367_2;
    wire c367;
    assign in367_1 = {c261};
    assign in367_2 = {c262};
    Half_Adder KS_367(s367, c367, in367_1, in367_2);
    wire[1:0] s368, in368_1, in368_2;
    wire c368;
    assign in368_1 = {c263,pp104[13]};
    assign in368_2 = {c264,pp105[12]};
    CLA_2 KS_368(s368, c368, in368_1, in368_2);
    wire[0:0] s369, in369_1, in369_2;
    wire c369;
    assign in369_1 = {c265};
    assign in369_2 = {c266};
    Half_Adder KS_369(s369, c369, in369_1, in369_2);
    wire[3:0] s370, in370_1, in370_2;
    wire c370;
    assign in370_1 = {c267,pp106[11],pp96[22],pp46[73]};
    assign in370_2 = {c268,pp107[10],pp97[21],pp47[72]};
    CLA_4 KS_370(s370, c370, in370_1, in370_2);
    wire[0:0] s371, in371_1, in371_2;
    wire c371;
    assign in371_1 = {c269};
    assign in371_2 = {c270};
    Half_Adder KS_371(s371, c371, in371_1, in371_2);
    wire[1:0] s372, in372_1, in372_2;
    wire c372;
    assign in372_1 = {c271,pp108[9]};
    assign in372_2 = {c272,pp109[8]};
    CLA_2 KS_372(s372, c372, in372_1, in372_2);
    wire[0:0] s373, in373_1, in373_2;
    wire c373;
    assign in373_1 = {c273};
    assign in373_2 = {c274};
    Half_Adder KS_373(s373, c373, in373_1, in373_2);
    wire[3:0] s374, in374_1, in374_2;
    wire c374;
    assign in374_1 = {c275,pp110[7],pp98[20],pp48[71]};
    assign in374_2 = {c276,pp111[6],pp99[19],pp49[70]};
    CLA_4 KS_374(s374, c374, in374_1, in374_2);
    wire[0:0] s375, in375_1, in375_2;
    wire c375;
    assign in375_1 = {c278};
    assign in375_2 = {c280};
    Full_Adder KS_375(s375, c375, in375_1, in375_2, c277);
    wire[3:0] s376, in376_1, in376_2;
    wire c376;
    assign in376_1 = {pp50[69],pp0[120],pp0[121],pp0[122]};
    assign in376_2 = {pp51[68],pp1[119],pp1[120],pp1[121]};
    CLA_4 KS_376(s376, c376, in376_1, in376_2);
    wire[3:0] s377, in377_1, in377_2;
    wire c377;
    assign in377_1 = {pp52[67],pp2[118],pp2[119],pp2[120]};
    assign in377_2 = {pp53[66],pp3[117],pp3[118],pp3[119]};
    CLA_4 KS_377(s377, c377, in377_1, in377_2);
    wire[3:0] s378, in378_1, in378_2;
    wire c378;
    assign in378_1 = {pp54[65],pp4[116],pp4[117],pp4[118]};
    assign in378_2 = {pp55[64],pp5[115],pp5[116],pp5[117]};
    CLA_4 KS_378(s378, c378, in378_1, in378_2);
    wire[3:0] s379, in379_1, in379_2;
    wire c379;
    assign in379_1 = {pp56[63],pp6[114],pp6[115],pp6[116]};
    assign in379_2 = {pp57[62],pp7[113],pp7[114],pp7[115]};
    CLA_4 KS_379(s379, c379, in379_1, in379_2);
    wire[3:0] s380, in380_1, in380_2;
    wire c380;
    assign in380_1 = {pp58[61],pp8[112],pp8[113],pp8[114]};
    assign in380_2 = {pp59[60],pp9[111],pp9[112],pp9[113]};
    CLA_4 KS_380(s380, c380, in380_1, in380_2);
    wire[3:0] s381, in381_1, in381_2;
    wire c381;
    assign in381_1 = {pp60[59],pp10[110],pp10[111],pp10[112]};
    assign in381_2 = {pp61[58],pp11[109],pp11[110],pp11[111]};
    CLA_4 KS_381(s381, c381, in381_1, in381_2);
    wire[3:0] s382, in382_1, in382_2;
    wire c382;
    assign in382_1 = {pp62[57],pp12[108],pp12[109],pp12[110]};
    assign in382_2 = {pp63[56],pp13[107],pp13[108],pp13[109]};
    CLA_4 KS_382(s382, c382, in382_1, in382_2);
    wire[3:0] s383, in383_1, in383_2;
    wire c383;
    assign in383_1 = {pp64[55],pp14[106],pp14[107],pp14[108]};
    assign in383_2 = {pp65[54],pp15[105],pp15[106],pp15[107]};
    CLA_4 KS_383(s383, c383, in383_1, in383_2);
    wire[3:0] s384, in384_1, in384_2;
    wire c384;
    assign in384_1 = {pp66[53],pp16[104],pp16[105],pp16[106]};
    assign in384_2 = {pp67[52],pp17[103],pp17[104],pp17[105]};
    CLA_4 KS_384(s384, c384, in384_1, in384_2);
    wire[3:0] s385, in385_1, in385_2;
    wire c385;
    assign in385_1 = {pp68[51],pp18[102],pp18[103],pp18[104]};
    assign in385_2 = {pp69[50],pp19[101],pp19[102],pp19[103]};
    CLA_4 KS_385(s385, c385, in385_1, in385_2);
    wire[3:0] s386, in386_1, in386_2;
    wire c386;
    assign in386_1 = {pp70[49],pp20[100],pp20[101],pp20[102]};
    assign in386_2 = {pp71[48],pp21[99],pp21[100],pp21[101]};
    CLA_4 KS_386(s386, c386, in386_1, in386_2);
    wire[3:0] s387, in387_1, in387_2;
    wire c387;
    assign in387_1 = {pp72[47],pp22[98],pp22[99],pp22[100]};
    assign in387_2 = {pp73[46],pp23[97],pp23[98],pp23[99]};
    CLA_4 KS_387(s387, c387, in387_1, in387_2);
    wire[3:0] s388, in388_1, in388_2;
    wire c388;
    assign in388_1 = {pp74[45],pp24[96],pp24[97],pp24[98]};
    assign in388_2 = {pp75[44],pp25[95],pp25[96],pp25[97]};
    CLA_4 KS_388(s388, c388, in388_1, in388_2);
    wire[3:0] s389, in389_1, in389_2;
    wire c389;
    assign in389_1 = {pp76[43],pp26[94],pp26[95],pp26[96]};
    assign in389_2 = {pp77[42],pp27[93],pp27[94],pp27[95]};
    CLA_4 KS_389(s389, c389, in389_1, in389_2);
    wire[3:0] s390, in390_1, in390_2;
    wire c390;
    assign in390_1 = {pp78[41],pp28[92],pp28[93],pp28[94]};
    assign in390_2 = {pp79[40],pp29[91],pp29[92],pp29[93]};
    CLA_4 KS_390(s390, c390, in390_1, in390_2);
    wire[3:0] s391, in391_1, in391_2;
    wire c391;
    assign in391_1 = {pp80[39],pp30[90],pp30[91],pp30[92]};
    assign in391_2 = {pp81[38],pp31[89],pp31[90],pp31[91]};
    CLA_4 KS_391(s391, c391, in391_1, in391_2);
    wire[3:0] s392, in392_1, in392_2;
    wire c392;
    assign in392_1 = {pp82[37],pp32[88],pp32[89],pp32[90]};
    assign in392_2 = {pp83[36],pp33[87],pp33[88],pp33[89]};
    CLA_4 KS_392(s392, c392, in392_1, in392_2);
    wire[3:0] s393, in393_1, in393_2;
    wire c393;
    assign in393_1 = {pp84[35],pp34[86],pp34[87],pp34[88]};
    assign in393_2 = {pp85[34],pp35[85],pp35[86],pp35[87]};
    CLA_4 KS_393(s393, c393, in393_1, in393_2);
    wire[3:0] s394, in394_1, in394_2;
    wire c394;
    assign in394_1 = {pp86[33],pp36[84],pp36[85],pp36[86]};
    assign in394_2 = {pp87[32],pp37[83],pp37[84],pp37[85]};
    CLA_4 KS_394(s394, c394, in394_1, in394_2);
    wire[3:0] s395, in395_1, in395_2;
    wire c395;
    assign in395_1 = {pp88[31],pp38[82],pp38[83],pp38[84]};
    assign in395_2 = {pp89[30],pp39[81],pp39[82],pp39[83]};
    CLA_4 KS_395(s395, c395, in395_1, in395_2);
    wire[3:0] s396, in396_1, in396_2;
    wire c396;
    assign in396_1 = {pp90[29],pp40[80],pp40[81],pp40[82]};
    assign in396_2 = {pp91[28],pp41[79],pp41[80],pp41[81]};
    CLA_4 KS_396(s396, c396, in396_1, in396_2);
    wire[3:0] s397, in397_1, in397_2;
    wire c397;
    assign in397_1 = {pp92[27],pp42[78],pp42[79],pp42[80]};
    assign in397_2 = {pp93[26],pp43[77],pp43[78],pp43[79]};
    CLA_4 KS_397(s397, c397, in397_1, in397_2);
    wire[3:0] s398, in398_1, in398_2;
    wire c398;
    assign in398_1 = {pp94[25],pp44[76],pp44[77],pp44[78]};
    assign in398_2 = {pp95[24],pp45[75],pp45[76],pp45[77]};
    CLA_4 KS_398(s398, c398, in398_1, in398_2);
    wire[3:0] s399, in399_1, in399_2;
    wire c399;
    assign in399_1 = {pp96[23],pp46[74],pp46[75],pp46[76]};
    assign in399_2 = {pp97[22],pp47[73],pp47[74],pp47[75]};
    CLA_4 KS_399(s399, c399, in399_1, in399_2);
    wire[3:0] s400, in400_1, in400_2;
    wire c400;
    assign in400_1 = {pp98[21],pp48[72],pp48[73],pp48[74]};
    assign in400_2 = {pp99[20],pp49[71],pp49[72],pp49[73]};
    CLA_4 KS_400(s400, c400, in400_1, in400_2);
    wire[3:0] s401, in401_1, in401_2;
    wire c401;
    assign in401_1 = {pp100[19],pp50[70],pp50[71],pp50[72]};
    assign in401_2 = {pp101[18],pp51[69],pp51[70],pp51[71]};
    CLA_4 KS_401(s401, c401, in401_1, in401_2);
    wire[3:0] s402, in402_1, in402_2;
    wire c402;
    assign in402_1 = {pp102[17],pp52[68],pp52[69],pp52[70]};
    assign in402_2 = {pp103[16],pp53[67],pp53[68],pp53[69]};
    CLA_4 KS_402(s402, c402, in402_1, in402_2);
    wire[3:0] s403, in403_1, in403_2;
    wire c403;
    assign in403_1 = {pp104[15],pp54[66],pp54[67],pp54[68]};
    assign in403_2 = {pp105[14],pp55[65],pp55[66],pp55[67]};
    CLA_4 KS_403(s403, c403, in403_1, in403_2);
    wire[3:0] s404, in404_1, in404_2;
    wire c404;
    assign in404_1 = {pp106[13],pp56[64],pp56[65],pp56[66]};
    assign in404_2 = {pp107[12],pp57[63],pp57[64],pp57[65]};
    CLA_4 KS_404(s404, c404, in404_1, in404_2);
    wire[3:0] s405, in405_1, in405_2;
    wire c405;
    assign in405_1 = {pp108[11],pp58[62],pp58[63],pp58[64]};
    assign in405_2 = {pp109[10],pp59[61],pp59[62],pp59[63]};
    CLA_4 KS_405(s405, c405, in405_1, in405_2);
    wire[3:0] s406, in406_1, in406_2;
    wire c406;
    assign in406_1 = {pp110[9],pp60[60],pp60[61],pp60[62]};
    assign in406_2 = {pp111[8],pp61[59],pp61[60],pp61[61]};
    CLA_4 KS_406(s406, c406, in406_1, in406_2);
    wire[3:0] s407, in407_1, in407_2;
    wire c407;
    assign in407_1 = {pp112[7],pp62[58],pp62[59],pp62[60]};
    assign in407_2 = {pp113[6],pp63[57],pp63[58],pp63[59]};
    CLA_4 KS_407(s407, c407, in407_1, in407_2);
    wire[3:0] s408, in408_1, in408_2;
    wire c408;
    assign in408_1 = {pp114[5],pp64[56],pp64[57],pp64[58]};
    assign in408_2 = {pp115[4],pp65[55],pp65[56],pp65[57]};
    CLA_4 KS_408(s408, c408, in408_1, in408_2);
    wire[3:0] s409, in409_1, in409_2;
    wire c409;
    assign in409_1 = {pp116[3],pp66[54],pp66[55],pp66[56]};
    assign in409_2 = {pp117[2],pp67[53],pp67[54],pp67[55]};
    CLA_4 KS_409(s409, c409, in409_1, in409_2);
    wire[3:0] s410, in410_1, in410_2;
    wire c410;
    assign in410_1 = {pp118[1],pp68[52],pp68[53],pp68[54]};
    assign in410_2 = {pp119[0],pp69[51],pp69[52],pp69[53]};
    CLA_4 KS_410(s410, c410, in410_1, in410_2);
    wire[3:0] s411, in411_1, in411_2;
    wire c411;
    assign in411_1 = {c306,pp70[50],pp70[51],pp70[52]};
    assign in411_2 = {c307,pp71[49],pp71[50],pp71[51]};
    CLA_4 KS_411(s411, c411, in411_1, in411_2);
    wire[3:0] s412, in412_1, in412_2;
    wire c412;
    assign in412_1 = {c308,pp72[48],pp72[49],pp72[50]};
    assign in412_2 = {c309,pp73[47],pp73[48],pp73[49]};
    CLA_4 KS_412(s412, c412, in412_1, in412_2);
    wire[3:0] s413, in413_1, in413_2;
    wire c413;
    assign in413_1 = {c310,pp74[46],pp74[47],pp74[48]};
    assign in413_2 = {c311,pp75[45],pp75[46],pp75[47]};
    CLA_4 KS_413(s413, c413, in413_1, in413_2);
    wire[3:0] s414, in414_1, in414_2;
    wire c414;
    assign in414_1 = {c312,pp76[44],pp76[45],pp76[46]};
    assign in414_2 = {c313,pp77[43],pp77[44],pp77[45]};
    CLA_4 KS_414(s414, c414, in414_1, in414_2);
    wire[3:0] s415, in415_1, in415_2;
    wire c415;
    assign in415_1 = {c314,pp78[42],pp78[43],pp78[44]};
    assign in415_2 = {c315,pp79[41],pp79[42],pp79[43]};
    CLA_4 KS_415(s415, c415, in415_1, in415_2);
    wire[3:0] s416, in416_1, in416_2;
    wire c416;
    assign in416_1 = {c316,pp80[40],pp80[41],pp80[42]};
    assign in416_2 = {c317,pp81[39],pp81[40],pp81[41]};
    CLA_4 KS_416(s416, c416, in416_1, in416_2);
    wire[3:0] s417, in417_1, in417_2;
    wire c417;
    assign in417_1 = {c318,pp82[38],pp82[39],pp82[40]};
    assign in417_2 = {c319,pp83[37],pp83[38],pp83[39]};
    CLA_4 KS_417(s417, c417, in417_1, in417_2);
    wire[3:0] s418, in418_1, in418_2;
    wire c418;
    assign in418_1 = {c321,pp84[36],pp84[37],pp84[38]};
    assign in418_2 = {c322,pp85[35],pp85[36],pp85[37]};
    CLA_4_c KS_418(s418, c418, in418_1, in418_2, c320);
    wire[3:0] s419, in419_1, in419_2;
    wire c419;
    assign in419_1 = {pp86[34],pp86[35],pp86[36],pp0[123]};
    assign in419_2 = {pp87[33],pp87[34],pp87[35],pp1[122]};
    CLA_4 KS_419(s419, c419, in419_1, in419_2);
    wire[3:0] s420, in420_1, in420_2;
    wire c420;
    assign in420_1 = {pp88[32],pp88[33],pp88[34],pp2[121]};
    assign in420_2 = {pp89[31],pp89[32],pp89[33],pp3[120]};
    CLA_4 KS_420(s420, c420, in420_1, in420_2);
    wire[3:0] s421, in421_1, in421_2;
    wire c421;
    assign in421_1 = {pp90[30],pp90[31],pp90[32],pp4[119]};
    assign in421_2 = {pp91[29],pp91[30],pp91[31],pp5[118]};
    CLA_4 KS_421(s421, c421, in421_1, in421_2);
    wire[3:0] s422, in422_1, in422_2;
    wire c422;
    assign in422_1 = {pp92[28],pp92[29],pp92[30],pp6[117]};
    assign in422_2 = {pp93[27],pp93[28],pp93[29],pp7[116]};
    CLA_4 KS_422(s422, c422, in422_1, in422_2);
    wire[0:0] s423, in423_1, in423_2;
    wire c423;
    assign in423_1 = {pp94[26]};
    assign in423_2 = {pp95[25]};
    Half_Adder KS_423(s423, c423, in423_1, in423_2);
    wire[3:0] s424, in424_1, in424_2;
    wire c424;
    assign in424_1 = {pp96[24],pp94[27],pp94[28],pp8[115]};
    assign in424_2 = {pp97[23],pp95[26],pp95[27],pp9[114]};
    CLA_4 KS_424(s424, c424, in424_1, in424_2);
    wire[0:0] s425, in425_1, in425_2;
    wire c425;
    assign in425_1 = {pp98[22]};
    assign in425_2 = {pp99[21]};
    Half_Adder KS_425(s425, c425, in425_1, in425_2);
    wire[1:0] s426, in426_1, in426_2;
    wire c426;
    assign in426_1 = {pp100[20],pp96[25]};
    assign in426_2 = {pp101[19],pp97[24]};
    CLA_2 KS_426(s426, c426, in426_1, in426_2);
    wire[0:0] s427, in427_1, in427_2;
    wire c427;
    assign in427_1 = {pp102[18]};
    assign in427_2 = {pp103[17]};
    Half_Adder KS_427(s427, c427, in427_1, in427_2);
    wire[3:0] s428, in428_1, in428_2;
    wire c428;
    assign in428_1 = {pp104[16],pp98[23],pp96[26],pp10[113]};
    assign in428_2 = {pp105[15],pp99[22],pp97[25],pp11[112]};
    CLA_4 KS_428(s428, c428, in428_1, in428_2);
    wire[0:0] s429, in429_1, in429_2;
    wire c429;
    assign in429_1 = {pp106[14]};
    assign in429_2 = {pp107[13]};
    Half_Adder KS_429(s429, c429, in429_1, in429_2);
    wire[1:0] s430, in430_1, in430_2;
    wire c430;
    assign in430_1 = {pp108[12],pp100[21]};
    assign in430_2 = {pp109[11],pp101[20]};
    CLA_2 KS_430(s430, c430, in430_1, in430_2);
    wire[0:0] s431, in431_1, in431_2;
    wire c431;
    assign in431_1 = {pp110[10]};
    assign in431_2 = {pp111[9]};
    Half_Adder KS_431(s431, c431, in431_1, in431_2);
    wire[3:0] s432, in432_1, in432_2;
    wire c432;
    assign in432_1 = {pp112[8],pp102[19],pp98[24],pp12[111]};
    assign in432_2 = {pp113[7],pp103[18],pp99[23],pp13[110]};
    CLA_4 KS_432(s432, c432, in432_1, in432_2);
    wire[0:0] s433, in433_1, in433_2;
    wire c433;
    assign in433_1 = {pp114[6]};
    assign in433_2 = {pp115[5]};
    Half_Adder KS_433(s433, c433, in433_1, in433_2);
    wire[1:0] s434, in434_1, in434_2;
    wire c434;
    assign in434_1 = {pp116[4],pp104[17]};
    assign in434_2 = {pp117[3],pp105[16]};
    CLA_2 KS_434(s434, c434, in434_1, in434_2);
    wire[0:0] s435, in435_1, in435_2;
    wire c435;
    assign in435_1 = {pp118[2]};
    assign in435_2 = {pp119[1]};
    Half_Adder KS_435(s435, c435, in435_1, in435_2);
    wire[3:0] s436, in436_1, in436_2;
    wire c436;
    assign in436_1 = {pp120[0],pp106[15],pp100[22],pp14[109]};
    assign in436_2 = {c331,pp107[14],pp101[21],pp15[108]};
    CLA_4 KS_436(s436, c436, in436_1, in436_2);
    wire[0:0] s437, in437_1, in437_2;
    wire c437;
    assign in437_1 = {c332};
    assign in437_2 = {c333};
    Half_Adder KS_437(s437, c437, in437_1, in437_2);
    wire[1:0] s438, in438_1, in438_2;
    wire c438;
    assign in438_1 = {c334,pp108[13]};
    assign in438_2 = {c335,pp109[12]};
    CLA_2 KS_438(s438, c438, in438_1, in438_2);
    wire[0:0] s439, in439_1, in439_2;
    wire c439;
    assign in439_1 = {c336};
    assign in439_2 = {c337};
    Half_Adder KS_439(s439, c439, in439_1, in439_2);
    wire[3:0] s440, in440_1, in440_2;
    wire c440;
    assign in440_1 = {c338,pp110[11],pp102[20],pp16[107]};
    assign in440_2 = {c339,pp111[10],pp103[19],pp17[106]};
    CLA_4 KS_440(s440, c440, in440_1, in440_2);
    wire[0:0] s441, in441_1, in441_2;
    wire c441;
    assign in441_1 = {c340};
    assign in441_2 = {c341};
    Half_Adder KS_441(s441, c441, in441_1, in441_2);
    wire[1:0] s442, in442_1, in442_2;
    wire c442;
    assign in442_1 = {c342,pp112[9]};
    assign in442_2 = {c343,pp113[8]};
    CLA_2 KS_442(s442, c442, in442_1, in442_2);
    wire[0:0] s443, in443_1, in443_2;
    wire c443;
    assign in443_1 = {c344};
    assign in443_2 = {c345};
    Half_Adder KS_443(s443, c443, in443_1, in443_2);
    wire[3:0] s444, in444_1, in444_2;
    wire c444;
    assign in444_1 = {c347,pp114[7],pp104[18],pp18[105]};
    assign in444_2 = {c348,pp115[6],pp105[17],pp19[104]};
    CLA_4_c KS_444(s444, c444, in444_1, in444_2, c346);
    wire[3:0] s445, in445_1, in445_2;
    wire c445;
    assign in445_1 = {pp20[103],pp0[124],pp0[125],pp0[126]};
    assign in445_2 = {pp21[102],pp1[123],pp1[124],pp1[125]};
    CLA_4 KS_445(s445, c445, in445_1, in445_2);
    wire[3:0] s446, in446_1, in446_2;
    wire c446;
    assign in446_1 = {pp22[101],pp2[122],pp2[123],pp2[124]};
    assign in446_2 = {pp23[100],pp3[121],pp3[122],pp3[123]};
    CLA_4 KS_446(s446, c446, in446_1, in446_2);
    wire[3:0] s447, in447_1, in447_2;
    wire c447;
    assign in447_1 = {pp24[99],pp4[120],pp4[121],pp4[122]};
    assign in447_2 = {pp25[98],pp5[119],pp5[120],pp5[121]};
    CLA_4 KS_447(s447, c447, in447_1, in447_2);
    wire[3:0] s448, in448_1, in448_2;
    wire c448;
    assign in448_1 = {pp26[97],pp6[118],pp6[119],pp6[120]};
    assign in448_2 = {pp27[96],pp7[117],pp7[118],pp7[119]};
    CLA_4 KS_448(s448, c448, in448_1, in448_2);
    wire[3:0] s449, in449_1, in449_2;
    wire c449;
    assign in449_1 = {pp28[95],pp8[116],pp8[117],pp8[118]};
    assign in449_2 = {pp29[94],pp9[115],pp9[116],pp9[117]};
    CLA_4 KS_449(s449, c449, in449_1, in449_2);
    wire[3:0] s450, in450_1, in450_2;
    wire c450;
    assign in450_1 = {pp30[93],pp10[114],pp10[115],pp10[116]};
    assign in450_2 = {pp31[92],pp11[113],pp11[114],pp11[115]};
    CLA_4 KS_450(s450, c450, in450_1, in450_2);
    wire[3:0] s451, in451_1, in451_2;
    wire c451;
    assign in451_1 = {pp32[91],pp12[112],pp12[113],pp12[114]};
    assign in451_2 = {pp33[90],pp13[111],pp13[112],pp13[113]};
    CLA_4 KS_451(s451, c451, in451_1, in451_2);
    wire[3:0] s452, in452_1, in452_2;
    wire c452;
    assign in452_1 = {pp34[89],pp14[110],pp14[111],pp14[112]};
    assign in452_2 = {pp35[88],pp15[109],pp15[110],pp15[111]};
    CLA_4 KS_452(s452, c452, in452_1, in452_2);
    wire[3:0] s453, in453_1, in453_2;
    wire c453;
    assign in453_1 = {pp36[87],pp16[108],pp16[109],pp16[110]};
    assign in453_2 = {pp37[86],pp17[107],pp17[108],pp17[109]};
    CLA_4 KS_453(s453, c453, in453_1, in453_2);
    wire[3:0] s454, in454_1, in454_2;
    wire c454;
    assign in454_1 = {pp38[85],pp18[106],pp18[107],pp18[108]};
    assign in454_2 = {pp39[84],pp19[105],pp19[106],pp19[107]};
    CLA_4 KS_454(s454, c454, in454_1, in454_2);
    wire[3:0] s455, in455_1, in455_2;
    wire c455;
    assign in455_1 = {pp40[83],pp20[104],pp20[105],pp20[106]};
    assign in455_2 = {pp41[82],pp21[103],pp21[104],pp21[105]};
    CLA_4 KS_455(s455, c455, in455_1, in455_2);
    wire[3:0] s456, in456_1, in456_2;
    wire c456;
    assign in456_1 = {pp42[81],pp22[102],pp22[103],pp22[104]};
    assign in456_2 = {pp43[80],pp23[101],pp23[102],pp23[103]};
    CLA_4 KS_456(s456, c456, in456_1, in456_2);
    wire[3:0] s457, in457_1, in457_2;
    wire c457;
    assign in457_1 = {pp44[79],pp24[100],pp24[101],pp24[102]};
    assign in457_2 = {pp45[78],pp25[99],pp25[100],pp25[101]};
    CLA_4 KS_457(s457, c457, in457_1, in457_2);
    wire[3:0] s458, in458_1, in458_2;
    wire c458;
    assign in458_1 = {pp46[77],pp26[98],pp26[99],pp26[100]};
    assign in458_2 = {pp47[76],pp27[97],pp27[98],pp27[99]};
    CLA_4 KS_458(s458, c458, in458_1, in458_2);
    wire[3:0] s459, in459_1, in459_2;
    wire c459;
    assign in459_1 = {pp48[75],pp28[96],pp28[97],pp28[98]};
    assign in459_2 = {pp49[74],pp29[95],pp29[96],pp29[97]};
    CLA_4 KS_459(s459, c459, in459_1, in459_2);
    wire[3:0] s460, in460_1, in460_2;
    wire c460;
    assign in460_1 = {pp50[73],pp30[94],pp30[95],pp30[96]};
    assign in460_2 = {pp51[72],pp31[93],pp31[94],pp31[95]};
    CLA_4 KS_460(s460, c460, in460_1, in460_2);
    wire[3:0] s461, in461_1, in461_2;
    wire c461;
    assign in461_1 = {pp52[71],pp32[92],pp32[93],pp32[94]};
    assign in461_2 = {pp53[70],pp33[91],pp33[92],pp33[93]};
    CLA_4 KS_461(s461, c461, in461_1, in461_2);
    wire[3:0] s462, in462_1, in462_2;
    wire c462;
    assign in462_1 = {pp54[69],pp34[90],pp34[91],pp34[92]};
    assign in462_2 = {pp55[68],pp35[89],pp35[90],pp35[91]};
    CLA_4 KS_462(s462, c462, in462_1, in462_2);
    wire[3:0] s463, in463_1, in463_2;
    wire c463;
    assign in463_1 = {pp56[67],pp36[88],pp36[89],pp36[90]};
    assign in463_2 = {pp57[66],pp37[87],pp37[88],pp37[89]};
    CLA_4 KS_463(s463, c463, in463_1, in463_2);
    wire[3:0] s464, in464_1, in464_2;
    wire c464;
    assign in464_1 = {pp58[65],pp38[86],pp38[87],pp38[88]};
    assign in464_2 = {pp59[64],pp39[85],pp39[86],pp39[87]};
    CLA_4 KS_464(s464, c464, in464_1, in464_2);
    wire[3:0] s465, in465_1, in465_2;
    wire c465;
    assign in465_1 = {pp60[63],pp40[84],pp40[85],pp40[86]};
    assign in465_2 = {pp61[62],pp41[83],pp41[84],pp41[85]};
    CLA_4 KS_465(s465, c465, in465_1, in465_2);
    wire[3:0] s466, in466_1, in466_2;
    wire c466;
    assign in466_1 = {pp62[61],pp42[82],pp42[83],pp42[84]};
    assign in466_2 = {pp63[60],pp43[81],pp43[82],pp43[83]};
    CLA_4 KS_466(s466, c466, in466_1, in466_2);
    wire[3:0] s467, in467_1, in467_2;
    wire c467;
    assign in467_1 = {pp64[59],pp44[80],pp44[81],pp44[82]};
    assign in467_2 = {pp65[58],pp45[79],pp45[80],pp45[81]};
    CLA_4 KS_467(s467, c467, in467_1, in467_2);
    wire[3:0] s468, in468_1, in468_2;
    wire c468;
    assign in468_1 = {pp66[57],pp46[78],pp46[79],pp46[80]};
    assign in468_2 = {pp67[56],pp47[77],pp47[78],pp47[79]};
    CLA_4 KS_468(s468, c468, in468_1, in468_2);
    wire[3:0] s469, in469_1, in469_2;
    wire c469;
    assign in469_1 = {pp68[55],pp48[76],pp48[77],pp48[78]};
    assign in469_2 = {pp69[54],pp49[75],pp49[76],pp49[77]};
    CLA_4 KS_469(s469, c469, in469_1, in469_2);
    wire[3:0] s470, in470_1, in470_2;
    wire c470;
    assign in470_1 = {pp70[53],pp50[74],pp50[75],pp50[76]};
    assign in470_2 = {pp71[52],pp51[73],pp51[74],pp51[75]};
    CLA_4 KS_470(s470, c470, in470_1, in470_2);
    wire[3:0] s471, in471_1, in471_2;
    wire c471;
    assign in471_1 = {pp72[51],pp52[72],pp52[73],pp52[74]};
    assign in471_2 = {pp73[50],pp53[71],pp53[72],pp53[73]};
    CLA_4 KS_471(s471, c471, in471_1, in471_2);
    wire[3:0] s472, in472_1, in472_2;
    wire c472;
    assign in472_1 = {pp74[49],pp54[70],pp54[71],pp54[72]};
    assign in472_2 = {pp75[48],pp55[69],pp55[70],pp55[71]};
    CLA_4 KS_472(s472, c472, in472_1, in472_2);
    wire[3:0] s473, in473_1, in473_2;
    wire c473;
    assign in473_1 = {pp76[47],pp56[68],pp56[69],pp56[70]};
    assign in473_2 = {pp77[46],pp57[67],pp57[68],pp57[69]};
    CLA_4 KS_473(s473, c473, in473_1, in473_2);
    wire[3:0] s474, in474_1, in474_2;
    wire c474;
    assign in474_1 = {pp78[45],pp58[66],pp58[67],pp58[68]};
    assign in474_2 = {pp79[44],pp59[65],pp59[66],pp59[67]};
    CLA_4 KS_474(s474, c474, in474_1, in474_2);
    wire[3:0] s475, in475_1, in475_2;
    wire c475;
    assign in475_1 = {pp80[43],pp60[64],pp60[65],pp60[66]};
    assign in475_2 = {pp81[42],pp61[63],pp61[64],pp61[65]};
    CLA_4 KS_475(s475, c475, in475_1, in475_2);
    wire[3:0] s476, in476_1, in476_2;
    wire c476;
    assign in476_1 = {pp82[41],pp62[62],pp62[63],pp62[64]};
    assign in476_2 = {pp83[40],pp63[61],pp63[62],pp63[63]};
    CLA_4 KS_476(s476, c476, in476_1, in476_2);
    wire[3:0] s477, in477_1, in477_2;
    wire c477;
    assign in477_1 = {pp84[39],pp64[60],pp64[61],pp64[62]};
    assign in477_2 = {pp85[38],pp65[59],pp65[60],pp65[61]};
    CLA_4 KS_477(s477, c477, in477_1, in477_2);
    wire[3:0] s478, in478_1, in478_2;
    wire c478;
    assign in478_1 = {pp86[37],pp66[58],pp66[59],pp66[60]};
    assign in478_2 = {pp87[36],pp67[57],pp67[58],pp67[59]};
    CLA_4 KS_478(s478, c478, in478_1, in478_2);
    wire[3:0] s479, in479_1, in479_2;
    wire c479;
    assign in479_1 = {pp88[35],pp68[56],pp68[57],pp68[58]};
    assign in479_2 = {pp89[34],pp69[55],pp69[56],pp69[57]};
    CLA_4 KS_479(s479, c479, in479_1, in479_2);
    wire[3:0] s480, in480_1, in480_2;
    wire c480;
    assign in480_1 = {pp90[33],pp70[54],pp70[55],pp70[56]};
    assign in480_2 = {pp91[32],pp71[53],pp71[54],pp71[55]};
    CLA_4 KS_480(s480, c480, in480_1, in480_2);
    wire[3:0] s481, in481_1, in481_2;
    wire c481;
    assign in481_1 = {pp92[31],pp72[52],pp72[53],pp72[54]};
    assign in481_2 = {pp93[30],pp73[51],pp73[52],pp73[53]};
    CLA_4 KS_481(s481, c481, in481_1, in481_2);
    wire[3:0] s482, in482_1, in482_2;
    wire c482;
    assign in482_1 = {pp94[29],pp74[50],pp74[51],pp74[52]};
    assign in482_2 = {pp95[28],pp75[49],pp75[50],pp75[51]};
    CLA_4 KS_482(s482, c482, in482_1, in482_2);
    wire[3:0] s483, in483_1, in483_2;
    wire c483;
    assign in483_1 = {pp96[27],pp76[48],pp76[49],pp76[50]};
    assign in483_2 = {pp97[26],pp77[47],pp77[48],pp77[49]};
    CLA_4 KS_483(s483, c483, in483_1, in483_2);
    wire[3:0] s484, in484_1, in484_2;
    wire c484;
    assign in484_1 = {pp98[25],pp78[46],pp78[47],pp78[48]};
    assign in484_2 = {pp99[24],pp79[45],pp79[46],pp79[47]};
    CLA_4 KS_484(s484, c484, in484_1, in484_2);
    wire[3:0] s485, in485_1, in485_2;
    wire c485;
    assign in485_1 = {pp100[23],pp80[44],pp80[45],pp80[46]};
    assign in485_2 = {pp101[22],pp81[43],pp81[44],pp81[45]};
    CLA_4 KS_485(s485, c485, in485_1, in485_2);
    wire[3:0] s486, in486_1, in486_2;
    wire c486;
    assign in486_1 = {pp102[21],pp82[42],pp82[43],pp82[44]};
    assign in486_2 = {pp103[20],pp83[41],pp83[42],pp83[43]};
    CLA_4 KS_486(s486, c486, in486_1, in486_2);
    wire[3:0] s487, in487_1, in487_2;
    wire c487;
    assign in487_1 = {pp104[19],pp84[40],pp84[41],pp84[42]};
    assign in487_2 = {pp105[18],pp85[39],pp85[40],pp85[41]};
    CLA_4 KS_487(s487, c487, in487_1, in487_2);
    wire[3:0] s488, in488_1, in488_2;
    wire c488;
    assign in488_1 = {pp106[17],pp86[38],pp86[39],pp86[40]};
    assign in488_2 = {pp107[16],pp87[37],pp87[38],pp87[39]};
    CLA_4 KS_488(s488, c488, in488_1, in488_2);
    wire[3:0] s489, in489_1, in489_2;
    wire c489;
    assign in489_1 = {pp108[15],pp88[36],pp88[37],pp88[38]};
    assign in489_2 = {pp109[14],pp89[35],pp89[36],pp89[37]};
    CLA_4 KS_489(s489, c489, in489_1, in489_2);
    wire[3:0] s490, in490_1, in490_2;
    wire c490;
    assign in490_1 = {pp110[13],pp90[34],pp90[35],pp90[36]};
    assign in490_2 = {pp111[12],pp91[33],pp91[34],pp91[35]};
    CLA_4 KS_490(s490, c490, in490_1, in490_2);
    wire[3:0] s491, in491_1, in491_2;
    wire c491;
    assign in491_1 = {pp112[11],pp92[32],pp92[33],pp92[34]};
    assign in491_2 = {pp113[10],pp93[31],pp93[32],pp93[33]};
    CLA_4 KS_491(s491, c491, in491_1, in491_2);
    wire[3:0] s492, in492_1, in492_2;
    wire c492;
    assign in492_1 = {pp114[9],pp94[30],pp94[31],pp94[32]};
    assign in492_2 = {pp115[8],pp95[29],pp95[30],pp95[31]};
    CLA_4 KS_492(s492, c492, in492_1, in492_2);
    wire[3:0] s493, in493_1, in493_2;
    wire c493;
    assign in493_1 = {pp116[7],pp96[28],pp96[29],pp96[30]};
    assign in493_2 = {pp117[6],pp97[27],pp97[28],pp97[29]};
    CLA_4 KS_493(s493, c493, in493_1, in493_2);
    wire[3:0] s494, in494_1, in494_2;
    wire c494;
    assign in494_1 = {pp118[5],pp98[26],pp98[27],pp98[28]};
    assign in494_2 = {pp119[4],pp99[25],pp99[26],pp99[27]};
    CLA_4 KS_494(s494, c494, in494_1, in494_2);
    wire[3:0] s495, in495_1, in495_2;
    wire c495;
    assign in495_1 = {pp120[3],pp100[24],pp100[25],pp100[26]};
    assign in495_2 = {pp121[2],pp101[23],pp101[24],pp101[25]};
    CLA_4 KS_495(s495, c495, in495_1, in495_2);
    wire[1:0] s496, in496_1, in496_2;
    wire c496;
    assign in496_1 = {pp122[1],pp102[22]};
    assign in496_2 = {pp123[0],pp103[21]};
    CLA_2 KS_496(s496, c496, in496_1, in496_2);
    wire[3:0] s497, in497_1, in497_2;
    wire c497;
    assign in497_1 = {c376,pp104[20],pp102[23],pp102[24]};
    assign in497_2 = {c377,pp105[19],pp103[22],pp103[23]};
    CLA_4 KS_497(s497, c497, in497_1, in497_2);
    wire[1:0] s498, in498_1, in498_2;
    wire c498;
    assign in498_1 = {c378,pp106[18]};
    assign in498_2 = {c379,pp107[17]};
    CLA_2 KS_498(s498, c498, in498_1, in498_2);
    wire[2:0] s499, in499_1, in499_2;
    wire c499;
    assign in499_1 = {c380,pp108[16],pp104[21]};
    assign in499_2 = {c381,pp109[15],pp105[20]};
    CLA_3 KS_499(s499, c499, in499_1, in499_2);
    wire[1:0] s500, in500_1, in500_2;
    wire c500;
    assign in500_1 = {c382,pp110[14]};
    assign in500_2 = {c383,pp111[13]};
    CLA_2 KS_500(s500, c500, in500_1, in500_2);
    wire[3:0] s501, in501_1, in501_2;
    wire c501;
    assign in501_1 = {c384,pp112[12],pp106[19],pp104[22]};
    assign in501_2 = {c385,pp113[11],pp107[18],pp105[21]};
    CLA_4 KS_501(s501, c501, in501_1, in501_2);
    wire[1:0] s502, in502_1, in502_2;
    wire c502;
    assign in502_1 = {c386,pp114[10]};
    assign in502_2 = {c387,pp115[9]};
    CLA_2 KS_502(s502, c502, in502_1, in502_2);
    wire[2:0] s503, in503_1, in503_2;
    wire c503;
    assign in503_1 = {c388,pp116[8],pp108[17]};
    assign in503_2 = {c389,pp117[7],pp109[16]};
    CLA_3 KS_503(s503, c503, in503_1, in503_2);
    wire[1:0] s504, in504_1, in504_2;
    wire c504;
    assign in504_1 = {c390,pp118[6]};
    assign in504_2 = {c391,pp119[5]};
    CLA_2 KS_504(s504, c504, in504_1, in504_2);
    wire[0:0] s505, in505_1, in505_2;
    wire c505;
    assign in505_1 = {c392};
    assign in505_2 = {c393};
    Half_Adder KS_505(s505, c505, in505_1, in505_2);
    wire[3:0] s506, in506_1, in506_2;
    wire c506;
    assign in506_1 = {c394,pp120[4],pp110[15],pp106[20]};
    assign in506_2 = {c395,pp121[3],pp111[14],pp107[19]};
    CLA_4 KS_506(s506, c506, in506_1, in506_2);
    wire[0:0] s507, in507_1, in507_2;
    wire c507;
    assign in507_1 = {c396};
    assign in507_2 = {c397};
    Half_Adder KS_507(s507, c507, in507_1, in507_2);
    wire[1:0] s508, in508_1, in508_2;
    wire c508;
    assign in508_1 = {c398,pp122[2]};
    assign in508_2 = {c399,pp123[1]};
    CLA_2 KS_508(s508, c508, in508_1, in508_2);
    wire[0:0] s509, in509_1, in509_2;
    wire c509;
    assign in509_1 = {c400};
    assign in509_2 = {c401};
    Half_Adder KS_509(s509, c509, in509_1, in509_2);
    wire[2:0] s510, in510_1, in510_2;
    wire c510;
    assign in510_1 = {c402,pp124[0],pp112[13]};
    assign in510_2 = {c403,c419,pp113[12]};
    CLA_3 KS_510(s510, c510, in510_1, in510_2);
    wire[0:0] s511, in511_1, in511_2;
    wire c511;
    assign in511_1 = {c404};
    assign in511_2 = {c405};
    Half_Adder KS_511(s511, c511, in511_1, in511_2);
    wire[1:0] s512, in512_1, in512_2;
    wire c512;
    assign in512_1 = {c406,c420};
    assign in512_2 = {c407,c421};
    CLA_2 KS_512(s512, c512, in512_1, in512_2);
    wire[0:0] s513, in513_1, in513_2;
    wire c513;
    assign in513_1 = {c408};
    assign in513_2 = {c409};
    Half_Adder KS_513(s513, c513, in513_1, in513_2);
    wire[3:0] s514, in514_1, in514_2;
    wire c514;
    assign in514_1 = {c410,c422,pp114[11],pp108[18]};
    assign in514_2 = {c411,c424,pp115[10],pp109[17]};
    CLA_4 KS_514(s514, c514, in514_1, in514_2);
    wire[0:0] s515, in515_1, in515_2;
    wire c515;
    assign in515_1 = {c412};
    assign in515_2 = {c413};
    Half_Adder KS_515(s515, c515, in515_1, in515_2);
    wire[1:0] s516, in516_1, in516_2;
    wire c516;
    assign in516_1 = {c414,c428};
    assign in516_2 = {c415,c432};
    CLA_2 KS_516(s516, c516, in516_1, in516_2);
    wire[0:0] s517, in517_1, in517_2;
    wire c517;
    assign in517_1 = {c416};
    assign in517_2 = {c417};
    Half_Adder KS_517(s517, c517, in517_1, in517_2);
    wire[2:0] s518, in518_1, in518_2;
    wire c518;
    assign in518_1 = {c418,c436,pp116[9]};
    assign in518_2 = {s419[3],c440,pp117[8]};
    CLA_3 KS_518(s518, c518, in518_1, in518_2);
    wire[0:0] s519, in519_1, in519_2;
    wire c519;
    assign in519_1 = {s420[3]};
    assign in519_2 = {s421[3]};
    Half_Adder KS_519(s519, c519, in519_1, in519_2);
    wire[1:0] s520, in520_1, in520_2;
    wire c520;
    assign in520_1 = {s422[3],c444};
    assign in520_2 = {s424[3],s445[1]};
    CLA_2 KS_520(s520, c520, in520_1, in520_2);
    wire[0:0] s521, in521_1, in521_2;
    wire c521;
    assign in521_1 = {s428[3]};
    assign in521_2 = {s432[3]};
    Half_Adder KS_521(s521, c521, in521_1, in521_2);
    wire[3:0] s522, in522_1, in522_2;
    wire c522;
    assign in522_1 = {s436[3],s446[1],pp118[7],pp110[16]};
    assign in522_2 = {s440[3],s447[1],pp119[6],pp111[15]};
    CLA_4 KS_522(s522, c522, in522_1, in522_2);
    wire[0:0] s523, in523_1, in523_2;
    wire c523;
    assign in523_1 = {s444[3]};
    assign in523_2 = {s445[0]};
    Half_Adder KS_523(s523, c523, in523_1, in523_2);
    wire[1:0] s524, in524_1, in524_2;
    wire c524;
    assign in524_1 = {s447[0],s448[1]};
    assign in524_2 = {s448[0],s449[1]};
    CLA_2_c KS_524(s524, c524, in524_1, in524_2, s446[0]);
    wire[3:0] s525, in525_1, in525_2;
    wire c525;
    assign in525_1 = {pp0[127],pp1[127],pp2[127],pp3[127]};
    assign in525_2 = {pp1[126],pp2[126],pp3[126],pp4[126]};
    CLA_4 KS_525(s525, c525, in525_1, in525_2);
    wire[3:0] s526, in526_1, in526_2;
    wire c526;
    assign in526_1 = {pp2[125],pp3[125],pp4[125],pp5[125]};
    assign in526_2 = {pp3[124],pp4[124],pp5[124],pp6[124]};
    CLA_4 KS_526(s526, c526, in526_1, in526_2);
    wire[3:0] s527, in527_1, in527_2;
    wire c527;
    assign in527_1 = {pp4[123],pp5[123],pp6[123],pp7[123]};
    assign in527_2 = {pp5[122],pp6[122],pp7[122],pp8[122]};
    CLA_4 KS_527(s527, c527, in527_1, in527_2);
    wire[3:0] s528, in528_1, in528_2;
    wire c528;
    assign in528_1 = {pp6[121],pp7[121],pp8[121],pp9[121]};
    assign in528_2 = {pp7[120],pp8[120],pp9[120],pp10[120]};
    CLA_4 KS_528(s528, c528, in528_1, in528_2);
    wire[3:0] s529, in529_1, in529_2;
    wire c529;
    assign in529_1 = {pp8[119],pp9[119],pp10[119],pp11[119]};
    assign in529_2 = {pp9[118],pp10[118],pp11[118],pp12[118]};
    CLA_4 KS_529(s529, c529, in529_1, in529_2);
    wire[3:0] s530, in530_1, in530_2;
    wire c530;
    assign in530_1 = {pp10[117],pp11[117],pp12[117],pp13[117]};
    assign in530_2 = {pp11[116],pp12[116],pp13[116],pp14[116]};
    CLA_4 KS_530(s530, c530, in530_1, in530_2);
    wire[3:0] s531, in531_1, in531_2;
    wire c531;
    assign in531_1 = {pp12[115],pp13[115],pp14[115],pp15[115]};
    assign in531_2 = {pp13[114],pp14[114],pp15[114],pp16[114]};
    CLA_4 KS_531(s531, c531, in531_1, in531_2);
    wire[3:0] s532, in532_1, in532_2;
    wire c532;
    assign in532_1 = {pp14[113],pp15[113],pp16[113],pp17[113]};
    assign in532_2 = {pp15[112],pp16[112],pp17[112],pp18[112]};
    CLA_4 KS_532(s532, c532, in532_1, in532_2);
    wire[3:0] s533, in533_1, in533_2;
    wire c533;
    assign in533_1 = {pp16[111],pp17[111],pp18[111],pp19[111]};
    assign in533_2 = {pp17[110],pp18[110],pp19[110],pp20[110]};
    CLA_4 KS_533(s533, c533, in533_1, in533_2);
    wire[3:0] s534, in534_1, in534_2;
    wire c534;
    assign in534_1 = {pp18[109],pp19[109],pp20[109],pp21[109]};
    assign in534_2 = {pp19[108],pp20[108],pp21[108],pp22[108]};
    CLA_4 KS_534(s534, c534, in534_1, in534_2);
    wire[3:0] s535, in535_1, in535_2;
    wire c535;
    assign in535_1 = {pp20[107],pp21[107],pp22[107],pp23[107]};
    assign in535_2 = {pp21[106],pp22[106],pp23[106],pp24[106]};
    CLA_4 KS_535(s535, c535, in535_1, in535_2);
    wire[3:0] s536, in536_1, in536_2;
    wire c536;
    assign in536_1 = {pp22[105],pp23[105],pp24[105],pp25[105]};
    assign in536_2 = {pp23[104],pp24[104],pp25[104],pp26[104]};
    CLA_4 KS_536(s536, c536, in536_1, in536_2);
    wire[3:0] s537, in537_1, in537_2;
    wire c537;
    assign in537_1 = {pp24[103],pp25[103],pp26[103],pp27[103]};
    assign in537_2 = {pp25[102],pp26[102],pp27[102],pp28[102]};
    CLA_4 KS_537(s537, c537, in537_1, in537_2);
    wire[3:0] s538, in538_1, in538_2;
    wire c538;
    assign in538_1 = {pp26[101],pp27[101],pp28[101],pp29[101]};
    assign in538_2 = {pp27[100],pp28[100],pp29[100],pp30[100]};
    CLA_4 KS_538(s538, c538, in538_1, in538_2);
    wire[3:0] s539, in539_1, in539_2;
    wire c539;
    assign in539_1 = {pp28[99],pp29[99],pp30[99],pp31[99]};
    assign in539_2 = {pp29[98],pp30[98],pp31[98],pp32[98]};
    CLA_4 KS_539(s539, c539, in539_1, in539_2);
    wire[3:0] s540, in540_1, in540_2;
    wire c540;
    assign in540_1 = {pp30[97],pp31[97],pp32[97],pp33[97]};
    assign in540_2 = {pp31[96],pp32[96],pp33[96],pp34[96]};
    CLA_4 KS_540(s540, c540, in540_1, in540_2);
    wire[3:0] s541, in541_1, in541_2;
    wire c541;
    assign in541_1 = {pp32[95],pp33[95],pp34[95],pp35[95]};
    assign in541_2 = {pp33[94],pp34[94],pp35[94],pp36[94]};
    CLA_4 KS_541(s541, c541, in541_1, in541_2);
    wire[3:0] s542, in542_1, in542_2;
    wire c542;
    assign in542_1 = {pp34[93],pp35[93],pp36[93],pp37[93]};
    assign in542_2 = {pp35[92],pp36[92],pp37[92],pp38[92]};
    CLA_4 KS_542(s542, c542, in542_1, in542_2);
    wire[3:0] s543, in543_1, in543_2;
    wire c543;
    assign in543_1 = {pp36[91],pp37[91],pp38[91],pp39[91]};
    assign in543_2 = {pp37[90],pp38[90],pp39[90],pp40[90]};
    CLA_4 KS_543(s543, c543, in543_1, in543_2);
    wire[3:0] s544, in544_1, in544_2;
    wire c544;
    assign in544_1 = {pp38[89],pp39[89],pp40[89],pp41[89]};
    assign in544_2 = {pp39[88],pp40[88],pp41[88],pp42[88]};
    CLA_4 KS_544(s544, c544, in544_1, in544_2);
    wire[3:0] s545, in545_1, in545_2;
    wire c545;
    assign in545_1 = {pp40[87],pp41[87],pp42[87],pp43[87]};
    assign in545_2 = {pp41[86],pp42[86],pp43[86],pp44[86]};
    CLA_4 KS_545(s545, c545, in545_1, in545_2);
    wire[3:0] s546, in546_1, in546_2;
    wire c546;
    assign in546_1 = {pp42[85],pp43[85],pp44[85],pp45[85]};
    assign in546_2 = {pp43[84],pp44[84],pp45[84],pp46[84]};
    CLA_4 KS_546(s546, c546, in546_1, in546_2);
    wire[3:0] s547, in547_1, in547_2;
    wire c547;
    assign in547_1 = {pp44[83],pp45[83],pp46[83],pp47[83]};
    assign in547_2 = {pp45[82],pp46[82],pp47[82],pp48[82]};
    CLA_4 KS_547(s547, c547, in547_1, in547_2);
    wire[3:0] s548, in548_1, in548_2;
    wire c548;
    assign in548_1 = {pp46[81],pp47[81],pp48[81],pp49[81]};
    assign in548_2 = {pp47[80],pp48[80],pp49[80],pp50[80]};
    CLA_4 KS_548(s548, c548, in548_1, in548_2);
    wire[3:0] s549, in549_1, in549_2;
    wire c549;
    assign in549_1 = {pp48[79],pp49[79],pp50[79],pp51[79]};
    assign in549_2 = {pp49[78],pp50[78],pp51[78],pp52[78]};
    CLA_4 KS_549(s549, c549, in549_1, in549_2);
    wire[3:0] s550, in550_1, in550_2;
    wire c550;
    assign in550_1 = {pp50[77],pp51[77],pp52[77],pp53[77]};
    assign in550_2 = {pp51[76],pp52[76],pp53[76],pp54[76]};
    CLA_4 KS_550(s550, c550, in550_1, in550_2);
    wire[3:0] s551, in551_1, in551_2;
    wire c551;
    assign in551_1 = {pp52[75],pp53[75],pp54[75],pp55[75]};
    assign in551_2 = {pp53[74],pp54[74],pp55[74],pp56[74]};
    CLA_4 KS_551(s551, c551, in551_1, in551_2);
    wire[3:0] s552, in552_1, in552_2;
    wire c552;
    assign in552_1 = {pp54[73],pp55[73],pp56[73],pp57[73]};
    assign in552_2 = {pp55[72],pp56[72],pp57[72],pp58[72]};
    CLA_4 KS_552(s552, c552, in552_1, in552_2);
    wire[3:0] s553, in553_1, in553_2;
    wire c553;
    assign in553_1 = {pp56[71],pp57[71],pp58[71],pp59[71]};
    assign in553_2 = {pp57[70],pp58[70],pp59[70],pp60[70]};
    CLA_4 KS_553(s553, c553, in553_1, in553_2);
    wire[3:0] s554, in554_1, in554_2;
    wire c554;
    assign in554_1 = {pp58[69],pp59[69],pp60[69],pp61[69]};
    assign in554_2 = {pp59[68],pp60[68],pp61[68],pp62[68]};
    CLA_4 KS_554(s554, c554, in554_1, in554_2);
    wire[3:0] s555, in555_1, in555_2;
    wire c555;
    assign in555_1 = {pp60[67],pp61[67],pp62[67],pp63[67]};
    assign in555_2 = {pp61[66],pp62[66],pp63[66],pp64[66]};
    CLA_4 KS_555(s555, c555, in555_1, in555_2);
    wire[3:0] s556, in556_1, in556_2;
    wire c556;
    assign in556_1 = {pp62[65],pp63[65],pp64[65],pp65[65]};
    assign in556_2 = {pp63[64],pp64[64],pp65[64],pp66[64]};
    CLA_4 KS_556(s556, c556, in556_1, in556_2);
    wire[3:0] s557, in557_1, in557_2;
    wire c557;
    assign in557_1 = {pp64[63],pp65[63],pp66[63],pp67[63]};
    assign in557_2 = {pp65[62],pp66[62],pp67[62],pp68[62]};
    CLA_4 KS_557(s557, c557, in557_1, in557_2);
    wire[3:0] s558, in558_1, in558_2;
    wire c558;
    assign in558_1 = {pp66[61],pp67[61],pp68[61],pp69[61]};
    assign in558_2 = {pp67[60],pp68[60],pp69[60],pp70[60]};
    CLA_4 KS_558(s558, c558, in558_1, in558_2);
    wire[3:0] s559, in559_1, in559_2;
    wire c559;
    assign in559_1 = {pp68[59],pp69[59],pp70[59],pp71[59]};
    assign in559_2 = {pp69[58],pp70[58],pp71[58],pp72[58]};
    CLA_4 KS_559(s559, c559, in559_1, in559_2);
    wire[3:0] s560, in560_1, in560_2;
    wire c560;
    assign in560_1 = {pp70[57],pp71[57],pp72[57],pp73[57]};
    assign in560_2 = {pp71[56],pp72[56],pp73[56],pp74[56]};
    CLA_4 KS_560(s560, c560, in560_1, in560_2);
    wire[3:0] s561, in561_1, in561_2;
    wire c561;
    assign in561_1 = {pp72[55],pp73[55],pp74[55],pp75[55]};
    assign in561_2 = {pp73[54],pp74[54],pp75[54],pp76[54]};
    CLA_4 KS_561(s561, c561, in561_1, in561_2);
    wire[3:0] s562, in562_1, in562_2;
    wire c562;
    assign in562_1 = {pp74[53],pp75[53],pp76[53],pp77[53]};
    assign in562_2 = {pp75[52],pp76[52],pp77[52],pp78[52]};
    CLA_4 KS_562(s562, c562, in562_1, in562_2);
    wire[3:0] s563, in563_1, in563_2;
    wire c563;
    assign in563_1 = {pp76[51],pp77[51],pp78[51],pp79[51]};
    assign in563_2 = {pp77[50],pp78[50],pp79[50],pp80[50]};
    CLA_4 KS_563(s563, c563, in563_1, in563_2);
    wire[3:0] s564, in564_1, in564_2;
    wire c564;
    assign in564_1 = {pp78[49],pp79[49],pp80[49],pp81[49]};
    assign in564_2 = {pp79[48],pp80[48],pp81[48],pp82[48]};
    CLA_4 KS_564(s564, c564, in564_1, in564_2);
    wire[3:0] s565, in565_1, in565_2;
    wire c565;
    assign in565_1 = {pp80[47],pp81[47],pp82[47],pp83[47]};
    assign in565_2 = {pp81[46],pp82[46],pp83[46],pp84[46]};
    CLA_4 KS_565(s565, c565, in565_1, in565_2);
    wire[3:0] s566, in566_1, in566_2;
    wire c566;
    assign in566_1 = {pp82[45],pp83[45],pp84[45],pp85[45]};
    assign in566_2 = {pp83[44],pp84[44],pp85[44],pp86[44]};
    CLA_4 KS_566(s566, c566, in566_1, in566_2);
    wire[3:0] s567, in567_1, in567_2;
    wire c567;
    assign in567_1 = {pp84[43],pp85[43],pp86[43],pp87[43]};
    assign in567_2 = {pp85[42],pp86[42],pp87[42],pp88[42]};
    CLA_4 KS_567(s567, c567, in567_1, in567_2);
    wire[3:0] s568, in568_1, in568_2;
    wire c568;
    assign in568_1 = {pp86[41],pp87[41],pp88[41],pp89[41]};
    assign in568_2 = {pp87[40],pp88[40],pp89[40],pp90[40]};
    CLA_4 KS_568(s568, c568, in568_1, in568_2);
    wire[3:0] s569, in569_1, in569_2;
    wire c569;
    assign in569_1 = {pp88[39],pp89[39],pp90[39],pp91[39]};
    assign in569_2 = {pp89[38],pp90[38],pp91[38],pp92[38]};
    CLA_4 KS_569(s569, c569, in569_1, in569_2);
    wire[3:0] s570, in570_1, in570_2;
    wire c570;
    assign in570_1 = {pp90[37],pp91[37],pp92[37],pp93[37]};
    assign in570_2 = {pp91[36],pp92[36],pp93[36],pp94[36]};
    CLA_4 KS_570(s570, c570, in570_1, in570_2);
    wire[3:0] s571, in571_1, in571_2;
    wire c571;
    assign in571_1 = {pp92[35],pp93[35],pp94[35],pp95[35]};
    assign in571_2 = {pp93[34],pp94[34],pp95[34],pp96[34]};
    CLA_4 KS_571(s571, c571, in571_1, in571_2);
    wire[3:0] s572, in572_1, in572_2;
    wire c572;
    assign in572_1 = {pp94[33],pp95[33],pp96[33],pp97[33]};
    assign in572_2 = {pp95[32],pp96[32],pp97[32],pp98[32]};
    CLA_4 KS_572(s572, c572, in572_1, in572_2);
    wire[3:0] s573, in573_1, in573_2;
    wire c573;
    assign in573_1 = {pp96[31],pp97[31],pp98[31],pp99[31]};
    assign in573_2 = {pp97[30],pp98[30],pp99[30],pp100[30]};
    CLA_4 KS_573(s573, c573, in573_1, in573_2);
    wire[3:0] s574, in574_1, in574_2;
    wire c574;
    assign in574_1 = {pp98[29],pp99[29],pp100[29],pp101[29]};
    assign in574_2 = {pp99[28],pp100[28],pp101[28],pp102[28]};
    CLA_4 KS_574(s574, c574, in574_1, in574_2);
    wire[2:0] s575, in575_1, in575_2;
    wire c575;
    assign in575_1 = {pp100[27],pp101[27],pp102[27]};
    assign in575_2 = {pp101[26],pp102[26],pp103[26]};
    CLA_3 KS_575(s575, c575, in575_1, in575_2);
    wire[1:0] s576, in576_1, in576_2;
    wire c576;
    assign in576_1 = {pp102[25],pp103[25]};
    assign in576_2 = {pp103[24],pp104[24]};
    CLA_2 KS_576(s576, c576, in576_1, in576_2);
    wire[3:0] s577, in577_1, in577_2;
    wire c577;
    assign in577_1 = {pp104[23],pp105[23],pp104[25],pp103[27]};
    assign in577_2 = {pp105[22],pp106[22],pp105[24],pp104[26]};
    CLA_4 KS_577(s577, c577, in577_1, in577_2);
    wire[0:0] s578, in578_1, in578_2;
    wire c578;
    assign in578_1 = {pp106[21]};
    assign in578_2 = {pp107[20]};
    Half_Adder KS_578(s578, c578, in578_1, in578_2);
    wire[1:0] s579, in579_1, in579_2;
    wire c579;
    assign in579_1 = {pp108[19],pp107[21]};
    assign in579_2 = {pp109[18],pp108[20]};
    CLA_2 KS_579(s579, c579, in579_1, in579_2);
    wire[0:0] s580, in580_1, in580_2;
    wire c580;
    assign in580_1 = {pp110[17]};
    assign in580_2 = {pp111[16]};
    Half_Adder KS_580(s580, c580, in580_1, in580_2);
    wire[2:0] s581, in581_1, in581_2;
    wire c581;
    assign in581_1 = {pp112[15],pp109[19],pp106[23]};
    assign in581_2 = {pp113[14],pp110[18],pp107[22]};
    CLA_3 KS_581(s581, c581, in581_1, in581_2);
    wire[0:0] s582, in582_1, in582_2;
    wire c582;
    assign in582_1 = {pp114[13]};
    assign in582_2 = {pp115[12]};
    Half_Adder KS_582(s582, c582, in582_1, in582_2);
    wire[1:0] s583, in583_1, in583_2;
    wire c583;
    assign in583_1 = {pp116[11],pp111[17]};
    assign in583_2 = {pp117[10],pp112[16]};
    CLA_2 KS_583(s583, c583, in583_1, in583_2);
    wire[0:0] s584, in584_1, in584_2;
    wire c584;
    assign in584_1 = {pp118[9]};
    assign in584_2 = {pp119[8]};
    Half_Adder KS_584(s584, c584, in584_1, in584_2);
    wire[3:0] s585, in585_1, in585_2;
    wire c585;
    assign in585_1 = {pp120[7],pp113[15],pp108[21],pp105[25]};
    assign in585_2 = {pp121[6],pp114[14],pp109[20],pp106[24]};
    CLA_4 KS_585(s585, c585, in585_1, in585_2);
    wire[0:0] s586, in586_1, in586_2;
    wire c586;
    assign in586_1 = {pp122[5]};
    assign in586_2 = {pp123[4]};
    Half_Adder KS_586(s586, c586, in586_1, in586_2);
    wire[1:0] s587, in587_1, in587_2;
    wire c587;
    assign in587_1 = {pp124[3],pp115[13]};
    assign in587_2 = {pp125[2],pp116[12]};
    CLA_2 KS_587(s587, c587, in587_1, in587_2);
    wire[0:0] s588, in588_1, in588_2;
    wire c588;
    assign in588_1 = {pp126[1]};
    assign in588_2 = {pp127[0]};
    Half_Adder KS_588(s588, c588, in588_1, in588_2);
    wire[2:0] s589, in589_1, in589_2;
    wire c589;
    assign in589_1 = {c445,pp117[11],pp110[19]};
    assign in589_2 = {c446,pp118[10],pp111[18]};
    CLA_3 KS_589(s589, c589, in589_1, in589_2);
    wire[0:0] s590, in590_1, in590_2;
    wire c590;
    assign in590_1 = {c447};
    assign in590_2 = {c448};
    Half_Adder KS_590(s590, c590, in590_1, in590_2);
    wire[1:0] s591, in591_1, in591_2;
    wire c591;
    assign in591_1 = {c449,pp119[9]};
    assign in591_2 = {c450,pp120[8]};
    CLA_2 KS_591(s591, c591, in591_1, in591_2);
    wire[0:0] s592, in592_1, in592_2;
    wire c592;
    assign in592_1 = {c451};
    assign in592_2 = {c452};
    Half_Adder KS_592(s592, c592, in592_1, in592_2);
    wire[3:0] s593, in593_1, in593_2;
    wire c593;
    assign in593_1 = {c453,pp121[7],pp112[17],pp107[23]};
    assign in593_2 = {c454,pp122[6],pp113[16],pp108[22]};
    CLA_4 KS_593(s593, c593, in593_1, in593_2);
    wire[0:0] s594, in594_1, in594_2;
    wire c594;
    assign in594_1 = {c455};
    assign in594_2 = {c456};
    Half_Adder KS_594(s594, c594, in594_1, in594_2);
    wire[1:0] s595, in595_1, in595_2;
    wire c595;
    assign in595_1 = {c457,pp123[5]};
    assign in595_2 = {c458,pp124[4]};
    CLA_2 KS_595(s595, c595, in595_1, in595_2);
    wire[0:0] s596, in596_1, in596_2;
    wire c596;
    assign in596_1 = {c459};
    assign in596_2 = {c460};
    Half_Adder KS_596(s596, c596, in596_1, in596_2);
    wire[2:0] s597, in597_1, in597_2;
    wire c597;
    assign in597_1 = {c461,pp125[3],pp114[15]};
    assign in597_2 = {c462,pp126[2],pp115[14]};
    CLA_3 KS_597(s597, c597, in597_1, in597_2);
    wire[0:0] s598, in598_1, in598_2;
    wire c598;
    assign in598_1 = {c463};
    assign in598_2 = {c464};
    Half_Adder KS_598(s598, c598, in598_1, in598_2);
    wire[1:0] s599, in599_1, in599_2;
    wire c599;
    assign in599_1 = {c465,pp127[1]};
    assign in599_2 = {c466,1'b0};
    CLA_2 KS_599(s599, c599, in599_1, in599_2);
    wire[0:0] s600, in600_1, in600_2;
    wire c600;
    assign in600_1 = {c467};
    assign in600_2 = {c468};
    Half_Adder KS_600(s600, c600, in600_1, in600_2);
    wire[3:0] s601, in601_1, in601_2;
    wire c601;
    assign in601_1 = {c469,s525[1],pp116[13],pp109[21]};
    assign in601_2 = {c470,s526[1],pp117[12],pp110[20]};
    CLA_4 KS_601(s601, c601, in601_1, in601_2);
    wire[0:0] s602, in602_1, in602_2;
    wire c602;
    assign in602_1 = {c471};
    assign in602_2 = {c472};
    Half_Adder KS_602(s602, c602, in602_1, in602_2);
    wire[1:0] s603, in603_1, in603_2;
    wire c603;
    assign in603_1 = {c473,s527[1]};
    assign in603_2 = {c474,s528[1]};
    CLA_2 KS_603(s603, c603, in603_1, in603_2);
    wire[0:0] s604, in604_1, in604_2;
    wire c604;
    assign in604_1 = {c475};
    assign in604_2 = {c476};
    Half_Adder KS_604(s604, c604, in604_1, in604_2);
    wire[2:0] s605, in605_1, in605_2;
    wire c605;
    assign in605_1 = {c477,s529[1],pp118[11]};
    assign in605_2 = {c478,s530[1],pp119[10]};
    CLA_3 KS_605(s605, c605, in605_1, in605_2);
    wire[0:0] s606, in606_1, in606_2;
    wire c606;
    assign in606_1 = {c479};
    assign in606_2 = {c480};
    Half_Adder KS_606(s606, c606, in606_1, in606_2);
    wire[1:0] s607, in607_1, in607_2;
    wire c607;
    assign in607_1 = {c481,s531[1]};
    assign in607_2 = {c482,s532[1]};
    CLA_2 KS_607(s607, c607, in607_1, in607_2);
    wire[0:0] s608, in608_1, in608_2;
    wire c608;
    assign in608_1 = {c483};
    assign in608_2 = {c484};
    Half_Adder KS_608(s608, c608, in608_1, in608_2);
    wire[3:0] s609, in609_1, in609_2;
    wire c609;
    assign in609_1 = {c485,s533[1],pp120[9],pp111[19]};
    assign in609_2 = {c486,s534[1],pp121[8],pp112[18]};
    CLA_4 KS_609(s609, c609, in609_1, in609_2);
    wire[0:0] s610, in610_1, in610_2;
    wire c610;
    assign in610_1 = {c487};
    assign in610_2 = {c488};
    Half_Adder KS_610(s610, c610, in610_1, in610_2);
    wire[1:0] s611, in611_1, in611_2;
    wire c611;
    assign in611_1 = {c489,s535[1]};
    assign in611_2 = {c490,s536[1]};
    CLA_2 KS_611(s611, c611, in611_1, in611_2);
    wire[0:0] s612, in612_1, in612_2;
    wire c612;
    assign in612_1 = {c491};
    assign in612_2 = {c492};
    Half_Adder KS_612(s612, c612, in612_1, in612_2);
    wire[2:0] s613, in613_1, in613_2;
    wire c613;
    assign in613_1 = {c493,s537[1],pp122[7]};
    assign in613_2 = {c494,s538[1],pp123[6]};
    CLA_3 KS_613(s613, c613, in613_1, in613_2);
    wire[0:0] s614, in614_1, in614_2;
    wire c614;
    assign in614_1 = {c495};
    assign in614_2 = {c497};
    Half_Adder KS_614(s614, c614, in614_1, in614_2);
    wire[1:0] s615, in615_1, in615_2;
    wire c615;
    assign in615_1 = {c501,s539[1]};
    assign in615_2 = {c506,s540[1]};
    CLA_2 KS_615(s615, c615, in615_1, in615_2);
    wire[0:0] s616, in616_1, in616_2;
    wire c616;
    assign in616_1 = {c514};
    assign in616_2 = {c522};
    Half_Adder KS_616(s616, c616, in616_1, in616_2);
    wire[3:0] s617, in617_1, in617_2;
    wire c617;
    assign in617_1 = {s525[0],s541[1],pp124[5],pp113[17]};
    assign in617_2 = {s526[0],s542[1],pp125[4],pp114[16]};
    CLA_4 KS_617(s617, c617, in617_1, in617_2);
    wire[0:0] s618, in618_1, in618_2;
    wire c618;
    assign in618_1 = {s527[0]};
    assign in618_2 = {s528[0]};
    Half_Adder KS_618(s618, c618, in618_1, in618_2);
    wire[1:0] s619, in619_1, in619_2;
    wire c619;
    assign in619_1 = {s529[0],s543[1]};
    assign in619_2 = {s530[0],s544[1]};
    CLA_2 KS_619(s619, c619, in619_1, in619_2);
    wire[0:0] s620, in620_1, in620_2;
    wire c620;
    assign in620_1 = {s531[0]};
    assign in620_2 = {s532[0]};
    Half_Adder KS_620(s620, c620, in620_1, in620_2);
    wire[2:0] s621, in621_1, in621_2;
    wire c621;
    assign in621_1 = {s533[0],s545[1],pp126[3]};
    assign in621_2 = {s534[0],s546[1],pp127[2]};
    CLA_3 KS_621(s621, c621, in621_1, in621_2);
    wire[0:0] s622, in622_1, in622_2;
    wire c622;
    assign in622_1 = {s535[0]};
    assign in622_2 = {s536[0]};
    Half_Adder KS_622(s622, c622, in622_1, in622_2);
    wire[1:0] s623, in623_1, in623_2;
    wire c623;
    assign in623_1 = {s537[0],s547[1]};
    assign in623_2 = {s538[0],s548[1]};
    CLA_2 KS_623(s623, c623, in623_1, in623_2);
    wire[0:0] s624, in624_1, in624_2;
    wire c624;
    assign in624_1 = {s539[0]};
    assign in624_2 = {s540[0]};
    Half_Adder KS_624(s624, c624, in624_1, in624_2);
    wire[3:0] s625, in625_1, in625_2;
    wire c625;
    assign in625_1 = {s541[0],s549[1],s525[2],pp115[15]};
    assign in625_2 = {s542[0],s550[1],s526[2],pp116[14]};
    CLA_4 KS_625(s625, c625, in625_1, in625_2);
    wire[0:0] s626, in626_1, in626_2;
    wire c626;
    assign in626_1 = {s543[0]};
    assign in626_2 = {s544[0]};
    Half_Adder KS_626(s626, c626, in626_1, in626_2);
    wire[1:0] s627, in627_1, in627_2;
    wire c627;
    assign in627_1 = {s545[0],s551[1]};
    assign in627_2 = {s546[0],s552[1]};
    CLA_2 KS_627(s627, c627, in627_1, in627_2);
    wire[0:0] s628, in628_1, in628_2;
    wire c628;
    assign in628_1 = {s547[0]};
    assign in628_2 = {s548[0]};
    Half_Adder KS_628(s628, c628, in628_1, in628_2);
    wire[2:0] s629, in629_1, in629_2;
    wire c629;
    assign in629_1 = {s549[0],s553[1],s527[2]};
    assign in629_2 = {s550[0],s554[1],s528[2]};
    CLA_3 KS_629(s629, c629, in629_1, in629_2);
    wire[0:0] s630, in630_1, in630_2;
    wire c630;
    assign in630_1 = {s551[0]};
    assign in630_2 = {s552[0]};
    Half_Adder KS_630(s630, c630, in630_1, in630_2);
    wire[1:0] s631, in631_1, in631_2;
    wire c631;
    assign in631_1 = {s554[0],s555[1]};
    assign in631_2 = {s555[0],s556[1]};
    CLA_2_c KS_631(s631, c631, in631_1, in631_2, s553[0]);
    wire[3:0] s632, in632_1, in632_2;
    wire c632;
    assign in632_1 = {pp4[127],pp5[127],pp6[127],pp7[127]};
    assign in632_2 = {pp5[126],pp6[126],pp7[126],pp8[126]};
    CLA_4 KS_632(s632, c632, in632_1, in632_2);
    wire[3:0] s633, in633_1, in633_2;
    wire c633;
    assign in633_1 = {pp6[125],pp7[125],pp8[125],pp9[125]};
    assign in633_2 = {pp7[124],pp8[124],pp9[124],pp10[124]};
    CLA_4 KS_633(s633, c633, in633_1, in633_2);
    wire[3:0] s634, in634_1, in634_2;
    wire c634;
    assign in634_1 = {pp8[123],pp9[123],pp10[123],pp11[123]};
    assign in634_2 = {pp9[122],pp10[122],pp11[122],pp12[122]};
    CLA_4 KS_634(s634, c634, in634_1, in634_2);
    wire[3:0] s635, in635_1, in635_2;
    wire c635;
    assign in635_1 = {pp10[121],pp11[121],pp12[121],pp13[121]};
    assign in635_2 = {pp11[120],pp12[120],pp13[120],pp14[120]};
    CLA_4 KS_635(s635, c635, in635_1, in635_2);
    wire[3:0] s636, in636_1, in636_2;
    wire c636;
    assign in636_1 = {pp12[119],pp13[119],pp14[119],pp15[119]};
    assign in636_2 = {pp13[118],pp14[118],pp15[118],pp16[118]};
    CLA_4 KS_636(s636, c636, in636_1, in636_2);
    wire[3:0] s637, in637_1, in637_2;
    wire c637;
    assign in637_1 = {pp14[117],pp15[117],pp16[117],pp17[117]};
    assign in637_2 = {pp15[116],pp16[116],pp17[116],pp18[116]};
    CLA_4 KS_637(s637, c637, in637_1, in637_2);
    wire[3:0] s638, in638_1, in638_2;
    wire c638;
    assign in638_1 = {pp16[115],pp17[115],pp18[115],pp19[115]};
    assign in638_2 = {pp17[114],pp18[114],pp19[114],pp20[114]};
    CLA_4 KS_638(s638, c638, in638_1, in638_2);
    wire[3:0] s639, in639_1, in639_2;
    wire c639;
    assign in639_1 = {pp18[113],pp19[113],pp20[113],pp21[113]};
    assign in639_2 = {pp19[112],pp20[112],pp21[112],pp22[112]};
    CLA_4 KS_639(s639, c639, in639_1, in639_2);
    wire[3:0] s640, in640_1, in640_2;
    wire c640;
    assign in640_1 = {pp20[111],pp21[111],pp22[111],pp23[111]};
    assign in640_2 = {pp21[110],pp22[110],pp23[110],pp24[110]};
    CLA_4 KS_640(s640, c640, in640_1, in640_2);
    wire[3:0] s641, in641_1, in641_2;
    wire c641;
    assign in641_1 = {pp22[109],pp23[109],pp24[109],pp25[109]};
    assign in641_2 = {pp23[108],pp24[108],pp25[108],pp26[108]};
    CLA_4 KS_641(s641, c641, in641_1, in641_2);
    wire[3:0] s642, in642_1, in642_2;
    wire c642;
    assign in642_1 = {pp24[107],pp25[107],pp26[107],pp27[107]};
    assign in642_2 = {pp25[106],pp26[106],pp27[106],pp28[106]};
    CLA_4 KS_642(s642, c642, in642_1, in642_2);
    wire[3:0] s643, in643_1, in643_2;
    wire c643;
    assign in643_1 = {pp26[105],pp27[105],pp28[105],pp29[105]};
    assign in643_2 = {pp27[104],pp28[104],pp29[104],pp30[104]};
    CLA_4 KS_643(s643, c643, in643_1, in643_2);
    wire[3:0] s644, in644_1, in644_2;
    wire c644;
    assign in644_1 = {pp28[103],pp29[103],pp30[103],pp31[103]};
    assign in644_2 = {pp29[102],pp30[102],pp31[102],pp32[102]};
    CLA_4 KS_644(s644, c644, in644_1, in644_2);
    wire[3:0] s645, in645_1, in645_2;
    wire c645;
    assign in645_1 = {pp30[101],pp31[101],pp32[101],pp33[101]};
    assign in645_2 = {pp31[100],pp32[100],pp33[100],pp34[100]};
    CLA_4 KS_645(s645, c645, in645_1, in645_2);
    wire[3:0] s646, in646_1, in646_2;
    wire c646;
    assign in646_1 = {pp32[99],pp33[99],pp34[99],pp35[99]};
    assign in646_2 = {pp33[98],pp34[98],pp35[98],pp36[98]};
    CLA_4 KS_646(s646, c646, in646_1, in646_2);
    wire[3:0] s647, in647_1, in647_2;
    wire c647;
    assign in647_1 = {pp34[97],pp35[97],pp36[97],pp37[97]};
    assign in647_2 = {pp35[96],pp36[96],pp37[96],pp38[96]};
    CLA_4 KS_647(s647, c647, in647_1, in647_2);
    wire[3:0] s648, in648_1, in648_2;
    wire c648;
    assign in648_1 = {pp36[95],pp37[95],pp38[95],pp39[95]};
    assign in648_2 = {pp37[94],pp38[94],pp39[94],pp40[94]};
    CLA_4 KS_648(s648, c648, in648_1, in648_2);
    wire[3:0] s649, in649_1, in649_2;
    wire c649;
    assign in649_1 = {pp38[93],pp39[93],pp40[93],pp41[93]};
    assign in649_2 = {pp39[92],pp40[92],pp41[92],pp42[92]};
    CLA_4 KS_649(s649, c649, in649_1, in649_2);
    wire[3:0] s650, in650_1, in650_2;
    wire c650;
    assign in650_1 = {pp40[91],pp41[91],pp42[91],pp43[91]};
    assign in650_2 = {pp41[90],pp42[90],pp43[90],pp44[90]};
    CLA_4 KS_650(s650, c650, in650_1, in650_2);
    wire[3:0] s651, in651_1, in651_2;
    wire c651;
    assign in651_1 = {pp42[89],pp43[89],pp44[89],pp45[89]};
    assign in651_2 = {pp43[88],pp44[88],pp45[88],pp46[88]};
    CLA_4 KS_651(s651, c651, in651_1, in651_2);
    wire[3:0] s652, in652_1, in652_2;
    wire c652;
    assign in652_1 = {pp44[87],pp45[87],pp46[87],pp47[87]};
    assign in652_2 = {pp45[86],pp46[86],pp47[86],pp48[86]};
    CLA_4 KS_652(s652, c652, in652_1, in652_2);
    wire[3:0] s653, in653_1, in653_2;
    wire c653;
    assign in653_1 = {pp46[85],pp47[85],pp48[85],pp49[85]};
    assign in653_2 = {pp47[84],pp48[84],pp49[84],pp50[84]};
    CLA_4 KS_653(s653, c653, in653_1, in653_2);
    wire[3:0] s654, in654_1, in654_2;
    wire c654;
    assign in654_1 = {pp48[83],pp49[83],pp50[83],pp51[83]};
    assign in654_2 = {pp49[82],pp50[82],pp51[82],pp52[82]};
    CLA_4 KS_654(s654, c654, in654_1, in654_2);
    wire[3:0] s655, in655_1, in655_2;
    wire c655;
    assign in655_1 = {pp50[81],pp51[81],pp52[81],pp53[81]};
    assign in655_2 = {pp51[80],pp52[80],pp53[80],pp54[80]};
    CLA_4 KS_655(s655, c655, in655_1, in655_2);
    wire[3:0] s656, in656_1, in656_2;
    wire c656;
    assign in656_1 = {pp52[79],pp53[79],pp54[79],pp55[79]};
    assign in656_2 = {pp53[78],pp54[78],pp55[78],pp56[78]};
    CLA_4 KS_656(s656, c656, in656_1, in656_2);
    wire[3:0] s657, in657_1, in657_2;
    wire c657;
    assign in657_1 = {pp54[77],pp55[77],pp56[77],pp57[77]};
    assign in657_2 = {pp55[76],pp56[76],pp57[76],pp58[76]};
    CLA_4 KS_657(s657, c657, in657_1, in657_2);
    wire[3:0] s658, in658_1, in658_2;
    wire c658;
    assign in658_1 = {pp56[75],pp57[75],pp58[75],pp59[75]};
    assign in658_2 = {pp57[74],pp58[74],pp59[74],pp60[74]};
    CLA_4 KS_658(s658, c658, in658_1, in658_2);
    wire[3:0] s659, in659_1, in659_2;
    wire c659;
    assign in659_1 = {pp58[73],pp59[73],pp60[73],pp61[73]};
    assign in659_2 = {pp59[72],pp60[72],pp61[72],pp62[72]};
    CLA_4 KS_659(s659, c659, in659_1, in659_2);
    wire[3:0] s660, in660_1, in660_2;
    wire c660;
    assign in660_1 = {pp60[71],pp61[71],pp62[71],pp63[71]};
    assign in660_2 = {pp61[70],pp62[70],pp63[70],pp64[70]};
    CLA_4 KS_660(s660, c660, in660_1, in660_2);
    wire[3:0] s661, in661_1, in661_2;
    wire c661;
    assign in661_1 = {pp62[69],pp63[69],pp64[69],pp65[69]};
    assign in661_2 = {pp63[68],pp64[68],pp65[68],pp66[68]};
    CLA_4 KS_661(s661, c661, in661_1, in661_2);
    wire[3:0] s662, in662_1, in662_2;
    wire c662;
    assign in662_1 = {pp64[67],pp65[67],pp66[67],pp67[67]};
    assign in662_2 = {pp65[66],pp66[66],pp67[66],pp68[66]};
    CLA_4 KS_662(s662, c662, in662_1, in662_2);
    wire[3:0] s663, in663_1, in663_2;
    wire c663;
    assign in663_1 = {pp66[65],pp67[65],pp68[65],pp69[65]};
    assign in663_2 = {pp67[64],pp68[64],pp69[64],pp70[64]};
    CLA_4 KS_663(s663, c663, in663_1, in663_2);
    wire[3:0] s664, in664_1, in664_2;
    wire c664;
    assign in664_1 = {pp68[63],pp69[63],pp70[63],pp71[63]};
    assign in664_2 = {pp69[62],pp70[62],pp71[62],pp72[62]};
    CLA_4 KS_664(s664, c664, in664_1, in664_2);
    wire[3:0] s665, in665_1, in665_2;
    wire c665;
    assign in665_1 = {pp70[61],pp71[61],pp72[61],pp73[61]};
    assign in665_2 = {pp71[60],pp72[60],pp73[60],pp74[60]};
    CLA_4 KS_665(s665, c665, in665_1, in665_2);
    wire[3:0] s666, in666_1, in666_2;
    wire c666;
    assign in666_1 = {pp72[59],pp73[59],pp74[59],pp75[59]};
    assign in666_2 = {pp73[58],pp74[58],pp75[58],pp76[58]};
    CLA_4 KS_666(s666, c666, in666_1, in666_2);
    wire[3:0] s667, in667_1, in667_2;
    wire c667;
    assign in667_1 = {pp74[57],pp75[57],pp76[57],pp77[57]};
    assign in667_2 = {pp75[56],pp76[56],pp77[56],pp78[56]};
    CLA_4 KS_667(s667, c667, in667_1, in667_2);
    wire[3:0] s668, in668_1, in668_2;
    wire c668;
    assign in668_1 = {pp76[55],pp77[55],pp78[55],pp79[55]};
    assign in668_2 = {pp77[54],pp78[54],pp79[54],pp80[54]};
    CLA_4 KS_668(s668, c668, in668_1, in668_2);
    wire[3:0] s669, in669_1, in669_2;
    wire c669;
    assign in669_1 = {pp78[53],pp79[53],pp80[53],pp81[53]};
    assign in669_2 = {pp79[52],pp80[52],pp81[52],pp82[52]};
    CLA_4 KS_669(s669, c669, in669_1, in669_2);
    wire[3:0] s670, in670_1, in670_2;
    wire c670;
    assign in670_1 = {pp80[51],pp81[51],pp82[51],pp83[51]};
    assign in670_2 = {pp81[50],pp82[50],pp83[50],pp84[50]};
    CLA_4 KS_670(s670, c670, in670_1, in670_2);
    wire[3:0] s671, in671_1, in671_2;
    wire c671;
    assign in671_1 = {pp82[49],pp83[49],pp84[49],pp85[49]};
    assign in671_2 = {pp83[48],pp84[48],pp85[48],pp86[48]};
    CLA_4 KS_671(s671, c671, in671_1, in671_2);
    wire[3:0] s672, in672_1, in672_2;
    wire c672;
    assign in672_1 = {pp84[47],pp85[47],pp86[47],pp87[47]};
    assign in672_2 = {pp85[46],pp86[46],pp87[46],pp88[46]};
    CLA_4 KS_672(s672, c672, in672_1, in672_2);
    wire[3:0] s673, in673_1, in673_2;
    wire c673;
    assign in673_1 = {pp86[45],pp87[45],pp88[45],pp89[45]};
    assign in673_2 = {pp87[44],pp88[44],pp89[44],pp90[44]};
    CLA_4 KS_673(s673, c673, in673_1, in673_2);
    wire[3:0] s674, in674_1, in674_2;
    wire c674;
    assign in674_1 = {pp88[43],pp89[43],pp90[43],pp91[43]};
    assign in674_2 = {pp89[42],pp90[42],pp91[42],pp92[42]};
    CLA_4 KS_674(s674, c674, in674_1, in674_2);
    wire[3:0] s675, in675_1, in675_2;
    wire c675;
    assign in675_1 = {pp90[41],pp91[41],pp92[41],pp93[41]};
    assign in675_2 = {pp91[40],pp92[40],pp93[40],pp94[40]};
    CLA_4 KS_675(s675, c675, in675_1, in675_2);
    wire[3:0] s676, in676_1, in676_2;
    wire c676;
    assign in676_1 = {pp92[39],pp93[39],pp94[39],pp95[39]};
    assign in676_2 = {pp93[38],pp94[38],pp95[38],pp96[38]};
    CLA_4 KS_676(s676, c676, in676_1, in676_2);
    wire[3:0] s677, in677_1, in677_2;
    wire c677;
    assign in677_1 = {pp94[37],pp95[37],pp96[37],pp97[37]};
    assign in677_2 = {pp95[36],pp96[36],pp97[36],pp98[36]};
    CLA_4 KS_677(s677, c677, in677_1, in677_2);
    wire[2:0] s678, in678_1, in678_2;
    wire c678;
    assign in678_1 = {pp96[35],pp97[35],pp98[35]};
    assign in678_2 = {pp97[34],pp98[34],pp99[34]};
    CLA_3 KS_678(s678, c678, in678_1, in678_2);
    wire[1:0] s679, in679_1, in679_2;
    wire c679;
    assign in679_1 = {pp98[33],pp99[33]};
    assign in679_2 = {pp99[32],pp100[32]};
    CLA_2 KS_679(s679, c679, in679_1, in679_2);
    wire[0:0] s680, in680_1, in680_2;
    wire c680;
    assign in680_1 = {pp100[31]};
    assign in680_2 = {pp101[30]};
    Half_Adder KS_680(s680, c680, in680_1, in680_2);
    wire[3:0] s681, in681_1, in681_2;
    wire c681;
    assign in681_1 = {pp102[29],pp101[31],pp100[33],pp99[35]};
    assign in681_2 = {pp103[28],pp102[30],pp101[32],pp100[34]};
    CLA_4 KS_681(s681, c681, in681_1, in681_2);
    wire[0:0] s682, in682_1, in682_2;
    wire c682;
    assign in682_1 = {pp104[27]};
    assign in682_2 = {pp105[26]};
    Half_Adder KS_682(s682, c682, in682_1, in682_2);
    wire[1:0] s683, in683_1, in683_2;
    wire c683;
    assign in683_1 = {pp106[25],pp103[29]};
    assign in683_2 = {pp107[24],pp104[28]};
    CLA_2 KS_683(s683, c683, in683_1, in683_2);
    wire[0:0] s684, in684_1, in684_2;
    wire c684;
    assign in684_1 = {pp108[23]};
    assign in684_2 = {pp109[22]};
    Half_Adder KS_684(s684, c684, in684_1, in684_2);
    wire[2:0] s685, in685_1, in685_2;
    wire c685;
    assign in685_1 = {pp110[21],pp105[27],pp102[31]};
    assign in685_2 = {pp111[20],pp106[26],pp103[30]};
    CLA_3 KS_685(s685, c685, in685_1, in685_2);
    wire[0:0] s686, in686_1, in686_2;
    wire c686;
    assign in686_1 = {pp112[19]};
    assign in686_2 = {pp113[18]};
    Half_Adder KS_686(s686, c686, in686_1, in686_2);
    wire[1:0] s687, in687_1, in687_2;
    wire c687;
    assign in687_1 = {pp114[17],pp107[25]};
    assign in687_2 = {pp115[16],pp108[24]};
    CLA_2 KS_687(s687, c687, in687_1, in687_2);
    wire[0:0] s688, in688_1, in688_2;
    wire c688;
    assign in688_1 = {pp116[15]};
    assign in688_2 = {pp117[14]};
    Half_Adder KS_688(s688, c688, in688_1, in688_2);
    wire[3:0] s689, in689_1, in689_2;
    wire c689;
    assign in689_1 = {pp118[13],pp109[23],pp104[29],pp101[33]};
    assign in689_2 = {pp119[12],pp110[22],pp105[28],pp102[32]};
    CLA_4 KS_689(s689, c689, in689_1, in689_2);
    wire[0:0] s690, in690_1, in690_2;
    wire c690;
    assign in690_1 = {pp120[11]};
    assign in690_2 = {pp121[10]};
    Half_Adder KS_690(s690, c690, in690_1, in690_2);
    wire[1:0] s691, in691_1, in691_2;
    wire c691;
    assign in691_1 = {pp122[9],pp111[21]};
    assign in691_2 = {pp123[8],pp112[20]};
    CLA_2 KS_691(s691, c691, in691_1, in691_2);
    wire[0:0] s692, in692_1, in692_2;
    wire c692;
    assign in692_1 = {pp124[7]};
    assign in692_2 = {pp125[6]};
    Half_Adder KS_692(s692, c692, in692_1, in692_2);
    wire[2:0] s693, in693_1, in693_2;
    wire c693;
    assign in693_1 = {pp126[5],pp113[19],pp106[27]};
    assign in693_2 = {pp127[4],pp114[18],pp107[26]};
    CLA_3 KS_693(s693, c693, in693_1, in693_2);
    wire[0:0] s694, in694_1, in694_2;
    wire c694;
    assign in694_1 = {c525};
    assign in694_2 = {c526};
    Half_Adder KS_694(s694, c694, in694_1, in694_2);
    wire[1:0] s695, in695_1, in695_2;
    wire c695;
    assign in695_1 = {c527,pp115[17]};
    assign in695_2 = {c528,pp116[16]};
    CLA_2 KS_695(s695, c695, in695_1, in695_2);
    wire[0:0] s696, in696_1, in696_2;
    wire c696;
    assign in696_1 = {c529};
    assign in696_2 = {c530};
    Half_Adder KS_696(s696, c696, in696_1, in696_2);
    wire[3:0] s697, in697_1, in697_2;
    wire c697;
    assign in697_1 = {c531,pp117[15],pp108[25],pp103[31]};
    assign in697_2 = {c532,pp118[14],pp109[24],pp104[30]};
    CLA_4 KS_697(s697, c697, in697_1, in697_2);
    wire[0:0] s698, in698_1, in698_2;
    wire c698;
    assign in698_1 = {c533};
    assign in698_2 = {c534};
    Half_Adder KS_698(s698, c698, in698_1, in698_2);
    wire[1:0] s699, in699_1, in699_2;
    wire c699;
    assign in699_1 = {c535,pp119[13]};
    assign in699_2 = {c536,pp120[12]};
    CLA_2 KS_699(s699, c699, in699_1, in699_2);
    wire[0:0] s700, in700_1, in700_2;
    wire c700;
    assign in700_1 = {c537};
    assign in700_2 = {c538};
    Half_Adder KS_700(s700, c700, in700_1, in700_2);
    wire[2:0] s701, in701_1, in701_2;
    wire c701;
    assign in701_1 = {c539,pp121[11],pp110[23]};
    assign in701_2 = {c540,pp122[10],pp111[22]};
    CLA_3 KS_701(s701, c701, in701_1, in701_2);
    wire[0:0] s702, in702_1, in702_2;
    wire c702;
    assign in702_1 = {c541};
    assign in702_2 = {c542};
    Half_Adder KS_702(s702, c702, in702_1, in702_2);
    wire[1:0] s703, in703_1, in703_2;
    wire c703;
    assign in703_1 = {c543,pp123[9]};
    assign in703_2 = {c544,pp124[8]};
    CLA_2 KS_703(s703, c703, in703_1, in703_2);
    wire[0:0] s704, in704_1, in704_2;
    wire c704;
    assign in704_1 = {c545};
    assign in704_2 = {c546};
    Half_Adder KS_704(s704, c704, in704_1, in704_2);
    wire[3:0] s705, in705_1, in705_2;
    wire c705;
    assign in705_1 = {c547,pp125[7],pp112[21],pp105[29]};
    assign in705_2 = {c548,pp126[6],pp113[20],pp106[28]};
    CLA_4 KS_705(s705, c705, in705_1, in705_2);
    wire[0:0] s706, in706_1, in706_2;
    wire c706;
    assign in706_1 = {c549};
    assign in706_2 = {c550};
    Half_Adder KS_706(s706, c706, in706_1, in706_2);
    wire[1:0] s707, in707_1, in707_2;
    wire c707;
    assign in707_1 = {c551,pp127[5]};
    assign in707_2 = {c552,s632[1]};
    CLA_2 KS_707(s707, c707, in707_1, in707_2);
    wire[0:0] s708, in708_1, in708_2;
    wire c708;
    assign in708_1 = {c553};
    assign in708_2 = {c554};
    Half_Adder KS_708(s708, c708, in708_1, in708_2);
    wire[2:0] s709, in709_1, in709_2;
    wire c709;
    assign in709_1 = {c555,s633[1],pp114[19]};
    assign in709_2 = {c556,s634[1],pp115[18]};
    CLA_3 KS_709(s709, c709, in709_1, in709_2);
    wire[0:0] s710, in710_1, in710_2;
    wire c710;
    assign in710_1 = {c557};
    assign in710_2 = {c558};
    Half_Adder KS_710(s710, c710, in710_1, in710_2);
    wire[1:0] s711, in711_1, in711_2;
    wire c711;
    assign in711_1 = {c559,s635[1]};
    assign in711_2 = {c560,s636[1]};
    CLA_2 KS_711(s711, c711, in711_1, in711_2);
    wire[0:0] s712, in712_1, in712_2;
    wire c712;
    assign in712_1 = {c561};
    assign in712_2 = {c562};
    Half_Adder KS_712(s712, c712, in712_1, in712_2);
    wire[3:0] s713, in713_1, in713_2;
    wire c713;
    assign in713_1 = {c563,s637[1],pp116[17],pp107[27]};
    assign in713_2 = {c564,s638[1],pp117[16],pp108[26]};
    CLA_4 KS_713(s713, c713, in713_1, in713_2);
    wire[0:0] s714, in714_1, in714_2;
    wire c714;
    assign in714_1 = {c565};
    assign in714_2 = {c566};
    Half_Adder KS_714(s714, c714, in714_1, in714_2);
    wire[1:0] s715, in715_1, in715_2;
    wire c715;
    assign in715_1 = {c567,s639[1]};
    assign in715_2 = {c568,s640[1]};
    CLA_2 KS_715(s715, c715, in715_1, in715_2);
    wire[0:0] s716, in716_1, in716_2;
    wire c716;
    assign in716_1 = {c569};
    assign in716_2 = {c570};
    Half_Adder KS_716(s716, c716, in716_1, in716_2);
    wire[2:0] s717, in717_1, in717_2;
    wire c717;
    assign in717_1 = {c571,s641[1],pp118[15]};
    assign in717_2 = {c572,s642[1],pp119[14]};
    CLA_3 KS_717(s717, c717, in717_1, in717_2);
    wire[0:0] s718, in718_1, in718_2;
    wire c718;
    assign in718_1 = {c573};
    assign in718_2 = {c574};
    Half_Adder KS_718(s718, c718, in718_1, in718_2);
    wire[1:0] s719, in719_1, in719_2;
    wire c719;
    assign in719_1 = {c577,s643[1]};
    assign in719_2 = {c585,s644[1]};
    CLA_2 KS_719(s719, c719, in719_1, in719_2);
    wire[0:0] s720, in720_1, in720_2;
    wire c720;
    assign in720_1 = {c593};
    assign in720_2 = {c601};
    Half_Adder KS_720(s720, c720, in720_1, in720_2);
    wire[3:0] s721, in721_1, in721_2;
    wire c721;
    assign in721_1 = {c609,s645[1],pp120[13],pp109[25]};
    assign in721_2 = {c617,s646[1],pp121[12],pp110[24]};
    CLA_4 KS_721(s721, c721, in721_1, in721_2);
    wire[0:0] s722, in722_1, in722_2;
    wire c722;
    assign in722_1 = {c625};
    assign in722_2 = {s632[0]};
    Half_Adder KS_722(s722, c722, in722_1, in722_2);
    wire[1:0] s723, in723_1, in723_2;
    wire c723;
    assign in723_1 = {s633[0],s647[1]};
    assign in723_2 = {s634[0],s648[1]};
    CLA_2 KS_723(s723, c723, in723_1, in723_2);
    wire[0:0] s724, in724_1, in724_2;
    wire c724;
    assign in724_1 = {s635[0]};
    assign in724_2 = {s636[0]};
    Half_Adder KS_724(s724, c724, in724_1, in724_2);
    wire[2:0] s725, in725_1, in725_2;
    wire c725;
    assign in725_1 = {s637[0],s649[1],pp122[11]};
    assign in725_2 = {s638[0],s650[1],pp123[10]};
    CLA_3 KS_725(s725, c725, in725_1, in725_2);
    wire[0:0] s726, in726_1, in726_2;
    wire c726;
    assign in726_1 = {s639[0]};
    assign in726_2 = {s640[0]};
    Half_Adder KS_726(s726, c726, in726_1, in726_2);
    wire[1:0] s727, in727_1, in727_2;
    wire c727;
    assign in727_1 = {s641[0],s651[1]};
    assign in727_2 = {s642[0],s652[1]};
    CLA_2 KS_727(s727, c727, in727_1, in727_2);
    wire[0:0] s728, in728_1, in728_2;
    wire c728;
    assign in728_1 = {s643[0]};
    assign in728_2 = {s644[0]};
    Half_Adder KS_728(s728, c728, in728_1, in728_2);
    wire[3:0] s729, in729_1, in729_2;
    wire c729;
    assign in729_1 = {s645[0],s653[1],pp124[9],pp111[23]};
    assign in729_2 = {s646[0],s654[1],pp125[8],pp112[22]};
    CLA_4 KS_729(s729, c729, in729_1, in729_2);
    wire[0:0] s730, in730_1, in730_2;
    wire c730;
    assign in730_1 = {s647[0]};
    assign in730_2 = {s648[0]};
    Half_Adder KS_730(s730, c730, in730_1, in730_2);
    wire[1:0] s731, in731_1, in731_2;
    wire c731;
    assign in731_1 = {s649[0],s655[1]};
    assign in731_2 = {s650[0],s656[1]};
    CLA_2 KS_731(s731, c731, in731_1, in731_2);
    wire[0:0] s732, in732_1, in732_2;
    wire c732;
    assign in732_1 = {s651[0]};
    assign in732_2 = {s652[0]};
    Half_Adder KS_732(s732, c732, in732_1, in732_2);
    wire[2:0] s733, in733_1, in733_2;
    wire c733;
    assign in733_1 = {s653[0],s657[1],pp126[7]};
    assign in733_2 = {s654[0],s658[1],pp127[6]};
    CLA_3 KS_733(s733, c733, in733_1, in733_2);
    wire[0:0] s734, in734_1, in734_2;
    wire c734;
    assign in734_1 = {s655[0]};
    assign in734_2 = {s656[0]};
    Half_Adder KS_734(s734, c734, in734_1, in734_2);
    wire[1:0] s735, in735_1, in735_2;
    wire c735;
    assign in735_1 = {s658[0],s659[1]};
    assign in735_2 = {s659[0],s660[1]};
    CLA_2_c KS_735(s735, c735, in735_1, in735_2, s657[0]);
    wire[3:0] s736, in736_1, in736_2;
    wire c736;
    assign in736_1 = {pp8[127],pp9[127],pp10[127],pp11[127]};
    assign in736_2 = {pp9[126],pp10[126],pp11[126],pp12[126]};
    CLA_4 KS_736(s736, c736, in736_1, in736_2);
    wire[3:0] s737, in737_1, in737_2;
    wire c737;
    assign in737_1 = {pp10[125],pp11[125],pp12[125],pp13[125]};
    assign in737_2 = {pp11[124],pp12[124],pp13[124],pp14[124]};
    CLA_4 KS_737(s737, c737, in737_1, in737_2);
    wire[3:0] s738, in738_1, in738_2;
    wire c738;
    assign in738_1 = {pp12[123],pp13[123],pp14[123],pp15[123]};
    assign in738_2 = {pp13[122],pp14[122],pp15[122],pp16[122]};
    CLA_4 KS_738(s738, c738, in738_1, in738_2);
    wire[3:0] s739, in739_1, in739_2;
    wire c739;
    assign in739_1 = {pp14[121],pp15[121],pp16[121],pp17[121]};
    assign in739_2 = {pp15[120],pp16[120],pp17[120],pp18[120]};
    CLA_4 KS_739(s739, c739, in739_1, in739_2);
    wire[3:0] s740, in740_1, in740_2;
    wire c740;
    assign in740_1 = {pp16[119],pp17[119],pp18[119],pp19[119]};
    assign in740_2 = {pp17[118],pp18[118],pp19[118],pp20[118]};
    CLA_4 KS_740(s740, c740, in740_1, in740_2);
    wire[3:0] s741, in741_1, in741_2;
    wire c741;
    assign in741_1 = {pp18[117],pp19[117],pp20[117],pp21[117]};
    assign in741_2 = {pp19[116],pp20[116],pp21[116],pp22[116]};
    CLA_4 KS_741(s741, c741, in741_1, in741_2);
    wire[3:0] s742, in742_1, in742_2;
    wire c742;
    assign in742_1 = {pp20[115],pp21[115],pp22[115],pp23[115]};
    assign in742_2 = {pp21[114],pp22[114],pp23[114],pp24[114]};
    CLA_4 KS_742(s742, c742, in742_1, in742_2);
    wire[3:0] s743, in743_1, in743_2;
    wire c743;
    assign in743_1 = {pp22[113],pp23[113],pp24[113],pp25[113]};
    assign in743_2 = {pp23[112],pp24[112],pp25[112],pp26[112]};
    CLA_4 KS_743(s743, c743, in743_1, in743_2);
    wire[3:0] s744, in744_1, in744_2;
    wire c744;
    assign in744_1 = {pp24[111],pp25[111],pp26[111],pp27[111]};
    assign in744_2 = {pp25[110],pp26[110],pp27[110],pp28[110]};
    CLA_4 KS_744(s744, c744, in744_1, in744_2);
    wire[3:0] s745, in745_1, in745_2;
    wire c745;
    assign in745_1 = {pp26[109],pp27[109],pp28[109],pp29[109]};
    assign in745_2 = {pp27[108],pp28[108],pp29[108],pp30[108]};
    CLA_4 KS_745(s745, c745, in745_1, in745_2);
    wire[3:0] s746, in746_1, in746_2;
    wire c746;
    assign in746_1 = {pp28[107],pp29[107],pp30[107],pp31[107]};
    assign in746_2 = {pp29[106],pp30[106],pp31[106],pp32[106]};
    CLA_4 KS_746(s746, c746, in746_1, in746_2);
    wire[3:0] s747, in747_1, in747_2;
    wire c747;
    assign in747_1 = {pp30[105],pp31[105],pp32[105],pp33[105]};
    assign in747_2 = {pp31[104],pp32[104],pp33[104],pp34[104]};
    CLA_4 KS_747(s747, c747, in747_1, in747_2);
    wire[3:0] s748, in748_1, in748_2;
    wire c748;
    assign in748_1 = {pp32[103],pp33[103],pp34[103],pp35[103]};
    assign in748_2 = {pp33[102],pp34[102],pp35[102],pp36[102]};
    CLA_4 KS_748(s748, c748, in748_1, in748_2);
    wire[3:0] s749, in749_1, in749_2;
    wire c749;
    assign in749_1 = {pp34[101],pp35[101],pp36[101],pp37[101]};
    assign in749_2 = {pp35[100],pp36[100],pp37[100],pp38[100]};
    CLA_4 KS_749(s749, c749, in749_1, in749_2);
    wire[3:0] s750, in750_1, in750_2;
    wire c750;
    assign in750_1 = {pp36[99],pp37[99],pp38[99],pp39[99]};
    assign in750_2 = {pp37[98],pp38[98],pp39[98],pp40[98]};
    CLA_4 KS_750(s750, c750, in750_1, in750_2);
    wire[3:0] s751, in751_1, in751_2;
    wire c751;
    assign in751_1 = {pp38[97],pp39[97],pp40[97],pp41[97]};
    assign in751_2 = {pp39[96],pp40[96],pp41[96],pp42[96]};
    CLA_4 KS_751(s751, c751, in751_1, in751_2);
    wire[3:0] s752, in752_1, in752_2;
    wire c752;
    assign in752_1 = {pp40[95],pp41[95],pp42[95],pp43[95]};
    assign in752_2 = {pp41[94],pp42[94],pp43[94],pp44[94]};
    CLA_4 KS_752(s752, c752, in752_1, in752_2);
    wire[3:0] s753, in753_1, in753_2;
    wire c753;
    assign in753_1 = {pp42[93],pp43[93],pp44[93],pp45[93]};
    assign in753_2 = {pp43[92],pp44[92],pp45[92],pp46[92]};
    CLA_4 KS_753(s753, c753, in753_1, in753_2);
    wire[3:0] s754, in754_1, in754_2;
    wire c754;
    assign in754_1 = {pp44[91],pp45[91],pp46[91],pp47[91]};
    assign in754_2 = {pp45[90],pp46[90],pp47[90],pp48[90]};
    CLA_4 KS_754(s754, c754, in754_1, in754_2);
    wire[3:0] s755, in755_1, in755_2;
    wire c755;
    assign in755_1 = {pp46[89],pp47[89],pp48[89],pp49[89]};
    assign in755_2 = {pp47[88],pp48[88],pp49[88],pp50[88]};
    CLA_4 KS_755(s755, c755, in755_1, in755_2);
    wire[3:0] s756, in756_1, in756_2;
    wire c756;
    assign in756_1 = {pp48[87],pp49[87],pp50[87],pp51[87]};
    assign in756_2 = {pp49[86],pp50[86],pp51[86],pp52[86]};
    CLA_4 KS_756(s756, c756, in756_1, in756_2);
    wire[3:0] s757, in757_1, in757_2;
    wire c757;
    assign in757_1 = {pp50[85],pp51[85],pp52[85],pp53[85]};
    assign in757_2 = {pp51[84],pp52[84],pp53[84],pp54[84]};
    CLA_4 KS_757(s757, c757, in757_1, in757_2);
    wire[3:0] s758, in758_1, in758_2;
    wire c758;
    assign in758_1 = {pp52[83],pp53[83],pp54[83],pp55[83]};
    assign in758_2 = {pp53[82],pp54[82],pp55[82],pp56[82]};
    CLA_4 KS_758(s758, c758, in758_1, in758_2);
    wire[3:0] s759, in759_1, in759_2;
    wire c759;
    assign in759_1 = {pp54[81],pp55[81],pp56[81],pp57[81]};
    assign in759_2 = {pp55[80],pp56[80],pp57[80],pp58[80]};
    CLA_4 KS_759(s759, c759, in759_1, in759_2);
    wire[3:0] s760, in760_1, in760_2;
    wire c760;
    assign in760_1 = {pp56[79],pp57[79],pp58[79],pp59[79]};
    assign in760_2 = {pp57[78],pp58[78],pp59[78],pp60[78]};
    CLA_4 KS_760(s760, c760, in760_1, in760_2);
    wire[3:0] s761, in761_1, in761_2;
    wire c761;
    assign in761_1 = {pp58[77],pp59[77],pp60[77],pp61[77]};
    assign in761_2 = {pp59[76],pp60[76],pp61[76],pp62[76]};
    CLA_4 KS_761(s761, c761, in761_1, in761_2);
    wire[3:0] s762, in762_1, in762_2;
    wire c762;
    assign in762_1 = {pp60[75],pp61[75],pp62[75],pp63[75]};
    assign in762_2 = {pp61[74],pp62[74],pp63[74],pp64[74]};
    CLA_4 KS_762(s762, c762, in762_1, in762_2);
    wire[3:0] s763, in763_1, in763_2;
    wire c763;
    assign in763_1 = {pp62[73],pp63[73],pp64[73],pp65[73]};
    assign in763_2 = {pp63[72],pp64[72],pp65[72],pp66[72]};
    CLA_4 KS_763(s763, c763, in763_1, in763_2);
    wire[3:0] s764, in764_1, in764_2;
    wire c764;
    assign in764_1 = {pp64[71],pp65[71],pp66[71],pp67[71]};
    assign in764_2 = {pp65[70],pp66[70],pp67[70],pp68[70]};
    CLA_4 KS_764(s764, c764, in764_1, in764_2);
    wire[3:0] s765, in765_1, in765_2;
    wire c765;
    assign in765_1 = {pp66[69],pp67[69],pp68[69],pp69[69]};
    assign in765_2 = {pp67[68],pp68[68],pp69[68],pp70[68]};
    CLA_4 KS_765(s765, c765, in765_1, in765_2);
    wire[3:0] s766, in766_1, in766_2;
    wire c766;
    assign in766_1 = {pp68[67],pp69[67],pp70[67],pp71[67]};
    assign in766_2 = {pp69[66],pp70[66],pp71[66],pp72[66]};
    CLA_4 KS_766(s766, c766, in766_1, in766_2);
    wire[3:0] s767, in767_1, in767_2;
    wire c767;
    assign in767_1 = {pp70[65],pp71[65],pp72[65],pp73[65]};
    assign in767_2 = {pp71[64],pp72[64],pp73[64],pp74[64]};
    CLA_4 KS_767(s767, c767, in767_1, in767_2);
    wire[3:0] s768, in768_1, in768_2;
    wire c768;
    assign in768_1 = {pp72[63],pp73[63],pp74[63],pp75[63]};
    assign in768_2 = {pp73[62],pp74[62],pp75[62],pp76[62]};
    CLA_4 KS_768(s768, c768, in768_1, in768_2);
    wire[3:0] s769, in769_1, in769_2;
    wire c769;
    assign in769_1 = {pp74[61],pp75[61],pp76[61],pp77[61]};
    assign in769_2 = {pp75[60],pp76[60],pp77[60],pp78[60]};
    CLA_4 KS_769(s769, c769, in769_1, in769_2);
    wire[3:0] s770, in770_1, in770_2;
    wire c770;
    assign in770_1 = {pp76[59],pp77[59],pp78[59],pp79[59]};
    assign in770_2 = {pp77[58],pp78[58],pp79[58],pp80[58]};
    CLA_4 KS_770(s770, c770, in770_1, in770_2);
    wire[3:0] s771, in771_1, in771_2;
    wire c771;
    assign in771_1 = {pp78[57],pp79[57],pp80[57],pp81[57]};
    assign in771_2 = {pp79[56],pp80[56],pp81[56],pp82[56]};
    CLA_4 KS_771(s771, c771, in771_1, in771_2);
    wire[3:0] s772, in772_1, in772_2;
    wire c772;
    assign in772_1 = {pp80[55],pp81[55],pp82[55],pp83[55]};
    assign in772_2 = {pp81[54],pp82[54],pp83[54],pp84[54]};
    CLA_4 KS_772(s772, c772, in772_1, in772_2);
    wire[3:0] s773, in773_1, in773_2;
    wire c773;
    assign in773_1 = {pp82[53],pp83[53],pp84[53],pp85[53]};
    assign in773_2 = {pp83[52],pp84[52],pp85[52],pp86[52]};
    CLA_4 KS_773(s773, c773, in773_1, in773_2);
    wire[3:0] s774, in774_1, in774_2;
    wire c774;
    assign in774_1 = {pp84[51],pp85[51],pp86[51],pp87[51]};
    assign in774_2 = {pp85[50],pp86[50],pp87[50],pp88[50]};
    CLA_4 KS_774(s774, c774, in774_1, in774_2);
    wire[3:0] s775, in775_1, in775_2;
    wire c775;
    assign in775_1 = {pp86[49],pp87[49],pp88[49],pp89[49]};
    assign in775_2 = {pp87[48],pp88[48],pp89[48],pp90[48]};
    CLA_4 KS_775(s775, c775, in775_1, in775_2);
    wire[3:0] s776, in776_1, in776_2;
    wire c776;
    assign in776_1 = {pp88[47],pp89[47],pp90[47],pp91[47]};
    assign in776_2 = {pp89[46],pp90[46],pp91[46],pp92[46]};
    CLA_4 KS_776(s776, c776, in776_1, in776_2);
    wire[3:0] s777, in777_1, in777_2;
    wire c777;
    assign in777_1 = {pp90[45],pp91[45],pp92[45],pp93[45]};
    assign in777_2 = {pp91[44],pp92[44],pp93[44],pp94[44]};
    CLA_4 KS_777(s777, c777, in777_1, in777_2);
    wire[2:0] s778, in778_1, in778_2;
    wire c778;
    assign in778_1 = {pp92[43],pp93[43],pp94[43]};
    assign in778_2 = {pp93[42],pp94[42],pp95[42]};
    CLA_3 KS_778(s778, c778, in778_1, in778_2);
    wire[1:0] s779, in779_1, in779_2;
    wire c779;
    assign in779_1 = {pp94[41],pp95[41]};
    assign in779_2 = {pp95[40],pp96[40]};
    CLA_2 KS_779(s779, c779, in779_1, in779_2);
    wire[0:0] s780, in780_1, in780_2;
    wire c780;
    assign in780_1 = {pp96[39]};
    assign in780_2 = {pp97[38]};
    Half_Adder KS_780(s780, c780, in780_1, in780_2);
    wire[3:0] s781, in781_1, in781_2;
    wire c781;
    assign in781_1 = {pp98[37],pp97[39],pp96[41],pp95[43]};
    assign in781_2 = {pp99[36],pp98[38],pp97[40],pp96[42]};
    CLA_4 KS_781(s781, c781, in781_1, in781_2);
    wire[0:0] s782, in782_1, in782_2;
    wire c782;
    assign in782_1 = {pp100[35]};
    assign in782_2 = {pp101[34]};
    Half_Adder KS_782(s782, c782, in782_1, in782_2);
    wire[1:0] s783, in783_1, in783_2;
    wire c783;
    assign in783_1 = {pp102[33],pp99[37]};
    assign in783_2 = {pp103[32],pp100[36]};
    CLA_2 KS_783(s783, c783, in783_1, in783_2);
    wire[0:0] s784, in784_1, in784_2;
    wire c784;
    assign in784_1 = {pp104[31]};
    assign in784_2 = {pp105[30]};
    Half_Adder KS_784(s784, c784, in784_1, in784_2);
    wire[2:0] s785, in785_1, in785_2;
    wire c785;
    assign in785_1 = {pp106[29],pp101[35],pp98[39]};
    assign in785_2 = {pp107[28],pp102[34],pp99[38]};
    CLA_3 KS_785(s785, c785, in785_1, in785_2);
    wire[0:0] s786, in786_1, in786_2;
    wire c786;
    assign in786_1 = {pp108[27]};
    assign in786_2 = {pp109[26]};
    Half_Adder KS_786(s786, c786, in786_1, in786_2);
    wire[1:0] s787, in787_1, in787_2;
    wire c787;
    assign in787_1 = {pp110[25],pp103[33]};
    assign in787_2 = {pp111[24],pp104[32]};
    CLA_2 KS_787(s787, c787, in787_1, in787_2);
    wire[0:0] s788, in788_1, in788_2;
    wire c788;
    assign in788_1 = {pp112[23]};
    assign in788_2 = {pp113[22]};
    Half_Adder KS_788(s788, c788, in788_1, in788_2);
    wire[3:0] s789, in789_1, in789_2;
    wire c789;
    assign in789_1 = {pp114[21],pp105[31],pp100[37],pp97[41]};
    assign in789_2 = {pp115[20],pp106[30],pp101[36],pp98[40]};
    CLA_4 KS_789(s789, c789, in789_1, in789_2);
    wire[0:0] s790, in790_1, in790_2;
    wire c790;
    assign in790_1 = {pp116[19]};
    assign in790_2 = {pp117[18]};
    Half_Adder KS_790(s790, c790, in790_1, in790_2);
    wire[1:0] s791, in791_1, in791_2;
    wire c791;
    assign in791_1 = {pp118[17],pp107[29]};
    assign in791_2 = {pp119[16],pp108[28]};
    CLA_2 KS_791(s791, c791, in791_1, in791_2);
    wire[0:0] s792, in792_1, in792_2;
    wire c792;
    assign in792_1 = {pp120[15]};
    assign in792_2 = {pp121[14]};
    Half_Adder KS_792(s792, c792, in792_1, in792_2);
    wire[2:0] s793, in793_1, in793_2;
    wire c793;
    assign in793_1 = {pp122[13],pp109[27],pp102[35]};
    assign in793_2 = {pp123[12],pp110[26],pp103[34]};
    CLA_3 KS_793(s793, c793, in793_1, in793_2);
    wire[0:0] s794, in794_1, in794_2;
    wire c794;
    assign in794_1 = {pp124[11]};
    assign in794_2 = {pp125[10]};
    Half_Adder KS_794(s794, c794, in794_1, in794_2);
    wire[1:0] s795, in795_1, in795_2;
    wire c795;
    assign in795_1 = {pp126[9],pp111[25]};
    assign in795_2 = {pp127[8],pp112[24]};
    CLA_2 KS_795(s795, c795, in795_1, in795_2);
    wire[0:0] s796, in796_1, in796_2;
    wire c796;
    assign in796_1 = {c632};
    assign in796_2 = {c633};
    Half_Adder KS_796(s796, c796, in796_1, in796_2);
    wire[3:0] s797, in797_1, in797_2;
    wire c797;
    assign in797_1 = {c634,pp113[23],pp104[33],pp99[39]};
    assign in797_2 = {c635,pp114[22],pp105[32],pp100[38]};
    CLA_4 KS_797(s797, c797, in797_1, in797_2);
    wire[0:0] s798, in798_1, in798_2;
    wire c798;
    assign in798_1 = {c636};
    assign in798_2 = {c637};
    Half_Adder KS_798(s798, c798, in798_1, in798_2);
    wire[1:0] s799, in799_1, in799_2;
    wire c799;
    assign in799_1 = {c638,pp115[21]};
    assign in799_2 = {c639,pp116[20]};
    CLA_2 KS_799(s799, c799, in799_1, in799_2);
    wire[0:0] s800, in800_1, in800_2;
    wire c800;
    assign in800_1 = {c640};
    assign in800_2 = {c641};
    Half_Adder KS_800(s800, c800, in800_1, in800_2);
    wire[2:0] s801, in801_1, in801_2;
    wire c801;
    assign in801_1 = {c642,pp117[19],pp106[31]};
    assign in801_2 = {c643,pp118[18],pp107[30]};
    CLA_3 KS_801(s801, c801, in801_1, in801_2);
    wire[0:0] s802, in802_1, in802_2;
    wire c802;
    assign in802_1 = {c644};
    assign in802_2 = {c645};
    Half_Adder KS_802(s802, c802, in802_1, in802_2);
    wire[1:0] s803, in803_1, in803_2;
    wire c803;
    assign in803_1 = {c646,pp119[17]};
    assign in803_2 = {c647,pp120[16]};
    CLA_2 KS_803(s803, c803, in803_1, in803_2);
    wire[0:0] s804, in804_1, in804_2;
    wire c804;
    assign in804_1 = {c648};
    assign in804_2 = {c649};
    Half_Adder KS_804(s804, c804, in804_1, in804_2);
    wire[3:0] s805, in805_1, in805_2;
    wire c805;
    assign in805_1 = {c650,pp121[15],pp108[29],pp101[37]};
    assign in805_2 = {c651,pp122[14],pp109[28],pp102[36]};
    CLA_4 KS_805(s805, c805, in805_1, in805_2);
    wire[0:0] s806, in806_1, in806_2;
    wire c806;
    assign in806_1 = {c652};
    assign in806_2 = {c653};
    Half_Adder KS_806(s806, c806, in806_1, in806_2);
    wire[1:0] s807, in807_1, in807_2;
    wire c807;
    assign in807_1 = {c654,pp123[13]};
    assign in807_2 = {c655,pp124[12]};
    CLA_2 KS_807(s807, c807, in807_1, in807_2);
    wire[0:0] s808, in808_1, in808_2;
    wire c808;
    assign in808_1 = {c656};
    assign in808_2 = {c657};
    Half_Adder KS_808(s808, c808, in808_1, in808_2);
    wire[2:0] s809, in809_1, in809_2;
    wire c809;
    assign in809_1 = {c658,pp125[11],pp110[27]};
    assign in809_2 = {c659,pp126[10],pp111[26]};
    CLA_3 KS_809(s809, c809, in809_1, in809_2);
    wire[0:0] s810, in810_1, in810_2;
    wire c810;
    assign in810_1 = {c660};
    assign in810_2 = {c661};
    Half_Adder KS_810(s810, c810, in810_1, in810_2);
    wire[1:0] s811, in811_1, in811_2;
    wire c811;
    assign in811_1 = {c662,pp127[9]};
    assign in811_2 = {c663,s736[1]};
    CLA_2 KS_811(s811, c811, in811_1, in811_2);
    wire[0:0] s812, in812_1, in812_2;
    wire c812;
    assign in812_1 = {c664};
    assign in812_2 = {c665};
    Half_Adder KS_812(s812, c812, in812_1, in812_2);
    wire[3:0] s813, in813_1, in813_2;
    wire c813;
    assign in813_1 = {c666,s737[1],pp112[25],pp103[35]};
    assign in813_2 = {c667,s738[1],pp113[24],pp104[34]};
    CLA_4 KS_813(s813, c813, in813_1, in813_2);
    wire[0:0] s814, in814_1, in814_2;
    wire c814;
    assign in814_1 = {c668};
    assign in814_2 = {c669};
    Half_Adder KS_814(s814, c814, in814_1, in814_2);
    wire[1:0] s815, in815_1, in815_2;
    wire c815;
    assign in815_1 = {c670,s739[1]};
    assign in815_2 = {c671,s740[1]};
    CLA_2 KS_815(s815, c815, in815_1, in815_2);
    wire[0:0] s816, in816_1, in816_2;
    wire c816;
    assign in816_1 = {c672};
    assign in816_2 = {c673};
    Half_Adder KS_816(s816, c816, in816_1, in816_2);
    wire[2:0] s817, in817_1, in817_2;
    wire c817;
    assign in817_1 = {c674,s741[1],pp114[23]};
    assign in817_2 = {c675,s742[1],pp115[22]};
    CLA_3 KS_817(s817, c817, in817_1, in817_2);
    wire[0:0] s818, in818_1, in818_2;
    wire c818;
    assign in818_1 = {c676};
    assign in818_2 = {c677};
    Half_Adder KS_818(s818, c818, in818_1, in818_2);
    wire[1:0] s819, in819_1, in819_2;
    wire c819;
    assign in819_1 = {c681,s743[1]};
    assign in819_2 = {c689,s744[1]};
    CLA_2 KS_819(s819, c819, in819_1, in819_2);
    wire[0:0] s820, in820_1, in820_2;
    wire c820;
    assign in820_1 = {c697};
    assign in820_2 = {c705};
    Half_Adder KS_820(s820, c820, in820_1, in820_2);
    wire[3:0] s821, in821_1, in821_2;
    wire c821;
    assign in821_1 = {c713,s745[1],pp116[21],pp105[33]};
    assign in821_2 = {c721,s746[1],pp117[20],pp106[32]};
    CLA_4 KS_821(s821, c821, in821_1, in821_2);
    wire[0:0] s822, in822_1, in822_2;
    wire c822;
    assign in822_1 = {c729};
    assign in822_2 = {s736[0]};
    Half_Adder KS_822(s822, c822, in822_1, in822_2);
    wire[1:0] s823, in823_1, in823_2;
    wire c823;
    assign in823_1 = {s737[0],s747[1]};
    assign in823_2 = {s738[0],s748[1]};
    CLA_2 KS_823(s823, c823, in823_1, in823_2);
    wire[0:0] s824, in824_1, in824_2;
    wire c824;
    assign in824_1 = {s739[0]};
    assign in824_2 = {s740[0]};
    Half_Adder KS_824(s824, c824, in824_1, in824_2);
    wire[2:0] s825, in825_1, in825_2;
    wire c825;
    assign in825_1 = {s741[0],s749[1],pp118[19]};
    assign in825_2 = {s742[0],s750[1],pp119[18]};
    CLA_3 KS_825(s825, c825, in825_1, in825_2);
    wire[0:0] s826, in826_1, in826_2;
    wire c826;
    assign in826_1 = {s743[0]};
    assign in826_2 = {s744[0]};
    Half_Adder KS_826(s826, c826, in826_1, in826_2);
    wire[1:0] s827, in827_1, in827_2;
    wire c827;
    assign in827_1 = {s745[0],s751[1]};
    assign in827_2 = {s746[0],s752[1]};
    CLA_2 KS_827(s827, c827, in827_1, in827_2);
    wire[0:0] s828, in828_1, in828_2;
    wire c828;
    assign in828_1 = {s747[0]};
    assign in828_2 = {s748[0]};
    Half_Adder KS_828(s828, c828, in828_1, in828_2);
    wire[3:0] s829, in829_1, in829_2;
    wire c829;
    assign in829_1 = {s749[0],s753[1],pp120[17],pp107[31]};
    assign in829_2 = {s750[0],s754[1],pp121[16],pp108[30]};
    CLA_4 KS_829(s829, c829, in829_1, in829_2);
    wire[0:0] s830, in830_1, in830_2;
    wire c830;
    assign in830_1 = {s751[0]};
    assign in830_2 = {s752[0]};
    Half_Adder KS_830(s830, c830, in830_1, in830_2);
    wire[1:0] s831, in831_1, in831_2;
    wire c831;
    assign in831_1 = {s754[0],s755[1]};
    assign in831_2 = {s755[0],s756[1]};
    CLA_2_c KS_831(s831, c831, in831_1, in831_2, s753[0]);
    wire[3:0] s832, in832_1, in832_2;
    wire c832;
    assign in832_1 = {pp12[127],pp13[127],pp14[127],pp15[127]};
    assign in832_2 = {pp13[126],pp14[126],pp15[126],pp16[126]};
    CLA_4 KS_832(s832, c832, in832_1, in832_2);
    wire[3:0] s833, in833_1, in833_2;
    wire c833;
    assign in833_1 = {pp14[125],pp15[125],pp16[125],pp17[125]};
    assign in833_2 = {pp15[124],pp16[124],pp17[124],pp18[124]};
    CLA_4 KS_833(s833, c833, in833_1, in833_2);
    wire[3:0] s834, in834_1, in834_2;
    wire c834;
    assign in834_1 = {pp16[123],pp17[123],pp18[123],pp19[123]};
    assign in834_2 = {pp17[122],pp18[122],pp19[122],pp20[122]};
    CLA_4 KS_834(s834, c834, in834_1, in834_2);
    wire[3:0] s835, in835_1, in835_2;
    wire c835;
    assign in835_1 = {pp18[121],pp19[121],pp20[121],pp21[121]};
    assign in835_2 = {pp19[120],pp20[120],pp21[120],pp22[120]};
    CLA_4 KS_835(s835, c835, in835_1, in835_2);
    wire[3:0] s836, in836_1, in836_2;
    wire c836;
    assign in836_1 = {pp20[119],pp21[119],pp22[119],pp23[119]};
    assign in836_2 = {pp21[118],pp22[118],pp23[118],pp24[118]};
    CLA_4 KS_836(s836, c836, in836_1, in836_2);
    wire[3:0] s837, in837_1, in837_2;
    wire c837;
    assign in837_1 = {pp22[117],pp23[117],pp24[117],pp25[117]};
    assign in837_2 = {pp23[116],pp24[116],pp25[116],pp26[116]};
    CLA_4 KS_837(s837, c837, in837_1, in837_2);
    wire[3:0] s838, in838_1, in838_2;
    wire c838;
    assign in838_1 = {pp24[115],pp25[115],pp26[115],pp27[115]};
    assign in838_2 = {pp25[114],pp26[114],pp27[114],pp28[114]};
    CLA_4 KS_838(s838, c838, in838_1, in838_2);
    wire[3:0] s839, in839_1, in839_2;
    wire c839;
    assign in839_1 = {pp26[113],pp27[113],pp28[113],pp29[113]};
    assign in839_2 = {pp27[112],pp28[112],pp29[112],pp30[112]};
    CLA_4 KS_839(s839, c839, in839_1, in839_2);
    wire[3:0] s840, in840_1, in840_2;
    wire c840;
    assign in840_1 = {pp28[111],pp29[111],pp30[111],pp31[111]};
    assign in840_2 = {pp29[110],pp30[110],pp31[110],pp32[110]};
    CLA_4 KS_840(s840, c840, in840_1, in840_2);
    wire[3:0] s841, in841_1, in841_2;
    wire c841;
    assign in841_1 = {pp30[109],pp31[109],pp32[109],pp33[109]};
    assign in841_2 = {pp31[108],pp32[108],pp33[108],pp34[108]};
    CLA_4 KS_841(s841, c841, in841_1, in841_2);
    wire[3:0] s842, in842_1, in842_2;
    wire c842;
    assign in842_1 = {pp32[107],pp33[107],pp34[107],pp35[107]};
    assign in842_2 = {pp33[106],pp34[106],pp35[106],pp36[106]};
    CLA_4 KS_842(s842, c842, in842_1, in842_2);
    wire[3:0] s843, in843_1, in843_2;
    wire c843;
    assign in843_1 = {pp34[105],pp35[105],pp36[105],pp37[105]};
    assign in843_2 = {pp35[104],pp36[104],pp37[104],pp38[104]};
    CLA_4 KS_843(s843, c843, in843_1, in843_2);
    wire[3:0] s844, in844_1, in844_2;
    wire c844;
    assign in844_1 = {pp36[103],pp37[103],pp38[103],pp39[103]};
    assign in844_2 = {pp37[102],pp38[102],pp39[102],pp40[102]};
    CLA_4 KS_844(s844, c844, in844_1, in844_2);
    wire[3:0] s845, in845_1, in845_2;
    wire c845;
    assign in845_1 = {pp38[101],pp39[101],pp40[101],pp41[101]};
    assign in845_2 = {pp39[100],pp40[100],pp41[100],pp42[100]};
    CLA_4 KS_845(s845, c845, in845_1, in845_2);
    wire[3:0] s846, in846_1, in846_2;
    wire c846;
    assign in846_1 = {pp40[99],pp41[99],pp42[99],pp43[99]};
    assign in846_2 = {pp41[98],pp42[98],pp43[98],pp44[98]};
    CLA_4 KS_846(s846, c846, in846_1, in846_2);
    wire[3:0] s847, in847_1, in847_2;
    wire c847;
    assign in847_1 = {pp42[97],pp43[97],pp44[97],pp45[97]};
    assign in847_2 = {pp43[96],pp44[96],pp45[96],pp46[96]};
    CLA_4 KS_847(s847, c847, in847_1, in847_2);
    wire[3:0] s848, in848_1, in848_2;
    wire c848;
    assign in848_1 = {pp44[95],pp45[95],pp46[95],pp47[95]};
    assign in848_2 = {pp45[94],pp46[94],pp47[94],pp48[94]};
    CLA_4 KS_848(s848, c848, in848_1, in848_2);
    wire[3:0] s849, in849_1, in849_2;
    wire c849;
    assign in849_1 = {pp46[93],pp47[93],pp48[93],pp49[93]};
    assign in849_2 = {pp47[92],pp48[92],pp49[92],pp50[92]};
    CLA_4 KS_849(s849, c849, in849_1, in849_2);
    wire[3:0] s850, in850_1, in850_2;
    wire c850;
    assign in850_1 = {pp48[91],pp49[91],pp50[91],pp51[91]};
    assign in850_2 = {pp49[90],pp50[90],pp51[90],pp52[90]};
    CLA_4 KS_850(s850, c850, in850_1, in850_2);
    wire[3:0] s851, in851_1, in851_2;
    wire c851;
    assign in851_1 = {pp50[89],pp51[89],pp52[89],pp53[89]};
    assign in851_2 = {pp51[88],pp52[88],pp53[88],pp54[88]};
    CLA_4 KS_851(s851, c851, in851_1, in851_2);
    wire[3:0] s852, in852_1, in852_2;
    wire c852;
    assign in852_1 = {pp52[87],pp53[87],pp54[87],pp55[87]};
    assign in852_2 = {pp53[86],pp54[86],pp55[86],pp56[86]};
    CLA_4 KS_852(s852, c852, in852_1, in852_2);
    wire[3:0] s853, in853_1, in853_2;
    wire c853;
    assign in853_1 = {pp54[85],pp55[85],pp56[85],pp57[85]};
    assign in853_2 = {pp55[84],pp56[84],pp57[84],pp58[84]};
    CLA_4 KS_853(s853, c853, in853_1, in853_2);
    wire[3:0] s854, in854_1, in854_2;
    wire c854;
    assign in854_1 = {pp56[83],pp57[83],pp58[83],pp59[83]};
    assign in854_2 = {pp57[82],pp58[82],pp59[82],pp60[82]};
    CLA_4 KS_854(s854, c854, in854_1, in854_2);
    wire[3:0] s855, in855_1, in855_2;
    wire c855;
    assign in855_1 = {pp58[81],pp59[81],pp60[81],pp61[81]};
    assign in855_2 = {pp59[80],pp60[80],pp61[80],pp62[80]};
    CLA_4 KS_855(s855, c855, in855_1, in855_2);
    wire[3:0] s856, in856_1, in856_2;
    wire c856;
    assign in856_1 = {pp60[79],pp61[79],pp62[79],pp63[79]};
    assign in856_2 = {pp61[78],pp62[78],pp63[78],pp64[78]};
    CLA_4 KS_856(s856, c856, in856_1, in856_2);
    wire[3:0] s857, in857_1, in857_2;
    wire c857;
    assign in857_1 = {pp62[77],pp63[77],pp64[77],pp65[77]};
    assign in857_2 = {pp63[76],pp64[76],pp65[76],pp66[76]};
    CLA_4 KS_857(s857, c857, in857_1, in857_2);
    wire[3:0] s858, in858_1, in858_2;
    wire c858;
    assign in858_1 = {pp64[75],pp65[75],pp66[75],pp67[75]};
    assign in858_2 = {pp65[74],pp66[74],pp67[74],pp68[74]};
    CLA_4 KS_858(s858, c858, in858_1, in858_2);
    wire[3:0] s859, in859_1, in859_2;
    wire c859;
    assign in859_1 = {pp66[73],pp67[73],pp68[73],pp69[73]};
    assign in859_2 = {pp67[72],pp68[72],pp69[72],pp70[72]};
    CLA_4 KS_859(s859, c859, in859_1, in859_2);
    wire[3:0] s860, in860_1, in860_2;
    wire c860;
    assign in860_1 = {pp68[71],pp69[71],pp70[71],pp71[71]};
    assign in860_2 = {pp69[70],pp70[70],pp71[70],pp72[70]};
    CLA_4 KS_860(s860, c860, in860_1, in860_2);
    wire[3:0] s861, in861_1, in861_2;
    wire c861;
    assign in861_1 = {pp70[69],pp71[69],pp72[69],pp73[69]};
    assign in861_2 = {pp71[68],pp72[68],pp73[68],pp74[68]};
    CLA_4 KS_861(s861, c861, in861_1, in861_2);
    wire[3:0] s862, in862_1, in862_2;
    wire c862;
    assign in862_1 = {pp72[67],pp73[67],pp74[67],pp75[67]};
    assign in862_2 = {pp73[66],pp74[66],pp75[66],pp76[66]};
    CLA_4 KS_862(s862, c862, in862_1, in862_2);
    wire[3:0] s863, in863_1, in863_2;
    wire c863;
    assign in863_1 = {pp74[65],pp75[65],pp76[65],pp77[65]};
    assign in863_2 = {pp75[64],pp76[64],pp77[64],pp78[64]};
    CLA_4 KS_863(s863, c863, in863_1, in863_2);
    wire[3:0] s864, in864_1, in864_2;
    wire c864;
    assign in864_1 = {pp76[63],pp77[63],pp78[63],pp79[63]};
    assign in864_2 = {pp77[62],pp78[62],pp79[62],pp80[62]};
    CLA_4 KS_864(s864, c864, in864_1, in864_2);
    wire[3:0] s865, in865_1, in865_2;
    wire c865;
    assign in865_1 = {pp78[61],pp79[61],pp80[61],pp81[61]};
    assign in865_2 = {pp79[60],pp80[60],pp81[60],pp82[60]};
    CLA_4 KS_865(s865, c865, in865_1, in865_2);
    wire[3:0] s866, in866_1, in866_2;
    wire c866;
    assign in866_1 = {pp80[59],pp81[59],pp82[59],pp83[59]};
    assign in866_2 = {pp81[58],pp82[58],pp83[58],pp84[58]};
    CLA_4 KS_866(s866, c866, in866_1, in866_2);
    wire[3:0] s867, in867_1, in867_2;
    wire c867;
    assign in867_1 = {pp82[57],pp83[57],pp84[57],pp85[57]};
    assign in867_2 = {pp83[56],pp84[56],pp85[56],pp86[56]};
    CLA_4 KS_867(s867, c867, in867_1, in867_2);
    wire[3:0] s868, in868_1, in868_2;
    wire c868;
    assign in868_1 = {pp84[55],pp85[55],pp86[55],pp87[55]};
    assign in868_2 = {pp85[54],pp86[54],pp87[54],pp88[54]};
    CLA_4 KS_868(s868, c868, in868_1, in868_2);
    wire[3:0] s869, in869_1, in869_2;
    wire c869;
    assign in869_1 = {pp86[53],pp87[53],pp88[53],pp89[53]};
    assign in869_2 = {pp87[52],pp88[52],pp89[52],pp90[52]};
    CLA_4 KS_869(s869, c869, in869_1, in869_2);
    wire[2:0] s870, in870_1, in870_2;
    wire c870;
    assign in870_1 = {pp88[51],pp89[51],pp90[51]};
    assign in870_2 = {pp89[50],pp90[50],pp91[50]};
    CLA_3 KS_870(s870, c870, in870_1, in870_2);
    wire[1:0] s871, in871_1, in871_2;
    wire c871;
    assign in871_1 = {pp90[49],pp91[49]};
    assign in871_2 = {pp91[48],pp92[48]};
    CLA_2 KS_871(s871, c871, in871_1, in871_2);
    wire[0:0] s872, in872_1, in872_2;
    wire c872;
    assign in872_1 = {pp92[47]};
    assign in872_2 = {pp93[46]};
    Half_Adder KS_872(s872, c872, in872_1, in872_2);
    wire[3:0] s873, in873_1, in873_2;
    wire c873;
    assign in873_1 = {pp94[45],pp93[47],pp92[49],pp91[51]};
    assign in873_2 = {pp95[44],pp94[46],pp93[48],pp92[50]};
    CLA_4 KS_873(s873, c873, in873_1, in873_2);
    wire[0:0] s874, in874_1, in874_2;
    wire c874;
    assign in874_1 = {pp96[43]};
    assign in874_2 = {pp97[42]};
    Half_Adder KS_874(s874, c874, in874_1, in874_2);
    wire[1:0] s875, in875_1, in875_2;
    wire c875;
    assign in875_1 = {pp98[41],pp95[45]};
    assign in875_2 = {pp99[40],pp96[44]};
    CLA_2 KS_875(s875, c875, in875_1, in875_2);
    wire[0:0] s876, in876_1, in876_2;
    wire c876;
    assign in876_1 = {pp100[39]};
    assign in876_2 = {pp101[38]};
    Half_Adder KS_876(s876, c876, in876_1, in876_2);
    wire[2:0] s877, in877_1, in877_2;
    wire c877;
    assign in877_1 = {pp102[37],pp97[43],pp94[47]};
    assign in877_2 = {pp103[36],pp98[42],pp95[46]};
    CLA_3 KS_877(s877, c877, in877_1, in877_2);
    wire[0:0] s878, in878_1, in878_2;
    wire c878;
    assign in878_1 = {pp104[35]};
    assign in878_2 = {pp105[34]};
    Half_Adder KS_878(s878, c878, in878_1, in878_2);
    wire[1:0] s879, in879_1, in879_2;
    wire c879;
    assign in879_1 = {pp106[33],pp99[41]};
    assign in879_2 = {pp107[32],pp100[40]};
    CLA_2 KS_879(s879, c879, in879_1, in879_2);
    wire[0:0] s880, in880_1, in880_2;
    wire c880;
    assign in880_1 = {pp108[31]};
    assign in880_2 = {pp109[30]};
    Half_Adder KS_880(s880, c880, in880_1, in880_2);
    wire[3:0] s881, in881_1, in881_2;
    wire c881;
    assign in881_1 = {pp110[29],pp101[39],pp96[45],pp93[49]};
    assign in881_2 = {pp111[28],pp102[38],pp97[44],pp94[48]};
    CLA_4 KS_881(s881, c881, in881_1, in881_2);
    wire[0:0] s882, in882_1, in882_2;
    wire c882;
    assign in882_1 = {pp112[27]};
    assign in882_2 = {pp113[26]};
    Half_Adder KS_882(s882, c882, in882_1, in882_2);
    wire[1:0] s883, in883_1, in883_2;
    wire c883;
    assign in883_1 = {pp114[25],pp103[37]};
    assign in883_2 = {pp115[24],pp104[36]};
    CLA_2 KS_883(s883, c883, in883_1, in883_2);
    wire[0:0] s884, in884_1, in884_2;
    wire c884;
    assign in884_1 = {pp116[23]};
    assign in884_2 = {pp117[22]};
    Half_Adder KS_884(s884, c884, in884_1, in884_2);
    wire[2:0] s885, in885_1, in885_2;
    wire c885;
    assign in885_1 = {pp118[21],pp105[35],pp98[43]};
    assign in885_2 = {pp119[20],pp106[34],pp99[42]};
    CLA_3 KS_885(s885, c885, in885_1, in885_2);
    wire[0:0] s886, in886_1, in886_2;
    wire c886;
    assign in886_1 = {pp120[19]};
    assign in886_2 = {pp121[18]};
    Half_Adder KS_886(s886, c886, in886_1, in886_2);
    wire[1:0] s887, in887_1, in887_2;
    wire c887;
    assign in887_1 = {pp122[17],pp107[33]};
    assign in887_2 = {pp123[16],pp108[32]};
    CLA_2 KS_887(s887, c887, in887_1, in887_2);
    wire[0:0] s888, in888_1, in888_2;
    wire c888;
    assign in888_1 = {pp124[15]};
    assign in888_2 = {pp125[14]};
    Half_Adder KS_888(s888, c888, in888_1, in888_2);
    wire[3:0] s889, in889_1, in889_2;
    wire c889;
    assign in889_1 = {pp126[13],pp109[31],pp100[41],pp95[47]};
    assign in889_2 = {pp127[12],pp110[30],pp101[40],pp96[46]};
    CLA_4 KS_889(s889, c889, in889_1, in889_2);
    wire[0:0] s890, in890_1, in890_2;
    wire c890;
    assign in890_1 = {c736};
    assign in890_2 = {c737};
    Half_Adder KS_890(s890, c890, in890_1, in890_2);
    wire[1:0] s891, in891_1, in891_2;
    wire c891;
    assign in891_1 = {c738,pp111[29]};
    assign in891_2 = {c739,pp112[28]};
    CLA_2 KS_891(s891, c891, in891_1, in891_2);
    wire[0:0] s892, in892_1, in892_2;
    wire c892;
    assign in892_1 = {c740};
    assign in892_2 = {c741};
    Half_Adder KS_892(s892, c892, in892_1, in892_2);
    wire[2:0] s893, in893_1, in893_2;
    wire c893;
    assign in893_1 = {c742,pp113[27],pp102[39]};
    assign in893_2 = {c743,pp114[26],pp103[38]};
    CLA_3 KS_893(s893, c893, in893_1, in893_2);
    wire[0:0] s894, in894_1, in894_2;
    wire c894;
    assign in894_1 = {c744};
    assign in894_2 = {c745};
    Half_Adder KS_894(s894, c894, in894_1, in894_2);
    wire[1:0] s895, in895_1, in895_2;
    wire c895;
    assign in895_1 = {c746,pp115[25]};
    assign in895_2 = {c747,pp116[24]};
    CLA_2 KS_895(s895, c895, in895_1, in895_2);
    wire[0:0] s896, in896_1, in896_2;
    wire c896;
    assign in896_1 = {c748};
    assign in896_2 = {c749};
    Half_Adder KS_896(s896, c896, in896_1, in896_2);
    wire[3:0] s897, in897_1, in897_2;
    wire c897;
    assign in897_1 = {c750,pp117[23],pp104[37],pp97[45]};
    assign in897_2 = {c751,pp118[22],pp105[36],pp98[44]};
    CLA_4 KS_897(s897, c897, in897_1, in897_2);
    wire[0:0] s898, in898_1, in898_2;
    wire c898;
    assign in898_1 = {c752};
    assign in898_2 = {c753};
    Half_Adder KS_898(s898, c898, in898_1, in898_2);
    wire[1:0] s899, in899_1, in899_2;
    wire c899;
    assign in899_1 = {c754,pp119[21]};
    assign in899_2 = {c755,pp120[20]};
    CLA_2 KS_899(s899, c899, in899_1, in899_2);
    wire[0:0] s900, in900_1, in900_2;
    wire c900;
    assign in900_1 = {c756};
    assign in900_2 = {c757};
    Half_Adder KS_900(s900, c900, in900_1, in900_2);
    wire[2:0] s901, in901_1, in901_2;
    wire c901;
    assign in901_1 = {c758,pp121[19],pp106[35]};
    assign in901_2 = {c759,pp122[18],pp107[34]};
    CLA_3 KS_901(s901, c901, in901_1, in901_2);
    wire[0:0] s902, in902_1, in902_2;
    wire c902;
    assign in902_1 = {c760};
    assign in902_2 = {c761};
    Half_Adder KS_902(s902, c902, in902_1, in902_2);
    wire[1:0] s903, in903_1, in903_2;
    wire c903;
    assign in903_1 = {c762,pp123[17]};
    assign in903_2 = {c763,pp124[16]};
    CLA_2 KS_903(s903, c903, in903_1, in903_2);
    wire[0:0] s904, in904_1, in904_2;
    wire c904;
    assign in904_1 = {c764};
    assign in904_2 = {c765};
    Half_Adder KS_904(s904, c904, in904_1, in904_2);
    wire[3:0] s905, in905_1, in905_2;
    wire c905;
    assign in905_1 = {c766,pp125[15],pp108[33],pp99[43]};
    assign in905_2 = {c767,pp126[14],pp109[32],pp100[42]};
    CLA_4 KS_905(s905, c905, in905_1, in905_2);
    wire[0:0] s906, in906_1, in906_2;
    wire c906;
    assign in906_1 = {c768};
    assign in906_2 = {c769};
    Half_Adder KS_906(s906, c906, in906_1, in906_2);
    wire[1:0] s907, in907_1, in907_2;
    wire c907;
    assign in907_1 = {c770,pp127[13]};
    assign in907_2 = {c771,s832[1]};
    CLA_2 KS_907(s907, c907, in907_1, in907_2);
    wire[0:0] s908, in908_1, in908_2;
    wire c908;
    assign in908_1 = {c772};
    assign in908_2 = {c773};
    Half_Adder KS_908(s908, c908, in908_1, in908_2);
    wire[2:0] s909, in909_1, in909_2;
    wire c909;
    assign in909_1 = {c774,s833[1],pp110[31]};
    assign in909_2 = {c775,s834[1],pp111[30]};
    CLA_3 KS_909(s909, c909, in909_1, in909_2);
    wire[0:0] s910, in910_1, in910_2;
    wire c910;
    assign in910_1 = {c776};
    assign in910_2 = {c777};
    Half_Adder KS_910(s910, c910, in910_1, in910_2);
    wire[1:0] s911, in911_1, in911_2;
    wire c911;
    assign in911_1 = {c781,s835[1]};
    assign in911_2 = {c789,s836[1]};
    CLA_2 KS_911(s911, c911, in911_1, in911_2);
    wire[0:0] s912, in912_1, in912_2;
    wire c912;
    assign in912_1 = {c797};
    assign in912_2 = {c805};
    Half_Adder KS_912(s912, c912, in912_1, in912_2);
    wire[3:0] s913, in913_1, in913_2;
    wire c913;
    assign in913_1 = {c813,s837[1],pp112[29],pp101[41]};
    assign in913_2 = {c821,s838[1],pp113[28],pp102[40]};
    CLA_4 KS_913(s913, c913, in913_1, in913_2);
    wire[0:0] s914, in914_1, in914_2;
    wire c914;
    assign in914_1 = {c829};
    assign in914_2 = {s832[0]};
    Half_Adder KS_914(s914, c914, in914_1, in914_2);
    wire[1:0] s915, in915_1, in915_2;
    wire c915;
    assign in915_1 = {s833[0],s839[1]};
    assign in915_2 = {s834[0],s840[1]};
    CLA_2 KS_915(s915, c915, in915_1, in915_2);
    wire[0:0] s916, in916_1, in916_2;
    wire c916;
    assign in916_1 = {s835[0]};
    assign in916_2 = {s836[0]};
    Half_Adder KS_916(s916, c916, in916_1, in916_2);
    wire[2:0] s917, in917_1, in917_2;
    wire c917;
    assign in917_1 = {s837[0],s841[1],pp114[27]};
    assign in917_2 = {s838[0],s842[1],pp115[26]};
    CLA_3 KS_917(s917, c917, in917_1, in917_2);
    wire[0:0] s918, in918_1, in918_2;
    wire c918;
    assign in918_1 = {s839[0]};
    assign in918_2 = {s840[0]};
    Half_Adder KS_918(s918, c918, in918_1, in918_2);
    wire[1:0] s919, in919_1, in919_2;
    wire c919;
    assign in919_1 = {s842[0],s843[1]};
    assign in919_2 = {s843[0],s844[1]};
    CLA_2_c KS_919(s919, c919, in919_1, in919_2, s841[0]);
    wire[3:0] s920, in920_1, in920_2;
    wire c920;
    assign in920_1 = {pp16[127],pp17[127],pp18[127],pp19[127]};
    assign in920_2 = {pp17[126],pp18[126],pp19[126],pp20[126]};
    CLA_4 KS_920(s920, c920, in920_1, in920_2);
    wire[3:0] s921, in921_1, in921_2;
    wire c921;
    assign in921_1 = {pp18[125],pp19[125],pp20[125],pp21[125]};
    assign in921_2 = {pp19[124],pp20[124],pp21[124],pp22[124]};
    CLA_4 KS_921(s921, c921, in921_1, in921_2);
    wire[3:0] s922, in922_1, in922_2;
    wire c922;
    assign in922_1 = {pp20[123],pp21[123],pp22[123],pp23[123]};
    assign in922_2 = {pp21[122],pp22[122],pp23[122],pp24[122]};
    CLA_4 KS_922(s922, c922, in922_1, in922_2);
    wire[3:0] s923, in923_1, in923_2;
    wire c923;
    assign in923_1 = {pp22[121],pp23[121],pp24[121],pp25[121]};
    assign in923_2 = {pp23[120],pp24[120],pp25[120],pp26[120]};
    CLA_4 KS_923(s923, c923, in923_1, in923_2);
    wire[3:0] s924, in924_1, in924_2;
    wire c924;
    assign in924_1 = {pp24[119],pp25[119],pp26[119],pp27[119]};
    assign in924_2 = {pp25[118],pp26[118],pp27[118],pp28[118]};
    CLA_4 KS_924(s924, c924, in924_1, in924_2);
    wire[3:0] s925, in925_1, in925_2;
    wire c925;
    assign in925_1 = {pp26[117],pp27[117],pp28[117],pp29[117]};
    assign in925_2 = {pp27[116],pp28[116],pp29[116],pp30[116]};
    CLA_4 KS_925(s925, c925, in925_1, in925_2);
    wire[3:0] s926, in926_1, in926_2;
    wire c926;
    assign in926_1 = {pp28[115],pp29[115],pp30[115],pp31[115]};
    assign in926_2 = {pp29[114],pp30[114],pp31[114],pp32[114]};
    CLA_4 KS_926(s926, c926, in926_1, in926_2);
    wire[3:0] s927, in927_1, in927_2;
    wire c927;
    assign in927_1 = {pp30[113],pp31[113],pp32[113],pp33[113]};
    assign in927_2 = {pp31[112],pp32[112],pp33[112],pp34[112]};
    CLA_4 KS_927(s927, c927, in927_1, in927_2);
    wire[3:0] s928, in928_1, in928_2;
    wire c928;
    assign in928_1 = {pp32[111],pp33[111],pp34[111],pp35[111]};
    assign in928_2 = {pp33[110],pp34[110],pp35[110],pp36[110]};
    CLA_4 KS_928(s928, c928, in928_1, in928_2);
    wire[3:0] s929, in929_1, in929_2;
    wire c929;
    assign in929_1 = {pp34[109],pp35[109],pp36[109],pp37[109]};
    assign in929_2 = {pp35[108],pp36[108],pp37[108],pp38[108]};
    CLA_4 KS_929(s929, c929, in929_1, in929_2);
    wire[3:0] s930, in930_1, in930_2;
    wire c930;
    assign in930_1 = {pp36[107],pp37[107],pp38[107],pp39[107]};
    assign in930_2 = {pp37[106],pp38[106],pp39[106],pp40[106]};
    CLA_4 KS_930(s930, c930, in930_1, in930_2);
    wire[3:0] s931, in931_1, in931_2;
    wire c931;
    assign in931_1 = {pp38[105],pp39[105],pp40[105],pp41[105]};
    assign in931_2 = {pp39[104],pp40[104],pp41[104],pp42[104]};
    CLA_4 KS_931(s931, c931, in931_1, in931_2);
    wire[3:0] s932, in932_1, in932_2;
    wire c932;
    assign in932_1 = {pp40[103],pp41[103],pp42[103],pp43[103]};
    assign in932_2 = {pp41[102],pp42[102],pp43[102],pp44[102]};
    CLA_4 KS_932(s932, c932, in932_1, in932_2);
    wire[3:0] s933, in933_1, in933_2;
    wire c933;
    assign in933_1 = {pp42[101],pp43[101],pp44[101],pp45[101]};
    assign in933_2 = {pp43[100],pp44[100],pp45[100],pp46[100]};
    CLA_4 KS_933(s933, c933, in933_1, in933_2);
    wire[3:0] s934, in934_1, in934_2;
    wire c934;
    assign in934_1 = {pp44[99],pp45[99],pp46[99],pp47[99]};
    assign in934_2 = {pp45[98],pp46[98],pp47[98],pp48[98]};
    CLA_4 KS_934(s934, c934, in934_1, in934_2);
    wire[3:0] s935, in935_1, in935_2;
    wire c935;
    assign in935_1 = {pp46[97],pp47[97],pp48[97],pp49[97]};
    assign in935_2 = {pp47[96],pp48[96],pp49[96],pp50[96]};
    CLA_4 KS_935(s935, c935, in935_1, in935_2);
    wire[3:0] s936, in936_1, in936_2;
    wire c936;
    assign in936_1 = {pp48[95],pp49[95],pp50[95],pp51[95]};
    assign in936_2 = {pp49[94],pp50[94],pp51[94],pp52[94]};
    CLA_4 KS_936(s936, c936, in936_1, in936_2);
    wire[3:0] s937, in937_1, in937_2;
    wire c937;
    assign in937_1 = {pp50[93],pp51[93],pp52[93],pp53[93]};
    assign in937_2 = {pp51[92],pp52[92],pp53[92],pp54[92]};
    CLA_4 KS_937(s937, c937, in937_1, in937_2);
    wire[3:0] s938, in938_1, in938_2;
    wire c938;
    assign in938_1 = {pp52[91],pp53[91],pp54[91],pp55[91]};
    assign in938_2 = {pp53[90],pp54[90],pp55[90],pp56[90]};
    CLA_4 KS_938(s938, c938, in938_1, in938_2);
    wire[3:0] s939, in939_1, in939_2;
    wire c939;
    assign in939_1 = {pp54[89],pp55[89],pp56[89],pp57[89]};
    assign in939_2 = {pp55[88],pp56[88],pp57[88],pp58[88]};
    CLA_4 KS_939(s939, c939, in939_1, in939_2);
    wire[3:0] s940, in940_1, in940_2;
    wire c940;
    assign in940_1 = {pp56[87],pp57[87],pp58[87],pp59[87]};
    assign in940_2 = {pp57[86],pp58[86],pp59[86],pp60[86]};
    CLA_4 KS_940(s940, c940, in940_1, in940_2);
    wire[3:0] s941, in941_1, in941_2;
    wire c941;
    assign in941_1 = {pp58[85],pp59[85],pp60[85],pp61[85]};
    assign in941_2 = {pp59[84],pp60[84],pp61[84],pp62[84]};
    CLA_4 KS_941(s941, c941, in941_1, in941_2);
    wire[3:0] s942, in942_1, in942_2;
    wire c942;
    assign in942_1 = {pp60[83],pp61[83],pp62[83],pp63[83]};
    assign in942_2 = {pp61[82],pp62[82],pp63[82],pp64[82]};
    CLA_4 KS_942(s942, c942, in942_1, in942_2);
    wire[3:0] s943, in943_1, in943_2;
    wire c943;
    assign in943_1 = {pp62[81],pp63[81],pp64[81],pp65[81]};
    assign in943_2 = {pp63[80],pp64[80],pp65[80],pp66[80]};
    CLA_4 KS_943(s943, c943, in943_1, in943_2);
    wire[3:0] s944, in944_1, in944_2;
    wire c944;
    assign in944_1 = {pp64[79],pp65[79],pp66[79],pp67[79]};
    assign in944_2 = {pp65[78],pp66[78],pp67[78],pp68[78]};
    CLA_4 KS_944(s944, c944, in944_1, in944_2);
    wire[3:0] s945, in945_1, in945_2;
    wire c945;
    assign in945_1 = {pp66[77],pp67[77],pp68[77],pp69[77]};
    assign in945_2 = {pp67[76],pp68[76],pp69[76],pp70[76]};
    CLA_4 KS_945(s945, c945, in945_1, in945_2);
    wire[3:0] s946, in946_1, in946_2;
    wire c946;
    assign in946_1 = {pp68[75],pp69[75],pp70[75],pp71[75]};
    assign in946_2 = {pp69[74],pp70[74],pp71[74],pp72[74]};
    CLA_4 KS_946(s946, c946, in946_1, in946_2);
    wire[3:0] s947, in947_1, in947_2;
    wire c947;
    assign in947_1 = {pp70[73],pp71[73],pp72[73],pp73[73]};
    assign in947_2 = {pp71[72],pp72[72],pp73[72],pp74[72]};
    CLA_4 KS_947(s947, c947, in947_1, in947_2);
    wire[3:0] s948, in948_1, in948_2;
    wire c948;
    assign in948_1 = {pp72[71],pp73[71],pp74[71],pp75[71]};
    assign in948_2 = {pp73[70],pp74[70],pp75[70],pp76[70]};
    CLA_4 KS_948(s948, c948, in948_1, in948_2);
    wire[3:0] s949, in949_1, in949_2;
    wire c949;
    assign in949_1 = {pp74[69],pp75[69],pp76[69],pp77[69]};
    assign in949_2 = {pp75[68],pp76[68],pp77[68],pp78[68]};
    CLA_4 KS_949(s949, c949, in949_1, in949_2);
    wire[3:0] s950, in950_1, in950_2;
    wire c950;
    assign in950_1 = {pp76[67],pp77[67],pp78[67],pp79[67]};
    assign in950_2 = {pp77[66],pp78[66],pp79[66],pp80[66]};
    CLA_4 KS_950(s950, c950, in950_1, in950_2);
    wire[3:0] s951, in951_1, in951_2;
    wire c951;
    assign in951_1 = {pp78[65],pp79[65],pp80[65],pp81[65]};
    assign in951_2 = {pp79[64],pp80[64],pp81[64],pp82[64]};
    CLA_4 KS_951(s951, c951, in951_1, in951_2);
    wire[3:0] s952, in952_1, in952_2;
    wire c952;
    assign in952_1 = {pp80[63],pp81[63],pp82[63],pp83[63]};
    assign in952_2 = {pp81[62],pp82[62],pp83[62],pp84[62]};
    CLA_4 KS_952(s952, c952, in952_1, in952_2);
    wire[3:0] s953, in953_1, in953_2;
    wire c953;
    assign in953_1 = {pp82[61],pp83[61],pp84[61],pp85[61]};
    assign in953_2 = {pp83[60],pp84[60],pp85[60],pp86[60]};
    CLA_4 KS_953(s953, c953, in953_1, in953_2);
    wire[2:0] s954, in954_1, in954_2;
    wire c954;
    assign in954_1 = {pp84[59],pp85[59],pp86[59]};
    assign in954_2 = {pp85[58],pp86[58],pp87[58]};
    CLA_3 KS_954(s954, c954, in954_1, in954_2);
    wire[1:0] s955, in955_1, in955_2;
    wire c955;
    assign in955_1 = {pp86[57],pp87[57]};
    assign in955_2 = {pp87[56],pp88[56]};
    CLA_2 KS_955(s955, c955, in955_1, in955_2);
    wire[0:0] s956, in956_1, in956_2;
    wire c956;
    assign in956_1 = {pp88[55]};
    assign in956_2 = {pp89[54]};
    Half_Adder KS_956(s956, c956, in956_1, in956_2);
    wire[3:0] s957, in957_1, in957_2;
    wire c957;
    assign in957_1 = {pp90[53],pp89[55],pp88[57],pp87[59]};
    assign in957_2 = {pp91[52],pp90[54],pp89[56],pp88[58]};
    CLA_4 KS_957(s957, c957, in957_1, in957_2);
    wire[0:0] s958, in958_1, in958_2;
    wire c958;
    assign in958_1 = {pp92[51]};
    assign in958_2 = {pp93[50]};
    Half_Adder KS_958(s958, c958, in958_1, in958_2);
    wire[1:0] s959, in959_1, in959_2;
    wire c959;
    assign in959_1 = {pp94[49],pp91[53]};
    assign in959_2 = {pp95[48],pp92[52]};
    CLA_2 KS_959(s959, c959, in959_1, in959_2);
    wire[0:0] s960, in960_1, in960_2;
    wire c960;
    assign in960_1 = {pp96[47]};
    assign in960_2 = {pp97[46]};
    Half_Adder KS_960(s960, c960, in960_1, in960_2);
    wire[2:0] s961, in961_1, in961_2;
    wire c961;
    assign in961_1 = {pp98[45],pp93[51],pp90[55]};
    assign in961_2 = {pp99[44],pp94[50],pp91[54]};
    CLA_3 KS_961(s961, c961, in961_1, in961_2);
    wire[0:0] s962, in962_1, in962_2;
    wire c962;
    assign in962_1 = {pp100[43]};
    assign in962_2 = {pp101[42]};
    Half_Adder KS_962(s962, c962, in962_1, in962_2);
    wire[1:0] s963, in963_1, in963_2;
    wire c963;
    assign in963_1 = {pp102[41],pp95[49]};
    assign in963_2 = {pp103[40],pp96[48]};
    CLA_2 KS_963(s963, c963, in963_1, in963_2);
    wire[0:0] s964, in964_1, in964_2;
    wire c964;
    assign in964_1 = {pp104[39]};
    assign in964_2 = {pp105[38]};
    Half_Adder KS_964(s964, c964, in964_1, in964_2);
    wire[3:0] s965, in965_1, in965_2;
    wire c965;
    assign in965_1 = {pp106[37],pp97[47],pp92[53],pp89[57]};
    assign in965_2 = {pp107[36],pp98[46],pp93[52],pp90[56]};
    CLA_4 KS_965(s965, c965, in965_1, in965_2);
    wire[0:0] s966, in966_1, in966_2;
    wire c966;
    assign in966_1 = {pp108[35]};
    assign in966_2 = {pp109[34]};
    Half_Adder KS_966(s966, c966, in966_1, in966_2);
    wire[1:0] s967, in967_1, in967_2;
    wire c967;
    assign in967_1 = {pp110[33],pp99[45]};
    assign in967_2 = {pp111[32],pp100[44]};
    CLA_2 KS_967(s967, c967, in967_1, in967_2);
    wire[0:0] s968, in968_1, in968_2;
    wire c968;
    assign in968_1 = {pp112[31]};
    assign in968_2 = {pp113[30]};
    Half_Adder KS_968(s968, c968, in968_1, in968_2);
    wire[2:0] s969, in969_1, in969_2;
    wire c969;
    assign in969_1 = {pp114[29],pp101[43],pp94[51]};
    assign in969_2 = {pp115[28],pp102[42],pp95[50]};
    CLA_3 KS_969(s969, c969, in969_1, in969_2);
    wire[0:0] s970, in970_1, in970_2;
    wire c970;
    assign in970_1 = {pp116[27]};
    assign in970_2 = {pp117[26]};
    Half_Adder KS_970(s970, c970, in970_1, in970_2);
    wire[1:0] s971, in971_1, in971_2;
    wire c971;
    assign in971_1 = {pp118[25],pp103[41]};
    assign in971_2 = {pp119[24],pp104[40]};
    CLA_2 KS_971(s971, c971, in971_1, in971_2);
    wire[0:0] s972, in972_1, in972_2;
    wire c972;
    assign in972_1 = {pp120[23]};
    assign in972_2 = {pp121[22]};
    Half_Adder KS_972(s972, c972, in972_1, in972_2);
    wire[3:0] s973, in973_1, in973_2;
    wire c973;
    assign in973_1 = {pp122[21],pp105[39],pp96[49],pp91[55]};
    assign in973_2 = {pp123[20],pp106[38],pp97[48],pp92[54]};
    CLA_4 KS_973(s973, c973, in973_1, in973_2);
    wire[0:0] s974, in974_1, in974_2;
    wire c974;
    assign in974_1 = {pp124[19]};
    assign in974_2 = {pp125[18]};
    Half_Adder KS_974(s974, c974, in974_1, in974_2);
    wire[1:0] s975, in975_1, in975_2;
    wire c975;
    assign in975_1 = {pp126[17],pp107[37]};
    assign in975_2 = {pp127[16],pp108[36]};
    CLA_2 KS_975(s975, c975, in975_1, in975_2);
    wire[0:0] s976, in976_1, in976_2;
    wire c976;
    assign in976_1 = {c832};
    assign in976_2 = {c833};
    Half_Adder KS_976(s976, c976, in976_1, in976_2);
    wire[2:0] s977, in977_1, in977_2;
    wire c977;
    assign in977_1 = {c834,pp109[35],pp98[47]};
    assign in977_2 = {c835,pp110[34],pp99[46]};
    CLA_3 KS_977(s977, c977, in977_1, in977_2);
    wire[0:0] s978, in978_1, in978_2;
    wire c978;
    assign in978_1 = {c836};
    assign in978_2 = {c837};
    Half_Adder KS_978(s978, c978, in978_1, in978_2);
    wire[1:0] s979, in979_1, in979_2;
    wire c979;
    assign in979_1 = {c838,pp111[33]};
    assign in979_2 = {c839,pp112[32]};
    CLA_2 KS_979(s979, c979, in979_1, in979_2);
    wire[0:0] s980, in980_1, in980_2;
    wire c980;
    assign in980_1 = {c840};
    assign in980_2 = {c841};
    Half_Adder KS_980(s980, c980, in980_1, in980_2);
    wire[3:0] s981, in981_1, in981_2;
    wire c981;
    assign in981_1 = {c842,pp113[31],pp100[45],pp93[53]};
    assign in981_2 = {c843,pp114[30],pp101[44],pp94[52]};
    CLA_4 KS_981(s981, c981, in981_1, in981_2);
    wire[0:0] s982, in982_1, in982_2;
    wire c982;
    assign in982_1 = {c844};
    assign in982_2 = {c845};
    Half_Adder KS_982(s982, c982, in982_1, in982_2);
    wire[1:0] s983, in983_1, in983_2;
    wire c983;
    assign in983_1 = {c846,pp115[29]};
    assign in983_2 = {c847,pp116[28]};
    CLA_2 KS_983(s983, c983, in983_1, in983_2);
    wire[0:0] s984, in984_1, in984_2;
    wire c984;
    assign in984_1 = {c848};
    assign in984_2 = {c849};
    Half_Adder KS_984(s984, c984, in984_1, in984_2);
    wire[2:0] s985, in985_1, in985_2;
    wire c985;
    assign in985_1 = {c850,pp117[27],pp102[43]};
    assign in985_2 = {c851,pp118[26],pp103[42]};
    CLA_3 KS_985(s985, c985, in985_1, in985_2);
    wire[0:0] s986, in986_1, in986_2;
    wire c986;
    assign in986_1 = {c852};
    assign in986_2 = {c853};
    Half_Adder KS_986(s986, c986, in986_1, in986_2);
    wire[1:0] s987, in987_1, in987_2;
    wire c987;
    assign in987_1 = {c854,pp119[25]};
    assign in987_2 = {c855,pp120[24]};
    CLA_2 KS_987(s987, c987, in987_1, in987_2);
    wire[0:0] s988, in988_1, in988_2;
    wire c988;
    assign in988_1 = {c856};
    assign in988_2 = {c857};
    Half_Adder KS_988(s988, c988, in988_1, in988_2);
    wire[3:0] s989, in989_1, in989_2;
    wire c989;
    assign in989_1 = {c858,pp121[23],pp104[41],pp95[51]};
    assign in989_2 = {c859,pp122[22],pp105[40],pp96[50]};
    CLA_4 KS_989(s989, c989, in989_1, in989_2);
    wire[0:0] s990, in990_1, in990_2;
    wire c990;
    assign in990_1 = {c860};
    assign in990_2 = {c861};
    Half_Adder KS_990(s990, c990, in990_1, in990_2);
    wire[1:0] s991, in991_1, in991_2;
    wire c991;
    assign in991_1 = {c862,pp123[21]};
    assign in991_2 = {c863,pp124[20]};
    CLA_2 KS_991(s991, c991, in991_1, in991_2);
    wire[0:0] s992, in992_1, in992_2;
    wire c992;
    assign in992_1 = {c864};
    assign in992_2 = {c865};
    Half_Adder KS_992(s992, c992, in992_1, in992_2);
    wire[2:0] s993, in993_1, in993_2;
    wire c993;
    assign in993_1 = {c866,pp125[19],pp106[39]};
    assign in993_2 = {c867,pp126[18],pp107[38]};
    CLA_3 KS_993(s993, c993, in993_1, in993_2);
    wire[0:0] s994, in994_1, in994_2;
    wire c994;
    assign in994_1 = {c868};
    assign in994_2 = {c869};
    Half_Adder KS_994(s994, c994, in994_1, in994_2);
    wire[1:0] s995, in995_1, in995_2;
    wire c995;
    assign in995_1 = {c873,pp127[17]};
    assign in995_2 = {c881,s920[1]};
    CLA_2 KS_995(s995, c995, in995_1, in995_2);
    wire[0:0] s996, in996_1, in996_2;
    wire c996;
    assign in996_1 = {c889};
    assign in996_2 = {c897};
    Half_Adder KS_996(s996, c996, in996_1, in996_2);
    wire[3:0] s997, in997_1, in997_2;
    wire c997;
    assign in997_1 = {c905,s921[1],pp108[37],pp97[49]};
    assign in997_2 = {c913,s922[1],pp109[36],pp98[48]};
    CLA_4 KS_997(s997, c997, in997_1, in997_2);
    wire[0:0] s998, in998_1, in998_2;
    wire c998;
    assign in998_1 = {s921[0]};
    assign in998_2 = {s922[0]};
    Full_Adder KS_998(s998, c998, in998_1, in998_2, s920[0]);
    wire[3:0] s999, in999_1, in999_2;
    wire c999;
    assign in999_1 = {pp20[127],pp21[127],pp22[127],pp23[127]};
    assign in999_2 = {pp21[126],pp22[126],pp23[126],pp24[126]};
    CLA_4 KS_999(s999, c999, in999_1, in999_2);
    wire[3:0] s1000, in1000_1, in1000_2;
    wire c1000;
    assign in1000_1 = {pp22[125],pp23[125],pp24[125],pp25[125]};
    assign in1000_2 = {pp23[124],pp24[124],pp25[124],pp26[124]};
    CLA_4 KS_1000(s1000, c1000, in1000_1, in1000_2);
    wire[3:0] s1001, in1001_1, in1001_2;
    wire c1001;
    assign in1001_1 = {pp24[123],pp25[123],pp26[123],pp27[123]};
    assign in1001_2 = {pp25[122],pp26[122],pp27[122],pp28[122]};
    CLA_4 KS_1001(s1001, c1001, in1001_1, in1001_2);
    wire[3:0] s1002, in1002_1, in1002_2;
    wire c1002;
    assign in1002_1 = {pp26[121],pp27[121],pp28[121],pp29[121]};
    assign in1002_2 = {pp27[120],pp28[120],pp29[120],pp30[120]};
    CLA_4 KS_1002(s1002, c1002, in1002_1, in1002_2);
    wire[3:0] s1003, in1003_1, in1003_2;
    wire c1003;
    assign in1003_1 = {pp28[119],pp29[119],pp30[119],pp31[119]};
    assign in1003_2 = {pp29[118],pp30[118],pp31[118],pp32[118]};
    CLA_4 KS_1003(s1003, c1003, in1003_1, in1003_2);
    wire[3:0] s1004, in1004_1, in1004_2;
    wire c1004;
    assign in1004_1 = {pp30[117],pp31[117],pp32[117],pp33[117]};
    assign in1004_2 = {pp31[116],pp32[116],pp33[116],pp34[116]};
    CLA_4 KS_1004(s1004, c1004, in1004_1, in1004_2);
    wire[3:0] s1005, in1005_1, in1005_2;
    wire c1005;
    assign in1005_1 = {pp32[115],pp33[115],pp34[115],pp35[115]};
    assign in1005_2 = {pp33[114],pp34[114],pp35[114],pp36[114]};
    CLA_4 KS_1005(s1005, c1005, in1005_1, in1005_2);
    wire[3:0] s1006, in1006_1, in1006_2;
    wire c1006;
    assign in1006_1 = {pp34[113],pp35[113],pp36[113],pp37[113]};
    assign in1006_2 = {pp35[112],pp36[112],pp37[112],pp38[112]};
    CLA_4 KS_1006(s1006, c1006, in1006_1, in1006_2);
    wire[3:0] s1007, in1007_1, in1007_2;
    wire c1007;
    assign in1007_1 = {pp36[111],pp37[111],pp38[111],pp39[111]};
    assign in1007_2 = {pp37[110],pp38[110],pp39[110],pp40[110]};
    CLA_4 KS_1007(s1007, c1007, in1007_1, in1007_2);
    wire[3:0] s1008, in1008_1, in1008_2;
    wire c1008;
    assign in1008_1 = {pp38[109],pp39[109],pp40[109],pp41[109]};
    assign in1008_2 = {pp39[108],pp40[108],pp41[108],pp42[108]};
    CLA_4 KS_1008(s1008, c1008, in1008_1, in1008_2);
    wire[3:0] s1009, in1009_1, in1009_2;
    wire c1009;
    assign in1009_1 = {pp40[107],pp41[107],pp42[107],pp43[107]};
    assign in1009_2 = {pp41[106],pp42[106],pp43[106],pp44[106]};
    CLA_4 KS_1009(s1009, c1009, in1009_1, in1009_2);
    wire[3:0] s1010, in1010_1, in1010_2;
    wire c1010;
    assign in1010_1 = {pp42[105],pp43[105],pp44[105],pp45[105]};
    assign in1010_2 = {pp43[104],pp44[104],pp45[104],pp46[104]};
    CLA_4 KS_1010(s1010, c1010, in1010_1, in1010_2);
    wire[3:0] s1011, in1011_1, in1011_2;
    wire c1011;
    assign in1011_1 = {pp44[103],pp45[103],pp46[103],pp47[103]};
    assign in1011_2 = {pp45[102],pp46[102],pp47[102],pp48[102]};
    CLA_4 KS_1011(s1011, c1011, in1011_1, in1011_2);
    wire[3:0] s1012, in1012_1, in1012_2;
    wire c1012;
    assign in1012_1 = {pp46[101],pp47[101],pp48[101],pp49[101]};
    assign in1012_2 = {pp47[100],pp48[100],pp49[100],pp50[100]};
    CLA_4 KS_1012(s1012, c1012, in1012_1, in1012_2);
    wire[3:0] s1013, in1013_1, in1013_2;
    wire c1013;
    assign in1013_1 = {pp48[99],pp49[99],pp50[99],pp51[99]};
    assign in1013_2 = {pp49[98],pp50[98],pp51[98],pp52[98]};
    CLA_4 KS_1013(s1013, c1013, in1013_1, in1013_2);
    wire[3:0] s1014, in1014_1, in1014_2;
    wire c1014;
    assign in1014_1 = {pp50[97],pp51[97],pp52[97],pp53[97]};
    assign in1014_2 = {pp51[96],pp52[96],pp53[96],pp54[96]};
    CLA_4 KS_1014(s1014, c1014, in1014_1, in1014_2);
    wire[3:0] s1015, in1015_1, in1015_2;
    wire c1015;
    assign in1015_1 = {pp52[95],pp53[95],pp54[95],pp55[95]};
    assign in1015_2 = {pp53[94],pp54[94],pp55[94],pp56[94]};
    CLA_4 KS_1015(s1015, c1015, in1015_1, in1015_2);
    wire[3:0] s1016, in1016_1, in1016_2;
    wire c1016;
    assign in1016_1 = {pp54[93],pp55[93],pp56[93],pp57[93]};
    assign in1016_2 = {pp55[92],pp56[92],pp57[92],pp58[92]};
    CLA_4 KS_1016(s1016, c1016, in1016_1, in1016_2);
    wire[3:0] s1017, in1017_1, in1017_2;
    wire c1017;
    assign in1017_1 = {pp56[91],pp57[91],pp58[91],pp59[91]};
    assign in1017_2 = {pp57[90],pp58[90],pp59[90],pp60[90]};
    CLA_4 KS_1017(s1017, c1017, in1017_1, in1017_2);
    wire[3:0] s1018, in1018_1, in1018_2;
    wire c1018;
    assign in1018_1 = {pp58[89],pp59[89],pp60[89],pp61[89]};
    assign in1018_2 = {pp59[88],pp60[88],pp61[88],pp62[88]};
    CLA_4 KS_1018(s1018, c1018, in1018_1, in1018_2);
    wire[3:0] s1019, in1019_1, in1019_2;
    wire c1019;
    assign in1019_1 = {pp60[87],pp61[87],pp62[87],pp63[87]};
    assign in1019_2 = {pp61[86],pp62[86],pp63[86],pp64[86]};
    CLA_4 KS_1019(s1019, c1019, in1019_1, in1019_2);
    wire[3:0] s1020, in1020_1, in1020_2;
    wire c1020;
    assign in1020_1 = {pp62[85],pp63[85],pp64[85],pp65[85]};
    assign in1020_2 = {pp63[84],pp64[84],pp65[84],pp66[84]};
    CLA_4 KS_1020(s1020, c1020, in1020_1, in1020_2);
    wire[3:0] s1021, in1021_1, in1021_2;
    wire c1021;
    assign in1021_1 = {pp64[83],pp65[83],pp66[83],pp67[83]};
    assign in1021_2 = {pp65[82],pp66[82],pp67[82],pp68[82]};
    CLA_4 KS_1021(s1021, c1021, in1021_1, in1021_2);
    wire[3:0] s1022, in1022_1, in1022_2;
    wire c1022;
    assign in1022_1 = {pp66[81],pp67[81],pp68[81],pp69[81]};
    assign in1022_2 = {pp67[80],pp68[80],pp69[80],pp70[80]};
    CLA_4 KS_1022(s1022, c1022, in1022_1, in1022_2);
    wire[3:0] s1023, in1023_1, in1023_2;
    wire c1023;
    assign in1023_1 = {pp68[79],pp69[79],pp70[79],pp71[79]};
    assign in1023_2 = {pp69[78],pp70[78],pp71[78],pp72[78]};
    CLA_4 KS_1023(s1023, c1023, in1023_1, in1023_2);
    wire[3:0] s1024, in1024_1, in1024_2;
    wire c1024;
    assign in1024_1 = {pp70[77],pp71[77],pp72[77],pp73[77]};
    assign in1024_2 = {pp71[76],pp72[76],pp73[76],pp74[76]};
    CLA_4 KS_1024(s1024, c1024, in1024_1, in1024_2);
    wire[3:0] s1025, in1025_1, in1025_2;
    wire c1025;
    assign in1025_1 = {pp72[75],pp73[75],pp74[75],pp75[75]};
    assign in1025_2 = {pp73[74],pp74[74],pp75[74],pp76[74]};
    CLA_4 KS_1025(s1025, c1025, in1025_1, in1025_2);
    wire[3:0] s1026, in1026_1, in1026_2;
    wire c1026;
    assign in1026_1 = {pp74[73],pp75[73],pp76[73],pp77[73]};
    assign in1026_2 = {pp75[72],pp76[72],pp77[72],pp78[72]};
    CLA_4 KS_1026(s1026, c1026, in1026_1, in1026_2);
    wire[3:0] s1027, in1027_1, in1027_2;
    wire c1027;
    assign in1027_1 = {pp76[71],pp77[71],pp78[71],pp79[71]};
    assign in1027_2 = {pp77[70],pp78[70],pp79[70],pp80[70]};
    CLA_4 KS_1027(s1027, c1027, in1027_1, in1027_2);
    wire[3:0] s1028, in1028_1, in1028_2;
    wire c1028;
    assign in1028_1 = {pp78[69],pp79[69],pp80[69],pp81[69]};
    assign in1028_2 = {pp79[68],pp80[68],pp81[68],pp82[68]};
    CLA_4 KS_1028(s1028, c1028, in1028_1, in1028_2);
    wire[2:0] s1029, in1029_1, in1029_2;
    wire c1029;
    assign in1029_1 = {pp80[67],pp81[67],pp82[67]};
    assign in1029_2 = {pp81[66],pp82[66],pp83[66]};
    CLA_3 KS_1029(s1029, c1029, in1029_1, in1029_2);
    wire[1:0] s1030, in1030_1, in1030_2;
    wire c1030;
    assign in1030_1 = {pp82[65],pp83[65]};
    assign in1030_2 = {pp83[64],pp84[64]};
    CLA_2 KS_1030(s1030, c1030, in1030_1, in1030_2);
    wire[0:0] s1031, in1031_1, in1031_2;
    wire c1031;
    assign in1031_1 = {pp84[63]};
    assign in1031_2 = {pp85[62]};
    Half_Adder KS_1031(s1031, c1031, in1031_1, in1031_2);
    wire[3:0] s1032, in1032_1, in1032_2;
    wire c1032;
    assign in1032_1 = {pp86[61],pp85[63],pp84[65],pp83[67]};
    assign in1032_2 = {pp87[60],pp86[62],pp85[64],pp84[66]};
    CLA_4 KS_1032(s1032, c1032, in1032_1, in1032_2);
    wire[0:0] s1033, in1033_1, in1033_2;
    wire c1033;
    assign in1033_1 = {pp88[59]};
    assign in1033_2 = {pp89[58]};
    Half_Adder KS_1033(s1033, c1033, in1033_1, in1033_2);
    wire[1:0] s1034, in1034_1, in1034_2;
    wire c1034;
    assign in1034_1 = {pp90[57],pp87[61]};
    assign in1034_2 = {pp91[56],pp88[60]};
    CLA_2 KS_1034(s1034, c1034, in1034_1, in1034_2);
    wire[0:0] s1035, in1035_1, in1035_2;
    wire c1035;
    assign in1035_1 = {pp92[55]};
    assign in1035_2 = {pp93[54]};
    Half_Adder KS_1035(s1035, c1035, in1035_1, in1035_2);
    wire[2:0] s1036, in1036_1, in1036_2;
    wire c1036;
    assign in1036_1 = {pp94[53],pp89[59],pp86[63]};
    assign in1036_2 = {pp95[52],pp90[58],pp87[62]};
    CLA_3 KS_1036(s1036, c1036, in1036_1, in1036_2);
    wire[0:0] s1037, in1037_1, in1037_2;
    wire c1037;
    assign in1037_1 = {pp96[51]};
    assign in1037_2 = {pp97[50]};
    Half_Adder KS_1037(s1037, c1037, in1037_1, in1037_2);
    wire[1:0] s1038, in1038_1, in1038_2;
    wire c1038;
    assign in1038_1 = {pp98[49],pp91[57]};
    assign in1038_2 = {pp99[48],pp92[56]};
    CLA_2 KS_1038(s1038, c1038, in1038_1, in1038_2);
    wire[0:0] s1039, in1039_1, in1039_2;
    wire c1039;
    assign in1039_1 = {pp100[47]};
    assign in1039_2 = {pp101[46]};
    Half_Adder KS_1039(s1039, c1039, in1039_1, in1039_2);
    wire[3:0] s1040, in1040_1, in1040_2;
    wire c1040;
    assign in1040_1 = {pp102[45],pp93[55],pp88[61],pp85[65]};
    assign in1040_2 = {pp103[44],pp94[54],pp89[60],pp86[64]};
    CLA_4 KS_1040(s1040, c1040, in1040_1, in1040_2);
    wire[0:0] s1041, in1041_1, in1041_2;
    wire c1041;
    assign in1041_1 = {pp104[43]};
    assign in1041_2 = {pp105[42]};
    Half_Adder KS_1041(s1041, c1041, in1041_1, in1041_2);
    wire[1:0] s1042, in1042_1, in1042_2;
    wire c1042;
    assign in1042_1 = {pp106[41],pp95[53]};
    assign in1042_2 = {pp107[40],pp96[52]};
    CLA_2 KS_1042(s1042, c1042, in1042_1, in1042_2);
    wire[0:0] s1043, in1043_1, in1043_2;
    wire c1043;
    assign in1043_1 = {pp108[39]};
    assign in1043_2 = {pp109[38]};
    Half_Adder KS_1043(s1043, c1043, in1043_1, in1043_2);
    wire[2:0] s1044, in1044_1, in1044_2;
    wire c1044;
    assign in1044_1 = {pp110[37],pp97[51],pp90[59]};
    assign in1044_2 = {pp111[36],pp98[50],pp91[58]};
    CLA_3 KS_1044(s1044, c1044, in1044_1, in1044_2);
    wire[0:0] s1045, in1045_1, in1045_2;
    wire c1045;
    assign in1045_1 = {pp112[35]};
    assign in1045_2 = {pp113[34]};
    Half_Adder KS_1045(s1045, c1045, in1045_1, in1045_2);
    wire[1:0] s1046, in1046_1, in1046_2;
    wire c1046;
    assign in1046_1 = {pp114[33],pp99[49]};
    assign in1046_2 = {pp115[32],pp100[48]};
    CLA_2 KS_1046(s1046, c1046, in1046_1, in1046_2);
    wire[0:0] s1047, in1047_1, in1047_2;
    wire c1047;
    assign in1047_1 = {pp116[31]};
    assign in1047_2 = {pp117[30]};
    Half_Adder KS_1047(s1047, c1047, in1047_1, in1047_2);
    wire[3:0] s1048, in1048_1, in1048_2;
    wire c1048;
    assign in1048_1 = {pp118[29],pp101[47],pp92[57],pp87[63]};
    assign in1048_2 = {pp119[28],pp102[46],pp93[56],pp88[62]};
    CLA_4 KS_1048(s1048, c1048, in1048_1, in1048_2);
    wire[0:0] s1049, in1049_1, in1049_2;
    wire c1049;
    assign in1049_1 = {pp120[27]};
    assign in1049_2 = {pp121[26]};
    Half_Adder KS_1049(s1049, c1049, in1049_1, in1049_2);
    wire[1:0] s1050, in1050_1, in1050_2;
    wire c1050;
    assign in1050_1 = {pp122[25],pp103[45]};
    assign in1050_2 = {pp123[24],pp104[44]};
    CLA_2 KS_1050(s1050, c1050, in1050_1, in1050_2);
    wire[0:0] s1051, in1051_1, in1051_2;
    wire c1051;
    assign in1051_1 = {pp124[23]};
    assign in1051_2 = {pp125[22]};
    Half_Adder KS_1051(s1051, c1051, in1051_1, in1051_2);
    wire[2:0] s1052, in1052_1, in1052_2;
    wire c1052;
    assign in1052_1 = {pp126[21],pp105[43],pp94[55]};
    assign in1052_2 = {pp127[20],pp106[42],pp95[54]};
    CLA_3 KS_1052(s1052, c1052, in1052_1, in1052_2);
    wire[0:0] s1053, in1053_1, in1053_2;
    wire c1053;
    assign in1053_1 = {c920};
    assign in1053_2 = {c921};
    Half_Adder KS_1053(s1053, c1053, in1053_1, in1053_2);
    wire[1:0] s1054, in1054_1, in1054_2;
    wire c1054;
    assign in1054_1 = {c922,pp107[41]};
    assign in1054_2 = {c923,pp108[40]};
    CLA_2 KS_1054(s1054, c1054, in1054_1, in1054_2);
    wire[0:0] s1055, in1055_1, in1055_2;
    wire c1055;
    assign in1055_1 = {c924};
    assign in1055_2 = {c925};
    Half_Adder KS_1055(s1055, c1055, in1055_1, in1055_2);
    wire[3:0] s1056, in1056_1, in1056_2;
    wire c1056;
    assign in1056_1 = {c926,pp109[39],pp96[53],pp89[61]};
    assign in1056_2 = {c927,pp110[38],pp97[52],pp90[60]};
    CLA_4 KS_1056(s1056, c1056, in1056_1, in1056_2);
    wire[0:0] s1057, in1057_1, in1057_2;
    wire c1057;
    assign in1057_1 = {c928};
    assign in1057_2 = {c929};
    Half_Adder KS_1057(s1057, c1057, in1057_1, in1057_2);
    wire[1:0] s1058, in1058_1, in1058_2;
    wire c1058;
    assign in1058_1 = {c930,pp111[37]};
    assign in1058_2 = {c931,pp112[36]};
    CLA_2 KS_1058(s1058, c1058, in1058_1, in1058_2);
    wire[0:0] s1059, in1059_1, in1059_2;
    wire c1059;
    assign in1059_1 = {c932};
    assign in1059_2 = {c933};
    Half_Adder KS_1059(s1059, c1059, in1059_1, in1059_2);
    wire[2:0] s1060, in1060_1, in1060_2;
    wire c1060;
    assign in1060_1 = {c934,pp113[35],pp98[51]};
    assign in1060_2 = {c935,pp114[34],pp99[50]};
    CLA_3 KS_1060(s1060, c1060, in1060_1, in1060_2);
    wire[0:0] s1061, in1061_1, in1061_2;
    wire c1061;
    assign in1061_1 = {c936};
    assign in1061_2 = {c937};
    Half_Adder KS_1061(s1061, c1061, in1061_1, in1061_2);
    wire[1:0] s1062, in1062_1, in1062_2;
    wire c1062;
    assign in1062_1 = {c938,pp115[33]};
    assign in1062_2 = {c939,pp116[32]};
    CLA_2 KS_1062(s1062, c1062, in1062_1, in1062_2);
    wire[0:0] s1063, in1063_1, in1063_2;
    wire c1063;
    assign in1063_1 = {c940};
    assign in1063_2 = {c941};
    Half_Adder KS_1063(s1063, c1063, in1063_1, in1063_2);
    wire[3:0] s1064, in1064_1, in1064_2;
    wire c1064;
    assign in1064_1 = {c942,pp117[31],pp100[49],pp91[59]};
    assign in1064_2 = {c943,pp118[30],pp101[48],pp92[58]};
    CLA_4 KS_1064(s1064, c1064, in1064_1, in1064_2);
    wire[0:0] s1065, in1065_1, in1065_2;
    wire c1065;
    assign in1065_1 = {c944};
    assign in1065_2 = {c945};
    Half_Adder KS_1065(s1065, c1065, in1065_1, in1065_2);
    wire[1:0] s1066, in1066_1, in1066_2;
    wire c1066;
    assign in1066_1 = {c946,pp119[29]};
    assign in1066_2 = {c947,pp120[28]};
    CLA_2 KS_1066(s1066, c1066, in1066_1, in1066_2);
    wire[0:0] s1067, in1067_1, in1067_2;
    wire c1067;
    assign in1067_1 = {c948};
    assign in1067_2 = {c949};
    Half_Adder KS_1067(s1067, c1067, in1067_1, in1067_2);
    wire[2:0] s1068, in1068_1, in1068_2;
    wire c1068;
    assign in1068_1 = {c950,pp121[27],pp102[47]};
    assign in1068_2 = {c951,pp122[26],pp103[46]};
    CLA_3 KS_1068(s1068, c1068, in1068_1, in1068_2);
    wire[0:0] s1069, in1069_1, in1069_2;
    wire c1069;
    assign in1069_1 = {c953};
    assign in1069_2 = {c957};
    Full_Adder KS_1069(s1069, c1069, in1069_1, in1069_2, c952);
    wire[3:0] s1070, in1070_1, in1070_2;
    wire c1070;
    assign in1070_1 = {pp24[127],pp25[127],pp26[127],pp27[127]};
    assign in1070_2 = {pp25[126],pp26[126],pp27[126],pp28[126]};
    CLA_4 KS_1070(s1070, c1070, in1070_1, in1070_2);
    wire[3:0] s1071, in1071_1, in1071_2;
    wire c1071;
    assign in1071_1 = {pp26[125],pp27[125],pp28[125],pp29[125]};
    assign in1071_2 = {pp27[124],pp28[124],pp29[124],pp30[124]};
    CLA_4 KS_1071(s1071, c1071, in1071_1, in1071_2);
    wire[3:0] s1072, in1072_1, in1072_2;
    wire c1072;
    assign in1072_1 = {pp28[123],pp29[123],pp30[123],pp31[123]};
    assign in1072_2 = {pp29[122],pp30[122],pp31[122],pp32[122]};
    CLA_4 KS_1072(s1072, c1072, in1072_1, in1072_2);
    wire[3:0] s1073, in1073_1, in1073_2;
    wire c1073;
    assign in1073_1 = {pp30[121],pp31[121],pp32[121],pp33[121]};
    assign in1073_2 = {pp31[120],pp32[120],pp33[120],pp34[120]};
    CLA_4 KS_1073(s1073, c1073, in1073_1, in1073_2);
    wire[3:0] s1074, in1074_1, in1074_2;
    wire c1074;
    assign in1074_1 = {pp32[119],pp33[119],pp34[119],pp35[119]};
    assign in1074_2 = {pp33[118],pp34[118],pp35[118],pp36[118]};
    CLA_4 KS_1074(s1074, c1074, in1074_1, in1074_2);
    wire[3:0] s1075, in1075_1, in1075_2;
    wire c1075;
    assign in1075_1 = {pp34[117],pp35[117],pp36[117],pp37[117]};
    assign in1075_2 = {pp35[116],pp36[116],pp37[116],pp38[116]};
    CLA_4 KS_1075(s1075, c1075, in1075_1, in1075_2);
    wire[3:0] s1076, in1076_1, in1076_2;
    wire c1076;
    assign in1076_1 = {pp36[115],pp37[115],pp38[115],pp39[115]};
    assign in1076_2 = {pp37[114],pp38[114],pp39[114],pp40[114]};
    CLA_4 KS_1076(s1076, c1076, in1076_1, in1076_2);
    wire[3:0] s1077, in1077_1, in1077_2;
    wire c1077;
    assign in1077_1 = {pp38[113],pp39[113],pp40[113],pp41[113]};
    assign in1077_2 = {pp39[112],pp40[112],pp41[112],pp42[112]};
    CLA_4 KS_1077(s1077, c1077, in1077_1, in1077_2);
    wire[3:0] s1078, in1078_1, in1078_2;
    wire c1078;
    assign in1078_1 = {pp40[111],pp41[111],pp42[111],pp43[111]};
    assign in1078_2 = {pp41[110],pp42[110],pp43[110],pp44[110]};
    CLA_4 KS_1078(s1078, c1078, in1078_1, in1078_2);
    wire[3:0] s1079, in1079_1, in1079_2;
    wire c1079;
    assign in1079_1 = {pp42[109],pp43[109],pp44[109],pp45[109]};
    assign in1079_2 = {pp43[108],pp44[108],pp45[108],pp46[108]};
    CLA_4 KS_1079(s1079, c1079, in1079_1, in1079_2);
    wire[3:0] s1080, in1080_1, in1080_2;
    wire c1080;
    assign in1080_1 = {pp44[107],pp45[107],pp46[107],pp47[107]};
    assign in1080_2 = {pp45[106],pp46[106],pp47[106],pp48[106]};
    CLA_4 KS_1080(s1080, c1080, in1080_1, in1080_2);
    wire[3:0] s1081, in1081_1, in1081_2;
    wire c1081;
    assign in1081_1 = {pp46[105],pp47[105],pp48[105],pp49[105]};
    assign in1081_2 = {pp47[104],pp48[104],pp49[104],pp50[104]};
    CLA_4 KS_1081(s1081, c1081, in1081_1, in1081_2);
    wire[3:0] s1082, in1082_1, in1082_2;
    wire c1082;
    assign in1082_1 = {pp48[103],pp49[103],pp50[103],pp51[103]};
    assign in1082_2 = {pp49[102],pp50[102],pp51[102],pp52[102]};
    CLA_4 KS_1082(s1082, c1082, in1082_1, in1082_2);
    wire[3:0] s1083, in1083_1, in1083_2;
    wire c1083;
    assign in1083_1 = {pp50[101],pp51[101],pp52[101],pp53[101]};
    assign in1083_2 = {pp51[100],pp52[100],pp53[100],pp54[100]};
    CLA_4 KS_1083(s1083, c1083, in1083_1, in1083_2);
    wire[3:0] s1084, in1084_1, in1084_2;
    wire c1084;
    assign in1084_1 = {pp52[99],pp53[99],pp54[99],pp55[99]};
    assign in1084_2 = {pp53[98],pp54[98],pp55[98],pp56[98]};
    CLA_4 KS_1084(s1084, c1084, in1084_1, in1084_2);
    wire[3:0] s1085, in1085_1, in1085_2;
    wire c1085;
    assign in1085_1 = {pp54[97],pp55[97],pp56[97],pp57[97]};
    assign in1085_2 = {pp55[96],pp56[96],pp57[96],pp58[96]};
    CLA_4 KS_1085(s1085, c1085, in1085_1, in1085_2);
    wire[3:0] s1086, in1086_1, in1086_2;
    wire c1086;
    assign in1086_1 = {pp56[95],pp57[95],pp58[95],pp59[95]};
    assign in1086_2 = {pp57[94],pp58[94],pp59[94],pp60[94]};
    CLA_4 KS_1086(s1086, c1086, in1086_1, in1086_2);
    wire[3:0] s1087, in1087_1, in1087_2;
    wire c1087;
    assign in1087_1 = {pp58[93],pp59[93],pp60[93],pp61[93]};
    assign in1087_2 = {pp59[92],pp60[92],pp61[92],pp62[92]};
    CLA_4 KS_1087(s1087, c1087, in1087_1, in1087_2);
    wire[3:0] s1088, in1088_1, in1088_2;
    wire c1088;
    assign in1088_1 = {pp60[91],pp61[91],pp62[91],pp63[91]};
    assign in1088_2 = {pp61[90],pp62[90],pp63[90],pp64[90]};
    CLA_4 KS_1088(s1088, c1088, in1088_1, in1088_2);
    wire[3:0] s1089, in1089_1, in1089_2;
    wire c1089;
    assign in1089_1 = {pp62[89],pp63[89],pp64[89],pp65[89]};
    assign in1089_2 = {pp63[88],pp64[88],pp65[88],pp66[88]};
    CLA_4 KS_1089(s1089, c1089, in1089_1, in1089_2);
    wire[3:0] s1090, in1090_1, in1090_2;
    wire c1090;
    assign in1090_1 = {pp64[87],pp65[87],pp66[87],pp67[87]};
    assign in1090_2 = {pp65[86],pp66[86],pp67[86],pp68[86]};
    CLA_4 KS_1090(s1090, c1090, in1090_1, in1090_2);
    wire[3:0] s1091, in1091_1, in1091_2;
    wire c1091;
    assign in1091_1 = {pp66[85],pp67[85],pp68[85],pp69[85]};
    assign in1091_2 = {pp67[84],pp68[84],pp69[84],pp70[84]};
    CLA_4 KS_1091(s1091, c1091, in1091_1, in1091_2);
    wire[3:0] s1092, in1092_1, in1092_2;
    wire c1092;
    assign in1092_1 = {pp68[83],pp69[83],pp70[83],pp71[83]};
    assign in1092_2 = {pp69[82],pp70[82],pp71[82],pp72[82]};
    CLA_4 KS_1092(s1092, c1092, in1092_1, in1092_2);
    wire[3:0] s1093, in1093_1, in1093_2;
    wire c1093;
    assign in1093_1 = {pp70[81],pp71[81],pp72[81],pp73[81]};
    assign in1093_2 = {pp71[80],pp72[80],pp73[80],pp74[80]};
    CLA_4 KS_1093(s1093, c1093, in1093_1, in1093_2);
    wire[3:0] s1094, in1094_1, in1094_2;
    wire c1094;
    assign in1094_1 = {pp72[79],pp73[79],pp74[79],pp75[79]};
    assign in1094_2 = {pp73[78],pp74[78],pp75[78],pp76[78]};
    CLA_4 KS_1094(s1094, c1094, in1094_1, in1094_2);
    wire[3:0] s1095, in1095_1, in1095_2;
    wire c1095;
    assign in1095_1 = {pp74[77],pp75[77],pp76[77],pp77[77]};
    assign in1095_2 = {pp75[76],pp76[76],pp77[76],pp78[76]};
    CLA_4 KS_1095(s1095, c1095, in1095_1, in1095_2);
    wire[2:0] s1096, in1096_1, in1096_2;
    wire c1096;
    assign in1096_1 = {pp76[75],pp77[75],pp78[75]};
    assign in1096_2 = {pp77[74],pp78[74],pp79[74]};
    CLA_3 KS_1096(s1096, c1096, in1096_1, in1096_2);
    wire[1:0] s1097, in1097_1, in1097_2;
    wire c1097;
    assign in1097_1 = {pp78[73],pp79[73]};
    assign in1097_2 = {pp79[72],pp80[72]};
    CLA_2 KS_1097(s1097, c1097, in1097_1, in1097_2);
    wire[0:0] s1098, in1098_1, in1098_2;
    wire c1098;
    assign in1098_1 = {pp80[71]};
    assign in1098_2 = {pp81[70]};
    Half_Adder KS_1098(s1098, c1098, in1098_1, in1098_2);
    wire[3:0] s1099, in1099_1, in1099_2;
    wire c1099;
    assign in1099_1 = {pp82[69],pp81[71],pp80[73],pp79[75]};
    assign in1099_2 = {pp83[68],pp82[70],pp81[72],pp80[74]};
    CLA_4 KS_1099(s1099, c1099, in1099_1, in1099_2);
    wire[0:0] s1100, in1100_1, in1100_2;
    wire c1100;
    assign in1100_1 = {pp84[67]};
    assign in1100_2 = {pp85[66]};
    Half_Adder KS_1100(s1100, c1100, in1100_1, in1100_2);
    wire[1:0] s1101, in1101_1, in1101_2;
    wire c1101;
    assign in1101_1 = {pp86[65],pp83[69]};
    assign in1101_2 = {pp87[64],pp84[68]};
    CLA_2 KS_1101(s1101, c1101, in1101_1, in1101_2);
    wire[0:0] s1102, in1102_1, in1102_2;
    wire c1102;
    assign in1102_1 = {pp88[63]};
    assign in1102_2 = {pp89[62]};
    Half_Adder KS_1102(s1102, c1102, in1102_1, in1102_2);
    wire[2:0] s1103, in1103_1, in1103_2;
    wire c1103;
    assign in1103_1 = {pp90[61],pp85[67],pp82[71]};
    assign in1103_2 = {pp91[60],pp86[66],pp83[70]};
    CLA_3 KS_1103(s1103, c1103, in1103_1, in1103_2);
    wire[0:0] s1104, in1104_1, in1104_2;
    wire c1104;
    assign in1104_1 = {pp92[59]};
    assign in1104_2 = {pp93[58]};
    Half_Adder KS_1104(s1104, c1104, in1104_1, in1104_2);
    wire[1:0] s1105, in1105_1, in1105_2;
    wire c1105;
    assign in1105_1 = {pp94[57],pp87[65]};
    assign in1105_2 = {pp95[56],pp88[64]};
    CLA_2 KS_1105(s1105, c1105, in1105_1, in1105_2);
    wire[0:0] s1106, in1106_1, in1106_2;
    wire c1106;
    assign in1106_1 = {pp96[55]};
    assign in1106_2 = {pp97[54]};
    Half_Adder KS_1106(s1106, c1106, in1106_1, in1106_2);
    wire[3:0] s1107, in1107_1, in1107_2;
    wire c1107;
    assign in1107_1 = {pp98[53],pp89[63],pp84[69],pp81[73]};
    assign in1107_2 = {pp99[52],pp90[62],pp85[68],pp82[72]};
    CLA_4 KS_1107(s1107, c1107, in1107_1, in1107_2);
    wire[0:0] s1108, in1108_1, in1108_2;
    wire c1108;
    assign in1108_1 = {pp100[51]};
    assign in1108_2 = {pp101[50]};
    Half_Adder KS_1108(s1108, c1108, in1108_1, in1108_2);
    wire[1:0] s1109, in1109_1, in1109_2;
    wire c1109;
    assign in1109_1 = {pp102[49],pp91[61]};
    assign in1109_2 = {pp103[48],pp92[60]};
    CLA_2 KS_1109(s1109, c1109, in1109_1, in1109_2);
    wire[0:0] s1110, in1110_1, in1110_2;
    wire c1110;
    assign in1110_1 = {pp104[47]};
    assign in1110_2 = {pp105[46]};
    Half_Adder KS_1110(s1110, c1110, in1110_1, in1110_2);
    wire[2:0] s1111, in1111_1, in1111_2;
    wire c1111;
    assign in1111_1 = {pp106[45],pp93[59],pp86[67]};
    assign in1111_2 = {pp107[44],pp94[58],pp87[66]};
    CLA_3 KS_1111(s1111, c1111, in1111_1, in1111_2);
    wire[0:0] s1112, in1112_1, in1112_2;
    wire c1112;
    assign in1112_1 = {pp108[43]};
    assign in1112_2 = {pp109[42]};
    Half_Adder KS_1112(s1112, c1112, in1112_1, in1112_2);
    wire[1:0] s1113, in1113_1, in1113_2;
    wire c1113;
    assign in1113_1 = {pp110[41],pp95[57]};
    assign in1113_2 = {pp111[40],pp96[56]};
    CLA_2 KS_1113(s1113, c1113, in1113_1, in1113_2);
    wire[0:0] s1114, in1114_1, in1114_2;
    wire c1114;
    assign in1114_1 = {pp112[39]};
    assign in1114_2 = {pp113[38]};
    Half_Adder KS_1114(s1114, c1114, in1114_1, in1114_2);
    wire[3:0] s1115, in1115_1, in1115_2;
    wire c1115;
    assign in1115_1 = {pp114[37],pp97[55],pp88[65],pp83[71]};
    assign in1115_2 = {pp115[36],pp98[54],pp89[64],pp84[70]};
    CLA_4 KS_1115(s1115, c1115, in1115_1, in1115_2);
    wire[0:0] s1116, in1116_1, in1116_2;
    wire c1116;
    assign in1116_1 = {pp116[35]};
    assign in1116_2 = {pp117[34]};
    Half_Adder KS_1116(s1116, c1116, in1116_1, in1116_2);
    wire[1:0] s1117, in1117_1, in1117_2;
    wire c1117;
    assign in1117_1 = {pp118[33],pp99[53]};
    assign in1117_2 = {pp119[32],pp100[52]};
    CLA_2 KS_1117(s1117, c1117, in1117_1, in1117_2);
    wire[0:0] s1118, in1118_1, in1118_2;
    wire c1118;
    assign in1118_1 = {pp120[31]};
    assign in1118_2 = {pp121[30]};
    Half_Adder KS_1118(s1118, c1118, in1118_1, in1118_2);
    wire[2:0] s1119, in1119_1, in1119_2;
    wire c1119;
    assign in1119_1 = {pp122[29],pp101[51],pp90[63]};
    assign in1119_2 = {pp123[28],pp102[50],pp91[62]};
    CLA_3 KS_1119(s1119, c1119, in1119_1, in1119_2);
    wire[0:0] s1120, in1120_1, in1120_2;
    wire c1120;
    assign in1120_1 = {pp124[27]};
    assign in1120_2 = {pp125[26]};
    Half_Adder KS_1120(s1120, c1120, in1120_1, in1120_2);
    wire[1:0] s1121, in1121_1, in1121_2;
    wire c1121;
    assign in1121_1 = {pp126[25],pp103[49]};
    assign in1121_2 = {pp127[24],pp104[48]};
    CLA_2 KS_1121(s1121, c1121, in1121_1, in1121_2);
    wire[0:0] s1122, in1122_1, in1122_2;
    wire c1122;
    assign in1122_1 = {c999};
    assign in1122_2 = {c1000};
    Half_Adder KS_1122(s1122, c1122, in1122_1, in1122_2);
    wire[3:0] s1123, in1123_1, in1123_2;
    wire c1123;
    assign in1123_1 = {c1001,pp105[47],pp92[61],pp85[69]};
    assign in1123_2 = {c1002,pp106[46],pp93[60],pp86[68]};
    CLA_4 KS_1123(s1123, c1123, in1123_1, in1123_2);
    wire[0:0] s1124, in1124_1, in1124_2;
    wire c1124;
    assign in1124_1 = {c1003};
    assign in1124_2 = {c1004};
    Half_Adder KS_1124(s1124, c1124, in1124_1, in1124_2);
    wire[1:0] s1125, in1125_1, in1125_2;
    wire c1125;
    assign in1125_1 = {c1005,pp107[45]};
    assign in1125_2 = {c1006,pp108[44]};
    CLA_2 KS_1125(s1125, c1125, in1125_1, in1125_2);
    wire[0:0] s1126, in1126_1, in1126_2;
    wire c1126;
    assign in1126_1 = {c1007};
    assign in1126_2 = {c1008};
    Half_Adder KS_1126(s1126, c1126, in1126_1, in1126_2);
    wire[2:0] s1127, in1127_1, in1127_2;
    wire c1127;
    assign in1127_1 = {c1009,pp109[43],pp94[59]};
    assign in1127_2 = {c1010,pp110[42],pp95[58]};
    CLA_3 KS_1127(s1127, c1127, in1127_1, in1127_2);
    wire[0:0] s1128, in1128_1, in1128_2;
    wire c1128;
    assign in1128_1 = {c1011};
    assign in1128_2 = {c1012};
    Half_Adder KS_1128(s1128, c1128, in1128_1, in1128_2);
    wire[1:0] s1129, in1129_1, in1129_2;
    wire c1129;
    assign in1129_1 = {c1013,pp111[41]};
    assign in1129_2 = {c1014,pp112[40]};
    CLA_2 KS_1129(s1129, c1129, in1129_1, in1129_2);
    wire[0:0] s1130, in1130_1, in1130_2;
    wire c1130;
    assign in1130_1 = {c1015};
    assign in1130_2 = {c1016};
    Half_Adder KS_1130(s1130, c1130, in1130_1, in1130_2);
    wire[3:0] s1131, in1131_1, in1131_2;
    wire c1131;
    assign in1131_1 = {c1018,pp113[39],pp96[57],pp87[67]};
    assign in1131_2 = {c1019,pp114[38],pp97[56],pp88[66]};
    CLA_4_c KS_1131(s1131, c1131, in1131_1, in1131_2, c1017);
    wire[3:0] s1132, in1132_1, in1132_2;
    wire c1132;
    assign in1132_1 = {pp28[127],pp29[127],pp30[127],pp31[127]};
    assign in1132_2 = {pp29[126],pp30[126],pp31[126],pp32[126]};
    CLA_4 KS_1132(s1132, c1132, in1132_1, in1132_2);
    wire[3:0] s1133, in1133_1, in1133_2;
    wire c1133;
    assign in1133_1 = {pp30[125],pp31[125],pp32[125],pp33[125]};
    assign in1133_2 = {pp31[124],pp32[124],pp33[124],pp34[124]};
    CLA_4 KS_1133(s1133, c1133, in1133_1, in1133_2);
    wire[3:0] s1134, in1134_1, in1134_2;
    wire c1134;
    assign in1134_1 = {pp32[123],pp33[123],pp34[123],pp35[123]};
    assign in1134_2 = {pp33[122],pp34[122],pp35[122],pp36[122]};
    CLA_4 KS_1134(s1134, c1134, in1134_1, in1134_2);
    wire[3:0] s1135, in1135_1, in1135_2;
    wire c1135;
    assign in1135_1 = {pp34[121],pp35[121],pp36[121],pp37[121]};
    assign in1135_2 = {pp35[120],pp36[120],pp37[120],pp38[120]};
    CLA_4 KS_1135(s1135, c1135, in1135_1, in1135_2);
    wire[3:0] s1136, in1136_1, in1136_2;
    wire c1136;
    assign in1136_1 = {pp36[119],pp37[119],pp38[119],pp39[119]};
    assign in1136_2 = {pp37[118],pp38[118],pp39[118],pp40[118]};
    CLA_4 KS_1136(s1136, c1136, in1136_1, in1136_2);
    wire[3:0] s1137, in1137_1, in1137_2;
    wire c1137;
    assign in1137_1 = {pp38[117],pp39[117],pp40[117],pp41[117]};
    assign in1137_2 = {pp39[116],pp40[116],pp41[116],pp42[116]};
    CLA_4 KS_1137(s1137, c1137, in1137_1, in1137_2);
    wire[3:0] s1138, in1138_1, in1138_2;
    wire c1138;
    assign in1138_1 = {pp40[115],pp41[115],pp42[115],pp43[115]};
    assign in1138_2 = {pp41[114],pp42[114],pp43[114],pp44[114]};
    CLA_4 KS_1138(s1138, c1138, in1138_1, in1138_2);
    wire[3:0] s1139, in1139_1, in1139_2;
    wire c1139;
    assign in1139_1 = {pp42[113],pp43[113],pp44[113],pp45[113]};
    assign in1139_2 = {pp43[112],pp44[112],pp45[112],pp46[112]};
    CLA_4 KS_1139(s1139, c1139, in1139_1, in1139_2);
    wire[3:0] s1140, in1140_1, in1140_2;
    wire c1140;
    assign in1140_1 = {pp44[111],pp45[111],pp46[111],pp47[111]};
    assign in1140_2 = {pp45[110],pp46[110],pp47[110],pp48[110]};
    CLA_4 KS_1140(s1140, c1140, in1140_1, in1140_2);
    wire[3:0] s1141, in1141_1, in1141_2;
    wire c1141;
    assign in1141_1 = {pp46[109],pp47[109],pp48[109],pp49[109]};
    assign in1141_2 = {pp47[108],pp48[108],pp49[108],pp50[108]};
    CLA_4 KS_1141(s1141, c1141, in1141_1, in1141_2);
    wire[3:0] s1142, in1142_1, in1142_2;
    wire c1142;
    assign in1142_1 = {pp48[107],pp49[107],pp50[107],pp51[107]};
    assign in1142_2 = {pp49[106],pp50[106],pp51[106],pp52[106]};
    CLA_4 KS_1142(s1142, c1142, in1142_1, in1142_2);
    wire[3:0] s1143, in1143_1, in1143_2;
    wire c1143;
    assign in1143_1 = {pp50[105],pp51[105],pp52[105],pp53[105]};
    assign in1143_2 = {pp51[104],pp52[104],pp53[104],pp54[104]};
    CLA_4 KS_1143(s1143, c1143, in1143_1, in1143_2);
    wire[3:0] s1144, in1144_1, in1144_2;
    wire c1144;
    assign in1144_1 = {pp52[103],pp53[103],pp54[103],pp55[103]};
    assign in1144_2 = {pp53[102],pp54[102],pp55[102],pp56[102]};
    CLA_4 KS_1144(s1144, c1144, in1144_1, in1144_2);
    wire[3:0] s1145, in1145_1, in1145_2;
    wire c1145;
    assign in1145_1 = {pp54[101],pp55[101],pp56[101],pp57[101]};
    assign in1145_2 = {pp55[100],pp56[100],pp57[100],pp58[100]};
    CLA_4 KS_1145(s1145, c1145, in1145_1, in1145_2);
    wire[3:0] s1146, in1146_1, in1146_2;
    wire c1146;
    assign in1146_1 = {pp56[99],pp57[99],pp58[99],pp59[99]};
    assign in1146_2 = {pp57[98],pp58[98],pp59[98],pp60[98]};
    CLA_4 KS_1146(s1146, c1146, in1146_1, in1146_2);
    wire[3:0] s1147, in1147_1, in1147_2;
    wire c1147;
    assign in1147_1 = {pp58[97],pp59[97],pp60[97],pp61[97]};
    assign in1147_2 = {pp59[96],pp60[96],pp61[96],pp62[96]};
    CLA_4 KS_1147(s1147, c1147, in1147_1, in1147_2);
    wire[3:0] s1148, in1148_1, in1148_2;
    wire c1148;
    assign in1148_1 = {pp60[95],pp61[95],pp62[95],pp63[95]};
    assign in1148_2 = {pp61[94],pp62[94],pp63[94],pp64[94]};
    CLA_4 KS_1148(s1148, c1148, in1148_1, in1148_2);
    wire[3:0] s1149, in1149_1, in1149_2;
    wire c1149;
    assign in1149_1 = {pp62[93],pp63[93],pp64[93],pp65[93]};
    assign in1149_2 = {pp63[92],pp64[92],pp65[92],pp66[92]};
    CLA_4 KS_1149(s1149, c1149, in1149_1, in1149_2);
    wire[3:0] s1150, in1150_1, in1150_2;
    wire c1150;
    assign in1150_1 = {pp64[91],pp65[91],pp66[91],pp67[91]};
    assign in1150_2 = {pp65[90],pp66[90],pp67[90],pp68[90]};
    CLA_4 KS_1150(s1150, c1150, in1150_1, in1150_2);
    wire[3:0] s1151, in1151_1, in1151_2;
    wire c1151;
    assign in1151_1 = {pp66[89],pp67[89],pp68[89],pp69[89]};
    assign in1151_2 = {pp67[88],pp68[88],pp69[88],pp70[88]};
    CLA_4 KS_1151(s1151, c1151, in1151_1, in1151_2);
    wire[3:0] s1152, in1152_1, in1152_2;
    wire c1152;
    assign in1152_1 = {pp68[87],pp69[87],pp70[87],pp71[87]};
    assign in1152_2 = {pp69[86],pp70[86],pp71[86],pp72[86]};
    CLA_4 KS_1152(s1152, c1152, in1152_1, in1152_2);
    wire[3:0] s1153, in1153_1, in1153_2;
    wire c1153;
    assign in1153_1 = {pp70[85],pp71[85],pp72[85],pp73[85]};
    assign in1153_2 = {pp71[84],pp72[84],pp73[84],pp74[84]};
    CLA_4 KS_1153(s1153, c1153, in1153_1, in1153_2);
    wire[2:0] s1154, in1154_1, in1154_2;
    wire c1154;
    assign in1154_1 = {pp72[83],pp73[83],pp74[83]};
    assign in1154_2 = {pp73[82],pp74[82],pp75[82]};
    CLA_3 KS_1154(s1154, c1154, in1154_1, in1154_2);
    wire[1:0] s1155, in1155_1, in1155_2;
    wire c1155;
    assign in1155_1 = {pp74[81],pp75[81]};
    assign in1155_2 = {pp75[80],pp76[80]};
    CLA_2 KS_1155(s1155, c1155, in1155_1, in1155_2);
    wire[0:0] s1156, in1156_1, in1156_2;
    wire c1156;
    assign in1156_1 = {pp76[79]};
    assign in1156_2 = {pp77[78]};
    Half_Adder KS_1156(s1156, c1156, in1156_1, in1156_2);
    wire[3:0] s1157, in1157_1, in1157_2;
    wire c1157;
    assign in1157_1 = {pp78[77],pp77[79],pp76[81],pp75[83]};
    assign in1157_2 = {pp79[76],pp78[78],pp77[80],pp76[82]};
    CLA_4 KS_1157(s1157, c1157, in1157_1, in1157_2);
    wire[0:0] s1158, in1158_1, in1158_2;
    wire c1158;
    assign in1158_1 = {pp80[75]};
    assign in1158_2 = {pp81[74]};
    Half_Adder KS_1158(s1158, c1158, in1158_1, in1158_2);
    wire[1:0] s1159, in1159_1, in1159_2;
    wire c1159;
    assign in1159_1 = {pp82[73],pp79[77]};
    assign in1159_2 = {pp83[72],pp80[76]};
    CLA_2 KS_1159(s1159, c1159, in1159_1, in1159_2);
    wire[0:0] s1160, in1160_1, in1160_2;
    wire c1160;
    assign in1160_1 = {pp84[71]};
    assign in1160_2 = {pp85[70]};
    Half_Adder KS_1160(s1160, c1160, in1160_1, in1160_2);
    wire[2:0] s1161, in1161_1, in1161_2;
    wire c1161;
    assign in1161_1 = {pp86[69],pp81[75],pp78[79]};
    assign in1161_2 = {pp87[68],pp82[74],pp79[78]};
    CLA_3 KS_1161(s1161, c1161, in1161_1, in1161_2);
    wire[0:0] s1162, in1162_1, in1162_2;
    wire c1162;
    assign in1162_1 = {pp88[67]};
    assign in1162_2 = {pp89[66]};
    Half_Adder KS_1162(s1162, c1162, in1162_1, in1162_2);
    wire[1:0] s1163, in1163_1, in1163_2;
    wire c1163;
    assign in1163_1 = {pp90[65],pp83[73]};
    assign in1163_2 = {pp91[64],pp84[72]};
    CLA_2 KS_1163(s1163, c1163, in1163_1, in1163_2);
    wire[0:0] s1164, in1164_1, in1164_2;
    wire c1164;
    assign in1164_1 = {pp92[63]};
    assign in1164_2 = {pp93[62]};
    Half_Adder KS_1164(s1164, c1164, in1164_1, in1164_2);
    wire[3:0] s1165, in1165_1, in1165_2;
    wire c1165;
    assign in1165_1 = {pp94[61],pp85[71],pp80[77],pp77[81]};
    assign in1165_2 = {pp95[60],pp86[70],pp81[76],pp78[80]};
    CLA_4 KS_1165(s1165, c1165, in1165_1, in1165_2);
    wire[0:0] s1166, in1166_1, in1166_2;
    wire c1166;
    assign in1166_1 = {pp96[59]};
    assign in1166_2 = {pp97[58]};
    Half_Adder KS_1166(s1166, c1166, in1166_1, in1166_2);
    wire[1:0] s1167, in1167_1, in1167_2;
    wire c1167;
    assign in1167_1 = {pp98[57],pp87[69]};
    assign in1167_2 = {pp99[56],pp88[68]};
    CLA_2 KS_1167(s1167, c1167, in1167_1, in1167_2);
    wire[0:0] s1168, in1168_1, in1168_2;
    wire c1168;
    assign in1168_1 = {pp100[55]};
    assign in1168_2 = {pp101[54]};
    Half_Adder KS_1168(s1168, c1168, in1168_1, in1168_2);
    wire[2:0] s1169, in1169_1, in1169_2;
    wire c1169;
    assign in1169_1 = {pp102[53],pp89[67],pp82[75]};
    assign in1169_2 = {pp103[52],pp90[66],pp83[74]};
    CLA_3 KS_1169(s1169, c1169, in1169_1, in1169_2);
    wire[0:0] s1170, in1170_1, in1170_2;
    wire c1170;
    assign in1170_1 = {pp104[51]};
    assign in1170_2 = {pp105[50]};
    Half_Adder KS_1170(s1170, c1170, in1170_1, in1170_2);
    wire[1:0] s1171, in1171_1, in1171_2;
    wire c1171;
    assign in1171_1 = {pp106[49],pp91[65]};
    assign in1171_2 = {pp107[48],pp92[64]};
    CLA_2 KS_1171(s1171, c1171, in1171_1, in1171_2);
    wire[0:0] s1172, in1172_1, in1172_2;
    wire c1172;
    assign in1172_1 = {pp108[47]};
    assign in1172_2 = {pp109[46]};
    Half_Adder KS_1172(s1172, c1172, in1172_1, in1172_2);
    wire[3:0] s1173, in1173_1, in1173_2;
    wire c1173;
    assign in1173_1 = {pp110[45],pp93[63],pp84[73],pp79[79]};
    assign in1173_2 = {pp111[44],pp94[62],pp85[72],pp80[78]};
    CLA_4 KS_1173(s1173, c1173, in1173_1, in1173_2);
    wire[0:0] s1174, in1174_1, in1174_2;
    wire c1174;
    assign in1174_1 = {pp112[43]};
    assign in1174_2 = {pp113[42]};
    Half_Adder KS_1174(s1174, c1174, in1174_1, in1174_2);
    wire[1:0] s1175, in1175_1, in1175_2;
    wire c1175;
    assign in1175_1 = {pp114[41],pp95[61]};
    assign in1175_2 = {pp115[40],pp96[60]};
    CLA_2 KS_1175(s1175, c1175, in1175_1, in1175_2);
    wire[0:0] s1176, in1176_1, in1176_2;
    wire c1176;
    assign in1176_1 = {pp116[39]};
    assign in1176_2 = {pp117[38]};
    Half_Adder KS_1176(s1176, c1176, in1176_1, in1176_2);
    wire[2:0] s1177, in1177_1, in1177_2;
    wire c1177;
    assign in1177_1 = {pp118[37],pp97[59],pp86[71]};
    assign in1177_2 = {pp119[36],pp98[58],pp87[70]};
    CLA_3 KS_1177(s1177, c1177, in1177_1, in1177_2);
    wire[0:0] s1178, in1178_1, in1178_2;
    wire c1178;
    assign in1178_1 = {pp120[35]};
    assign in1178_2 = {pp121[34]};
    Half_Adder KS_1178(s1178, c1178, in1178_1, in1178_2);
    wire[1:0] s1179, in1179_1, in1179_2;
    wire c1179;
    assign in1179_1 = {pp122[33],pp99[57]};
    assign in1179_2 = {pp123[32],pp100[56]};
    CLA_2 KS_1179(s1179, c1179, in1179_1, in1179_2);
    wire[0:0] s1180, in1180_1, in1180_2;
    wire c1180;
    assign in1180_1 = {pp124[31]};
    assign in1180_2 = {pp125[30]};
    Half_Adder KS_1180(s1180, c1180, in1180_1, in1180_2);
    wire[3:0] s1181, in1181_1, in1181_2;
    wire c1181;
    assign in1181_1 = {pp126[29],pp101[55],pp88[69],pp81[77]};
    assign in1181_2 = {pp127[28],pp102[54],pp89[68],pp82[76]};
    CLA_4 KS_1181(s1181, c1181, in1181_1, in1181_2);
    wire[0:0] s1182, in1182_1, in1182_2;
    wire c1182;
    assign in1182_1 = {c1070};
    assign in1182_2 = {c1071};
    Half_Adder KS_1182(s1182, c1182, in1182_1, in1182_2);
    wire[1:0] s1183, in1183_1, in1183_2;
    wire c1183;
    assign in1183_1 = {c1072,pp103[53]};
    assign in1183_2 = {c1073,pp104[52]};
    CLA_2 KS_1183(s1183, c1183, in1183_1, in1183_2);
    wire[0:0] s1184, in1184_1, in1184_2;
    wire c1184;
    assign in1184_1 = {c1074};
    assign in1184_2 = {c1075};
    Half_Adder KS_1184(s1184, c1184, in1184_1, in1184_2);
    wire[2:0] s1185, in1185_1, in1185_2;
    wire c1185;
    assign in1185_1 = {c1077,pp105[51],pp90[67]};
    assign in1185_2 = {c1078,pp106[50],pp91[66]};
    CLA_3_c KS_1185(s1185, c1185, in1185_1, in1185_2, c1076);
    wire[3:0] s1186, in1186_1, in1186_2;
    wire c1186;
    assign in1186_1 = {pp32[127],pp33[127],pp34[127],pp35[127]};
    assign in1186_2 = {pp33[126],pp34[126],pp35[126],pp36[126]};
    CLA_4 KS_1186(s1186, c1186, in1186_1, in1186_2);
    wire[3:0] s1187, in1187_1, in1187_2;
    wire c1187;
    assign in1187_1 = {pp34[125],pp35[125],pp36[125],pp37[125]};
    assign in1187_2 = {pp35[124],pp36[124],pp37[124],pp38[124]};
    CLA_4 KS_1187(s1187, c1187, in1187_1, in1187_2);
    wire[3:0] s1188, in1188_1, in1188_2;
    wire c1188;
    assign in1188_1 = {pp36[123],pp37[123],pp38[123],pp39[123]};
    assign in1188_2 = {pp37[122],pp38[122],pp39[122],pp40[122]};
    CLA_4 KS_1188(s1188, c1188, in1188_1, in1188_2);
    wire[3:0] s1189, in1189_1, in1189_2;
    wire c1189;
    assign in1189_1 = {pp38[121],pp39[121],pp40[121],pp41[121]};
    assign in1189_2 = {pp39[120],pp40[120],pp41[120],pp42[120]};
    CLA_4 KS_1189(s1189, c1189, in1189_1, in1189_2);
    wire[3:0] s1190, in1190_1, in1190_2;
    wire c1190;
    assign in1190_1 = {pp40[119],pp41[119],pp42[119],pp43[119]};
    assign in1190_2 = {pp41[118],pp42[118],pp43[118],pp44[118]};
    CLA_4 KS_1190(s1190, c1190, in1190_1, in1190_2);
    wire[3:0] s1191, in1191_1, in1191_2;
    wire c1191;
    assign in1191_1 = {pp42[117],pp43[117],pp44[117],pp45[117]};
    assign in1191_2 = {pp43[116],pp44[116],pp45[116],pp46[116]};
    CLA_4 KS_1191(s1191, c1191, in1191_1, in1191_2);
    wire[3:0] s1192, in1192_1, in1192_2;
    wire c1192;
    assign in1192_1 = {pp44[115],pp45[115],pp46[115],pp47[115]};
    assign in1192_2 = {pp45[114],pp46[114],pp47[114],pp48[114]};
    CLA_4 KS_1192(s1192, c1192, in1192_1, in1192_2);
    wire[3:0] s1193, in1193_1, in1193_2;
    wire c1193;
    assign in1193_1 = {pp46[113],pp47[113],pp48[113],pp49[113]};
    assign in1193_2 = {pp47[112],pp48[112],pp49[112],pp50[112]};
    CLA_4 KS_1193(s1193, c1193, in1193_1, in1193_2);
    wire[3:0] s1194, in1194_1, in1194_2;
    wire c1194;
    assign in1194_1 = {pp48[111],pp49[111],pp50[111],pp51[111]};
    assign in1194_2 = {pp49[110],pp50[110],pp51[110],pp52[110]};
    CLA_4 KS_1194(s1194, c1194, in1194_1, in1194_2);
    wire[3:0] s1195, in1195_1, in1195_2;
    wire c1195;
    assign in1195_1 = {pp50[109],pp51[109],pp52[109],pp53[109]};
    assign in1195_2 = {pp51[108],pp52[108],pp53[108],pp54[108]};
    CLA_4 KS_1195(s1195, c1195, in1195_1, in1195_2);
    wire[3:0] s1196, in1196_1, in1196_2;
    wire c1196;
    assign in1196_1 = {pp52[107],pp53[107],pp54[107],pp55[107]};
    assign in1196_2 = {pp53[106],pp54[106],pp55[106],pp56[106]};
    CLA_4 KS_1196(s1196, c1196, in1196_1, in1196_2);
    wire[3:0] s1197, in1197_1, in1197_2;
    wire c1197;
    assign in1197_1 = {pp54[105],pp55[105],pp56[105],pp57[105]};
    assign in1197_2 = {pp55[104],pp56[104],pp57[104],pp58[104]};
    CLA_4 KS_1197(s1197, c1197, in1197_1, in1197_2);
    wire[3:0] s1198, in1198_1, in1198_2;
    wire c1198;
    assign in1198_1 = {pp56[103],pp57[103],pp58[103],pp59[103]};
    assign in1198_2 = {pp57[102],pp58[102],pp59[102],pp60[102]};
    CLA_4 KS_1198(s1198, c1198, in1198_1, in1198_2);
    wire[3:0] s1199, in1199_1, in1199_2;
    wire c1199;
    assign in1199_1 = {pp58[101],pp59[101],pp60[101],pp61[101]};
    assign in1199_2 = {pp59[100],pp60[100],pp61[100],pp62[100]};
    CLA_4 KS_1199(s1199, c1199, in1199_1, in1199_2);
    wire[3:0] s1200, in1200_1, in1200_2;
    wire c1200;
    assign in1200_1 = {pp60[99],pp61[99],pp62[99],pp63[99]};
    assign in1200_2 = {pp61[98],pp62[98],pp63[98],pp64[98]};
    CLA_4 KS_1200(s1200, c1200, in1200_1, in1200_2);
    wire[3:0] s1201, in1201_1, in1201_2;
    wire c1201;
    assign in1201_1 = {pp62[97],pp63[97],pp64[97],pp65[97]};
    assign in1201_2 = {pp63[96],pp64[96],pp65[96],pp66[96]};
    CLA_4 KS_1201(s1201, c1201, in1201_1, in1201_2);
    wire[3:0] s1202, in1202_1, in1202_2;
    wire c1202;
    assign in1202_1 = {pp64[95],pp65[95],pp66[95],pp67[95]};
    assign in1202_2 = {pp65[94],pp66[94],pp67[94],pp68[94]};
    CLA_4 KS_1202(s1202, c1202, in1202_1, in1202_2);
    wire[3:0] s1203, in1203_1, in1203_2;
    wire c1203;
    assign in1203_1 = {pp66[93],pp67[93],pp68[93],pp69[93]};
    assign in1203_2 = {pp67[92],pp68[92],pp69[92],pp70[92]};
    CLA_4 KS_1203(s1203, c1203, in1203_1, in1203_2);
    wire[2:0] s1204, in1204_1, in1204_2;
    wire c1204;
    assign in1204_1 = {pp68[91],pp69[91],pp70[91]};
    assign in1204_2 = {pp69[90],pp70[90],pp71[90]};
    CLA_3 KS_1204(s1204, c1204, in1204_1, in1204_2);
    wire[1:0] s1205, in1205_1, in1205_2;
    wire c1205;
    assign in1205_1 = {pp70[89],pp71[89]};
    assign in1205_2 = {pp71[88],pp72[88]};
    CLA_2 KS_1205(s1205, c1205, in1205_1, in1205_2);
    wire[0:0] s1206, in1206_1, in1206_2;
    wire c1206;
    assign in1206_1 = {pp72[87]};
    assign in1206_2 = {pp73[86]};
    Half_Adder KS_1206(s1206, c1206, in1206_1, in1206_2);
    wire[3:0] s1207, in1207_1, in1207_2;
    wire c1207;
    assign in1207_1 = {pp74[85],pp73[87],pp72[89],pp71[91]};
    assign in1207_2 = {pp75[84],pp74[86],pp73[88],pp72[90]};
    CLA_4 KS_1207(s1207, c1207, in1207_1, in1207_2);
    wire[0:0] s1208, in1208_1, in1208_2;
    wire c1208;
    assign in1208_1 = {pp76[83]};
    assign in1208_2 = {pp77[82]};
    Half_Adder KS_1208(s1208, c1208, in1208_1, in1208_2);
    wire[1:0] s1209, in1209_1, in1209_2;
    wire c1209;
    assign in1209_1 = {pp78[81],pp75[85]};
    assign in1209_2 = {pp79[80],pp76[84]};
    CLA_2 KS_1209(s1209, c1209, in1209_1, in1209_2);
    wire[0:0] s1210, in1210_1, in1210_2;
    wire c1210;
    assign in1210_1 = {pp80[79]};
    assign in1210_2 = {pp81[78]};
    Half_Adder KS_1210(s1210, c1210, in1210_1, in1210_2);
    wire[2:0] s1211, in1211_1, in1211_2;
    wire c1211;
    assign in1211_1 = {pp82[77],pp77[83],pp74[87]};
    assign in1211_2 = {pp83[76],pp78[82],pp75[86]};
    CLA_3 KS_1211(s1211, c1211, in1211_1, in1211_2);
    wire[0:0] s1212, in1212_1, in1212_2;
    wire c1212;
    assign in1212_1 = {pp84[75]};
    assign in1212_2 = {pp85[74]};
    Half_Adder KS_1212(s1212, c1212, in1212_1, in1212_2);
    wire[1:0] s1213, in1213_1, in1213_2;
    wire c1213;
    assign in1213_1 = {pp86[73],pp79[81]};
    assign in1213_2 = {pp87[72],pp80[80]};
    CLA_2 KS_1213(s1213, c1213, in1213_1, in1213_2);
    wire[0:0] s1214, in1214_1, in1214_2;
    wire c1214;
    assign in1214_1 = {pp88[71]};
    assign in1214_2 = {pp89[70]};
    Half_Adder KS_1214(s1214, c1214, in1214_1, in1214_2);
    wire[3:0] s1215, in1215_1, in1215_2;
    wire c1215;
    assign in1215_1 = {pp90[69],pp81[79],pp76[85],pp73[89]};
    assign in1215_2 = {pp91[68],pp82[78],pp77[84],pp74[88]};
    CLA_4 KS_1215(s1215, c1215, in1215_1, in1215_2);
    wire[0:0] s1216, in1216_1, in1216_2;
    wire c1216;
    assign in1216_1 = {pp92[67]};
    assign in1216_2 = {pp93[66]};
    Half_Adder KS_1216(s1216, c1216, in1216_1, in1216_2);
    wire[1:0] s1217, in1217_1, in1217_2;
    wire c1217;
    assign in1217_1 = {pp94[65],pp83[77]};
    assign in1217_2 = {pp95[64],pp84[76]};
    CLA_2 KS_1217(s1217, c1217, in1217_1, in1217_2);
    wire[0:0] s1218, in1218_1, in1218_2;
    wire c1218;
    assign in1218_1 = {pp96[63]};
    assign in1218_2 = {pp97[62]};
    Half_Adder KS_1218(s1218, c1218, in1218_1, in1218_2);
    wire[2:0] s1219, in1219_1, in1219_2;
    wire c1219;
    assign in1219_1 = {pp98[61],pp85[75],pp78[83]};
    assign in1219_2 = {pp99[60],pp86[74],pp79[82]};
    CLA_3 KS_1219(s1219, c1219, in1219_1, in1219_2);
    wire[0:0] s1220, in1220_1, in1220_2;
    wire c1220;
    assign in1220_1 = {pp100[59]};
    assign in1220_2 = {pp101[58]};
    Half_Adder KS_1220(s1220, c1220, in1220_1, in1220_2);
    wire[1:0] s1221, in1221_1, in1221_2;
    wire c1221;
    assign in1221_1 = {pp102[57],pp87[73]};
    assign in1221_2 = {pp103[56],pp88[72]};
    CLA_2 KS_1221(s1221, c1221, in1221_1, in1221_2);
    wire[0:0] s1222, in1222_1, in1222_2;
    wire c1222;
    assign in1222_1 = {pp104[55]};
    assign in1222_2 = {pp105[54]};
    Half_Adder KS_1222(s1222, c1222, in1222_1, in1222_2);
    wire[3:0] s1223, in1223_1, in1223_2;
    wire c1223;
    assign in1223_1 = {pp106[53],pp89[71],pp80[81],pp75[87]};
    assign in1223_2 = {pp107[52],pp90[70],pp81[80],pp76[86]};
    CLA_4 KS_1223(s1223, c1223, in1223_1, in1223_2);
    wire[0:0] s1224, in1224_1, in1224_2;
    wire c1224;
    assign in1224_1 = {pp108[51]};
    assign in1224_2 = {pp109[50]};
    Half_Adder KS_1224(s1224, c1224, in1224_1, in1224_2);
    wire[1:0] s1225, in1225_1, in1225_2;
    wire c1225;
    assign in1225_1 = {pp110[49],pp91[69]};
    assign in1225_2 = {pp111[48],pp92[68]};
    CLA_2 KS_1225(s1225, c1225, in1225_1, in1225_2);
    wire[0:0] s1226, in1226_1, in1226_2;
    wire c1226;
    assign in1226_1 = {pp112[47]};
    assign in1226_2 = {pp113[46]};
    Half_Adder KS_1226(s1226, c1226, in1226_1, in1226_2);
    wire[2:0] s1227, in1227_1, in1227_2;
    wire c1227;
    assign in1227_1 = {pp114[45],pp93[67],pp82[79]};
    assign in1227_2 = {pp115[44],pp94[66],pp83[78]};
    CLA_3 KS_1227(s1227, c1227, in1227_1, in1227_2);
    wire[0:0] s1228, in1228_1, in1228_2;
    wire c1228;
    assign in1228_1 = {pp116[43]};
    assign in1228_2 = {pp117[42]};
    Half_Adder KS_1228(s1228, c1228, in1228_1, in1228_2);
    wire[1:0] s1229, in1229_1, in1229_2;
    wire c1229;
    assign in1229_1 = {pp118[41],pp95[65]};
    assign in1229_2 = {pp119[40],pp96[64]};
    CLA_2 KS_1229(s1229, c1229, in1229_1, in1229_2);
    wire[0:0] s1230, in1230_1, in1230_2;
    wire c1230;
    assign in1230_1 = {pp121[38]};
    assign in1230_2 = {pp122[37]};
    Full_Adder KS_1230(s1230, c1230, in1230_1, in1230_2, pp120[39]);
    wire[3:0] s1231, in1231_1, in1231_2;
    wire c1231;
    assign in1231_1 = {pp36[127],pp37[127],pp38[127],pp39[127]};
    assign in1231_2 = {pp37[126],pp38[126],pp39[126],pp40[126]};
    CLA_4 KS_1231(s1231, c1231, in1231_1, in1231_2);
    wire[3:0] s1232, in1232_1, in1232_2;
    wire c1232;
    assign in1232_1 = {pp38[125],pp39[125],pp40[125],pp41[125]};
    assign in1232_2 = {pp39[124],pp40[124],pp41[124],pp42[124]};
    CLA_4 KS_1232(s1232, c1232, in1232_1, in1232_2);
    wire[3:0] s1233, in1233_1, in1233_2;
    wire c1233;
    assign in1233_1 = {pp40[123],pp41[123],pp42[123],pp43[123]};
    assign in1233_2 = {pp41[122],pp42[122],pp43[122],pp44[122]};
    CLA_4 KS_1233(s1233, c1233, in1233_1, in1233_2);
    wire[3:0] s1234, in1234_1, in1234_2;
    wire c1234;
    assign in1234_1 = {pp42[121],pp43[121],pp44[121],pp45[121]};
    assign in1234_2 = {pp43[120],pp44[120],pp45[120],pp46[120]};
    CLA_4 KS_1234(s1234, c1234, in1234_1, in1234_2);
    wire[3:0] s1235, in1235_1, in1235_2;
    wire c1235;
    assign in1235_1 = {pp44[119],pp45[119],pp46[119],pp47[119]};
    assign in1235_2 = {pp45[118],pp46[118],pp47[118],pp48[118]};
    CLA_4 KS_1235(s1235, c1235, in1235_1, in1235_2);
    wire[3:0] s1236, in1236_1, in1236_2;
    wire c1236;
    assign in1236_1 = {pp46[117],pp47[117],pp48[117],pp49[117]};
    assign in1236_2 = {pp47[116],pp48[116],pp49[116],pp50[116]};
    CLA_4 KS_1236(s1236, c1236, in1236_1, in1236_2);
    wire[3:0] s1237, in1237_1, in1237_2;
    wire c1237;
    assign in1237_1 = {pp48[115],pp49[115],pp50[115],pp51[115]};
    assign in1237_2 = {pp49[114],pp50[114],pp51[114],pp52[114]};
    CLA_4 KS_1237(s1237, c1237, in1237_1, in1237_2);
    wire[3:0] s1238, in1238_1, in1238_2;
    wire c1238;
    assign in1238_1 = {pp50[113],pp51[113],pp52[113],pp53[113]};
    assign in1238_2 = {pp51[112],pp52[112],pp53[112],pp54[112]};
    CLA_4 KS_1238(s1238, c1238, in1238_1, in1238_2);
    wire[3:0] s1239, in1239_1, in1239_2;
    wire c1239;
    assign in1239_1 = {pp52[111],pp53[111],pp54[111],pp55[111]};
    assign in1239_2 = {pp53[110],pp54[110],pp55[110],pp56[110]};
    CLA_4 KS_1239(s1239, c1239, in1239_1, in1239_2);
    wire[3:0] s1240, in1240_1, in1240_2;
    wire c1240;
    assign in1240_1 = {pp54[109],pp55[109],pp56[109],pp57[109]};
    assign in1240_2 = {pp55[108],pp56[108],pp57[108],pp58[108]};
    CLA_4 KS_1240(s1240, c1240, in1240_1, in1240_2);
    wire[3:0] s1241, in1241_1, in1241_2;
    wire c1241;
    assign in1241_1 = {pp56[107],pp57[107],pp58[107],pp59[107]};
    assign in1241_2 = {pp57[106],pp58[106],pp59[106],pp60[106]};
    CLA_4 KS_1241(s1241, c1241, in1241_1, in1241_2);
    wire[3:0] s1242, in1242_1, in1242_2;
    wire c1242;
    assign in1242_1 = {pp58[105],pp59[105],pp60[105],pp61[105]};
    assign in1242_2 = {pp59[104],pp60[104],pp61[104],pp62[104]};
    CLA_4 KS_1242(s1242, c1242, in1242_1, in1242_2);
    wire[3:0] s1243, in1243_1, in1243_2;
    wire c1243;
    assign in1243_1 = {pp60[103],pp61[103],pp62[103],pp63[103]};
    assign in1243_2 = {pp61[102],pp62[102],pp63[102],pp64[102]};
    CLA_4 KS_1243(s1243, c1243, in1243_1, in1243_2);
    wire[3:0] s1244, in1244_1, in1244_2;
    wire c1244;
    assign in1244_1 = {pp62[101],pp63[101],pp64[101],pp65[101]};
    assign in1244_2 = {pp63[100],pp64[100],pp65[100],pp66[100]};
    CLA_4 KS_1244(s1244, c1244, in1244_1, in1244_2);
    wire[2:0] s1245, in1245_1, in1245_2;
    wire c1245;
    assign in1245_1 = {pp64[99],pp65[99],pp66[99]};
    assign in1245_2 = {pp65[98],pp66[98],pp67[98]};
    CLA_3 KS_1245(s1245, c1245, in1245_1, in1245_2);
    wire[1:0] s1246, in1246_1, in1246_2;
    wire c1246;
    assign in1246_1 = {pp66[97],pp67[97]};
    assign in1246_2 = {pp67[96],pp68[96]};
    CLA_2 KS_1246(s1246, c1246, in1246_1, in1246_2);
    wire[0:0] s1247, in1247_1, in1247_2;
    wire c1247;
    assign in1247_1 = {pp68[95]};
    assign in1247_2 = {pp69[94]};
    Half_Adder KS_1247(s1247, c1247, in1247_1, in1247_2);
    wire[3:0] s1248, in1248_1, in1248_2;
    wire c1248;
    assign in1248_1 = {pp70[93],pp69[95],pp68[97],pp67[99]};
    assign in1248_2 = {pp71[92],pp70[94],pp69[96],pp68[98]};
    CLA_4 KS_1248(s1248, c1248, in1248_1, in1248_2);
    wire[0:0] s1249, in1249_1, in1249_2;
    wire c1249;
    assign in1249_1 = {pp72[91]};
    assign in1249_2 = {pp73[90]};
    Half_Adder KS_1249(s1249, c1249, in1249_1, in1249_2);
    wire[1:0] s1250, in1250_1, in1250_2;
    wire c1250;
    assign in1250_1 = {pp74[89],pp71[93]};
    assign in1250_2 = {pp75[88],pp72[92]};
    CLA_2 KS_1250(s1250, c1250, in1250_1, in1250_2);
    wire[0:0] s1251, in1251_1, in1251_2;
    wire c1251;
    assign in1251_1 = {pp76[87]};
    assign in1251_2 = {pp77[86]};
    Half_Adder KS_1251(s1251, c1251, in1251_1, in1251_2);
    wire[2:0] s1252, in1252_1, in1252_2;
    wire c1252;
    assign in1252_1 = {pp78[85],pp73[91],pp70[95]};
    assign in1252_2 = {pp79[84],pp74[90],pp71[94]};
    CLA_3 KS_1252(s1252, c1252, in1252_1, in1252_2);
    wire[0:0] s1253, in1253_1, in1253_2;
    wire c1253;
    assign in1253_1 = {pp80[83]};
    assign in1253_2 = {pp81[82]};
    Half_Adder KS_1253(s1253, c1253, in1253_1, in1253_2);
    wire[1:0] s1254, in1254_1, in1254_2;
    wire c1254;
    assign in1254_1 = {pp82[81],pp75[89]};
    assign in1254_2 = {pp83[80],pp76[88]};
    CLA_2 KS_1254(s1254, c1254, in1254_1, in1254_2);
    wire[0:0] s1255, in1255_1, in1255_2;
    wire c1255;
    assign in1255_1 = {pp84[79]};
    assign in1255_2 = {pp85[78]};
    Half_Adder KS_1255(s1255, c1255, in1255_1, in1255_2);
    wire[3:0] s1256, in1256_1, in1256_2;
    wire c1256;
    assign in1256_1 = {pp86[77],pp77[87],pp72[93],pp69[97]};
    assign in1256_2 = {pp87[76],pp78[86],pp73[92],pp70[96]};
    CLA_4 KS_1256(s1256, c1256, in1256_1, in1256_2);
    wire[0:0] s1257, in1257_1, in1257_2;
    wire c1257;
    assign in1257_1 = {pp88[75]};
    assign in1257_2 = {pp89[74]};
    Half_Adder KS_1257(s1257, c1257, in1257_1, in1257_2);
    wire[1:0] s1258, in1258_1, in1258_2;
    wire c1258;
    assign in1258_1 = {pp90[73],pp79[85]};
    assign in1258_2 = {pp91[72],pp80[84]};
    CLA_2 KS_1258(s1258, c1258, in1258_1, in1258_2);
    wire[0:0] s1259, in1259_1, in1259_2;
    wire c1259;
    assign in1259_1 = {pp92[71]};
    assign in1259_2 = {pp93[70]};
    Half_Adder KS_1259(s1259, c1259, in1259_1, in1259_2);
    wire[2:0] s1260, in1260_1, in1260_2;
    wire c1260;
    assign in1260_1 = {pp94[69],pp81[83],pp74[91]};
    assign in1260_2 = {pp95[68],pp82[82],pp75[90]};
    CLA_3 KS_1260(s1260, c1260, in1260_1, in1260_2);
    wire[0:0] s1261, in1261_1, in1261_2;
    wire c1261;
    assign in1261_1 = {pp96[67]};
    assign in1261_2 = {pp97[66]};
    Half_Adder KS_1261(s1261, c1261, in1261_1, in1261_2);
    wire[1:0] s1262, in1262_1, in1262_2;
    wire c1262;
    assign in1262_1 = {pp98[65],pp83[81]};
    assign in1262_2 = {pp99[64],pp84[80]};
    CLA_2 KS_1262(s1262, c1262, in1262_1, in1262_2);
    wire[0:0] s1263, in1263_1, in1263_2;
    wire c1263;
    assign in1263_1 = {pp100[63]};
    assign in1263_2 = {pp101[62]};
    Half_Adder KS_1263(s1263, c1263, in1263_1, in1263_2);
    wire[3:0] s1264, in1264_1, in1264_2;
    wire c1264;
    assign in1264_1 = {pp102[61],pp85[79],pp76[89],pp71[95]};
    assign in1264_2 = {pp103[60],pp86[78],pp77[88],pp72[94]};
    CLA_4 KS_1264(s1264, c1264, in1264_1, in1264_2);
    wire[0:0] s1265, in1265_1, in1265_2;
    wire c1265;
    assign in1265_1 = {pp104[59]};
    assign in1265_2 = {pp105[58]};
    Half_Adder KS_1265(s1265, c1265, in1265_1, in1265_2);
    wire[1:0] s1266, in1266_1, in1266_2;
    wire c1266;
    assign in1266_1 = {pp107[56],pp87[77]};
    assign in1266_2 = {pp108[55],pp88[76]};
    CLA_2_c KS_1266(s1266, c1266, in1266_1, in1266_2, pp106[57]);
    wire[3:0] s1267, in1267_1, in1267_2;
    wire c1267;
    assign in1267_1 = {pp40[127],pp41[127],pp42[127],pp43[127]};
    assign in1267_2 = {pp41[126],pp42[126],pp43[126],pp44[126]};
    CLA_4 KS_1267(s1267, c1267, in1267_1, in1267_2);
    wire[3:0] s1268, in1268_1, in1268_2;
    wire c1268;
    assign in1268_1 = {pp42[125],pp43[125],pp44[125],pp45[125]};
    assign in1268_2 = {pp43[124],pp44[124],pp45[124],pp46[124]};
    CLA_4 KS_1268(s1268, c1268, in1268_1, in1268_2);
    wire[3:0] s1269, in1269_1, in1269_2;
    wire c1269;
    assign in1269_1 = {pp44[123],pp45[123],pp46[123],pp47[123]};
    assign in1269_2 = {pp45[122],pp46[122],pp47[122],pp48[122]};
    CLA_4 KS_1269(s1269, c1269, in1269_1, in1269_2);
    wire[3:0] s1270, in1270_1, in1270_2;
    wire c1270;
    assign in1270_1 = {pp46[121],pp47[121],pp48[121],pp49[121]};
    assign in1270_2 = {pp47[120],pp48[120],pp49[120],pp50[120]};
    CLA_4 KS_1270(s1270, c1270, in1270_1, in1270_2);
    wire[3:0] s1271, in1271_1, in1271_2;
    wire c1271;
    assign in1271_1 = {pp48[119],pp49[119],pp50[119],pp51[119]};
    assign in1271_2 = {pp49[118],pp50[118],pp51[118],pp52[118]};
    CLA_4 KS_1271(s1271, c1271, in1271_1, in1271_2);
    wire[3:0] s1272, in1272_1, in1272_2;
    wire c1272;
    assign in1272_1 = {pp50[117],pp51[117],pp52[117],pp53[117]};
    assign in1272_2 = {pp51[116],pp52[116],pp53[116],pp54[116]};
    CLA_4 KS_1272(s1272, c1272, in1272_1, in1272_2);
    wire[3:0] s1273, in1273_1, in1273_2;
    wire c1273;
    assign in1273_1 = {pp52[115],pp53[115],pp54[115],pp55[115]};
    assign in1273_2 = {pp53[114],pp54[114],pp55[114],pp56[114]};
    CLA_4 KS_1273(s1273, c1273, in1273_1, in1273_2);
    wire[3:0] s1274, in1274_1, in1274_2;
    wire c1274;
    assign in1274_1 = {pp54[113],pp55[113],pp56[113],pp57[113]};
    assign in1274_2 = {pp55[112],pp56[112],pp57[112],pp58[112]};
    CLA_4 KS_1274(s1274, c1274, in1274_1, in1274_2);
    wire[3:0] s1275, in1275_1, in1275_2;
    wire c1275;
    assign in1275_1 = {pp56[111],pp57[111],pp58[111],pp59[111]};
    assign in1275_2 = {pp57[110],pp58[110],pp59[110],pp60[110]};
    CLA_4 KS_1275(s1275, c1275, in1275_1, in1275_2);
    wire[3:0] s1276, in1276_1, in1276_2;
    wire c1276;
    assign in1276_1 = {pp58[109],pp59[109],pp60[109],pp61[109]};
    assign in1276_2 = {pp59[108],pp60[108],pp61[108],pp62[108]};
    CLA_4 KS_1276(s1276, c1276, in1276_1, in1276_2);
    wire[2:0] s1277, in1277_1, in1277_2;
    wire c1277;
    assign in1277_1 = {pp60[107],pp61[107],pp62[107]};
    assign in1277_2 = {pp61[106],pp62[106],pp63[106]};
    CLA_3 KS_1277(s1277, c1277, in1277_1, in1277_2);
    wire[1:0] s1278, in1278_1, in1278_2;
    wire c1278;
    assign in1278_1 = {pp62[105],pp63[105]};
    assign in1278_2 = {pp63[104],pp64[104]};
    CLA_2 KS_1278(s1278, c1278, in1278_1, in1278_2);
    wire[0:0] s1279, in1279_1, in1279_2;
    wire c1279;
    assign in1279_1 = {pp64[103]};
    assign in1279_2 = {pp65[102]};
    Half_Adder KS_1279(s1279, c1279, in1279_1, in1279_2);
    wire[3:0] s1280, in1280_1, in1280_2;
    wire c1280;
    assign in1280_1 = {pp66[101],pp65[103],pp64[105],pp63[107]};
    assign in1280_2 = {pp67[100],pp66[102],pp65[104],pp64[106]};
    CLA_4 KS_1280(s1280, c1280, in1280_1, in1280_2);
    wire[0:0] s1281, in1281_1, in1281_2;
    wire c1281;
    assign in1281_1 = {pp68[99]};
    assign in1281_2 = {pp69[98]};
    Half_Adder KS_1281(s1281, c1281, in1281_1, in1281_2);
    wire[1:0] s1282, in1282_1, in1282_2;
    wire c1282;
    assign in1282_1 = {pp70[97],pp67[101]};
    assign in1282_2 = {pp71[96],pp68[100]};
    CLA_2 KS_1282(s1282, c1282, in1282_1, in1282_2);
    wire[0:0] s1283, in1283_1, in1283_2;
    wire c1283;
    assign in1283_1 = {pp72[95]};
    assign in1283_2 = {pp73[94]};
    Half_Adder KS_1283(s1283, c1283, in1283_1, in1283_2);
    wire[2:0] s1284, in1284_1, in1284_2;
    wire c1284;
    assign in1284_1 = {pp74[93],pp69[99],pp66[103]};
    assign in1284_2 = {pp75[92],pp70[98],pp67[102]};
    CLA_3 KS_1284(s1284, c1284, in1284_1, in1284_2);
    wire[0:0] s1285, in1285_1, in1285_2;
    wire c1285;
    assign in1285_1 = {pp76[91]};
    assign in1285_2 = {pp77[90]};
    Half_Adder KS_1285(s1285, c1285, in1285_1, in1285_2);
    wire[1:0] s1286, in1286_1, in1286_2;
    wire c1286;
    assign in1286_1 = {pp78[89],pp71[97]};
    assign in1286_2 = {pp79[88],pp72[96]};
    CLA_2 KS_1286(s1286, c1286, in1286_1, in1286_2);
    wire[0:0] s1287, in1287_1, in1287_2;
    wire c1287;
    assign in1287_1 = {pp80[87]};
    assign in1287_2 = {pp81[86]};
    Half_Adder KS_1287(s1287, c1287, in1287_1, in1287_2);
    wire[3:0] s1288, in1288_1, in1288_2;
    wire c1288;
    assign in1288_1 = {pp82[85],pp73[95],pp68[101],pp65[105]};
    assign in1288_2 = {pp83[84],pp74[94],pp69[100],pp66[104]};
    CLA_4 KS_1288(s1288, c1288, in1288_1, in1288_2);
    wire[0:0] s1289, in1289_1, in1289_2;
    wire c1289;
    assign in1289_1 = {pp84[83]};
    assign in1289_2 = {pp85[82]};
    Half_Adder KS_1289(s1289, c1289, in1289_1, in1289_2);
    wire[1:0] s1290, in1290_1, in1290_2;
    wire c1290;
    assign in1290_1 = {pp86[81],pp75[93]};
    assign in1290_2 = {pp87[80],pp76[92]};
    CLA_2 KS_1290(s1290, c1290, in1290_1, in1290_2);
    wire[0:0] s1291, in1291_1, in1291_2;
    wire c1291;
    assign in1291_1 = {pp88[79]};
    assign in1291_2 = {pp89[78]};
    Half_Adder KS_1291(s1291, c1291, in1291_1, in1291_2);
    wire[2:0] s1292, in1292_1, in1292_2;
    wire c1292;
    assign in1292_1 = {pp90[77],pp77[91],pp70[99]};
    assign in1292_2 = {pp91[76],pp78[90],pp71[98]};
    CLA_3 KS_1292(s1292, c1292, in1292_1, in1292_2);
    wire[0:0] s1293, in1293_1, in1293_2;
    wire c1293;
    assign in1293_1 = {pp92[75]};
    assign in1293_2 = {pp93[74]};
    Half_Adder KS_1293(s1293, c1293, in1293_1, in1293_2);
    wire[1:0] s1294, in1294_1, in1294_2;
    wire c1294;
    assign in1294_1 = {pp95[72],pp79[89]};
    assign in1294_2 = {pp96[71],pp80[88]};
    CLA_2_c KS_1294(s1294, c1294, in1294_1, in1294_2, pp94[73]);
    wire[3:0] s1295, in1295_1, in1295_2;
    wire c1295;
    assign in1295_1 = {pp44[127],pp45[127],pp46[127],pp47[127]};
    assign in1295_2 = {pp45[126],pp46[126],pp47[126],pp48[126]};
    CLA_4 KS_1295(s1295, c1295, in1295_1, in1295_2);
    wire[3:0] s1296, in1296_1, in1296_2;
    wire c1296;
    assign in1296_1 = {pp46[125],pp47[125],pp48[125],pp49[125]};
    assign in1296_2 = {pp47[124],pp48[124],pp49[124],pp50[124]};
    CLA_4 KS_1296(s1296, c1296, in1296_1, in1296_2);
    wire[3:0] s1297, in1297_1, in1297_2;
    wire c1297;
    assign in1297_1 = {pp48[123],pp49[123],pp50[123],pp51[123]};
    assign in1297_2 = {pp49[122],pp50[122],pp51[122],pp52[122]};
    CLA_4 KS_1297(s1297, c1297, in1297_1, in1297_2);
    wire[3:0] s1298, in1298_1, in1298_2;
    wire c1298;
    assign in1298_1 = {pp50[121],pp51[121],pp52[121],pp53[121]};
    assign in1298_2 = {pp51[120],pp52[120],pp53[120],pp54[120]};
    CLA_4 KS_1298(s1298, c1298, in1298_1, in1298_2);
    wire[3:0] s1299, in1299_1, in1299_2;
    wire c1299;
    assign in1299_1 = {pp52[119],pp53[119],pp54[119],pp55[119]};
    assign in1299_2 = {pp53[118],pp54[118],pp55[118],pp56[118]};
    CLA_4 KS_1299(s1299, c1299, in1299_1, in1299_2);
    wire[3:0] s1300, in1300_1, in1300_2;
    wire c1300;
    assign in1300_1 = {pp54[117],pp55[117],pp56[117],pp57[117]};
    assign in1300_2 = {pp55[116],pp56[116],pp57[116],pp58[116]};
    CLA_4 KS_1300(s1300, c1300, in1300_1, in1300_2);
    wire[2:0] s1301, in1301_1, in1301_2;
    wire c1301;
    assign in1301_1 = {pp56[115],pp57[115],pp58[115]};
    assign in1301_2 = {pp57[114],pp58[114],pp59[114]};
    CLA_3 KS_1301(s1301, c1301, in1301_1, in1301_2);
    wire[1:0] s1302, in1302_1, in1302_2;
    wire c1302;
    assign in1302_1 = {pp58[113],pp59[113]};
    assign in1302_2 = {pp59[112],pp60[112]};
    CLA_2 KS_1302(s1302, c1302, in1302_1, in1302_2);
    wire[0:0] s1303, in1303_1, in1303_2;
    wire c1303;
    assign in1303_1 = {pp60[111]};
    assign in1303_2 = {pp61[110]};
    Half_Adder KS_1303(s1303, c1303, in1303_1, in1303_2);
    wire[3:0] s1304, in1304_1, in1304_2;
    wire c1304;
    assign in1304_1 = {pp62[109],pp61[111],pp60[113],pp59[115]};
    assign in1304_2 = {pp63[108],pp62[110],pp61[112],pp60[114]};
    CLA_4 KS_1304(s1304, c1304, in1304_1, in1304_2);
    wire[0:0] s1305, in1305_1, in1305_2;
    wire c1305;
    assign in1305_1 = {pp64[107]};
    assign in1305_2 = {pp65[106]};
    Half_Adder KS_1305(s1305, c1305, in1305_1, in1305_2);
    wire[1:0] s1306, in1306_1, in1306_2;
    wire c1306;
    assign in1306_1 = {pp66[105],pp63[109]};
    assign in1306_2 = {pp67[104],pp64[108]};
    CLA_2 KS_1306(s1306, c1306, in1306_1, in1306_2);
    wire[0:0] s1307, in1307_1, in1307_2;
    wire c1307;
    assign in1307_1 = {pp68[103]};
    assign in1307_2 = {pp69[102]};
    Half_Adder KS_1307(s1307, c1307, in1307_1, in1307_2);
    wire[2:0] s1308, in1308_1, in1308_2;
    wire c1308;
    assign in1308_1 = {pp70[101],pp65[107],pp62[111]};
    assign in1308_2 = {pp71[100],pp66[106],pp63[110]};
    CLA_3 KS_1308(s1308, c1308, in1308_1, in1308_2);
    wire[0:0] s1309, in1309_1, in1309_2;
    wire c1309;
    assign in1309_1 = {pp72[99]};
    assign in1309_2 = {pp73[98]};
    Half_Adder KS_1309(s1309, c1309, in1309_1, in1309_2);
    wire[1:0] s1310, in1310_1, in1310_2;
    wire c1310;
    assign in1310_1 = {pp74[97],pp67[105]};
    assign in1310_2 = {pp75[96],pp68[104]};
    CLA_2 KS_1310(s1310, c1310, in1310_1, in1310_2);
    wire[0:0] s1311, in1311_1, in1311_2;
    wire c1311;
    assign in1311_1 = {pp76[95]};
    assign in1311_2 = {pp77[94]};
    Half_Adder KS_1311(s1311, c1311, in1311_1, in1311_2);
    wire[3:0] s1312, in1312_1, in1312_2;
    wire c1312;
    assign in1312_1 = {pp78[93],pp69[103],pp64[109],pp61[113]};
    assign in1312_2 = {pp79[92],pp70[102],pp65[108],pp62[112]};
    CLA_4 KS_1312(s1312, c1312, in1312_1, in1312_2);
    wire[0:0] s1313, in1313_1, in1313_2;
    wire c1313;
    assign in1313_1 = {pp81[90]};
    assign in1313_2 = {pp82[89]};
    Full_Adder KS_1313(s1313, c1313, in1313_1, in1313_2, pp80[91]);
    wire[3:0] s1314, in1314_1, in1314_2;
    wire c1314;
    assign in1314_1 = {pp48[127],pp49[127],pp50[127],pp51[127]};
    assign in1314_2 = {pp49[126],pp50[126],pp51[126],pp52[126]};
    CLA_4 KS_1314(s1314, c1314, in1314_1, in1314_2);
    wire[3:0] s1315, in1315_1, in1315_2;
    wire c1315;
    assign in1315_1 = {pp50[125],pp51[125],pp52[125],pp53[125]};
    assign in1315_2 = {pp51[124],pp52[124],pp53[124],pp54[124]};
    CLA_4 KS_1315(s1315, c1315, in1315_1, in1315_2);
    wire[2:0] s1316, in1316_1, in1316_2;
    wire c1316;
    assign in1316_1 = {pp52[123],pp53[123],pp54[123]};
    assign in1316_2 = {pp53[122],pp54[122],pp55[122]};
    CLA_3 KS_1316(s1316, c1316, in1316_1, in1316_2);
    wire[1:0] s1317, in1317_1, in1317_2;
    wire c1317;
    assign in1317_1 = {pp54[121],pp55[121]};
    assign in1317_2 = {pp55[120],pp56[120]};
    CLA_2 KS_1317(s1317, c1317, in1317_1, in1317_2);
    wire[0:0] s1318, in1318_1, in1318_2;
    wire c1318;
    assign in1318_1 = {pp56[119]};
    assign in1318_2 = {pp57[118]};
    Half_Adder KS_1318(s1318, c1318, in1318_1, in1318_2);
    wire[3:0] s1319, in1319_1, in1319_2;
    wire c1319;
    assign in1319_1 = {pp58[117],pp57[119],pp56[121],pp55[123]};
    assign in1319_2 = {pp59[116],pp58[118],pp57[120],pp56[122]};
    CLA_4 KS_1319(s1319, c1319, in1319_1, in1319_2);
    wire[0:0] s1320, in1320_1, in1320_2;
    wire c1320;
    assign in1320_1 = {pp60[115]};
    assign in1320_2 = {pp61[114]};
    Half_Adder KS_1320(s1320, c1320, in1320_1, in1320_2);
    wire[1:0] s1321, in1321_1, in1321_2;
    wire c1321;
    assign in1321_1 = {pp62[113],pp59[117]};
    assign in1321_2 = {pp63[112],pp60[116]};
    CLA_2 KS_1321(s1321, c1321, in1321_1, in1321_2);
    wire[0:0] s1322, in1322_1, in1322_2;
    wire c1322;
    assign in1322_1 = {pp64[111]};
    assign in1322_2 = {pp65[110]};
    Half_Adder KS_1322(s1322, c1322, in1322_1, in1322_2);
    wire[2:0] s1323, in1323_1, in1323_2;
    wire c1323;
    assign in1323_1 = {pp66[109],pp61[115],pp58[119]};
    assign in1323_2 = {pp67[108],pp62[114],pp59[118]};
    CLA_3 KS_1323(s1323, c1323, in1323_1, in1323_2);
    wire[0:0] s1324, in1324_1, in1324_2;
    wire c1324;
    assign in1324_1 = {pp69[106]};
    assign in1324_2 = {pp70[105]};
    Full_Adder KS_1324(s1324, c1324, in1324_1, in1324_2, pp68[107]);
    wire[0:0] s1325, in1325_1, in1325_2;
    wire c1325;
    assign in1325_1 = {pp52[127]};
    assign in1325_2 = {pp53[126]};
    Half_Adder KS_1325(s1325, c1325, in1325_1, in1325_2);
    wire[1:0] s1326, in1326_1, in1326_2;
    wire c1326;
    assign in1326_1 = {pp55[124],pp53[127]};
    assign in1326_2 = {pp56[123],pp54[126]};
    CLA_2_c KS_1326(s1326, c1326, in1326_1, in1326_2, pp54[125]);

    /*Stage 2*/
    wire[3:0] s1327, in1327_1, in1327_2;
    wire c1327;
    assign in1327_1 = {pp0[45],pp0[46],pp0[47],pp0[48]};
    assign in1327_2 = {pp1[44],pp1[45],pp1[46],pp1[47]};
    CLA_4 KS_1327(s1327, c1327, in1327_1, in1327_2);
    wire[3:0] s1328, in1328_1, in1328_2;
    wire c1328;
    assign in1328_1 = {pp2[44],pp2[45],pp2[46],pp0[49]};
    assign in1328_2 = {pp3[43],pp3[44],pp3[45],pp1[48]};
    CLA_4 KS_1328(s1328, c1328, in1328_1, in1328_2);
    wire[3:0] s1329, in1329_1, in1329_2;
    wire c1329;
    assign in1329_1 = {pp4[43],pp4[44],pp2[47],pp0[50]};
    assign in1329_2 = {pp5[42],pp5[43],pp3[46],pp1[49]};
    CLA_4 KS_1329(s1329, c1329, in1329_1, in1329_2);
    wire[3:0] s1330, in1330_1, in1330_2;
    wire c1330;
    assign in1330_1 = {pp6[42],pp4[45],pp2[48],pp0[51]};
    assign in1330_2 = {pp7[41],pp5[44],pp3[47],pp1[50]};
    CLA_4 KS_1330(s1330, c1330, in1330_1, in1330_2);
    wire[3:0] s1331, in1331_1, in1331_2;
    wire c1331;
    assign in1331_1 = {pp6[43],pp4[46],pp2[49],pp0[52]};
    assign in1331_2 = {pp7[42],pp5[45],pp3[48],pp1[51]};
    CLA_4 KS_1331(s1331, c1331, in1331_1, in1331_2);
    wire[3:0] s1332, in1332_1, in1332_2;
    wire c1332;
    assign in1332_1 = {pp9[40],pp6[44],pp4[47],pp2[50]};
    assign in1332_2 = {pp10[39],pp7[43],pp5[46],pp3[49]};
    CLA_4_c KS_1332(s1332, c1332, in1332_1, in1332_2, pp8[41]);
    wire[3:0] s1333, in1333_1, in1333_2;
    wire c1333;
    assign in1333_1 = {pp8[42],pp6[45],pp4[48],pp0[53]};
    assign in1333_2 = {pp9[41],pp7[44],pp5[47],pp1[52]};
    CLA_4 KS_1333(s1333, c1333, in1333_1, in1333_2);
    wire[3:0] s1334, in1334_1, in1334_2;
    wire c1334;
    assign in1334_1 = {pp11[39],pp8[43],pp6[46],pp2[51]};
    assign in1334_2 = {pp12[38],pp9[42],pp7[45],pp3[50]};
    CLA_4_c KS_1334(s1334, c1334, in1334_1, in1334_2, pp10[40]);
    wire[3:0] s1335, in1335_1, in1335_2;
    wire c1335;
    assign in1335_1 = {pp10[41],pp8[44],pp4[49],pp0[54]};
    assign in1335_2 = {pp11[40],pp9[43],pp5[48],pp1[53]};
    CLA_4 KS_1335(s1335, c1335, in1335_1, in1335_2);
    wire[3:0] s1336, in1336_1, in1336_2;
    wire c1336;
    assign in1336_1 = {pp13[38],pp10[42],pp6[47],pp2[52]};
    assign in1336_2 = {pp14[37],pp11[41],pp7[46],pp3[51]};
    CLA_4_c KS_1336(s1336, c1336, in1336_1, in1336_2, pp12[39]);
    wire[3:0] s1337, in1337_1, in1337_2;
    wire c1337;
    assign in1337_1 = {pp12[40],pp8[45],pp4[50],pp0[55]};
    assign in1337_2 = {pp13[39],pp9[44],pp5[49],pp1[54]};
    CLA_4 KS_1337(s1337, c1337, in1337_1, in1337_2);
    wire[3:0] s1338, in1338_1, in1338_2;
    wire c1338;
    assign in1338_1 = {pp15[37],pp10[43],pp6[48],pp2[53]};
    assign in1338_2 = {pp16[36],pp11[42],pp7[47],pp3[52]};
    CLA_4_c KS_1338(s1338, c1338, in1338_1, in1338_2, pp14[38]);
    wire[3:0] s1339, in1339_1, in1339_2;
    wire c1339;
    assign in1339_1 = {pp12[41],pp8[46],pp4[51],pp0[56]};
    assign in1339_2 = {pp13[40],pp9[45],pp5[50],pp1[55]};
    CLA_4 KS_1339(s1339, c1339, in1339_1, in1339_2);
    wire[3:0] s1340, in1340_1, in1340_2;
    wire c1340;
    assign in1340_1 = {pp14[39],pp10[44],pp6[49],pp2[54]};
    assign in1340_2 = {pp15[38],pp11[43],pp7[48],pp3[53]};
    CLA_4 KS_1340(s1340, c1340, in1340_1, in1340_2);
    wire[3:0] s1341, in1341_1, in1341_2;
    wire c1341;
    assign in1341_1 = {pp16[37],pp12[42],pp8[47],pp4[52]};
    assign in1341_2 = {pp17[36],pp13[41],pp9[46],pp5[51]};
    CLA_4 KS_1341(s1341, c1341, in1341_1, in1341_2);
    wire[3:0] s1342, in1342_1, in1342_2;
    wire c1342;
    assign in1342_1 = {pp19[34],pp14[40],pp10[45],pp6[50]};
    assign in1342_2 = {pp20[33],pp15[39],pp11[44],pp7[49]};
    CLA_4_c KS_1342(s1342, c1342, in1342_1, in1342_2, pp18[35]);
    wire[3:0] s1343, in1343_1, in1343_2;
    wire c1343;
    assign in1343_1 = {pp16[38],pp12[43],pp8[48],pp0[57]};
    assign in1343_2 = {pp17[37],pp13[42],pp9[47],pp1[56]};
    CLA_4 KS_1343(s1343, c1343, in1343_1, in1343_2);
    wire[3:0] s1344, in1344_1, in1344_2;
    wire c1344;
    assign in1344_1 = {pp18[36],pp14[41],pp10[46],pp2[55]};
    assign in1344_2 = {pp19[35],pp15[40],pp11[45],pp3[54]};
    CLA_4 KS_1344(s1344, c1344, in1344_1, in1344_2);
    wire[3:0] s1345, in1345_1, in1345_2;
    wire c1345;
    assign in1345_1 = {pp21[33],pp16[39],pp12[44],pp4[53]};
    assign in1345_2 = {pp22[32],pp17[38],pp13[43],pp5[52]};
    CLA_4_c KS_1345(s1345, c1345, in1345_1, in1345_2, pp20[34]);
    wire[3:0] s1346, in1346_1, in1346_2;
    wire c1346;
    assign in1346_1 = {pp18[37],pp14[42],pp6[51],pp0[58]};
    assign in1346_2 = {pp19[36],pp15[41],pp7[50],pp1[57]};
    CLA_4 KS_1346(s1346, c1346, in1346_1, in1346_2);
    wire[3:0] s1347, in1347_1, in1347_2;
    wire c1347;
    assign in1347_1 = {pp20[35],pp16[40],pp8[49],pp2[56]};
    assign in1347_2 = {pp21[34],pp17[39],pp9[48],pp3[55]};
    CLA_4 KS_1347(s1347, c1347, in1347_1, in1347_2);
    wire[3:0] s1348, in1348_1, in1348_2;
    wire c1348;
    assign in1348_1 = {pp23[32],pp18[38],pp10[47],pp4[54]};
    assign in1348_2 = {pp24[31],pp19[37],pp11[46],pp5[53]};
    CLA_4_c KS_1348(s1348, c1348, in1348_1, in1348_2, pp22[33]);
    wire[3:0] s1349, in1349_1, in1349_2;
    wire c1349;
    assign in1349_1 = {pp20[36],pp12[45],pp6[52],pp0[59]};
    assign in1349_2 = {pp21[35],pp13[44],pp7[51],pp1[58]};
    CLA_4 KS_1349(s1349, c1349, in1349_1, in1349_2);
    wire[3:0] s1350, in1350_1, in1350_2;
    wire c1350;
    assign in1350_1 = {pp22[34],pp14[43],pp8[50],pp2[57]};
    assign in1350_2 = {pp23[33],pp15[42],pp9[49],pp3[56]};
    CLA_4 KS_1350(s1350, c1350, in1350_1, in1350_2);
    wire[3:0] s1351, in1351_1, in1351_2;
    wire c1351;
    assign in1351_1 = {pp25[31],pp16[41],pp10[48],pp4[55]};
    assign in1351_2 = {pp26[30],pp17[40],pp11[47],pp5[54]};
    CLA_4_c KS_1351(s1351, c1351, in1351_1, in1351_2, pp24[32]);
    wire[3:0] s1352, in1352_1, in1352_2;
    wire c1352;
    assign in1352_1 = {pp18[39],pp12[46],pp6[53],pp0[60]};
    assign in1352_2 = {pp19[38],pp13[45],pp7[52],pp1[59]};
    CLA_4 KS_1352(s1352, c1352, in1352_1, in1352_2);
    wire[3:0] s1353, in1353_1, in1353_2;
    wire c1353;
    assign in1353_1 = {pp20[37],pp14[44],pp8[51],pp2[58]};
    assign in1353_2 = {pp21[36],pp15[43],pp9[50],pp3[57]};
    CLA_4 KS_1353(s1353, c1353, in1353_1, in1353_2);
    wire[3:0] s1354, in1354_1, in1354_2;
    wire c1354;
    assign in1354_1 = {pp22[35],pp16[42],pp10[49],pp4[56]};
    assign in1354_2 = {pp23[34],pp17[41],pp11[48],pp5[55]};
    CLA_4 KS_1354(s1354, c1354, in1354_1, in1354_2);
    wire[3:0] s1355, in1355_1, in1355_2;
    wire c1355;
    assign in1355_1 = {pp24[33],pp18[40],pp12[47],pp6[54]};
    assign in1355_2 = {pp25[32],pp19[39],pp13[46],pp7[53]};
    CLA_4 KS_1355(s1355, c1355, in1355_1, in1355_2);
    wire[3:0] s1356, in1356_1, in1356_2;
    wire c1356;
    assign in1356_1 = {pp26[31],pp20[38],pp14[45],pp8[52]};
    assign in1356_2 = {pp27[30],pp21[37],pp15[44],pp9[51]};
    CLA_4 KS_1356(s1356, c1356, in1356_1, in1356_2);
    wire[3:0] s1357, in1357_1, in1357_2;
    wire c1357;
    assign in1357_1 = {pp28[29],pp22[36],pp16[43],pp10[50]};
    assign in1357_2 = {pp29[28],pp23[35],pp17[42],pp11[49]};
    CLA_4 KS_1357(s1357, c1357, in1357_1, in1357_2);
    wire[3:0] s1358, in1358_1, in1358_2;
    wire c1358;
    assign in1358_1 = {pp31[26],pp24[34],pp18[41],pp12[48]};
    assign in1358_2 = {pp32[25],pp25[33],pp19[40],pp13[47]};
    CLA_4_c KS_1358(s1358, c1358, in1358_1, in1358_2, pp30[27]);
    wire[3:0] s1359, in1359_1, in1359_2;
    wire c1359;
    assign in1359_1 = {pp26[32],pp20[39],pp14[46],pp0[61]};
    assign in1359_2 = {pp27[31],pp21[38],pp15[45],pp1[60]};
    CLA_4 KS_1359(s1359, c1359, in1359_1, in1359_2);
    wire[3:0] s1360, in1360_1, in1360_2;
    wire c1360;
    assign in1360_1 = {pp28[30],pp22[37],pp16[44],pp2[59]};
    assign in1360_2 = {pp29[29],pp23[36],pp17[43],pp3[58]};
    CLA_4 KS_1360(s1360, c1360, in1360_1, in1360_2);
    wire[3:0] s1361, in1361_1, in1361_2;
    wire c1361;
    assign in1361_1 = {pp31[27],pp24[35],pp18[42],pp4[57]};
    assign in1361_2 = {pp32[26],pp25[34],pp19[41],pp5[56]};
    CLA_4_c KS_1361(s1361, c1361, in1361_1, in1361_2, pp30[28]);
    wire[3:0] s1362, in1362_1, in1362_2;
    wire c1362;
    assign in1362_1 = {pp26[33],pp20[40],pp6[55],pp0[62]};
    assign in1362_2 = {pp27[32],pp21[39],pp7[54],pp1[61]};
    CLA_4 KS_1362(s1362, c1362, in1362_1, in1362_2);
    wire[3:0] s1363, in1363_1, in1363_2;
    wire c1363;
    assign in1363_1 = {pp28[31],pp22[38],pp8[53],pp2[60]};
    assign in1363_2 = {pp29[30],pp23[37],pp9[52],pp3[59]};
    CLA_4 KS_1363(s1363, c1363, in1363_1, in1363_2);
    wire[3:0] s1364, in1364_1, in1364_2;
    wire c1364;
    assign in1364_1 = {pp30[29],pp24[36],pp10[51],pp4[58]};
    assign in1364_2 = {pp31[28],pp25[35],pp11[50],pp5[57]};
    CLA_4 KS_1364(s1364, c1364, in1364_1, in1364_2);
    wire[3:0] s1365, in1365_1, in1365_2;
    wire c1365;
    assign in1365_1 = {pp33[26],pp26[34],pp12[49],pp6[56]};
    assign in1365_2 = {pp34[25],pp27[33],pp13[48],pp7[55]};
    CLA_4_c KS_1365(s1365, c1365, in1365_1, in1365_2, pp32[27]);
    wire[3:0] s1366, in1366_1, in1366_2;
    wire c1366;
    assign in1366_1 = {pp28[32],pp14[47],pp8[54],pp0[63]};
    assign in1366_2 = {pp29[31],pp15[46],pp9[53],pp1[62]};
    CLA_4 KS_1366(s1366, c1366, in1366_1, in1366_2);
    wire[3:0] s1367, in1367_1, in1367_2;
    wire c1367;
    assign in1367_1 = {pp30[30],pp16[45],pp10[52],pp2[61]};
    assign in1367_2 = {pp31[29],pp17[44],pp11[51],pp3[60]};
    CLA_4 KS_1367(s1367, c1367, in1367_1, in1367_2);
    wire[3:0] s1368, in1368_1, in1368_2;
    wire c1368;
    assign in1368_1 = {pp32[28],pp18[43],pp12[50],pp4[59]};
    assign in1368_2 = {pp33[27],pp19[42],pp13[49],pp5[58]};
    CLA_4 KS_1368(s1368, c1368, in1368_1, in1368_2);
    wire[3:0] s1369, in1369_1, in1369_2;
    wire c1369;
    assign in1369_1 = {pp35[25],pp20[41],pp14[48],pp6[57]};
    assign in1369_2 = {pp36[24],pp21[40],pp15[47],pp7[56]};
    CLA_4_c KS_1369(s1369, c1369, in1369_1, in1369_2, pp34[26]);
    wire[3:0] s1370, in1370_1, in1370_2;
    wire c1370;
    assign in1370_1 = {pp22[39],pp16[46],pp8[55],pp0[64]};
    assign in1370_2 = {pp23[38],pp17[45],pp9[54],pp1[63]};
    CLA_4 KS_1370(s1370, c1370, in1370_1, in1370_2);
    wire[3:0] s1371, in1371_1, in1371_2;
    wire c1371;
    assign in1371_1 = {pp24[37],pp18[44],pp10[53],pp2[62]};
    assign in1371_2 = {pp25[36],pp19[43],pp11[52],pp3[61]};
    CLA_4 KS_1371(s1371, c1371, in1371_1, in1371_2);
    wire[3:0] s1372, in1372_1, in1372_2;
    wire c1372;
    assign in1372_1 = {pp26[35],pp20[42],pp12[51],pp4[60]};
    assign in1372_2 = {pp27[34],pp21[41],pp13[50],pp5[59]};
    CLA_4 KS_1372(s1372, c1372, in1372_1, in1372_2);
    wire[3:0] s1373, in1373_1, in1373_2;
    wire c1373;
    assign in1373_1 = {pp28[33],pp22[40],pp14[49],pp6[58]};
    assign in1373_2 = {pp29[32],pp23[39],pp15[48],pp7[57]};
    CLA_4 KS_1373(s1373, c1373, in1373_1, in1373_2);
    wire[3:0] s1374, in1374_1, in1374_2;
    wire c1374;
    assign in1374_1 = {pp30[31],pp24[38],pp16[47],pp8[56]};
    assign in1374_2 = {pp31[30],pp25[37],pp17[46],pp9[55]};
    CLA_4 KS_1374(s1374, c1374, in1374_1, in1374_2);
    wire[3:0] s1375, in1375_1, in1375_2;
    wire c1375;
    assign in1375_1 = {pp32[29],pp26[36],pp18[45],pp10[54]};
    assign in1375_2 = {pp33[28],pp27[35],pp19[44],pp11[53]};
    CLA_4 KS_1375(s1375, c1375, in1375_1, in1375_2);
    wire[3:0] s1376, in1376_1, in1376_2;
    wire c1376;
    assign in1376_1 = {pp34[27],pp28[34],pp20[43],pp12[52]};
    assign in1376_2 = {pp35[26],pp29[33],pp21[42],pp13[51]};
    CLA_4 KS_1376(s1376, c1376, in1376_1, in1376_2);
    wire[3:0] s1377, in1377_1, in1377_2;
    wire c1377;
    assign in1377_1 = {pp36[25],pp30[32],pp22[41],pp14[50]};
    assign in1377_2 = {pp37[24],pp31[31],pp23[40],pp15[49]};
    CLA_4 KS_1377(s1377, c1377, in1377_1, in1377_2);
    wire[3:0] s1378, in1378_1, in1378_2;
    wire c1378;
    assign in1378_1 = {pp38[23],pp32[30],pp24[39],pp16[48]};
    assign in1378_2 = {pp39[22],pp33[29],pp25[38],pp17[47]};
    CLA_4 KS_1378(s1378, c1378, in1378_1, in1378_2);
    wire[3:0] s1379, in1379_1, in1379_2;
    wire c1379;
    assign in1379_1 = {pp40[21],pp34[28],pp26[37],pp18[46]};
    assign in1379_2 = {pp41[20],pp35[27],pp27[36],pp19[45]};
    CLA_4 KS_1379(s1379, c1379, in1379_1, in1379_2);
    wire[3:0] s1380, in1380_1, in1380_2;
    wire c1380;
    assign in1380_1 = {pp42[19],pp36[26],pp28[35],pp20[44]};
    assign in1380_2 = {pp43[18],pp37[25],pp29[34],pp21[43]};
    CLA_4 KS_1380(s1380, c1380, in1380_1, in1380_2);
    wire[3:0] s1381, in1381_1, in1381_2;
    wire c1381;
    assign in1381_1 = {pp45[16],pp38[24],pp30[33],pp22[42]};
    assign in1381_2 = {pp46[15],pp39[23],pp31[32],pp23[41]};
    CLA_4_c KS_1381(s1381, c1381, in1381_1, in1381_2, pp44[17]);
    wire[3:0] s1382, in1382_1, in1382_2;
    wire c1382;
    assign in1382_1 = {pp40[22],pp32[31],pp24[40],pp0[65]};
    assign in1382_2 = {pp41[21],pp33[30],pp25[39],pp1[64]};
    CLA_4 KS_1382(s1382, c1382, in1382_1, in1382_2);
    wire[3:0] s1383, in1383_1, in1383_2;
    wire c1383;
    assign in1383_1 = {pp34[29],pp26[38],pp2[63],pp0[66]};
    assign in1383_2 = {pp35[28],pp27[37],pp3[62],pp1[65]};
    CLA_4 KS_1383(s1383, c1383, in1383_1, in1383_2);
    wire[3:0] s1384, in1384_1, in1384_2;
    wire c1384;
    assign in1384_1 = {pp36[27],pp28[36],pp4[61],pp2[64]};
    assign in1384_2 = {pp37[26],pp29[35],pp5[60],pp3[63]};
    CLA_4 KS_1384(s1384, c1384, in1384_1, in1384_2);
    wire[3:0] s1385, in1385_1, in1385_2;
    wire c1385;
    assign in1385_1 = {pp38[25],pp30[34],pp6[59],pp4[62]};
    assign in1385_2 = {pp39[24],pp31[33],pp7[58],pp5[61]};
    CLA_4 KS_1385(s1385, c1385, in1385_1, in1385_2);
    wire[3:0] s1386, in1386_1, in1386_2;
    wire c1386;
    assign in1386_1 = {pp40[23],pp32[32],pp8[57],pp6[60]};
    assign in1386_2 = {pp41[22],pp33[31],pp9[56],pp7[59]};
    CLA_4 KS_1386(s1386, c1386, in1386_1, in1386_2);
    wire[3:0] s1387, in1387_1, in1387_2;
    wire c1387;
    assign in1387_1 = {pp43[20],pp34[30],pp10[55],pp8[58]};
    assign in1387_2 = {pp44[19],pp35[29],pp11[54],pp9[57]};
    CLA_4_c KS_1387(s1387, c1387, in1387_1, in1387_2, pp42[21]);
    wire[3:0] s1388, in1388_1, in1388_2;
    wire c1388;
    assign in1388_1 = {pp36[28],pp12[53],pp10[56],pp0[67]};
    assign in1388_2 = {pp37[27],pp13[52],pp11[55],pp1[66]};
    CLA_4 KS_1388(s1388, c1388, in1388_1, in1388_2);
    wire[3:0] s1389, in1389_1, in1389_2;
    wire c1389;
    assign in1389_1 = {pp38[26],pp14[51],pp12[54],pp2[65]};
    assign in1389_2 = {pp39[25],pp15[50],pp13[53],pp3[64]};
    CLA_4 KS_1389(s1389, c1389, in1389_1, in1389_2);
    wire[3:0] s1390, in1390_1, in1390_2;
    wire c1390;
    assign in1390_1 = {pp40[24],pp16[49],pp14[52],pp4[63]};
    assign in1390_2 = {pp41[23],pp17[48],pp15[51],pp5[62]};
    CLA_4 KS_1390(s1390, c1390, in1390_1, in1390_2);
    wire[3:0] s1391, in1391_1, in1391_2;
    wire c1391;
    assign in1391_1 = {pp42[22],pp18[47],pp16[50],pp6[61]};
    assign in1391_2 = {pp43[21],pp19[46],pp17[49],pp7[60]};
    CLA_4 KS_1391(s1391, c1391, in1391_1, in1391_2);
    wire[3:0] s1392, in1392_1, in1392_2;
    wire c1392;
    assign in1392_1 = {pp45[19],pp20[45],pp18[48],pp8[59]};
    assign in1392_2 = {pp46[18],pp21[44],pp19[47],pp9[58]};
    CLA_4_c KS_1392(s1392, c1392, in1392_1, in1392_2, pp44[20]);
    wire[3:0] s1393, in1393_1, in1393_2;
    wire c1393;
    assign in1393_1 = {pp22[43],pp20[46],pp10[57],pp0[68]};
    assign in1393_2 = {pp23[42],pp21[45],pp11[56],pp1[67]};
    CLA_4 KS_1393(s1393, c1393, in1393_1, in1393_2);
    wire[3:0] s1394, in1394_1, in1394_2;
    wire c1394;
    assign in1394_1 = {pp24[41],pp22[44],pp12[55],pp2[66]};
    assign in1394_2 = {pp25[40],pp23[43],pp13[54],pp3[65]};
    CLA_4 KS_1394(s1394, c1394, in1394_1, in1394_2);
    wire[3:0] s1395, in1395_1, in1395_2;
    wire c1395;
    assign in1395_1 = {pp26[39],pp24[42],pp14[53],pp4[64]};
    assign in1395_2 = {pp27[38],pp25[41],pp15[52],pp5[63]};
    CLA_4 KS_1395(s1395, c1395, in1395_1, in1395_2);
    wire[3:0] s1396, in1396_1, in1396_2;
    wire c1396;
    assign in1396_1 = {pp28[37],pp26[40],pp16[51],pp6[62]};
    assign in1396_2 = {pp29[36],pp27[39],pp17[50],pp7[61]};
    CLA_4 KS_1396(s1396, c1396, in1396_1, in1396_2);
    wire[3:0] s1397, in1397_1, in1397_2;
    wire c1397;
    assign in1397_1 = {pp30[35],pp28[38],pp18[49],pp8[60]};
    assign in1397_2 = {pp31[34],pp29[37],pp19[48],pp9[59]};
    CLA_4 KS_1397(s1397, c1397, in1397_1, in1397_2);
    wire[3:0] s1398, in1398_1, in1398_2;
    wire c1398;
    assign in1398_1 = {pp32[33],pp30[36],pp20[47],pp10[58]};
    assign in1398_2 = {pp33[32],pp31[35],pp21[46],pp11[57]};
    CLA_4 KS_1398(s1398, c1398, in1398_1, in1398_2);
    wire[3:0] s1399, in1399_1, in1399_2;
    wire c1399;
    assign in1399_1 = {pp34[31],pp32[34],pp22[45],pp12[56]};
    assign in1399_2 = {pp35[30],pp33[33],pp23[44],pp13[55]};
    CLA_4 KS_1399(s1399, c1399, in1399_1, in1399_2);
    wire[3:0] s1400, in1400_1, in1400_2;
    wire c1400;
    assign in1400_1 = {pp36[29],pp34[32],pp24[43],pp14[54]};
    assign in1400_2 = {pp37[28],pp35[31],pp25[42],pp15[53]};
    CLA_4 KS_1400(s1400, c1400, in1400_1, in1400_2);
    wire[3:0] s1401, in1401_1, in1401_2;
    wire c1401;
    assign in1401_1 = {pp38[27],pp36[30],pp26[41],pp16[52]};
    assign in1401_2 = {pp39[26],pp37[29],pp27[40],pp17[51]};
    CLA_4 KS_1401(s1401, c1401, in1401_1, in1401_2);
    wire[3:0] s1402, in1402_1, in1402_2;
    wire c1402;
    assign in1402_1 = {pp40[25],pp38[28],pp28[39],pp18[50]};
    assign in1402_2 = {pp41[24],pp39[27],pp29[38],pp19[49]};
    CLA_4 KS_1402(s1402, c1402, in1402_1, in1402_2);
    wire[3:0] s1403, in1403_1, in1403_2;
    wire c1403;
    assign in1403_1 = {pp42[23],pp40[26],pp30[37],pp20[48]};
    assign in1403_2 = {pp43[22],pp41[25],pp31[36],pp21[47]};
    CLA_4 KS_1403(s1403, c1403, in1403_1, in1403_2);
    wire[3:0] s1404, in1404_1, in1404_2;
    wire c1404;
    assign in1404_1 = {pp44[21],pp42[24],pp32[35],pp22[46]};
    assign in1404_2 = {pp45[20],pp43[23],pp33[34],pp23[45]};
    CLA_4 KS_1404(s1404, c1404, in1404_1, in1404_2);
    wire[3:0] s1405, in1405_1, in1405_2;
    wire c1405;
    assign in1405_1 = {pp46[19],pp44[22],pp34[33],pp24[44]};
    assign in1405_2 = {pp47[18],pp45[21],pp35[32],pp25[43]};
    CLA_4 KS_1405(s1405, c1405, in1405_1, in1405_2);
    wire[3:0] s1406, in1406_1, in1406_2;
    wire c1406;
    assign in1406_1 = {pp48[17],pp46[20],pp36[31],pp26[42]};
    assign in1406_2 = {pp49[16],pp47[19],pp37[30],pp27[41]};
    CLA_4 KS_1406(s1406, c1406, in1406_1, in1406_2);
    wire[0:0] s1407, in1407_1, in1407_2;
    wire c1407;
    assign in1407_1 = {pp50[15]};
    assign in1407_2 = {pp51[14]};
    Half_Adder KS_1407(s1407, c1407, in1407_1, in1407_2);
    wire[3:0] s1408, in1408_1, in1408_2;
    wire c1408;
    assign in1408_1 = {pp52[13],pp48[18],pp38[29],pp28[40]};
    assign in1408_2 = {pp53[12],pp49[17],pp39[28],pp29[39]};
    CLA_4 KS_1408(s1408, c1408, in1408_1, in1408_2);
    wire[0:0] s1409, in1409_1, in1409_2;
    wire c1409;
    assign in1409_1 = {pp54[11]};
    assign in1409_2 = {pp55[10]};
    Half_Adder KS_1409(s1409, c1409, in1409_1, in1409_2);
    wire[3:0] s1410, in1410_1, in1410_2;
    wire c1410;
    assign in1410_1 = {pp56[9],pp50[16],pp40[27],pp30[38]};
    assign in1410_2 = {pp57[8],pp51[15],pp41[26],pp31[37]};
    CLA_4 KS_1410(s1410, c1410, in1410_1, in1410_2);
    wire[0:0] s1411, in1411_1, in1411_2;
    wire c1411;
    assign in1411_1 = {pp58[7]};
    assign in1411_2 = {pp59[6]};
    Half_Adder KS_1411(s1411, c1411, in1411_1, in1411_2);
    wire[3:0] s1412, in1412_1, in1412_2;
    wire c1412;
    assign in1412_1 = {pp60[5],pp52[14],pp42[25],pp32[36]};
    assign in1412_2 = {pp61[4],pp53[13],pp43[24],pp33[35]};
    CLA_4 KS_1412(s1412, c1412, in1412_1, in1412_2);
    wire[0:0] s1413, in1413_1, in1413_2;
    wire c1413;
    assign in1413_1 = {pp63[2]};
    assign in1413_2 = {pp64[1]};
    Full_Adder KS_1413(s1413, c1413, in1413_1, in1413_2, pp62[3]);
    wire[3:0] s1414, in1414_1, in1414_2;
    wire c1414;
    assign in1414_1 = {pp44[23],pp34[34],pp0[69],pp0[70]};
    assign in1414_2 = {pp45[22],pp35[33],pp1[68],pp1[69]};
    CLA_4 KS_1414(s1414, c1414, in1414_1, in1414_2);
    wire[3:0] s1415, in1415_1, in1415_2;
    wire c1415;
    assign in1415_1 = {pp46[21],pp36[32],pp2[67],pp2[68]};
    assign in1415_2 = {pp47[20],pp37[31],pp3[66],pp3[67]};
    CLA_4 KS_1415(s1415, c1415, in1415_1, in1415_2);
    wire[3:0] s1416, in1416_1, in1416_2;
    wire c1416;
    assign in1416_1 = {pp48[19],pp38[30],pp4[65],pp4[66]};
    assign in1416_2 = {pp49[18],pp39[29],pp5[64],pp5[65]};
    CLA_4 KS_1416(s1416, c1416, in1416_1, in1416_2);
    wire[3:0] s1417, in1417_1, in1417_2;
    wire c1417;
    assign in1417_1 = {pp50[17],pp40[28],pp6[63],pp6[64]};
    assign in1417_2 = {pp51[16],pp41[27],pp7[62],pp7[63]};
    CLA_4 KS_1417(s1417, c1417, in1417_1, in1417_2);
    wire[3:0] s1418, in1418_1, in1418_2;
    wire c1418;
    assign in1418_1 = {pp53[14],pp42[26],pp8[61],pp8[62]};
    assign in1418_2 = {pp54[13],pp43[25],pp9[60],pp9[61]};
    CLA_4_c KS_1418(s1418, c1418, in1418_1, in1418_2, pp52[15]);
    wire[3:0] s1419, in1419_1, in1419_2;
    wire c1419;
    assign in1419_1 = {pp44[24],pp10[59],pp10[60],pp0[71]};
    assign in1419_2 = {pp45[23],pp11[58],pp11[59],pp1[70]};
    CLA_4 KS_1419(s1419, c1419, in1419_1, in1419_2);
    wire[3:0] s1420, in1420_1, in1420_2;
    wire c1420;
    assign in1420_1 = {pp46[22],pp12[57],pp12[58],pp2[69]};
    assign in1420_2 = {pp47[21],pp13[56],pp13[57],pp3[68]};
    CLA_4 KS_1420(s1420, c1420, in1420_1, in1420_2);
    wire[3:0] s1421, in1421_1, in1421_2;
    wire c1421;
    assign in1421_1 = {pp48[20],pp14[55],pp14[56],pp4[67]};
    assign in1421_2 = {pp49[19],pp15[54],pp15[55],pp5[66]};
    CLA_4 KS_1421(s1421, c1421, in1421_1, in1421_2);
    wire[3:0] s1422, in1422_1, in1422_2;
    wire c1422;
    assign in1422_1 = {pp50[18],pp16[53],pp16[54],pp6[65]};
    assign in1422_2 = {pp51[17],pp17[52],pp17[53],pp7[64]};
    CLA_4 KS_1422(s1422, c1422, in1422_1, in1422_2);
    wire[3:0] s1423, in1423_1, in1423_2;
    wire c1423;
    assign in1423_1 = {pp52[16],pp18[51],pp18[52],pp8[63]};
    assign in1423_2 = {pp53[15],pp19[50],pp19[51],pp9[62]};
    CLA_4 KS_1423(s1423, c1423, in1423_1, in1423_2);
    wire[3:0] s1424, in1424_1, in1424_2;
    wire c1424;
    assign in1424_1 = {pp55[13],pp20[49],pp20[50],pp10[61]};
    assign in1424_2 = {pp56[12],pp21[48],pp21[49],pp11[60]};
    CLA_4_c KS_1424(s1424, c1424, in1424_1, in1424_2, pp54[14]);
    wire[3:0] s1425, in1425_1, in1425_2;
    wire c1425;
    assign in1425_1 = {pp22[47],pp22[48],pp12[59],pp0[72]};
    assign in1425_2 = {pp23[46],pp23[47],pp13[58],pp1[71]};
    CLA_4 KS_1425(s1425, c1425, in1425_1, in1425_2);
    wire[3:0] s1426, in1426_1, in1426_2;
    wire c1426;
    assign in1426_1 = {pp24[45],pp24[46],pp14[57],pp2[70]};
    assign in1426_2 = {pp25[44],pp25[45],pp15[56],pp3[69]};
    CLA_4 KS_1426(s1426, c1426, in1426_1, in1426_2);
    wire[3:0] s1427, in1427_1, in1427_2;
    wire c1427;
    assign in1427_1 = {pp26[43],pp26[44],pp16[55],pp4[68]};
    assign in1427_2 = {pp27[42],pp27[43],pp17[54],pp5[67]};
    CLA_4 KS_1427(s1427, c1427, in1427_1, in1427_2);
    wire[3:0] s1428, in1428_1, in1428_2;
    wire c1428;
    assign in1428_1 = {pp28[41],pp28[42],pp18[53],pp6[66]};
    assign in1428_2 = {pp29[40],pp29[41],pp19[52],pp7[65]};
    CLA_4 KS_1428(s1428, c1428, in1428_1, in1428_2);
    wire[3:0] s1429, in1429_1, in1429_2;
    wire c1429;
    assign in1429_1 = {pp30[39],pp30[40],pp20[51],pp8[64]};
    assign in1429_2 = {pp31[38],pp31[39],pp21[50],pp9[63]};
    CLA_4 KS_1429(s1429, c1429, in1429_1, in1429_2);
    wire[3:0] s1430, in1430_1, in1430_2;
    wire c1430;
    assign in1430_1 = {pp32[37],pp32[38],pp22[49],pp10[62]};
    assign in1430_2 = {pp33[36],pp33[37],pp23[48],pp11[61]};
    CLA_4 KS_1430(s1430, c1430, in1430_1, in1430_2);
    wire[3:0] s1431, in1431_1, in1431_2;
    wire c1431;
    assign in1431_1 = {pp34[35],pp34[36],pp24[47],pp12[60]};
    assign in1431_2 = {pp35[34],pp35[35],pp25[46],pp13[59]};
    CLA_4 KS_1431(s1431, c1431, in1431_1, in1431_2);
    wire[3:0] s1432, in1432_1, in1432_2;
    wire c1432;
    assign in1432_1 = {pp36[33],pp36[34],pp26[45],pp14[58]};
    assign in1432_2 = {pp37[32],pp37[33],pp27[44],pp15[57]};
    CLA_4 KS_1432(s1432, c1432, in1432_1, in1432_2);
    wire[3:0] s1433, in1433_1, in1433_2;
    wire c1433;
    assign in1433_1 = {pp38[31],pp38[32],pp28[43],pp16[56]};
    assign in1433_2 = {pp39[30],pp39[31],pp29[42],pp17[55]};
    CLA_4 KS_1433(s1433, c1433, in1433_1, in1433_2);
    wire[3:0] s1434, in1434_1, in1434_2;
    wire c1434;
    assign in1434_1 = {pp40[29],pp40[30],pp30[41],pp18[54]};
    assign in1434_2 = {pp41[28],pp41[29],pp31[40],pp19[53]};
    CLA_4 KS_1434(s1434, c1434, in1434_1, in1434_2);
    wire[3:0] s1435, in1435_1, in1435_2;
    wire c1435;
    assign in1435_1 = {pp42[27],pp42[28],pp32[39],pp20[52]};
    assign in1435_2 = {pp43[26],pp43[27],pp33[38],pp21[51]};
    CLA_4 KS_1435(s1435, c1435, in1435_1, in1435_2);
    wire[3:0] s1436, in1436_1, in1436_2;
    wire c1436;
    assign in1436_1 = {pp44[25],pp44[26],pp34[37],pp22[50]};
    assign in1436_2 = {pp45[24],pp45[25],pp35[36],pp23[49]};
    CLA_4 KS_1436(s1436, c1436, in1436_1, in1436_2);
    wire[3:0] s1437, in1437_1, in1437_2;
    wire c1437;
    assign in1437_1 = {pp46[23],pp46[24],pp36[35],pp24[48]};
    assign in1437_2 = {pp47[22],pp47[23],pp37[34],pp25[47]};
    CLA_4 KS_1437(s1437, c1437, in1437_1, in1437_2);
    wire[3:0] s1438, in1438_1, in1438_2;
    wire c1438;
    assign in1438_1 = {pp48[21],pp48[22],pp38[33],pp26[46]};
    assign in1438_2 = {pp49[20],pp49[21],pp39[32],pp27[45]};
    CLA_4 KS_1438(s1438, c1438, in1438_1, in1438_2);
    wire[3:0] s1439, in1439_1, in1439_2;
    wire c1439;
    assign in1439_1 = {pp50[19],pp50[20],pp40[31],pp28[44]};
    assign in1439_2 = {pp51[18],pp51[19],pp41[30],pp29[43]};
    CLA_4 KS_1439(s1439, c1439, in1439_1, in1439_2);
    wire[3:0] s1440, in1440_1, in1440_2;
    wire c1440;
    assign in1440_1 = {pp52[17],pp52[18],pp42[29],pp30[42]};
    assign in1440_2 = {pp53[16],pp53[17],pp43[28],pp31[41]};
    CLA_4 KS_1440(s1440, c1440, in1440_1, in1440_2);
    wire[0:0] s1441, in1441_1, in1441_2;
    wire c1441;
    assign in1441_1 = {pp54[15]};
    assign in1441_2 = {pp55[14]};
    Half_Adder KS_1441(s1441, c1441, in1441_1, in1441_2);
    wire[3:0] s1442, in1442_1, in1442_2;
    wire c1442;
    assign in1442_1 = {pp56[13],pp54[16],pp44[27],pp32[40]};
    assign in1442_2 = {pp57[12],pp55[15],pp45[26],pp33[39]};
    CLA_4 KS_1442(s1442, c1442, in1442_1, in1442_2);
    wire[0:0] s1443, in1443_1, in1443_2;
    wire c1443;
    assign in1443_1 = {pp58[11]};
    assign in1443_2 = {pp59[10]};
    Half_Adder KS_1443(s1443, c1443, in1443_1, in1443_2);
    wire[3:0] s1444, in1444_1, in1444_2;
    wire c1444;
    assign in1444_1 = {pp60[9],pp56[14],pp46[25],pp34[38]};
    assign in1444_2 = {pp61[8],pp57[13],pp47[24],pp35[37]};
    CLA_4 KS_1444(s1444, c1444, in1444_1, in1444_2);
    wire[0:0] s1445, in1445_1, in1445_2;
    wire c1445;
    assign in1445_1 = {pp62[7]};
    assign in1445_2 = {pp63[6]};
    Half_Adder KS_1445(s1445, c1445, in1445_1, in1445_2);
    wire[3:0] s1446, in1446_1, in1446_2;
    wire c1446;
    assign in1446_1 = {pp64[5],pp58[12],pp48[23],pp36[36]};
    assign in1446_2 = {pp65[4],pp59[11],pp49[22],pp37[35]};
    CLA_4 KS_1446(s1446, c1446, in1446_1, in1446_2);
    wire[0:0] s1447, in1447_1, in1447_2;
    wire c1447;
    assign in1447_1 = {pp66[3]};
    assign in1447_2 = {pp67[2]};
    Half_Adder KS_1447(s1447, c1447, in1447_1, in1447_2);
    wire[3:0] s1448, in1448_1, in1448_2;
    wire c1448;
    assign in1448_1 = {pp68[1],pp60[10],pp50[21],pp38[34]};
    assign in1448_2 = {pp69[0],pp61[9],pp51[20],pp39[33]};
    CLA_4 KS_1448(s1448, c1448, in1448_1, in1448_2);
    wire[0:0] s1449, in1449_1, in1449_2;
    wire c1449;
    assign in1449_1 = {c1393};
    assign in1449_2 = {c1394};
    Half_Adder KS_1449(s1449, c1449, in1449_1, in1449_2);
    wire[3:0] s1450, in1450_1, in1450_2;
    wire c1450;
    assign in1450_1 = {c1395,pp62[8],pp52[19],pp40[32]};
    assign in1450_2 = {c1396,pp63[7],pp53[18],pp41[31]};
    CLA_4 KS_1450(s1450, c1450, in1450_1, in1450_2);
    wire[0:0] s1451, in1451_1, in1451_2;
    wire c1451;
    assign in1451_1 = {c1397};
    assign in1451_2 = {c1398};
    Half_Adder KS_1451(s1451, c1451, in1451_1, in1451_2);
    wire[3:0] s1452, in1452_1, in1452_2;
    wire c1452;
    assign in1452_1 = {c1399,pp64[6],pp54[17],pp42[30]};
    assign in1452_2 = {c1400,pp65[5],pp55[16],pp43[29]};
    CLA_4 KS_1452(s1452, c1452, in1452_1, in1452_2);
    wire[0:0] s1453, in1453_1, in1453_2;
    wire c1453;
    assign in1453_1 = {c1401};
    assign in1453_2 = {c1402};
    Half_Adder KS_1453(s1453, c1453, in1453_1, in1453_2);
    wire[3:0] s1454, in1454_1, in1454_2;
    wire c1454;
    assign in1454_1 = {c1404,pp66[4],pp56[15],pp44[28]};
    assign in1454_2 = {c1405,pp67[3],pp57[14],pp45[27]};
    CLA_4_c KS_1454(s1454, c1454, in1454_1, in1454_2, c1403);
    wire[3:0] s1455, in1455_1, in1455_2;
    wire c1455;
    assign in1455_1 = {pp58[13],pp46[26],pp0[73],pp0[74]};
    assign in1455_2 = {pp59[12],pp47[25],pp1[72],pp1[73]};
    CLA_4 KS_1455(s1455, c1455, in1455_1, in1455_2);
    wire[3:0] s1456, in1456_1, in1456_2;
    wire c1456;
    assign in1456_1 = {pp61[10],pp48[24],pp2[71],pp2[72]};
    assign in1456_2 = {pp62[9],pp49[23],pp3[70],pp3[71]};
    CLA_4_c KS_1456(s1456, c1456, in1456_1, in1456_2, pp60[11]);
    wire[3:0] s1457, in1457_1, in1457_2;
    wire c1457;
    assign in1457_1 = {pp50[22],pp4[69],pp4[70],pp0[75]};
    assign in1457_2 = {pp51[21],pp5[68],pp5[69],pp1[74]};
    CLA_4 KS_1457(s1457, c1457, in1457_1, in1457_2);
    wire[3:0] s1458, in1458_1, in1458_2;
    wire c1458;
    assign in1458_1 = {pp52[20],pp6[67],pp6[68],pp2[73]};
    assign in1458_2 = {pp53[19],pp7[66],pp7[67],pp3[72]};
    CLA_4 KS_1458(s1458, c1458, in1458_1, in1458_2);
    wire[3:0] s1459, in1459_1, in1459_2;
    wire c1459;
    assign in1459_1 = {pp54[18],pp8[65],pp8[66],pp4[71]};
    assign in1459_2 = {pp55[17],pp9[64],pp9[65],pp5[70]};
    CLA_4 KS_1459(s1459, c1459, in1459_1, in1459_2);
    wire[3:0] s1460, in1460_1, in1460_2;
    wire c1460;
    assign in1460_1 = {pp56[16],pp10[63],pp10[64],pp6[69]};
    assign in1460_2 = {pp57[15],pp11[62],pp11[63],pp7[68]};
    CLA_4 KS_1460(s1460, c1460, in1460_1, in1460_2);
    wire[3:0] s1461, in1461_1, in1461_2;
    wire c1461;
    assign in1461_1 = {pp58[14],pp12[61],pp12[62],pp8[67]};
    assign in1461_2 = {pp59[13],pp13[60],pp13[61],pp9[66]};
    CLA_4 KS_1461(s1461, c1461, in1461_1, in1461_2);
    wire[3:0] s1462, in1462_1, in1462_2;
    wire c1462;
    assign in1462_1 = {pp60[12],pp14[59],pp14[60],pp10[65]};
    assign in1462_2 = {pp61[11],pp15[58],pp15[59],pp11[64]};
    CLA_4 KS_1462(s1462, c1462, in1462_1, in1462_2);
    wire[3:0] s1463, in1463_1, in1463_2;
    wire c1463;
    assign in1463_1 = {pp62[10],pp16[57],pp16[58],pp12[63]};
    assign in1463_2 = {pp63[9],pp17[56],pp17[57],pp13[62]};
    CLA_4 KS_1463(s1463, c1463, in1463_1, in1463_2);
    wire[3:0] s1464, in1464_1, in1464_2;
    wire c1464;
    assign in1464_1 = {pp65[7],pp18[55],pp18[56],pp14[61]};
    assign in1464_2 = {pp66[6],pp19[54],pp19[55],pp15[60]};
    CLA_4_c KS_1464(s1464, c1464, in1464_1, in1464_2, pp64[8]);
    wire[3:0] s1465, in1465_1, in1465_2;
    wire c1465;
    assign in1465_1 = {pp20[53],pp20[54],pp16[59],pp2[74]};
    assign in1465_2 = {pp21[52],pp21[53],pp17[58],pp3[73]};
    CLA_4 KS_1465(s1465, c1465, in1465_1, in1465_2);
    wire[3:0] s1466, in1466_1, in1466_2;
    wire c1466;
    assign in1466_1 = {pp22[51],pp22[52],pp18[57],pp4[72]};
    assign in1466_2 = {pp23[50],pp23[51],pp19[56],pp5[71]};
    CLA_4 KS_1466(s1466, c1466, in1466_1, in1466_2);
    wire[3:0] s1467, in1467_1, in1467_2;
    wire c1467;
    assign in1467_1 = {pp24[49],pp24[50],pp20[55],pp6[70]};
    assign in1467_2 = {pp25[48],pp25[49],pp21[54],pp7[69]};
    CLA_4 KS_1467(s1467, c1467, in1467_1, in1467_2);
    wire[3:0] s1468, in1468_1, in1468_2;
    wire c1468;
    assign in1468_1 = {pp26[47],pp26[48],pp22[53],pp8[68]};
    assign in1468_2 = {pp27[46],pp27[47],pp23[52],pp9[67]};
    CLA_4 KS_1468(s1468, c1468, in1468_1, in1468_2);
    wire[3:0] s1469, in1469_1, in1469_2;
    wire c1469;
    assign in1469_1 = {pp28[45],pp28[46],pp24[51],pp10[66]};
    assign in1469_2 = {pp29[44],pp29[45],pp25[50],pp11[65]};
    CLA_4 KS_1469(s1469, c1469, in1469_1, in1469_2);
    wire[3:0] s1470, in1470_1, in1470_2;
    wire c1470;
    assign in1470_1 = {pp30[43],pp30[44],pp26[49],pp12[64]};
    assign in1470_2 = {pp31[42],pp31[43],pp27[48],pp13[63]};
    CLA_4 KS_1470(s1470, c1470, in1470_1, in1470_2);
    wire[3:0] s1471, in1471_1, in1471_2;
    wire c1471;
    assign in1471_1 = {pp32[41],pp32[42],pp28[47],pp14[62]};
    assign in1471_2 = {pp33[40],pp33[41],pp29[46],pp15[61]};
    CLA_4 KS_1471(s1471, c1471, in1471_1, in1471_2);
    wire[3:0] s1472, in1472_1, in1472_2;
    wire c1472;
    assign in1472_1 = {pp34[39],pp34[40],pp30[45],pp16[60]};
    assign in1472_2 = {pp35[38],pp35[39],pp31[44],pp17[59]};
    CLA_4 KS_1472(s1472, c1472, in1472_1, in1472_2);
    wire[3:0] s1473, in1473_1, in1473_2;
    wire c1473;
    assign in1473_1 = {pp36[37],pp36[38],pp32[43],pp18[58]};
    assign in1473_2 = {pp37[36],pp37[37],pp33[42],pp19[57]};
    CLA_4 KS_1473(s1473, c1473, in1473_1, in1473_2);
    wire[3:0] s1474, in1474_1, in1474_2;
    wire c1474;
    assign in1474_1 = {pp38[35],pp38[36],pp34[41],pp20[56]};
    assign in1474_2 = {pp39[34],pp39[35],pp35[40],pp21[55]};
    CLA_4 KS_1474(s1474, c1474, in1474_1, in1474_2);
    wire[3:0] s1475, in1475_1, in1475_2;
    wire c1475;
    assign in1475_1 = {pp40[33],pp40[34],pp36[39],pp22[54]};
    assign in1475_2 = {pp41[32],pp41[33],pp37[38],pp23[53]};
    CLA_4 KS_1475(s1475, c1475, in1475_1, in1475_2);
    wire[3:0] s1476, in1476_1, in1476_2;
    wire c1476;
    assign in1476_1 = {pp42[31],pp42[32],pp38[37],pp24[52]};
    assign in1476_2 = {pp43[30],pp43[31],pp39[36],pp25[51]};
    CLA_4 KS_1476(s1476, c1476, in1476_1, in1476_2);
    wire[3:0] s1477, in1477_1, in1477_2;
    wire c1477;
    assign in1477_1 = {pp44[29],pp44[30],pp40[35],pp26[50]};
    assign in1477_2 = {pp45[28],pp45[29],pp41[34],pp27[49]};
    CLA_4 KS_1477(s1477, c1477, in1477_1, in1477_2);
    wire[3:0] s1478, in1478_1, in1478_2;
    wire c1478;
    assign in1478_1 = {pp46[27],pp46[28],pp42[33],pp28[48]};
    assign in1478_2 = {pp47[26],pp47[27],pp43[32],pp29[47]};
    CLA_4 KS_1478(s1478, c1478, in1478_1, in1478_2);
    wire[3:0] s1479, in1479_1, in1479_2;
    wire c1479;
    assign in1479_1 = {pp48[25],pp48[26],pp44[31],pp30[46]};
    assign in1479_2 = {pp49[24],pp49[25],pp45[30],pp31[45]};
    CLA_4 KS_1479(s1479, c1479, in1479_1, in1479_2);
    wire[3:0] s1480, in1480_1, in1480_2;
    wire c1480;
    assign in1480_1 = {pp50[23],pp50[24],pp46[29],pp32[44]};
    assign in1480_2 = {pp51[22],pp51[23],pp47[28],pp33[43]};
    CLA_4 KS_1480(s1480, c1480, in1480_1, in1480_2);
    wire[3:0] s1481, in1481_1, in1481_2;
    wire c1481;
    assign in1481_1 = {pp52[21],pp52[22],pp48[27],pp34[42]};
    assign in1481_2 = {pp53[20],pp53[21],pp49[26],pp35[41]};
    CLA_4 KS_1481(s1481, c1481, in1481_1, in1481_2);
    wire[3:0] s1482, in1482_1, in1482_2;
    wire c1482;
    assign in1482_1 = {pp54[19],pp54[20],pp50[25],pp36[40]};
    assign in1482_2 = {pp55[18],pp55[19],pp51[24],pp37[39]};
    CLA_4 KS_1482(s1482, c1482, in1482_1, in1482_2);
    wire[3:0] s1483, in1483_1, in1483_2;
    wire c1483;
    assign in1483_1 = {pp56[17],pp56[18],pp52[23],pp38[38]};
    assign in1483_2 = {pp57[16],pp57[17],pp53[22],pp39[37]};
    CLA_4 KS_1483(s1483, c1483, in1483_1, in1483_2);
    wire[3:0] s1484, in1484_1, in1484_2;
    wire c1484;
    assign in1484_1 = {pp58[15],pp58[16],pp54[21],pp40[36]};
    assign in1484_2 = {pp59[14],pp59[15],pp55[20],pp41[35]};
    CLA_4 KS_1484(s1484, c1484, in1484_1, in1484_2);
    wire[3:0] s1485, in1485_1, in1485_2;
    wire c1485;
    assign in1485_1 = {pp60[13],pp60[14],pp56[19],pp42[34]};
    assign in1485_2 = {pp61[12],pp61[13],pp57[18],pp43[33]};
    CLA_4 KS_1485(s1485, c1485, in1485_1, in1485_2);
    wire[0:0] s1486, in1486_1, in1486_2;
    wire c1486;
    assign in1486_1 = {pp62[11]};
    assign in1486_2 = {pp63[10]};
    Half_Adder KS_1486(s1486, c1486, in1486_1, in1486_2);
    wire[3:0] s1487, in1487_1, in1487_2;
    wire c1487;
    assign in1487_1 = {pp64[9],pp62[12],pp58[17],pp44[32]};
    assign in1487_2 = {pp65[8],pp63[11],pp59[16],pp45[31]};
    CLA_4 KS_1487(s1487, c1487, in1487_1, in1487_2);
    wire[0:0] s1488, in1488_1, in1488_2;
    wire c1488;
    assign in1488_1 = {pp66[7]};
    assign in1488_2 = {pp67[6]};
    Half_Adder KS_1488(s1488, c1488, in1488_1, in1488_2);
    wire[3:0] s1489, in1489_1, in1489_2;
    wire c1489;
    assign in1489_1 = {pp68[5],pp64[10],pp60[15],pp46[30]};
    assign in1489_2 = {pp69[4],pp65[9],pp61[14],pp47[29]};
    CLA_4 KS_1489(s1489, c1489, in1489_1, in1489_2);
    wire[0:0] s1490, in1490_1, in1490_2;
    wire c1490;
    assign in1490_1 = {pp70[3]};
    assign in1490_2 = {pp71[2]};
    Half_Adder KS_1490(s1490, c1490, in1490_1, in1490_2);
    wire[3:0] s1491, in1491_1, in1491_2;
    wire c1491;
    assign in1491_1 = {pp72[1],pp66[8],pp62[13],pp48[28]};
    assign in1491_2 = {pp73[0],pp67[7],pp63[12],pp49[27]};
    CLA_4 KS_1491(s1491, c1491, in1491_1, in1491_2);
    wire[0:0] s1492, in1492_1, in1492_2;
    wire c1492;
    assign in1492_1 = {c1425};
    assign in1492_2 = {c1426};
    Half_Adder KS_1492(s1492, c1492, in1492_1, in1492_2);
    wire[3:0] s1493, in1493_1, in1493_2;
    wire c1493;
    assign in1493_1 = {c1427,pp68[6],pp64[11],pp50[26]};
    assign in1493_2 = {c1428,pp69[5],pp65[10],pp51[25]};
    CLA_4 KS_1493(s1493, c1493, in1493_1, in1493_2);
    wire[0:0] s1494, in1494_1, in1494_2;
    wire c1494;
    assign in1494_1 = {c1429};
    assign in1494_2 = {c1430};
    Half_Adder KS_1494(s1494, c1494, in1494_1, in1494_2);
    wire[3:0] s1495, in1495_1, in1495_2;
    wire c1495;
    assign in1495_1 = {c1431,pp70[4],pp66[9],pp52[24]};
    assign in1495_2 = {c1432,pp71[3],pp67[8],pp53[23]};
    CLA_4 KS_1495(s1495, c1495, in1495_1, in1495_2);
    wire[0:0] s1496, in1496_1, in1496_2;
    wire c1496;
    assign in1496_1 = {c1433};
    assign in1496_2 = {c1434};
    Half_Adder KS_1496(s1496, c1496, in1496_1, in1496_2);
    wire[1:0] s1497, in1497_1, in1497_2;
    wire c1497;
    assign in1497_1 = {c1435,pp72[2]};
    assign in1497_2 = {c1436,pp73[1]};
    CLA_2 KS_1497(s1497, c1497, in1497_1, in1497_2);
    wire[0:0] s1498, in1498_1, in1498_2;
    wire c1498;
    assign in1498_1 = {c1437};
    assign in1498_2 = {c1438};
    Half_Adder KS_1498(s1498, c1498, in1498_1, in1498_2);
    wire[3:0] s1499, in1499_1, in1499_2;
    wire c1499;
    assign in1499_1 = {c1439,pp74[0],pp68[7],pp54[22]};
    assign in1499_2 = {c1440,s1455[3],pp69[6],pp55[21]};
    CLA_4 KS_1499(s1499, c1499, in1499_1, in1499_2);
    wire[0:0] s1500, in1500_1, in1500_2;
    wire c1500;
    assign in1500_1 = {c1442};
    assign in1500_2 = {c1444};
    Half_Adder KS_1500(s1500, c1500, in1500_1, in1500_2);
    wire[1:0] s1501, in1501_1, in1501_2;
    wire c1501;
    assign in1501_1 = {c1446,s1456[3]};
    assign in1501_2 = {c1448,s1457[2]};
    CLA_2 KS_1501(s1501, c1501, in1501_1, in1501_2);
    wire[0:0] s1502, in1502_1, in1502_2;
    wire c1502;
    assign in1502_1 = {c1450};
    assign in1502_2 = {c1452};
    Half_Adder KS_1502(s1502, c1502, in1502_1, in1502_2);
    wire[3:0] s1503, in1503_1, in1503_2;
    wire c1503;
    assign in1503_1 = {c1454,s1458[2],pp70[5],pp56[20]};
    assign in1503_2 = {s1455[2],s1459[2],pp71[4],pp57[19]};
    CLA_4 KS_1503(s1503, c1503, in1503_1, in1503_2);
    wire[0:0] s1504, in1504_1, in1504_2;
    wire c1504;
    assign in1504_1 = {s1456[2]};
    assign in1504_2 = {s1457[1]};
    Half_Adder KS_1504(s1504, c1504, in1504_1, in1504_2);
    wire[1:0] s1505, in1505_1, in1505_2;
    wire c1505;
    assign in1505_1 = {s1459[1],s1460[2]};
    assign in1505_2 = {s1460[1],s1461[2]};
    CLA_2_c KS_1505(s1505, c1505, in1505_1, in1505_2, s1458[1]);
    wire[3:0] s1506, in1506_1, in1506_2;
    wire c1506;
    assign in1506_1 = {pp58[18],pp4[73],pp6[72],pp8[71]};
    assign in1506_2 = {pp59[17],pp5[72],pp7[71],pp9[70]};
    CLA_4 KS_1506(s1506, c1506, in1506_1, in1506_2);
    wire[3:0] s1507, in1507_1, in1507_2;
    wire c1507;
    assign in1507_1 = {pp60[16],pp6[71],pp8[70],pp10[69]};
    assign in1507_2 = {pp61[15],pp7[70],pp9[69],pp11[68]};
    CLA_4 KS_1507(s1507, c1507, in1507_1, in1507_2);
    wire[3:0] s1508, in1508_1, in1508_2;
    wire c1508;
    assign in1508_1 = {pp62[14],pp8[69],pp10[68],pp12[67]};
    assign in1508_2 = {pp63[13],pp9[68],pp11[67],pp13[66]};
    CLA_4 KS_1508(s1508, c1508, in1508_1, in1508_2);
    wire[3:0] s1509, in1509_1, in1509_2;
    wire c1509;
    assign in1509_1 = {pp64[12],pp10[67],pp12[66],pp14[65]};
    assign in1509_2 = {pp65[11],pp11[66],pp13[65],pp15[64]};
    CLA_4 KS_1509(s1509, c1509, in1509_1, in1509_2);
    wire[3:0] s1510, in1510_1, in1510_2;
    wire c1510;
    assign in1510_1 = {pp66[10],pp12[65],pp14[64],pp16[63]};
    assign in1510_2 = {pp67[9],pp13[64],pp15[63],pp17[62]};
    CLA_4 KS_1510(s1510, c1510, in1510_1, in1510_2);
    wire[3:0] s1511, in1511_1, in1511_2;
    wire c1511;
    assign in1511_1 = {pp68[8],pp14[63],pp16[62],pp18[61]};
    assign in1511_2 = {pp69[7],pp15[62],pp17[61],pp19[60]};
    CLA_4 KS_1511(s1511, c1511, in1511_1, in1511_2);
    wire[3:0] s1512, in1512_1, in1512_2;
    wire c1512;
    assign in1512_1 = {pp70[6],pp16[61],pp18[60],pp20[59]};
    assign in1512_2 = {pp71[5],pp17[60],pp19[59],pp21[58]};
    CLA_4 KS_1512(s1512, c1512, in1512_1, in1512_2);
    wire[3:0] s1513, in1513_1, in1513_2;
    wire c1513;
    assign in1513_1 = {pp72[4],pp18[59],pp20[58],pp22[57]};
    assign in1513_2 = {pp73[3],pp19[58],pp21[57],pp23[56]};
    CLA_4 KS_1513(s1513, c1513, in1513_1, in1513_2);
    wire[3:0] s1514, in1514_1, in1514_2;
    wire c1514;
    assign in1514_1 = {pp74[2],pp20[57],pp22[56],pp24[55]};
    assign in1514_2 = {pp75[1],pp21[56],pp23[55],pp25[54]};
    CLA_4 KS_1514(s1514, c1514, in1514_1, in1514_2);
    wire[3:0] s1515, in1515_1, in1515_2;
    wire c1515;
    assign in1515_1 = {s1[0],pp22[55],pp24[54],pp26[53]};
    assign in1515_2 = {c1457,pp23[54],pp25[53],pp27[52]};
    CLA_4_c KS_1515(s1515, c1515, in1515_1, in1515_2, pp76[0]);
    wire[3:0] s1516, in1516_1, in1516_2;
    wire c1516;
    assign in1516_1 = {pp24[53],pp26[52],pp28[51],pp11[69]};
    assign in1516_2 = {pp25[52],pp27[51],pp29[50],pp12[68]};
    CLA_4 KS_1516(s1516, c1516, in1516_1, in1516_2);
    wire[3:0] s1517, in1517_1, in1517_2;
    wire c1517;
    assign in1517_1 = {pp26[51],pp28[50],pp30[49],pp13[67]};
    assign in1517_2 = {pp27[50],pp29[49],pp31[48],pp14[66]};
    CLA_4 KS_1517(s1517, c1517, in1517_1, in1517_2);
    wire[3:0] s1518, in1518_1, in1518_2;
    wire c1518;
    assign in1518_1 = {pp28[49],pp30[48],pp32[47],pp15[65]};
    assign in1518_2 = {pp29[48],pp31[47],pp33[46],pp16[64]};
    CLA_4 KS_1518(s1518, c1518, in1518_1, in1518_2);
    wire[3:0] s1519, in1519_1, in1519_2;
    wire c1519;
    assign in1519_1 = {pp30[47],pp32[46],pp34[45],pp17[63]};
    assign in1519_2 = {pp31[46],pp33[45],pp35[44],pp18[62]};
    CLA_4 KS_1519(s1519, c1519, in1519_1, in1519_2);
    wire[3:0] s1520, in1520_1, in1520_2;
    wire c1520;
    assign in1520_1 = {pp32[45],pp34[44],pp36[43],pp19[61]};
    assign in1520_2 = {pp33[44],pp35[43],pp37[42],pp20[60]};
    CLA_4 KS_1520(s1520, c1520, in1520_1, in1520_2);
    wire[3:0] s1521, in1521_1, in1521_2;
    wire c1521;
    assign in1521_1 = {pp34[43],pp36[42],pp38[41],pp21[59]};
    assign in1521_2 = {pp35[42],pp37[41],pp39[40],pp22[58]};
    CLA_4 KS_1521(s1521, c1521, in1521_1, in1521_2);
    wire[3:0] s1522, in1522_1, in1522_2;
    wire c1522;
    assign in1522_1 = {pp36[41],pp38[40],pp40[39],pp23[57]};
    assign in1522_2 = {pp37[40],pp39[39],pp41[38],pp24[56]};
    CLA_4 KS_1522(s1522, c1522, in1522_1, in1522_2);
    wire[3:0] s1523, in1523_1, in1523_2;
    wire c1523;
    assign in1523_1 = {pp38[39],pp40[38],pp42[37],pp25[55]};
    assign in1523_2 = {pp39[38],pp41[37],pp43[36],pp26[54]};
    CLA_4 KS_1523(s1523, c1523, in1523_1, in1523_2);
    wire[3:0] s1524, in1524_1, in1524_2;
    wire c1524;
    assign in1524_1 = {pp40[37],pp42[36],pp44[35],pp27[53]};
    assign in1524_2 = {pp41[36],pp43[35],pp45[34],pp28[52]};
    CLA_4 KS_1524(s1524, c1524, in1524_1, in1524_2);
    wire[3:0] s1525, in1525_1, in1525_2;
    wire c1525;
    assign in1525_1 = {pp42[35],pp44[34],pp46[33],pp29[51]};
    assign in1525_2 = {pp43[34],pp45[33],pp47[32],pp30[50]};
    CLA_4 KS_1525(s1525, c1525, in1525_1, in1525_2);
    wire[3:0] s1526, in1526_1, in1526_2;
    wire c1526;
    assign in1526_1 = {pp44[33],pp46[32],pp48[31],pp31[49]};
    assign in1526_2 = {pp45[32],pp47[31],pp49[30],pp32[48]};
    CLA_4 KS_1526(s1526, c1526, in1526_1, in1526_2);
    wire[3:0] s1527, in1527_1, in1527_2;
    wire c1527;
    assign in1527_1 = {pp46[31],pp48[30],pp50[29],pp33[47]};
    assign in1527_2 = {pp47[30],pp49[29],pp51[28],pp34[46]};
    CLA_4 KS_1527(s1527, c1527, in1527_1, in1527_2);
    wire[3:0] s1528, in1528_1, in1528_2;
    wire c1528;
    assign in1528_1 = {pp48[29],pp50[28],pp52[27],pp35[45]};
    assign in1528_2 = {pp49[28],pp51[27],pp53[26],pp36[44]};
    CLA_4 KS_1528(s1528, c1528, in1528_1, in1528_2);
    wire[3:0] s1529, in1529_1, in1529_2;
    wire c1529;
    assign in1529_1 = {pp50[27],pp52[26],pp54[25],pp37[43]};
    assign in1529_2 = {pp51[26],pp53[25],pp55[24],pp38[42]};
    CLA_4 KS_1529(s1529, c1529, in1529_1, in1529_2);
    wire[3:0] s1530, in1530_1, in1530_2;
    wire c1530;
    assign in1530_1 = {pp52[25],pp54[24],pp56[23],pp39[41]};
    assign in1530_2 = {pp53[24],pp55[23],pp57[22],pp40[40]};
    CLA_4 KS_1530(s1530, c1530, in1530_1, in1530_2);
    wire[3:0] s1531, in1531_1, in1531_2;
    wire c1531;
    assign in1531_1 = {pp54[23],pp56[22],pp58[21],pp41[39]};
    assign in1531_2 = {pp55[22],pp57[21],pp59[20],pp42[38]};
    CLA_4 KS_1531(s1531, c1531, in1531_1, in1531_2);
    wire[3:0] s1532, in1532_1, in1532_2;
    wire c1532;
    assign in1532_1 = {pp56[21],pp58[20],pp60[19],pp43[37]};
    assign in1532_2 = {pp57[20],pp59[19],pp61[18],pp44[36]};
    CLA_4 KS_1532(s1532, c1532, in1532_1, in1532_2);
    wire[3:0] s1533, in1533_1, in1533_2;
    wire c1533;
    assign in1533_1 = {pp58[19],pp60[18],pp62[17],pp45[35]};
    assign in1533_2 = {pp59[18],pp61[17],pp63[16],pp46[34]};
    CLA_4 KS_1533(s1533, c1533, in1533_1, in1533_2);
    wire[3:0] s1534, in1534_1, in1534_2;
    wire c1534;
    assign in1534_1 = {pp60[17],pp62[16],pp64[15],pp47[33]};
    assign in1534_2 = {pp61[16],pp63[15],pp65[14],pp48[32]};
    CLA_4 KS_1534(s1534, c1534, in1534_1, in1534_2);
    wire[3:0] s1535, in1535_1, in1535_2;
    wire c1535;
    assign in1535_1 = {pp62[15],pp64[14],pp66[13],pp49[31]};
    assign in1535_2 = {pp63[14],pp65[13],pp67[12],pp50[30]};
    CLA_4 KS_1535(s1535, c1535, in1535_1, in1535_2);
    wire[3:0] s1536, in1536_1, in1536_2;
    wire c1536;
    assign in1536_1 = {pp64[13],pp66[12],pp68[11],pp51[29]};
    assign in1536_2 = {pp65[12],pp67[11],pp69[10],pp52[28]};
    CLA_4 KS_1536(s1536, c1536, in1536_1, in1536_2);
    wire[3:0] s1537, in1537_1, in1537_2;
    wire c1537;
    assign in1537_1 = {pp66[11],pp68[10],pp70[9],pp53[27]};
    assign in1537_2 = {pp67[10],pp69[9],pp71[8],pp54[26]};
    CLA_4 KS_1537(s1537, c1537, in1537_1, in1537_2);
    wire[0:0] s1538, in1538_1, in1538_2;
    wire c1538;
    assign in1538_1 = {pp68[9]};
    assign in1538_2 = {pp69[8]};
    Half_Adder KS_1538(s1538, c1538, in1538_1, in1538_2);
    wire[1:0] s1539, in1539_1, in1539_2;
    wire c1539;
    assign in1539_1 = {pp70[7],pp70[8]};
    assign in1539_2 = {pp71[6],pp71[7]};
    CLA_2 KS_1539(s1539, c1539, in1539_1, in1539_2);
    wire[0:0] s1540, in1540_1, in1540_2;
    wire c1540;
    assign in1540_1 = {pp72[5]};
    assign in1540_2 = {pp73[4]};
    Half_Adder KS_1540(s1540, c1540, in1540_1, in1540_2);
    wire[3:0] s1541, in1541_1, in1541_2;
    wire c1541;
    assign in1541_1 = {pp74[3],pp72[6],pp72[7],pp55[25]};
    assign in1541_2 = {pp75[2],pp73[5],pp73[6],pp56[24]};
    CLA_4 KS_1541(s1541, c1541, in1541_1, in1541_2);
    wire[0:0] s1542, in1542_1, in1542_2;
    wire c1542;
    assign in1542_1 = {pp76[1]};
    assign in1542_2 = {pp77[0]};
    Half_Adder KS_1542(s1542, c1542, in1542_1, in1542_2);
    wire[1:0] s1543, in1543_1, in1543_2;
    wire c1543;
    assign in1543_1 = {s1[1],pp74[4]};
    assign in1543_2 = {s2[0],pp75[3]};
    CLA_2 KS_1543(s1543, c1543, in1543_1, in1543_2);
    wire[0:0] s1544, in1544_1, in1544_2;
    wire c1544;
    assign in1544_1 = {c1465};
    assign in1544_2 = {c1466};
    Half_Adder KS_1544(s1544, c1544, in1544_1, in1544_2);
    wire[3:0] s1545, in1545_1, in1545_2;
    wire c1545;
    assign in1545_1 = {c1467,pp76[2],pp74[5],pp57[23]};
    assign in1545_2 = {c1468,pp77[1],pp75[4],pp58[22]};
    CLA_4 KS_1545(s1545, c1545, in1545_1, in1545_2);
    wire[0:0] s1546, in1546_1, in1546_2;
    wire c1546;
    assign in1546_1 = {c1469};
    assign in1546_2 = {c1470};
    Half_Adder KS_1546(s1546, c1546, in1546_1, in1546_2);
    wire[1:0] s1547, in1547_1, in1547_2;
    wire c1547;
    assign in1547_1 = {c1471,pp78[0]};
    assign in1547_2 = {c1472,s1[2]};
    CLA_2 KS_1547(s1547, c1547, in1547_1, in1547_2);
    wire[0:0] s1548, in1548_1, in1548_2;
    wire c1548;
    assign in1548_1 = {c1473};
    assign in1548_2 = {c1474};
    Half_Adder KS_1548(s1548, c1548, in1548_1, in1548_2);
    wire[3:0] s1549, in1549_1, in1549_2;
    wire c1549;
    assign in1549_1 = {c1475,s2[1],pp76[3],pp59[21]};
    assign in1549_2 = {c1476,s3[0],pp77[2],pp60[20]};
    CLA_4 KS_1549(s1549, c1549, in1549_1, in1549_2);
    wire[0:0] s1550, in1550_1, in1550_2;
    wire c1550;
    assign in1550_1 = {c1477};
    assign in1550_2 = {c1478};
    Half_Adder KS_1550(s1550, c1550, in1550_1, in1550_2);
    wire[1:0] s1551, in1551_1, in1551_2;
    wire c1551;
    assign in1551_1 = {c1479,s1506[2]};
    assign in1551_2 = {c1480,s1507[2]};
    CLA_2 KS_1551(s1551, c1551, in1551_1, in1551_2);
    wire[0:0] s1552, in1552_1, in1552_2;
    wire c1552;
    assign in1552_1 = {c1481};
    assign in1552_2 = {c1482};
    Half_Adder KS_1552(s1552, c1552, in1552_1, in1552_2);
    wire[3:0] s1553, in1553_1, in1553_2;
    wire c1553;
    assign in1553_1 = {c1483,s1508[2],pp78[1],pp61[19]};
    assign in1553_2 = {c1484,s1509[2],pp79[0],pp62[18]};
    CLA_4 KS_1553(s1553, c1553, in1553_1, in1553_2);
    wire[0:0] s1554, in1554_1, in1554_2;
    wire c1554;
    assign in1554_1 = {c1485};
    assign in1554_2 = {c1487};
    Half_Adder KS_1554(s1554, c1554, in1554_1, in1554_2);
    wire[1:0] s1555, in1555_1, in1555_2;
    wire c1555;
    assign in1555_1 = {c1489,s1510[2]};
    assign in1555_2 = {c1491,s1511[2]};
    CLA_2 KS_1555(s1555, c1555, in1555_1, in1555_2);
    wire[0:0] s1556, in1556_1, in1556_2;
    wire c1556;
    assign in1556_1 = {c1493};
    assign in1556_2 = {c1495};
    Half_Adder KS_1556(s1556, c1556, in1556_1, in1556_2);
    wire[3:0] s1557, in1557_1, in1557_2;
    wire c1557;
    assign in1557_1 = {c1499,s1512[2],s1[3],pp63[17]};
    assign in1557_2 = {c1503,s1513[2],s2[2],pp64[16]};
    CLA_4 KS_1557(s1557, c1557, in1557_1, in1557_2);
    wire[0:0] s1558, in1558_1, in1558_2;
    wire c1558;
    assign in1558_1 = {s1506[1]};
    assign in1558_2 = {s1507[1]};
    Half_Adder KS_1558(s1558, c1558, in1558_1, in1558_2);
    wire[1:0] s1559, in1559_1, in1559_2;
    wire c1559;
    assign in1559_1 = {s1508[1],s1514[2]};
    assign in1559_2 = {s1509[1],s1515[2]};
    CLA_2 KS_1559(s1559, c1559, in1559_1, in1559_2);
    wire[0:0] s1560, in1560_1, in1560_2;
    wire c1560;
    assign in1560_1 = {s1510[1]};
    assign in1560_2 = {s1511[1]};
    Half_Adder KS_1560(s1560, c1560, in1560_1, in1560_2);
    wire[3:0] s1561, in1561_1, in1561_2;
    wire c1561;
    assign in1561_1 = {s1512[1],s1516[1],s3[1],pp65[15]};
    assign in1561_2 = {s1513[1],s1517[1],s4[0],pp66[14]};
    CLA_4 KS_1561(s1561, c1561, in1561_1, in1561_2);
    wire[0:0] s1562, in1562_1, in1562_2;
    wire c1562;
    assign in1562_1 = {s1514[1]};
    assign in1562_2 = {s1515[1]};
    Half_Adder KS_1562(s1562, c1562, in1562_1, in1562_2);
    wire[1:0] s1563, in1563_1, in1563_2;
    wire c1563;
    assign in1563_1 = {s1517[0],s1518[1]};
    assign in1563_2 = {s1518[0],s1519[1]};
    CLA_2_c KS_1563(s1563, c1563, in1563_1, in1563_2, s1516[0]);
    wire[3:0] s1564, in1564_1, in1564_2;
    wire c1564;
    assign in1564_1 = {pp67[13],pp13[68],pp15[67],pp17[66]};
    assign in1564_2 = {pp68[12],pp14[67],pp16[66],pp18[65]};
    CLA_4 KS_1564(s1564, c1564, in1564_1, in1564_2);
    wire[3:0] s1565, in1565_1, in1565_2;
    wire c1565;
    assign in1565_1 = {pp69[11],pp15[66],pp17[65],pp19[64]};
    assign in1565_2 = {pp70[10],pp16[65],pp18[64],pp20[63]};
    CLA_4 KS_1565(s1565, c1565, in1565_1, in1565_2);
    wire[3:0] s1566, in1566_1, in1566_2;
    wire c1566;
    assign in1566_1 = {pp71[9],pp17[64],pp19[63],pp21[62]};
    assign in1566_2 = {pp72[8],pp18[63],pp20[62],pp22[61]};
    CLA_4 KS_1566(s1566, c1566, in1566_1, in1566_2);
    wire[3:0] s1567, in1567_1, in1567_2;
    wire c1567;
    assign in1567_1 = {pp73[7],pp19[62],pp21[61],pp23[60]};
    assign in1567_2 = {pp74[6],pp20[61],pp22[60],pp24[59]};
    CLA_4 KS_1567(s1567, c1567, in1567_1, in1567_2);
    wire[3:0] s1568, in1568_1, in1568_2;
    wire c1568;
    assign in1568_1 = {pp75[5],pp21[60],pp23[59],pp25[58]};
    assign in1568_2 = {pp76[4],pp22[59],pp24[58],pp26[57]};
    CLA_4 KS_1568(s1568, c1568, in1568_1, in1568_2);
    wire[3:0] s1569, in1569_1, in1569_2;
    wire c1569;
    assign in1569_1 = {pp77[3],pp23[58],pp25[57],pp27[56]};
    assign in1569_2 = {pp78[2],pp24[57],pp26[56],pp28[55]};
    CLA_4 KS_1569(s1569, c1569, in1569_1, in1569_2);
    wire[3:0] s1570, in1570_1, in1570_2;
    wire c1570;
    assign in1570_1 = {pp79[1],pp25[56],pp27[55],pp29[54]};
    assign in1570_2 = {pp80[0],pp26[55],pp28[54],pp30[53]};
    CLA_4 KS_1570(s1570, c1570, in1570_1, in1570_2);
    wire[3:0] s1571, in1571_1, in1571_2;
    wire c1571;
    assign in1571_1 = {c1,pp27[54],pp29[53],pp31[52]};
    assign in1571_2 = {s2[3],pp28[53],pp30[52],pp32[51]};
    CLA_4 KS_1571(s1571, c1571, in1571_1, in1571_2);
    wire[3:0] s1572, in1572_1, in1572_2;
    wire c1572;
    assign in1572_1 = {s3[2],pp29[52],pp31[51],pp33[50]};
    assign in1572_2 = {s4[1],pp30[51],pp32[50],pp34[49]};
    CLA_4 KS_1572(s1572, c1572, in1572_1, in1572_2);
    wire[3:0] s1573, in1573_1, in1573_2;
    wire c1573;
    assign in1573_1 = {s5[0],pp31[50],pp33[49],pp35[48]};
    assign in1573_2 = {s6[0],pp32[49],pp34[48],pp36[47]};
    CLA_4 KS_1573(s1573, c1573, in1573_1, in1573_2);
    wire[3:0] s1574, in1574_1, in1574_2;
    wire c1574;
    assign in1574_1 = {c1506,pp33[48],pp35[47],pp37[46]};
    assign in1574_2 = {c1507,pp34[47],pp36[46],pp38[45]};
    CLA_4 KS_1574(s1574, c1574, in1574_1, in1574_2);
    wire[3:0] s1575, in1575_1, in1575_2;
    wire c1575;
    assign in1575_1 = {c1509,pp35[46],pp37[45],pp39[44]};
    assign in1575_2 = {c1510,pp36[45],pp38[44],pp40[43]};
    CLA_4_c KS_1575(s1575, c1575, in1575_1, in1575_2, c1508);
    wire[3:0] s1576, in1576_1, in1576_2;
    wire c1576;
    assign in1576_1 = {pp37[44],pp39[43],pp41[42],pp21[63]};
    assign in1576_2 = {pp38[43],pp40[42],pp42[41],pp22[62]};
    CLA_4 KS_1576(s1576, c1576, in1576_1, in1576_2);
    wire[3:0] s1577, in1577_1, in1577_2;
    wire c1577;
    assign in1577_1 = {pp39[42],pp41[41],pp43[40],pp23[61]};
    assign in1577_2 = {pp40[41],pp42[40],pp44[39],pp24[60]};
    CLA_4 KS_1577(s1577, c1577, in1577_1, in1577_2);
    wire[3:0] s1578, in1578_1, in1578_2;
    wire c1578;
    assign in1578_1 = {pp41[40],pp43[39],pp45[38],pp25[59]};
    assign in1578_2 = {pp42[39],pp44[38],pp46[37],pp26[58]};
    CLA_4 KS_1578(s1578, c1578, in1578_1, in1578_2);
    wire[3:0] s1579, in1579_1, in1579_2;
    wire c1579;
    assign in1579_1 = {pp43[38],pp45[37],pp47[36],pp27[57]};
    assign in1579_2 = {pp44[37],pp46[36],pp48[35],pp28[56]};
    CLA_4 KS_1579(s1579, c1579, in1579_1, in1579_2);
    wire[3:0] s1580, in1580_1, in1580_2;
    wire c1580;
    assign in1580_1 = {pp45[36],pp47[35],pp49[34],pp29[55]};
    assign in1580_2 = {pp46[35],pp48[34],pp50[33],pp30[54]};
    CLA_4 KS_1580(s1580, c1580, in1580_1, in1580_2);
    wire[3:0] s1581, in1581_1, in1581_2;
    wire c1581;
    assign in1581_1 = {pp47[34],pp49[33],pp51[32],pp31[53]};
    assign in1581_2 = {pp48[33],pp50[32],pp52[31],pp32[52]};
    CLA_4 KS_1581(s1581, c1581, in1581_1, in1581_2);
    wire[3:0] s1582, in1582_1, in1582_2;
    wire c1582;
    assign in1582_1 = {pp49[32],pp51[31],pp53[30],pp33[51]};
    assign in1582_2 = {pp50[31],pp52[30],pp54[29],pp34[50]};
    CLA_4 KS_1582(s1582, c1582, in1582_1, in1582_2);
    wire[3:0] s1583, in1583_1, in1583_2;
    wire c1583;
    assign in1583_1 = {pp51[30],pp53[29],pp55[28],pp35[49]};
    assign in1583_2 = {pp52[29],pp54[28],pp56[27],pp36[48]};
    CLA_4 KS_1583(s1583, c1583, in1583_1, in1583_2);
    wire[3:0] s1584, in1584_1, in1584_2;
    wire c1584;
    assign in1584_1 = {pp53[28],pp55[27],pp57[26],pp37[47]};
    assign in1584_2 = {pp54[27],pp56[26],pp58[25],pp38[46]};
    CLA_4 KS_1584(s1584, c1584, in1584_1, in1584_2);
    wire[3:0] s1585, in1585_1, in1585_2;
    wire c1585;
    assign in1585_1 = {pp55[26],pp57[25],pp59[24],pp39[45]};
    assign in1585_2 = {pp56[25],pp58[24],pp60[23],pp40[44]};
    CLA_4 KS_1585(s1585, c1585, in1585_1, in1585_2);
    wire[3:0] s1586, in1586_1, in1586_2;
    wire c1586;
    assign in1586_1 = {pp57[24],pp59[23],pp61[22],pp41[43]};
    assign in1586_2 = {pp58[23],pp60[22],pp62[21],pp42[42]};
    CLA_4 KS_1586(s1586, c1586, in1586_1, in1586_2);
    wire[3:0] s1587, in1587_1, in1587_2;
    wire c1587;
    assign in1587_1 = {pp59[22],pp61[21],pp63[20],pp43[41]};
    assign in1587_2 = {pp60[21],pp62[20],pp64[19],pp44[40]};
    CLA_4 KS_1587(s1587, c1587, in1587_1, in1587_2);
    wire[3:0] s1588, in1588_1, in1588_2;
    wire c1588;
    assign in1588_1 = {pp61[20],pp63[19],pp65[18],pp45[39]};
    assign in1588_2 = {pp62[19],pp64[18],pp66[17],pp46[38]};
    CLA_4 KS_1588(s1588, c1588, in1588_1, in1588_2);
    wire[3:0] s1589, in1589_1, in1589_2;
    wire c1589;
    assign in1589_1 = {pp63[18],pp65[17],pp67[16],pp47[37]};
    assign in1589_2 = {pp64[17],pp66[16],pp68[15],pp48[36]};
    CLA_4 KS_1589(s1589, c1589, in1589_1, in1589_2);
    wire[3:0] s1590, in1590_1, in1590_2;
    wire c1590;
    assign in1590_1 = {pp65[16],pp67[15],pp69[14],pp49[35]};
    assign in1590_2 = {pp66[15],pp68[14],pp70[13],pp50[34]};
    CLA_4 KS_1590(s1590, c1590, in1590_1, in1590_2);
    wire[3:0] s1591, in1591_1, in1591_2;
    wire c1591;
    assign in1591_1 = {pp67[14],pp69[13],pp71[12],pp51[33]};
    assign in1591_2 = {pp68[13],pp70[12],pp72[11],pp52[32]};
    CLA_4 KS_1591(s1591, c1591, in1591_1, in1591_2);
    wire[3:0] s1592, in1592_1, in1592_2;
    wire c1592;
    assign in1592_1 = {pp69[12],pp71[11],pp73[10],pp53[31]};
    assign in1592_2 = {pp70[11],pp72[10],pp74[9],pp54[30]};
    CLA_4 KS_1592(s1592, c1592, in1592_1, in1592_2);
    wire[3:0] s1593, in1593_1, in1593_2;
    wire c1593;
    assign in1593_1 = {pp71[10],pp73[9],pp75[8],pp55[29]};
    assign in1593_2 = {pp72[9],pp74[8],pp76[7],pp56[28]};
    CLA_4 KS_1593(s1593, c1593, in1593_1, in1593_2);
    wire[3:0] s1594, in1594_1, in1594_2;
    wire c1594;
    assign in1594_1 = {pp73[8],pp75[7],pp77[6],pp57[27]};
    assign in1594_2 = {pp74[7],pp76[6],pp78[5],pp58[26]};
    CLA_4 KS_1594(s1594, c1594, in1594_1, in1594_2);
    wire[3:0] s1595, in1595_1, in1595_2;
    wire c1595;
    assign in1595_1 = {pp75[6],pp77[5],pp79[4],pp59[25]};
    assign in1595_2 = {pp76[5],pp78[4],pp80[3],pp60[24]};
    CLA_4 KS_1595(s1595, c1595, in1595_1, in1595_2);
    wire[0:0] s1596, in1596_1, in1596_2;
    wire c1596;
    assign in1596_1 = {pp77[4]};
    assign in1596_2 = {pp78[3]};
    Half_Adder KS_1596(s1596, c1596, in1596_1, in1596_2);
    wire[1:0] s1597, in1597_1, in1597_2;
    wire c1597;
    assign in1597_1 = {pp79[2],pp79[3]};
    assign in1597_2 = {pp80[1],pp80[2]};
    CLA_2 KS_1597(s1597, c1597, in1597_1, in1597_2);
    wire[0:0] s1598, in1598_1, in1598_2;
    wire c1598;
    assign in1598_1 = {pp81[0]};
    assign in1598_2 = {c2};
    Half_Adder KS_1598(s1598, c1598, in1598_1, in1598_2);
    wire[3:0] s1599, in1599_1, in1599_2;
    wire c1599;
    assign in1599_1 = {s3[3],pp81[1],pp81[2],pp61[23]};
    assign in1599_2 = {s4[2],pp82[0],pp82[1],pp62[22]};
    CLA_4 KS_1599(s1599, c1599, in1599_1, in1599_2);
    wire[0:0] s1600, in1600_1, in1600_2;
    wire c1600;
    assign in1600_1 = {s5[1]};
    assign in1600_2 = {s6[1]};
    Half_Adder KS_1600(s1600, c1600, in1600_1, in1600_2);
    wire[1:0] s1601, in1601_1, in1601_2;
    wire c1601;
    assign in1601_1 = {s7[0],c3};
    assign in1601_2 = {s8[0],s4[3]};
    CLA_2 KS_1601(s1601, c1601, in1601_1, in1601_2);
    wire[0:0] s1602, in1602_1, in1602_2;
    wire c1602;
    assign in1602_1 = {c1516};
    assign in1602_2 = {c1517};
    Half_Adder KS_1602(s1602, c1602, in1602_1, in1602_2);
    wire[3:0] s1603, in1603_1, in1603_2;
    wire c1603;
    assign in1603_1 = {c1518,s5[2],pp83[0],pp63[21]};
    assign in1603_2 = {c1519,s6[2],c4,pp64[20]};
    CLA_4 KS_1603(s1603, c1603, in1603_1, in1603_2);
    wire[0:0] s1604, in1604_1, in1604_2;
    wire c1604;
    assign in1604_1 = {c1520};
    assign in1604_2 = {c1521};
    Half_Adder KS_1604(s1604, c1604, in1604_1, in1604_2);
    wire[1:0] s1605, in1605_1, in1605_2;
    wire c1605;
    assign in1605_1 = {c1522,s7[1]};
    assign in1605_2 = {c1523,s8[1]};
    CLA_2 KS_1605(s1605, c1605, in1605_1, in1605_2);
    wire[0:0] s1606, in1606_1, in1606_2;
    wire c1606;
    assign in1606_1 = {c1524};
    assign in1606_2 = {c1525};
    Half_Adder KS_1606(s1606, c1606, in1606_1, in1606_2);
    wire[3:0] s1607, in1607_1, in1607_2;
    wire c1607;
    assign in1607_1 = {c1526,s9[0],s5[3],pp65[19]};
    assign in1607_2 = {c1527,s10[0],s6[3],pp66[18]};
    CLA_4 KS_1607(s1607, c1607, in1607_1, in1607_2);
    wire[0:0] s1608, in1608_1, in1608_2;
    wire c1608;
    assign in1608_1 = {c1528};
    assign in1608_2 = {c1529};
    Half_Adder KS_1608(s1608, c1608, in1608_1, in1608_2);
    wire[1:0] s1609, in1609_1, in1609_2;
    wire c1609;
    assign in1609_1 = {c1530,s1564[2]};
    assign in1609_2 = {c1531,s1565[2]};
    CLA_2 KS_1609(s1609, c1609, in1609_1, in1609_2);
    wire[0:0] s1610, in1610_1, in1610_2;
    wire c1610;
    assign in1610_1 = {c1532};
    assign in1610_2 = {c1533};
    Half_Adder KS_1610(s1610, c1610, in1610_1, in1610_2);
    wire[3:0] s1611, in1611_1, in1611_2;
    wire c1611;
    assign in1611_1 = {c1534,s1566[2],s7[2],pp67[17]};
    assign in1611_2 = {c1535,s1567[2],s8[2],pp68[16]};
    CLA_4 KS_1611(s1611, c1611, in1611_1, in1611_2);
    wire[0:0] s1612, in1612_1, in1612_2;
    wire c1612;
    assign in1612_1 = {c1536};
    assign in1612_2 = {c1537};
    Half_Adder KS_1612(s1612, c1612, in1612_1, in1612_2);
    wire[1:0] s1613, in1613_1, in1613_2;
    wire c1613;
    assign in1613_1 = {c1541,s1568[2]};
    assign in1613_2 = {c1545,s1569[2]};
    CLA_2 KS_1613(s1613, c1613, in1613_1, in1613_2);
    wire[0:0] s1614, in1614_1, in1614_2;
    wire c1614;
    assign in1614_1 = {c1549};
    assign in1614_2 = {c1553};
    Half_Adder KS_1614(s1614, c1614, in1614_1, in1614_2);
    wire[3:0] s1615, in1615_1, in1615_2;
    wire c1615;
    assign in1615_1 = {c1557,s1570[2],s9[1],pp69[15]};
    assign in1615_2 = {c1561,s1571[2],s10[1],pp70[14]};
    CLA_4 KS_1615(s1615, c1615, in1615_1, in1615_2);
    wire[0:0] s1616, in1616_1, in1616_2;
    wire c1616;
    assign in1616_1 = {s1564[1]};
    assign in1616_2 = {s1565[1]};
    Half_Adder KS_1616(s1616, c1616, in1616_1, in1616_2);
    wire[1:0] s1617, in1617_1, in1617_2;
    wire c1617;
    assign in1617_1 = {s1566[1],s1572[2]};
    assign in1617_2 = {s1567[1],s1573[2]};
    CLA_2 KS_1617(s1617, c1617, in1617_1, in1617_2);
    wire[0:0] s1618, in1618_1, in1618_2;
    wire c1618;
    assign in1618_1 = {s1568[1]};
    assign in1618_2 = {s1569[1]};
    Half_Adder KS_1618(s1618, c1618, in1618_1, in1618_2);
    wire[3:0] s1619, in1619_1, in1619_2;
    wire c1619;
    assign in1619_1 = {s1570[1],s1574[2],s11[0],pp71[13]};
    assign in1619_2 = {s1571[1],s1575[2],s12[0],pp72[12]};
    CLA_4 KS_1619(s1619, c1619, in1619_1, in1619_2);
    wire[0:0] s1620, in1620_1, in1620_2;
    wire c1620;
    assign in1620_1 = {s1572[1]};
    assign in1620_2 = {s1573[1]};
    Half_Adder KS_1620(s1620, c1620, in1620_1, in1620_2);
    wire[1:0] s1621, in1621_1, in1621_2;
    wire c1621;
    assign in1621_1 = {s1575[1],s1576[1]};
    assign in1621_2 = {s1576[0],s1577[1]};
    CLA_2_c KS_1621(s1621, c1621, in1621_1, in1621_2, s1574[1]);
    wire[3:0] s1622, in1622_1, in1622_2;
    wire c1622;
    assign in1622_1 = {pp73[11],pp23[62],pp25[61],pp27[60]};
    assign in1622_2 = {pp74[10],pp24[61],pp26[60],pp28[59]};
    CLA_4 KS_1622(s1622, c1622, in1622_1, in1622_2);
    wire[3:0] s1623, in1623_1, in1623_2;
    wire c1623;
    assign in1623_1 = {pp75[9],pp25[60],pp27[59],pp29[58]};
    assign in1623_2 = {pp76[8],pp26[59],pp28[58],pp30[57]};
    CLA_4 KS_1623(s1623, c1623, in1623_1, in1623_2);
    wire[3:0] s1624, in1624_1, in1624_2;
    wire c1624;
    assign in1624_1 = {pp77[7],pp27[58],pp29[57],pp31[56]};
    assign in1624_2 = {pp78[6],pp28[57],pp30[56],pp32[55]};
    CLA_4 KS_1624(s1624, c1624, in1624_1, in1624_2);
    wire[3:0] s1625, in1625_1, in1625_2;
    wire c1625;
    assign in1625_1 = {pp79[5],pp29[56],pp31[55],pp33[54]};
    assign in1625_2 = {pp80[4],pp30[55],pp32[54],pp34[53]};
    CLA_4 KS_1625(s1625, c1625, in1625_1, in1625_2);
    wire[3:0] s1626, in1626_1, in1626_2;
    wire c1626;
    assign in1626_1 = {pp81[3],pp31[54],pp33[53],pp35[52]};
    assign in1626_2 = {pp82[2],pp32[53],pp34[52],pp36[51]};
    CLA_4 KS_1626(s1626, c1626, in1626_1, in1626_2);
    wire[3:0] s1627, in1627_1, in1627_2;
    wire c1627;
    assign in1627_1 = {pp83[1],pp33[52],pp35[51],pp37[50]};
    assign in1627_2 = {pp84[0],pp34[51],pp36[50],pp38[49]};
    CLA_4 KS_1627(s1627, c1627, in1627_1, in1627_2);
    wire[3:0] s1628, in1628_1, in1628_2;
    wire c1628;
    assign in1628_1 = {c5,pp35[50],pp37[49],pp39[48]};
    assign in1628_2 = {c6,pp36[49],pp38[48],pp40[47]};
    CLA_4 KS_1628(s1628, c1628, in1628_1, in1628_2);
    wire[3:0] s1629, in1629_1, in1629_2;
    wire c1629;
    assign in1629_1 = {s7[3],pp37[48],pp39[47],pp41[46]};
    assign in1629_2 = {s8[3],pp38[47],pp40[46],pp42[45]};
    CLA_4 KS_1629(s1629, c1629, in1629_1, in1629_2);
    wire[3:0] s1630, in1630_1, in1630_2;
    wire c1630;
    assign in1630_1 = {s9[2],pp39[46],pp41[45],pp43[44]};
    assign in1630_2 = {s10[2],pp40[45],pp42[44],pp44[43]};
    CLA_4 KS_1630(s1630, c1630, in1630_1, in1630_2);
    wire[3:0] s1631, in1631_1, in1631_2;
    wire c1631;
    assign in1631_1 = {s11[1],pp41[44],pp43[43],pp45[42]};
    assign in1631_2 = {s12[1],pp42[43],pp44[42],pp46[41]};
    CLA_4 KS_1631(s1631, c1631, in1631_1, in1631_2);
    wire[3:0] s1632, in1632_1, in1632_2;
    wire c1632;
    assign in1632_1 = {s13[0],pp43[42],pp45[41],pp47[40]};
    assign in1632_2 = {s14[0],pp44[41],pp46[40],pp48[39]};
    CLA_4 KS_1632(s1632, c1632, in1632_1, in1632_2);
    wire[3:0] s1633, in1633_1, in1633_2;
    wire c1633;
    assign in1633_1 = {s15[0],pp45[40],pp47[39],pp49[38]};
    assign in1633_2 = {s16[0],pp46[39],pp48[38],pp50[37]};
    CLA_4 KS_1633(s1633, c1633, in1633_1, in1633_2);
    wire[3:0] s1634, in1634_1, in1634_2;
    wire c1634;
    assign in1634_1 = {c1564,pp47[38],pp49[37],pp51[36]};
    assign in1634_2 = {c1565,pp48[37],pp50[36],pp52[35]};
    CLA_4 KS_1634(s1634, c1634, in1634_1, in1634_2);
    wire[3:0] s1635, in1635_1, in1635_2;
    wire c1635;
    assign in1635_1 = {c1566,pp49[36],pp51[35],pp53[34]};
    assign in1635_2 = {c1567,pp50[35],pp52[34],pp54[33]};
    CLA_4 KS_1635(s1635, c1635, in1635_1, in1635_2);
    wire[3:0] s1636, in1636_1, in1636_2;
    wire c1636;
    assign in1636_1 = {c1568,pp51[34],pp53[33],pp55[32]};
    assign in1636_2 = {c1569,pp52[33],pp54[32],pp56[31]};
    CLA_4 KS_1636(s1636, c1636, in1636_1, in1636_2);
    wire[3:0] s1637, in1637_1, in1637_2;
    wire c1637;
    assign in1637_1 = {c1571,pp53[32],pp55[31],pp57[30]};
    assign in1637_2 = {c1572,pp54[31],pp56[30],pp58[29]};
    CLA_4_c KS_1637(s1637, c1637, in1637_1, in1637_2, c1570);
    wire[3:0] s1638, in1638_1, in1638_2;
    wire c1638;
    assign in1638_1 = {pp55[30],pp57[29],pp59[28],pp33[55]};
    assign in1638_2 = {pp56[29],pp58[28],pp60[27],pp34[54]};
    CLA_4 KS_1638(s1638, c1638, in1638_1, in1638_2);
    wire[3:0] s1639, in1639_1, in1639_2;
    wire c1639;
    assign in1639_1 = {pp57[28],pp59[27],pp61[26],pp35[53]};
    assign in1639_2 = {pp58[27],pp60[26],pp62[25],pp36[52]};
    CLA_4 KS_1639(s1639, c1639, in1639_1, in1639_2);
    wire[3:0] s1640, in1640_1, in1640_2;
    wire c1640;
    assign in1640_1 = {pp59[26],pp61[25],pp63[24],pp37[51]};
    assign in1640_2 = {pp60[25],pp62[24],pp64[23],pp38[50]};
    CLA_4 KS_1640(s1640, c1640, in1640_1, in1640_2);
    wire[3:0] s1641, in1641_1, in1641_2;
    wire c1641;
    assign in1641_1 = {pp61[24],pp63[23],pp65[22],pp39[49]};
    assign in1641_2 = {pp62[23],pp64[22],pp66[21],pp40[48]};
    CLA_4 KS_1641(s1641, c1641, in1641_1, in1641_2);
    wire[3:0] s1642, in1642_1, in1642_2;
    wire c1642;
    assign in1642_1 = {pp63[22],pp65[21],pp67[20],pp41[47]};
    assign in1642_2 = {pp64[21],pp66[20],pp68[19],pp42[46]};
    CLA_4 KS_1642(s1642, c1642, in1642_1, in1642_2);
    wire[3:0] s1643, in1643_1, in1643_2;
    wire c1643;
    assign in1643_1 = {pp65[20],pp67[19],pp69[18],pp43[45]};
    assign in1643_2 = {pp66[19],pp68[18],pp70[17],pp44[44]};
    CLA_4 KS_1643(s1643, c1643, in1643_1, in1643_2);
    wire[3:0] s1644, in1644_1, in1644_2;
    wire c1644;
    assign in1644_1 = {pp67[18],pp69[17],pp71[16],pp45[43]};
    assign in1644_2 = {pp68[17],pp70[16],pp72[15],pp46[42]};
    CLA_4 KS_1644(s1644, c1644, in1644_1, in1644_2);
    wire[3:0] s1645, in1645_1, in1645_2;
    wire c1645;
    assign in1645_1 = {pp69[16],pp71[15],pp73[14],pp47[41]};
    assign in1645_2 = {pp70[15],pp72[14],pp74[13],pp48[40]};
    CLA_4 KS_1645(s1645, c1645, in1645_1, in1645_2);
    wire[3:0] s1646, in1646_1, in1646_2;
    wire c1646;
    assign in1646_1 = {pp71[14],pp73[13],pp75[12],pp49[39]};
    assign in1646_2 = {pp72[13],pp74[12],pp76[11],pp50[38]};
    CLA_4 KS_1646(s1646, c1646, in1646_1, in1646_2);
    wire[3:0] s1647, in1647_1, in1647_2;
    wire c1647;
    assign in1647_1 = {pp73[12],pp75[11],pp77[10],pp51[37]};
    assign in1647_2 = {pp74[11],pp76[10],pp78[9],pp52[36]};
    CLA_4 KS_1647(s1647, c1647, in1647_1, in1647_2);
    wire[3:0] s1648, in1648_1, in1648_2;
    wire c1648;
    assign in1648_1 = {pp75[10],pp77[9],pp79[8],pp53[35]};
    assign in1648_2 = {pp76[9],pp78[8],pp80[7],pp54[34]};
    CLA_4 KS_1648(s1648, c1648, in1648_1, in1648_2);
    wire[3:0] s1649, in1649_1, in1649_2;
    wire c1649;
    assign in1649_1 = {pp77[8],pp79[7],pp81[6],pp55[33]};
    assign in1649_2 = {pp78[7],pp80[6],pp82[5],pp56[32]};
    CLA_4 KS_1649(s1649, c1649, in1649_1, in1649_2);
    wire[3:0] s1650, in1650_1, in1650_2;
    wire c1650;
    assign in1650_1 = {pp79[6],pp81[5],pp83[4],pp57[31]};
    assign in1650_2 = {pp80[5],pp82[4],pp84[3],pp58[30]};
    CLA_4 KS_1650(s1650, c1650, in1650_1, in1650_2);
    wire[3:0] s1651, in1651_1, in1651_2;
    wire c1651;
    assign in1651_1 = {pp81[4],pp83[3],pp85[2],pp59[29]};
    assign in1651_2 = {pp82[3],pp84[2],pp86[1],pp60[28]};
    CLA_4 KS_1651(s1651, c1651, in1651_1, in1651_2);
    wire[3:0] s1652, in1652_1, in1652_2;
    wire c1652;
    assign in1652_1 = {pp83[2],pp85[1],pp87[0],pp61[27]};
    assign in1652_2 = {pp84[1],pp86[0],c11,pp62[26]};
    CLA_4 KS_1652(s1652, c1652, in1652_1, in1652_2);
    wire[3:0] s1653, in1653_1, in1653_2;
    wire c1653;
    assign in1653_1 = {pp85[0],c9,c12,pp63[25]};
    assign in1653_2 = {c7,c10,s13[3],pp64[24]};
    CLA_4 KS_1653(s1653, c1653, in1653_1, in1653_2);
    wire[0:0] s1654, in1654_1, in1654_2;
    wire c1654;
    assign in1654_1 = {c8};
    assign in1654_2 = {s9[3]};
    Half_Adder KS_1654(s1654, c1654, in1654_1, in1654_2);
    wire[1:0] s1655, in1655_1, in1655_2;
    wire c1655;
    assign in1655_1 = {s10[3],s11[3]};
    assign in1655_2 = {s11[2],s12[3]};
    CLA_2 KS_1655(s1655, c1655, in1655_1, in1655_2);
    wire[0:0] s1656, in1656_1, in1656_2;
    wire c1656;
    assign in1656_1 = {s12[2]};
    assign in1656_2 = {s13[1]};
    Half_Adder KS_1656(s1656, c1656, in1656_1, in1656_2);
    wire[3:0] s1657, in1657_1, in1657_2;
    wire c1657;
    assign in1657_1 = {s14[1],s13[2],s14[3],pp65[23]};
    assign in1657_2 = {s15[1],s14[2],s15[3],pp66[22]};
    CLA_4 KS_1657(s1657, c1657, in1657_1, in1657_2);
    wire[0:0] s1658, in1658_1, in1658_2;
    wire c1658;
    assign in1658_1 = {s16[1]};
    assign in1658_2 = {s17[0]};
    Half_Adder KS_1658(s1658, c1658, in1658_1, in1658_2);
    wire[1:0] s1659, in1659_1, in1659_2;
    wire c1659;
    assign in1659_1 = {s18[0],s15[2]};
    assign in1659_2 = {s19[0],s16[2]};
    CLA_2 KS_1659(s1659, c1659, in1659_1, in1659_2);
    wire[0:0] s1660, in1660_1, in1660_2;
    wire c1660;
    assign in1660_1 = {c1576};
    assign in1660_2 = {c1577};
    Half_Adder KS_1660(s1660, c1660, in1660_1, in1660_2);
    wire[3:0] s1661, in1661_1, in1661_2;
    wire c1661;
    assign in1661_1 = {c1578,s17[1],s16[3],pp67[21]};
    assign in1661_2 = {c1579,s18[1],s17[2],pp68[20]};
    CLA_4 KS_1661(s1661, c1661, in1661_1, in1661_2);
    wire[0:0] s1662, in1662_1, in1662_2;
    wire c1662;
    assign in1662_1 = {c1580};
    assign in1662_2 = {c1581};
    Half_Adder KS_1662(s1662, c1662, in1662_1, in1662_2);
    wire[1:0] s1663, in1663_1, in1663_2;
    wire c1663;
    assign in1663_1 = {c1582,s19[1]};
    assign in1663_2 = {c1583,s20[0]};
    CLA_2 KS_1663(s1663, c1663, in1663_1, in1663_2);
    wire[0:0] s1664, in1664_1, in1664_2;
    wire c1664;
    assign in1664_1 = {c1584};
    assign in1664_2 = {c1585};
    Half_Adder KS_1664(s1664, c1664, in1664_1, in1664_2);
    wire[3:0] s1665, in1665_1, in1665_2;
    wire c1665;
    assign in1665_1 = {c1586,s21[0],s18[2],pp69[19]};
    assign in1665_2 = {c1587,s22[0],s19[2],pp70[18]};
    CLA_4 KS_1665(s1665, c1665, in1665_1, in1665_2);
    wire[0:0] s1666, in1666_1, in1666_2;
    wire c1666;
    assign in1666_1 = {c1588};
    assign in1666_2 = {c1589};
    Half_Adder KS_1666(s1666, c1666, in1666_1, in1666_2);
    wire[1:0] s1667, in1667_1, in1667_2;
    wire c1667;
    assign in1667_1 = {c1590,s1622[2]};
    assign in1667_2 = {c1591,s1623[2]};
    CLA_2 KS_1667(s1667, c1667, in1667_1, in1667_2);
    wire[0:0] s1668, in1668_1, in1668_2;
    wire c1668;
    assign in1668_1 = {c1592};
    assign in1668_2 = {c1593};
    Half_Adder KS_1668(s1668, c1668, in1668_1, in1668_2);
    wire[3:0] s1669, in1669_1, in1669_2;
    wire c1669;
    assign in1669_1 = {c1594,s1624[2],s20[1],pp71[17]};
    assign in1669_2 = {c1595,s1625[2],s21[1],pp72[16]};
    CLA_4 KS_1669(s1669, c1669, in1669_1, in1669_2);
    wire[0:0] s1670, in1670_1, in1670_2;
    wire c1670;
    assign in1670_1 = {c1599};
    assign in1670_2 = {c1603};
    Half_Adder KS_1670(s1670, c1670, in1670_1, in1670_2);
    wire[1:0] s1671, in1671_1, in1671_2;
    wire c1671;
    assign in1671_1 = {c1607,s1626[2]};
    assign in1671_2 = {c1611,s1627[2]};
    CLA_2 KS_1671(s1671, c1671, in1671_1, in1671_2);
    wire[0:0] s1672, in1672_1, in1672_2;
    wire c1672;
    assign in1672_1 = {c1615};
    assign in1672_2 = {c1619};
    Half_Adder KS_1672(s1672, c1672, in1672_1, in1672_2);
    wire[3:0] s1673, in1673_1, in1673_2;
    wire c1673;
    assign in1673_1 = {s1622[1],s1628[2],s22[1],pp73[15]};
    assign in1673_2 = {s1623[1],s1629[2],s23[0],pp74[14]};
    CLA_4 KS_1673(s1673, c1673, in1673_1, in1673_2);
    wire[0:0] s1674, in1674_1, in1674_2;
    wire c1674;
    assign in1674_1 = {s1624[1]};
    assign in1674_2 = {s1625[1]};
    Half_Adder KS_1674(s1674, c1674, in1674_1, in1674_2);
    wire[1:0] s1675, in1675_1, in1675_2;
    wire c1675;
    assign in1675_1 = {s1626[1],s1630[2]};
    assign in1675_2 = {s1627[1],s1631[2]};
    CLA_2 KS_1675(s1675, c1675, in1675_1, in1675_2);
    wire[0:0] s1676, in1676_1, in1676_2;
    wire c1676;
    assign in1676_1 = {s1628[1]};
    assign in1676_2 = {s1629[1]};
    Half_Adder KS_1676(s1676, c1676, in1676_1, in1676_2);
    wire[3:0] s1677, in1677_1, in1677_2;
    wire c1677;
    assign in1677_1 = {s1631[1],s1632[2],s24[0],pp75[13]};
    assign in1677_2 = {s1632[1],s1633[2],s25[0],pp76[12]};
    CLA_4_c KS_1677(s1677, c1677, in1677_1, in1677_2, s1630[1]);
    wire[3:0] s1678, in1678_1, in1678_2;
    wire c1678;
    assign in1678_1 = {pp77[11],pp33[56],pp35[55],pp37[54]};
    assign in1678_2 = {pp78[10],pp34[55],pp36[54],pp38[53]};
    CLA_4 KS_1678(s1678, c1678, in1678_1, in1678_2);
    wire[3:0] s1679, in1679_1, in1679_2;
    wire c1679;
    assign in1679_1 = {pp79[9],pp35[54],pp37[53],pp39[52]};
    assign in1679_2 = {pp80[8],pp36[53],pp38[52],pp40[51]};
    CLA_4 KS_1679(s1679, c1679, in1679_1, in1679_2);
    wire[3:0] s1680, in1680_1, in1680_2;
    wire c1680;
    assign in1680_1 = {pp81[7],pp37[52],pp39[51],pp41[50]};
    assign in1680_2 = {pp82[6],pp38[51],pp40[50],pp42[49]};
    CLA_4 KS_1680(s1680, c1680, in1680_1, in1680_2);
    wire[3:0] s1681, in1681_1, in1681_2;
    wire c1681;
    assign in1681_1 = {pp83[5],pp39[50],pp41[49],pp43[48]};
    assign in1681_2 = {pp84[4],pp40[49],pp42[48],pp44[47]};
    CLA_4 KS_1681(s1681, c1681, in1681_1, in1681_2);
    wire[3:0] s1682, in1682_1, in1682_2;
    wire c1682;
    assign in1682_1 = {pp85[3],pp41[48],pp43[47],pp45[46]};
    assign in1682_2 = {pp86[2],pp42[47],pp44[46],pp46[45]};
    CLA_4 KS_1682(s1682, c1682, in1682_1, in1682_2);
    wire[3:0] s1683, in1683_1, in1683_2;
    wire c1683;
    assign in1683_1 = {pp87[1],pp43[46],pp45[45],pp47[44]};
    assign in1683_2 = {pp88[0],pp44[45],pp46[44],pp48[43]};
    CLA_4 KS_1683(s1683, c1683, in1683_1, in1683_2);
    wire[3:0] s1684, in1684_1, in1684_2;
    wire c1684;
    assign in1684_1 = {c13,pp45[44],pp47[43],pp49[42]};
    assign in1684_2 = {c14,pp46[43],pp48[42],pp50[41]};
    CLA_4 KS_1684(s1684, c1684, in1684_1, in1684_2);
    wire[3:0] s1685, in1685_1, in1685_2;
    wire c1685;
    assign in1685_1 = {c15,pp47[42],pp49[41],pp51[40]};
    assign in1685_2 = {c16,pp48[41],pp50[40],pp52[39]};
    CLA_4 KS_1685(s1685, c1685, in1685_1, in1685_2);
    wire[3:0] s1686, in1686_1, in1686_2;
    wire c1686;
    assign in1686_1 = {s17[3],pp49[40],pp51[39],pp53[38]};
    assign in1686_2 = {s18[3],pp50[39],pp52[38],pp54[37]};
    CLA_4 KS_1686(s1686, c1686, in1686_1, in1686_2);
    wire[3:0] s1687, in1687_1, in1687_2;
    wire c1687;
    assign in1687_1 = {s19[3],pp51[38],pp53[37],pp55[36]};
    assign in1687_2 = {s20[2],pp52[37],pp54[36],pp56[35]};
    CLA_4 KS_1687(s1687, c1687, in1687_1, in1687_2);
    wire[3:0] s1688, in1688_1, in1688_2;
    wire c1688;
    assign in1688_1 = {s21[2],pp53[36],pp55[35],pp57[34]};
    assign in1688_2 = {s22[2],pp54[35],pp56[34],pp58[33]};
    CLA_4 KS_1688(s1688, c1688, in1688_1, in1688_2);
    wire[3:0] s1689, in1689_1, in1689_2;
    wire c1689;
    assign in1689_1 = {s23[1],pp55[34],pp57[33],pp59[32]};
    assign in1689_2 = {s24[1],pp56[33],pp58[32],pp60[31]};
    CLA_4 KS_1689(s1689, c1689, in1689_1, in1689_2);
    wire[3:0] s1690, in1690_1, in1690_2;
    wire c1690;
    assign in1690_1 = {s25[1],pp57[32],pp59[31],pp61[30]};
    assign in1690_2 = {s26[0],pp58[31],pp60[30],pp62[29]};
    CLA_4 KS_1690(s1690, c1690, in1690_1, in1690_2);
    wire[3:0] s1691, in1691_1, in1691_2;
    wire c1691;
    assign in1691_1 = {s27[0],pp59[30],pp61[29],pp63[28]};
    assign in1691_2 = {s28[0],pp60[29],pp62[28],pp64[27]};
    CLA_4 KS_1691(s1691, c1691, in1691_1, in1691_2);
    wire[3:0] s1692, in1692_1, in1692_2;
    wire c1692;
    assign in1692_1 = {s29[0],pp61[28],pp63[27],pp65[26]};
    assign in1692_2 = {s30[0],pp62[27],pp64[26],pp66[25]};
    CLA_4 KS_1692(s1692, c1692, in1692_1, in1692_2);
    wire[3:0] s1693, in1693_1, in1693_2;
    wire c1693;
    assign in1693_1 = {s31[0],pp63[26],pp65[25],pp67[24]};
    assign in1693_2 = {s32[0],pp64[25],pp66[24],pp68[23]};
    CLA_4 KS_1693(s1693, c1693, in1693_1, in1693_2);
    wire[3:0] s1694, in1694_1, in1694_2;
    wire c1694;
    assign in1694_1 = {c1622,pp65[24],pp67[23],pp69[22]};
    assign in1694_2 = {c1623,pp66[23],pp68[22],pp70[21]};
    CLA_4 KS_1694(s1694, c1694, in1694_1, in1694_2);
    wire[3:0] s1695, in1695_1, in1695_2;
    wire c1695;
    assign in1695_1 = {c1624,pp67[22],pp69[21],pp71[20]};
    assign in1695_2 = {c1625,pp68[21],pp70[20],pp72[19]};
    CLA_4 KS_1695(s1695, c1695, in1695_1, in1695_2);
    wire[3:0] s1696, in1696_1, in1696_2;
    wire c1696;
    assign in1696_1 = {c1626,pp69[20],pp71[19],pp73[18]};
    assign in1696_2 = {c1627,pp70[19],pp72[18],pp74[17]};
    CLA_4 KS_1696(s1696, c1696, in1696_1, in1696_2);
    wire[3:0] s1697, in1697_1, in1697_2;
    wire c1697;
    assign in1697_1 = {c1628,pp71[18],pp73[17],pp75[16]};
    assign in1697_2 = {c1629,pp72[17],pp74[16],pp76[15]};
    CLA_4 KS_1697(s1697, c1697, in1697_1, in1697_2);
    wire[3:0] s1698, in1698_1, in1698_2;
    wire c1698;
    assign in1698_1 = {c1630,pp73[16],pp75[15],pp77[14]};
    assign in1698_2 = {c1631,pp74[15],pp76[14],pp78[13]};
    CLA_4 KS_1698(s1698, c1698, in1698_1, in1698_2);
    wire[3:0] s1699, in1699_1, in1699_2;
    wire c1699;
    assign in1699_1 = {c1632,pp75[14],pp77[13],pp79[12]};
    assign in1699_2 = {c1633,pp76[13],pp78[12],pp80[11]};
    CLA_4 KS_1699(s1699, c1699, in1699_1, in1699_2);
    wire[3:0] s1700, in1700_1, in1700_2;
    wire c1700;
    assign in1700_1 = {c1634,pp77[12],pp79[11],pp81[10]};
    assign in1700_2 = {c1635,pp78[11],pp80[10],pp82[9]};
    CLA_4 KS_1700(s1700, c1700, in1700_1, in1700_2);
    wire[3:0] s1701, in1701_1, in1701_2;
    wire c1701;
    assign in1701_1 = {c1637,pp79[10],pp81[9],pp83[8]};
    assign in1701_2 = {s1638[3],pp80[9],pp82[8],pp84[7]};
    CLA_4_c KS_1701(s1701, c1701, in1701_1, in1701_2, c1636);
    wire[3:0] s1702, in1702_1, in1702_2;
    wire c1702;
    assign in1702_1 = {pp81[8],pp83[7],pp85[6],pp47[45]};
    assign in1702_2 = {pp82[7],pp84[6],pp86[5],pp48[44]};
    CLA_4 KS_1702(s1702, c1702, in1702_1, in1702_2);
    wire[3:0] s1703, in1703_1, in1703_2;
    wire c1703;
    assign in1703_1 = {pp83[6],pp85[5],pp87[4],pp49[43]};
    assign in1703_2 = {pp84[5],pp86[4],pp88[3],pp50[42]};
    CLA_4 KS_1703(s1703, c1703, in1703_1, in1703_2);
    wire[3:0] s1704, in1704_1, in1704_2;
    wire c1704;
    assign in1704_1 = {pp85[4],pp87[3],pp89[2],pp51[41]};
    assign in1704_2 = {pp86[3],pp88[2],pp90[1],pp52[40]};
    CLA_4 KS_1704(s1704, c1704, in1704_1, in1704_2);
    wire[3:0] s1705, in1705_1, in1705_2;
    wire c1705;
    assign in1705_1 = {pp87[2],pp89[1],pp91[0],pp53[39]};
    assign in1705_2 = {pp88[1],pp90[0],c23,pp54[38]};
    CLA_4 KS_1705(s1705, c1705, in1705_1, in1705_2);
    wire[3:0] s1706, in1706_1, in1706_2;
    wire c1706;
    assign in1706_1 = {pp89[0],c20,c24,pp55[37]};
    assign in1706_2 = {c17,c21,c25,pp56[36]};
    CLA_4 KS_1706(s1706, c1706, in1706_1, in1706_2);
    wire[3:0] s1707, in1707_1, in1707_2;
    wire c1707;
    assign in1707_1 = {c18,c22,s26[3],pp57[35]};
    assign in1707_2 = {c19,s23[3],s27[3],pp58[34]};
    CLA_4 KS_1707(s1707, c1707, in1707_1, in1707_2);
    wire[3:0] s1708, in1708_1, in1708_2;
    wire c1708;
    assign in1708_1 = {s20[3],s24[3],s28[3],pp59[33]};
    assign in1708_2 = {s21[3],s25[3],s29[3],pp60[32]};
    CLA_4 KS_1708(s1708, c1708, in1708_1, in1708_2);
    wire[3:0] s1709, in1709_1, in1709_2;
    wire c1709;
    assign in1709_1 = {s22[3],s26[2],s30[3],pp61[31]};
    assign in1709_2 = {s23[2],s27[2],s31[3],pp62[30]};
    CLA_4 KS_1709(s1709, c1709, in1709_1, in1709_2);
    wire[0:0] s1710, in1710_1, in1710_2;
    wire c1710;
    assign in1710_1 = {s24[2]};
    assign in1710_2 = {s25[2]};
    Half_Adder KS_1710(s1710, c1710, in1710_1, in1710_2);
    wire[1:0] s1711, in1711_1, in1711_2;
    wire c1711;
    assign in1711_1 = {s26[1],s28[2]};
    assign in1711_2 = {s27[1],s29[2]};
    CLA_2 KS_1711(s1711, c1711, in1711_1, in1711_2);
    wire[0:0] s1712, in1712_1, in1712_2;
    wire c1712;
    assign in1712_1 = {s28[1]};
    assign in1712_2 = {s29[1]};
    Half_Adder KS_1712(s1712, c1712, in1712_1, in1712_2);
    wire[3:0] s1713, in1713_1, in1713_2;
    wire c1713;
    assign in1713_1 = {s30[1],s30[2],s32[3],pp63[29]};
    assign in1713_2 = {s31[1],s31[2],s33[2],pp64[28]};
    CLA_4 KS_1713(s1713, c1713, in1713_1, in1713_2);
    wire[0:0] s1714, in1714_1, in1714_2;
    wire c1714;
    assign in1714_1 = {s32[1]};
    assign in1714_2 = {s33[0]};
    Half_Adder KS_1714(s1714, c1714, in1714_1, in1714_2);
    wire[1:0] s1715, in1715_1, in1715_2;
    wire c1715;
    assign in1715_1 = {s34[0],s32[2]};
    assign in1715_2 = {s35[0],s33[1]};
    CLA_2 KS_1715(s1715, c1715, in1715_1, in1715_2);
    wire[0:0] s1716, in1716_1, in1716_2;
    wire c1716;
    assign in1716_1 = {c1638};
    assign in1716_2 = {c1639};
    Half_Adder KS_1716(s1716, c1716, in1716_1, in1716_2);
    wire[3:0] s1717, in1717_1, in1717_2;
    wire c1717;
    assign in1717_1 = {c1640,s34[1],s34[2],pp65[27]};
    assign in1717_2 = {c1641,s35[1],s35[2],pp66[26]};
    CLA_4 KS_1717(s1717, c1717, in1717_1, in1717_2);
    wire[0:0] s1718, in1718_1, in1718_2;
    wire c1718;
    assign in1718_1 = {c1642};
    assign in1718_2 = {c1643};
    Half_Adder KS_1718(s1718, c1718, in1718_1, in1718_2);
    wire[1:0] s1719, in1719_1, in1719_2;
    wire c1719;
    assign in1719_1 = {c1644,s36[0]};
    assign in1719_2 = {c1645,s37[0]};
    CLA_2 KS_1719(s1719, c1719, in1719_1, in1719_2);
    wire[0:0] s1720, in1720_1, in1720_2;
    wire c1720;
    assign in1720_1 = {c1646};
    assign in1720_2 = {c1647};
    Half_Adder KS_1720(s1720, c1720, in1720_1, in1720_2);
    wire[3:0] s1721, in1721_1, in1721_2;
    wire c1721;
    assign in1721_1 = {c1648,s38[0],s36[1],pp67[25]};
    assign in1721_2 = {c1649,s39[0],s37[1],pp68[24]};
    CLA_4 KS_1721(s1721, c1721, in1721_1, in1721_2);
    wire[0:0] s1722, in1722_1, in1722_2;
    wire c1722;
    assign in1722_1 = {c1650};
    assign in1722_2 = {c1651};
    Half_Adder KS_1722(s1722, c1722, in1722_1, in1722_2);
    wire[1:0] s1723, in1723_1, in1723_2;
    wire c1723;
    assign in1723_1 = {c1652,s1678[2]};
    assign in1723_2 = {c1653,s1679[2]};
    CLA_2 KS_1723(s1723, c1723, in1723_1, in1723_2);
    wire[0:0] s1724, in1724_1, in1724_2;
    wire c1724;
    assign in1724_1 = {c1657};
    assign in1724_2 = {c1661};
    Half_Adder KS_1724(s1724, c1724, in1724_1, in1724_2);
    wire[3:0] s1725, in1725_1, in1725_2;
    wire c1725;
    assign in1725_1 = {c1665,s1680[2],s38[1],pp69[23]};
    assign in1725_2 = {c1669,s1681[2],s39[1],pp70[22]};
    CLA_4 KS_1725(s1725, c1725, in1725_1, in1725_2);
    wire[0:0] s1726, in1726_1, in1726_2;
    wire c1726;
    assign in1726_1 = {c1673};
    assign in1726_2 = {c1677};
    Half_Adder KS_1726(s1726, c1726, in1726_1, in1726_2);
    wire[1:0] s1727, in1727_1, in1727_2;
    wire c1727;
    assign in1727_1 = {s1678[1],s1682[2]};
    assign in1727_2 = {s1679[1],s1683[2]};
    CLA_2 KS_1727(s1727, c1727, in1727_1, in1727_2);
    wire[0:0] s1728, in1728_1, in1728_2;
    wire c1728;
    assign in1728_1 = {s1680[1]};
    assign in1728_2 = {s1681[1]};
    Half_Adder KS_1728(s1728, c1728, in1728_1, in1728_2);
    wire[3:0] s1729, in1729_1, in1729_2;
    wire c1729;
    assign in1729_1 = {s1683[1],s1684[2],s40[0],pp71[21]};
    assign in1729_2 = {s1684[1],s1685[2],s41[0],pp72[20]};
    CLA_4_c KS_1729(s1729, c1729, in1729_1, in1729_2, s1682[1]);
    wire[3:0] s1730, in1730_1, in1730_2;
    wire c1730;
    assign in1730_1 = {pp73[19],pp42[51],pp45[49],pp47[48]};
    assign in1730_2 = {pp74[18],pp43[50],pp46[48],pp48[47]};
    CLA_4 KS_1730(s1730, c1730, in1730_1, in1730_2);
    wire[3:0] s1731, in1731_1, in1731_2;
    wire c1731;
    assign in1731_1 = {pp75[17],pp44[49],pp47[47],pp49[46]};
    assign in1731_2 = {pp76[16],pp45[48],pp48[46],pp50[45]};
    CLA_4 KS_1731(s1731, c1731, in1731_1, in1731_2);
    wire[3:0] s1732, in1732_1, in1732_2;
    wire c1732;
    assign in1732_1 = {pp77[15],pp46[47],pp49[45],pp51[44]};
    assign in1732_2 = {pp78[14],pp47[46],pp50[44],pp52[43]};
    CLA_4 KS_1732(s1732, c1732, in1732_1, in1732_2);
    wire[3:0] s1733, in1733_1, in1733_2;
    wire c1733;
    assign in1733_1 = {pp79[13],pp48[45],pp51[43],pp53[42]};
    assign in1733_2 = {pp80[12],pp49[44],pp52[42],pp54[41]};
    CLA_4 KS_1733(s1733, c1733, in1733_1, in1733_2);
    wire[3:0] s1734, in1734_1, in1734_2;
    wire c1734;
    assign in1734_1 = {pp81[11],pp50[43],pp53[41],pp55[40]};
    assign in1734_2 = {pp82[10],pp51[42],pp54[40],pp56[39]};
    CLA_4 KS_1734(s1734, c1734, in1734_1, in1734_2);
    wire[3:0] s1735, in1735_1, in1735_2;
    wire c1735;
    assign in1735_1 = {pp83[9],pp52[41],pp55[39],pp57[38]};
    assign in1735_2 = {pp84[8],pp53[40],pp56[38],pp58[37]};
    CLA_4 KS_1735(s1735, c1735, in1735_1, in1735_2);
    wire[3:0] s1736, in1736_1, in1736_2;
    wire c1736;
    assign in1736_1 = {pp85[7],pp54[39],pp57[37],pp59[36]};
    assign in1736_2 = {pp86[6],pp55[38],pp58[36],pp60[35]};
    CLA_4 KS_1736(s1736, c1736, in1736_1, in1736_2);
    wire[3:0] s1737, in1737_1, in1737_2;
    wire c1737;
    assign in1737_1 = {pp87[5],pp56[37],pp59[35],pp61[34]};
    assign in1737_2 = {pp88[4],pp57[36],pp60[34],pp62[33]};
    CLA_4 KS_1737(s1737, c1737, in1737_1, in1737_2);
    wire[3:0] s1738, in1738_1, in1738_2;
    wire c1738;
    assign in1738_1 = {pp89[3],pp58[35],pp61[33],pp63[32]};
    assign in1738_2 = {pp90[2],pp59[34],pp62[32],pp64[31]};
    CLA_4 KS_1738(s1738, c1738, in1738_1, in1738_2);
    wire[3:0] s1739, in1739_1, in1739_2;
    wire c1739;
    assign in1739_1 = {pp91[1],pp60[33],pp63[31],pp65[30]};
    assign in1739_2 = {pp92[0],pp61[32],pp64[30],pp66[29]};
    CLA_4 KS_1739(s1739, c1739, in1739_1, in1739_2);
    wire[3:0] s1740, in1740_1, in1740_2;
    wire c1740;
    assign in1740_1 = {c26,pp62[31],pp65[29],pp67[28]};
    assign in1740_2 = {c27,pp63[30],pp66[28],pp68[27]};
    CLA_4 KS_1740(s1740, c1740, in1740_1, in1740_2);
    wire[3:0] s1741, in1741_1, in1741_2;
    wire c1741;
    assign in1741_1 = {c28,pp64[29],pp67[27],pp69[26]};
    assign in1741_2 = {c29,pp65[28],pp68[26],pp70[25]};
    CLA_4 KS_1741(s1741, c1741, in1741_1, in1741_2);
    wire[3:0] s1742, in1742_1, in1742_2;
    wire c1742;
    assign in1742_1 = {c30,pp66[27],pp69[25],pp71[24]};
    assign in1742_2 = {c31,pp67[26],pp70[24],pp72[23]};
    CLA_4 KS_1742(s1742, c1742, in1742_1, in1742_2);
    wire[3:0] s1743, in1743_1, in1743_2;
    wire c1743;
    assign in1743_1 = {c32,pp68[25],pp71[23],pp73[22]};
    assign in1743_2 = {s33[3],pp69[24],pp72[22],pp74[21]};
    CLA_4 KS_1743(s1743, c1743, in1743_1, in1743_2);
    wire[3:0] s1744, in1744_1, in1744_2;
    wire c1744;
    assign in1744_1 = {s34[3],pp70[23],pp73[21],pp75[20]};
    assign in1744_2 = {s35[3],pp71[22],pp74[20],pp76[19]};
    CLA_4 KS_1744(s1744, c1744, in1744_1, in1744_2);
    wire[3:0] s1745, in1745_1, in1745_2;
    wire c1745;
    assign in1745_1 = {s36[2],pp72[21],pp75[19],pp77[18]};
    assign in1745_2 = {s37[2],pp73[20],pp76[18],pp78[17]};
    CLA_4 KS_1745(s1745, c1745, in1745_1, in1745_2);
    wire[3:0] s1746, in1746_1, in1746_2;
    wire c1746;
    assign in1746_1 = {s38[2],pp74[19],pp77[17],pp79[16]};
    assign in1746_2 = {s39[2],pp75[18],pp78[16],pp80[15]};
    CLA_4 KS_1746(s1746, c1746, in1746_1, in1746_2);
    wire[3:0] s1747, in1747_1, in1747_2;
    wire c1747;
    assign in1747_1 = {s40[1],pp76[17],pp79[15],pp81[14]};
    assign in1747_2 = {s41[1],pp77[16],pp80[14],pp82[13]};
    CLA_4 KS_1747(s1747, c1747, in1747_1, in1747_2);
    wire[3:0] s1748, in1748_1, in1748_2;
    wire c1748;
    assign in1748_1 = {s42[1],pp78[15],pp81[13],pp83[12]};
    assign in1748_2 = {s43[1],pp79[14],pp82[12],pp84[11]};
    CLA_4 KS_1748(s1748, c1748, in1748_1, in1748_2);
    wire[3:0] s1749, in1749_1, in1749_2;
    wire c1749;
    assign in1749_1 = {s44[0],pp80[13],pp83[11],pp85[10]};
    assign in1749_2 = {s45[0],pp81[12],pp84[10],pp86[9]};
    CLA_4 KS_1749(s1749, c1749, in1749_1, in1749_2);
    wire[3:0] s1750, in1750_1, in1750_2;
    wire c1750;
    assign in1750_1 = {s46[0],pp82[11],pp85[9],pp87[8]};
    assign in1750_2 = {s47[0],pp83[10],pp86[8],pp88[7]};
    CLA_4 KS_1750(s1750, c1750, in1750_1, in1750_2);
    wire[3:0] s1751, in1751_1, in1751_2;
    wire c1751;
    assign in1751_1 = {s48[0],pp84[9],pp87[7],pp89[6]};
    assign in1751_2 = {s49[0],pp85[8],pp88[6],pp90[5]};
    CLA_4 KS_1751(s1751, c1751, in1751_1, in1751_2);
    wire[3:0] s1752, in1752_1, in1752_2;
    wire c1752;
    assign in1752_1 = {s50[0],pp86[7],pp89[5],pp91[4]};
    assign in1752_2 = {s51[0],pp87[6],pp90[4],pp92[3]};
    CLA_4 KS_1752(s1752, c1752, in1752_1, in1752_2);
    wire[3:0] s1753, in1753_1, in1753_2;
    wire c1753;
    assign in1753_1 = {s52[0],pp88[5],pp91[3],pp93[2]};
    assign in1753_2 = {s53[0],pp89[4],pp92[2],pp94[1]};
    CLA_4 KS_1753(s1753, c1753, in1753_1, in1753_2);
    wire[3:0] s1754, in1754_1, in1754_2;
    wire c1754;
    assign in1754_1 = {s54[0],pp90[3],pp93[1],pp95[0]};
    assign in1754_2 = {s55[0],pp91[2],pp94[0],c40};
    CLA_4 KS_1754(s1754, c1754, in1754_1, in1754_2);
    wire[3:0] s1755, in1755_1, in1755_2;
    wire c1755;
    assign in1755_1 = {c1678,pp92[1],c36,c41};
    assign in1755_2 = {c1679,pp93[0],c37,c42};
    CLA_4 KS_1755(s1755, c1755, in1755_1, in1755_2);
    wire[3:0] s1756, in1756_1, in1756_2;
    wire c1756;
    assign in1756_1 = {c1680,c33,c38,c43};
    assign in1756_2 = {c1681,c34,c39,s44[3]};
    CLA_4 KS_1756(s1756, c1756, in1756_1, in1756_2);
    wire[3:0] s1757, in1757_1, in1757_2;
    wire c1757;
    assign in1757_1 = {c1682,c35,s40[3],s45[3]};
    assign in1757_2 = {c1683,s36[3],s41[3],s46[3]};
    CLA_4 KS_1757(s1757, c1757, in1757_1, in1757_2);
    wire[3:0] s1758, in1758_1, in1758_2;
    wire c1758;
    assign in1758_1 = {c1684,s37[3],s42[3],s47[3]};
    assign in1758_2 = {c1685,s38[3],s43[3],s48[3]};
    CLA_4 KS_1758(s1758, c1758, in1758_1, in1758_2);
    wire[3:0] s1759, in1759_1, in1759_2;
    wire c1759;
    assign in1759_1 = {c1686,s39[3],s44[2],s49[3]};
    assign in1759_2 = {c1687,s40[2],s45[2],s50[3]};
    CLA_4 KS_1759(s1759, c1759, in1759_1, in1759_2);
    wire[3:0] s1760, in1760_1, in1760_2;
    wire c1760;
    assign in1760_1 = {c1688,s41[2],s46[2],s51[3]};
    assign in1760_2 = {c1689,s42[2],s47[2],s52[3]};
    CLA_4 KS_1760(s1760, c1760, in1760_1, in1760_2);
    wire[3:0] s1761, in1761_1, in1761_2;
    wire c1761;
    assign in1761_1 = {c1690,s43[2],s48[2],s53[3]};
    assign in1761_2 = {c1691,s44[1],s49[2],s54[3]};
    CLA_4 KS_1761(s1761, c1761, in1761_1, in1761_2);
    wire[1:0] s1762, in1762_1, in1762_2;
    wire c1762;
    assign in1762_1 = {c1692,s45[1]};
    assign in1762_2 = {c1693,s46[1]};
    CLA_2 KS_1762(s1762, c1762, in1762_1, in1762_2);
    wire[2:0] s1763, in1763_1, in1763_2;
    wire c1763;
    assign in1763_1 = {c1694,s47[1],s50[2]};
    assign in1763_2 = {c1695,s48[1],s51[2]};
    CLA_3 KS_1763(s1763, c1763, in1763_1, in1763_2);
    wire[1:0] s1764, in1764_1, in1764_2;
    wire c1764;
    assign in1764_1 = {c1696,s49[1]};
    assign in1764_2 = {c1697,s50[1]};
    CLA_2 KS_1764(s1764, c1764, in1764_1, in1764_2);
    wire[3:0] s1765, in1765_1, in1765_2;
    wire c1765;
    assign in1765_1 = {c1698,s51[1],s52[2],s55[3]};
    assign in1765_2 = {c1699,s52[1],s53[2],s56[2]};
    CLA_4 KS_1765(s1765, c1765, in1765_1, in1765_2);
    wire[1:0] s1766, in1766_1, in1766_2;
    wire c1766;
    assign in1766_1 = {c1700,s53[1]};
    assign in1766_2 = {c1701,s54[1]};
    CLA_2 KS_1766(s1766, c1766, in1766_1, in1766_2);
    wire[2:0] s1767, in1767_1, in1767_2;
    wire c1767;
    assign in1767_1 = {s1702[3],s55[1],s54[2]};
    assign in1767_2 = {s1703[3],s56[0],s55[2]};
    CLA_3 KS_1767(s1767, c1767, in1767_1, in1767_2);
    wire[1:0] s1768, in1768_1, in1768_2;
    wire c1768;
    assign in1768_1 = {s1704[3],c1702};
    assign in1768_2 = {s1705[3],c1703};
    CLA_2 KS_1768(s1768, c1768, in1768_1, in1768_2);
    wire[3:0] s1769, in1769_1, in1769_2;
    wire c1769;
    assign in1769_1 = {s1706[3],c1704,s56[1],s57[1]};
    assign in1769_2 = {s1707[3],c1705,s57[0],s58[1]};
    CLA_4 KS_1769(s1769, c1769, in1769_1, in1769_2);
    wire[1:0] s1770, in1770_1, in1770_2;
    wire c1770;
    assign in1770_1 = {s1709[3],c1706};
    assign in1770_2 = {s1713[3],c1707};
    CLA_2_c KS_1770(s1770, c1770, in1770_1, in1770_2, s1708[3]);
    wire[1:0] s1771, in1771_1, in1771_2;
    wire c1771;
    assign in1771_1 = {c1708,s58[0]};
    assign in1771_2 = {c1709,s59[0]};
    CLA_2 KS_1771(s1771, c1771, in1771_1, in1771_2);
    wire[0:0] s1772, in1772_1, in1772_2;
    wire c1772;
    assign in1772_1 = {c1717};
    assign in1772_2 = {c1721};
    Full_Adder KS_1772(s1772, c1772, in1772_1, in1772_2, c1713);
    wire[3:0] s1773, in1773_1, in1773_2;
    wire c1773;
    assign in1773_1 = {pp65[31],pp54[43],pp55[43],pp57[42]};
    assign in1773_2 = {pp66[30],pp55[42],pp56[42],pp58[41]};
    CLA_4 KS_1773(s1773, c1773, in1773_1, in1773_2);
    wire[3:0] s1774, in1774_1, in1774_2;
    wire c1774;
    assign in1774_1 = {pp67[29],pp56[41],pp57[41],pp59[40]};
    assign in1774_2 = {pp68[28],pp57[40],pp58[40],pp60[39]};
    CLA_4 KS_1774(s1774, c1774, in1774_1, in1774_2);
    wire[3:0] s1775, in1775_1, in1775_2;
    wire c1775;
    assign in1775_1 = {pp69[27],pp58[39],pp59[39],pp61[38]};
    assign in1775_2 = {pp70[26],pp59[38],pp60[38],pp62[37]};
    CLA_4 KS_1775(s1775, c1775, in1775_1, in1775_2);
    wire[3:0] s1776, in1776_1, in1776_2;
    wire c1776;
    assign in1776_1 = {pp71[25],pp60[37],pp61[37],pp63[36]};
    assign in1776_2 = {pp72[24],pp61[36],pp62[36],pp64[35]};
    CLA_4 KS_1776(s1776, c1776, in1776_1, in1776_2);
    wire[3:0] s1777, in1777_1, in1777_2;
    wire c1777;
    assign in1777_1 = {pp73[23],pp62[35],pp63[35],pp65[34]};
    assign in1777_2 = {pp74[22],pp63[34],pp64[34],pp66[33]};
    CLA_4 KS_1777(s1777, c1777, in1777_1, in1777_2);
    wire[3:0] s1778, in1778_1, in1778_2;
    wire c1778;
    assign in1778_1 = {pp75[21],pp64[33],pp65[33],pp67[32]};
    assign in1778_2 = {pp76[20],pp65[32],pp66[32],pp68[31]};
    CLA_4 KS_1778(s1778, c1778, in1778_1, in1778_2);
    wire[3:0] s1779, in1779_1, in1779_2;
    wire c1779;
    assign in1779_1 = {pp77[19],pp66[31],pp67[31],pp69[30]};
    assign in1779_2 = {pp78[18],pp67[30],pp68[30],pp70[29]};
    CLA_4 KS_1779(s1779, c1779, in1779_1, in1779_2);
    wire[3:0] s1780, in1780_1, in1780_2;
    wire c1780;
    assign in1780_1 = {pp79[17],pp68[29],pp69[29],pp71[28]};
    assign in1780_2 = {pp80[16],pp69[28],pp70[28],pp72[27]};
    CLA_4 KS_1780(s1780, c1780, in1780_1, in1780_2);
    wire[3:0] s1781, in1781_1, in1781_2;
    wire c1781;
    assign in1781_1 = {pp81[15],pp70[27],pp71[27],pp73[26]};
    assign in1781_2 = {pp82[14],pp71[26],pp72[26],pp74[25]};
    CLA_4 KS_1781(s1781, c1781, in1781_1, in1781_2);
    wire[3:0] s1782, in1782_1, in1782_2;
    wire c1782;
    assign in1782_1 = {pp83[13],pp72[25],pp73[25],pp75[24]};
    assign in1782_2 = {pp84[12],pp73[24],pp74[24],pp76[23]};
    CLA_4 KS_1782(s1782, c1782, in1782_1, in1782_2);
    wire[3:0] s1783, in1783_1, in1783_2;
    wire c1783;
    assign in1783_1 = {pp85[11],pp74[23],pp75[23],pp77[22]};
    assign in1783_2 = {pp86[10],pp75[22],pp76[22],pp78[21]};
    CLA_4 KS_1783(s1783, c1783, in1783_1, in1783_2);
    wire[3:0] s1784, in1784_1, in1784_2;
    wire c1784;
    assign in1784_1 = {pp87[9],pp76[21],pp77[21],pp79[20]};
    assign in1784_2 = {pp88[8],pp77[20],pp78[20],pp80[19]};
    CLA_4 KS_1784(s1784, c1784, in1784_1, in1784_2);
    wire[3:0] s1785, in1785_1, in1785_2;
    wire c1785;
    assign in1785_1 = {pp89[7],pp78[19],pp79[19],pp81[18]};
    assign in1785_2 = {pp90[6],pp79[18],pp80[18],pp82[17]};
    CLA_4 KS_1785(s1785, c1785, in1785_1, in1785_2);
    wire[3:0] s1786, in1786_1, in1786_2;
    wire c1786;
    assign in1786_1 = {pp91[5],pp80[17],pp81[17],pp83[16]};
    assign in1786_2 = {pp92[4],pp81[16],pp82[16],pp84[15]};
    CLA_4 KS_1786(s1786, c1786, in1786_1, in1786_2);
    wire[3:0] s1787, in1787_1, in1787_2;
    wire c1787;
    assign in1787_1 = {pp93[3],pp82[15],pp83[15],pp85[14]};
    assign in1787_2 = {pp94[2],pp83[14],pp84[14],pp86[13]};
    CLA_4 KS_1787(s1787, c1787, in1787_1, in1787_2);
    wire[3:0] s1788, in1788_1, in1788_2;
    wire c1788;
    assign in1788_1 = {pp95[1],pp84[13],pp85[13],pp87[12]};
    assign in1788_2 = {pp96[0],pp85[12],pp86[12],pp88[11]};
    CLA_4 KS_1788(s1788, c1788, in1788_1, in1788_2);
    wire[3:0] s1789, in1789_1, in1789_2;
    wire c1789;
    assign in1789_1 = {c44,pp86[11],pp87[11],pp89[10]};
    assign in1789_2 = {c45,pp87[10],pp88[10],pp90[9]};
    CLA_4 KS_1789(s1789, c1789, in1789_1, in1789_2);
    wire[3:0] s1790, in1790_1, in1790_2;
    wire c1790;
    assign in1790_1 = {c46,pp88[9],pp89[9],pp91[8]};
    assign in1790_2 = {c47,pp89[8],pp90[8],pp92[7]};
    CLA_4 KS_1790(s1790, c1790, in1790_1, in1790_2);
    wire[3:0] s1791, in1791_1, in1791_2;
    wire c1791;
    assign in1791_1 = {c48,pp90[7],pp91[7],pp93[6]};
    assign in1791_2 = {c49,pp91[6],pp92[6],pp94[5]};
    CLA_4 KS_1791(s1791, c1791, in1791_1, in1791_2);
    wire[3:0] s1792, in1792_1, in1792_2;
    wire c1792;
    assign in1792_1 = {c50,pp92[5],pp93[5],pp95[4]};
    assign in1792_2 = {c51,pp93[4],pp94[4],pp96[3]};
    CLA_4 KS_1792(s1792, c1792, in1792_1, in1792_2);
    wire[3:0] s1793, in1793_1, in1793_2;
    wire c1793;
    assign in1793_1 = {c52,pp94[3],pp95[3],pp97[2]};
    assign in1793_2 = {c53,pp95[2],pp96[2],pp98[1]};
    CLA_4 KS_1793(s1793, c1793, in1793_1, in1793_2);
    wire[3:0] s1794, in1794_1, in1794_2;
    wire c1794;
    assign in1794_1 = {c54,pp96[1],pp97[1],pp99[0]};
    assign in1794_2 = {c55,pp97[0],pp98[0],c62};
    CLA_4 KS_1794(s1794, c1794, in1794_1, in1794_2);
    wire[3:0] s1795, in1795_1, in1795_2;
    wire c1795;
    assign in1795_1 = {s56[3],c56,c57,c63};
    assign in1795_2 = {s57[2],s57[3],c58,c64};
    CLA_4 KS_1795(s1795, c1795, in1795_1, in1795_2);
    wire[3:0] s1796, in1796_1, in1796_2;
    wire c1796;
    assign in1796_1 = {s58[2],s58[3],c59,c65};
    assign in1796_2 = {s59[2],s59[3],c60,c66};
    CLA_4 KS_1796(s1796, c1796, in1796_1, in1796_2);
    wire[3:0] s1797, in1797_1, in1797_2;
    wire c1797;
    assign in1797_1 = {s60[2],s60[3],c61,s67[3]};
    assign in1797_2 = {s61[2],s61[3],s62[3],s68[3]};
    CLA_4 KS_1797(s1797, c1797, in1797_1, in1797_2);
    wire[3:0] s1798, in1798_1, in1798_2;
    wire c1798;
    assign in1798_1 = {s62[1],s62[2],s63[3],s69[3]};
    assign in1798_2 = {s63[1],s63[2],s64[3],s70[3]};
    CLA_4 KS_1798(s1798, c1798, in1798_1, in1798_2);
    wire[3:0] s1799, in1799_1, in1799_2;
    wire c1799;
    assign in1799_1 = {s64[1],s64[2],s65[3],s71[3]};
    assign in1799_2 = {s65[1],s65[2],s66[3],s72[3]};
    CLA_4 KS_1799(s1799, c1799, in1799_1, in1799_2);
    wire[3:0] s1800, in1800_1, in1800_2;
    wire c1800;
    assign in1800_1 = {s66[1],s66[2],s67[2],s73[3]};
    assign in1800_2 = {s67[0],s67[1],s68[2],s74[3]};
    CLA_4 KS_1800(s1800, c1800, in1800_1, in1800_2);
    wire[3:0] s1801, in1801_1, in1801_2;
    wire c1801;
    assign in1801_1 = {s68[0],s68[1],s69[2],s75[3]};
    assign in1801_2 = {s69[0],s69[1],s70[2],s76[3]};
    CLA_4 KS_1801(s1801, c1801, in1801_1, in1801_2);
    wire[3:0] s1802, in1802_1, in1802_2;
    wire c1802;
    assign in1802_1 = {s70[0],s70[1],s71[2],s77[3]};
    assign in1802_2 = {s71[0],s71[1],s72[2],s78[3]};
    CLA_4 KS_1802(s1802, c1802, in1802_1, in1802_2);
    wire[3:0] s1803, in1803_1, in1803_2;
    wire c1803;
    assign in1803_1 = {s72[0],s72[1],s73[2],s79[3]};
    assign in1803_2 = {s73[0],s73[1],s74[2],s80[3]};
    CLA_4 KS_1803(s1803, c1803, in1803_1, in1803_2);
    wire[3:0] s1804, in1804_1, in1804_2;
    wire c1804;
    assign in1804_1 = {s74[0],s74[1],s75[2],s82[3]};
    assign in1804_2 = {s75[0],s75[1],s76[2],s84[3]};
    CLA_4 KS_1804(s1804, c1804, in1804_1, in1804_2);
    wire[0:0] s1805, in1805_1, in1805_2;
    wire c1805;
    assign in1805_1 = {s76[0]};
    assign in1805_2 = {s77[0]};
    Half_Adder KS_1805(s1805, c1805, in1805_1, in1805_2);
    wire[1:0] s1806, in1806_1, in1806_2;
    wire c1806;
    assign in1806_1 = {s78[0],s76[1]};
    assign in1806_2 = {s79[0],s77[1]};
    CLA_2 KS_1806(s1806, c1806, in1806_1, in1806_2);
    wire[0:0] s1807, in1807_1, in1807_2;
    wire c1807;
    assign in1807_1 = {s80[0]};
    assign in1807_2 = {s81[0]};
    Half_Adder KS_1807(s1807, c1807, in1807_1, in1807_2);
    wire[2:0] s1808, in1808_1, in1808_2;
    wire c1808;
    assign in1808_1 = {s82[0],s78[1],s77[2]};
    assign in1808_2 = {s83[0],s79[1],s78[2]};
    CLA_3 KS_1808(s1808, c1808, in1808_1, in1808_2);
    wire[0:0] s1809, in1809_1, in1809_2;
    wire c1809;
    assign in1809_1 = {s84[0]};
    assign in1809_2 = {s85[0]};
    Half_Adder KS_1809(s1809, c1809, in1809_1, in1809_2);
    wire[1:0] s1810, in1810_1, in1810_2;
    wire c1810;
    assign in1810_1 = {s86[0],s80[1]};
    assign in1810_2 = {s87[0],c81};
    CLA_2 KS_1810(s1810, c1810, in1810_1, in1810_2);
    wire[0:0] s1811, in1811_1, in1811_2;
    wire c1811;
    assign in1811_1 = {c1730};
    assign in1811_2 = {c1731};
    Half_Adder KS_1811(s1811, c1811, in1811_1, in1811_2);
    wire[3:0] s1812, in1812_1, in1812_2;
    wire c1812;
    assign in1812_1 = {c1732,s82[1],s79[2],s86[3]};
    assign in1812_2 = {c1733,c83,s80[2],s88[1]};
    CLA_4 KS_1812(s1812, c1812, in1812_1, in1812_2);
    wire[0:0] s1813, in1813_1, in1813_2;
    wire c1813;
    assign in1813_1 = {c1734};
    assign in1813_2 = {c1735};
    Half_Adder KS_1813(s1813, c1813, in1813_1, in1813_2);
    wire[1:0] s1814, in1814_1, in1814_2;
    wire c1814;
    assign in1814_1 = {c1736,s84[1]};
    assign in1814_2 = {c1737,c85};
    CLA_2 KS_1814(s1814, c1814, in1814_1, in1814_2);
    wire[0:0] s1815, in1815_1, in1815_2;
    wire c1815;
    assign in1815_1 = {c1738};
    assign in1815_2 = {c1739};
    Half_Adder KS_1815(s1815, c1815, in1815_1, in1815_2);
    wire[2:0] s1816, in1816_1, in1816_2;
    wire c1816;
    assign in1816_1 = {c1740,s86[1],s82[2]};
    assign in1816_2 = {c1741,c87,s84[2]};
    CLA_3 KS_1816(s1816, c1816, in1816_1, in1816_2);
    wire[0:0] s1817, in1817_1, in1817_2;
    wire c1817;
    assign in1817_1 = {c1742};
    assign in1817_2 = {c1743};
    Half_Adder KS_1817(s1817, c1817, in1817_1, in1817_2);
    wire[1:0] s1818, in1818_1, in1818_2;
    wire c1818;
    assign in1818_1 = {c1744,s1773[1]};
    assign in1818_2 = {c1745,s1774[1]};
    CLA_2 KS_1818(s1818, c1818, in1818_1, in1818_2);
    wire[0:0] s1819, in1819_1, in1819_2;
    wire c1819;
    assign in1819_1 = {c1746};
    assign in1819_2 = {c1747};
    Half_Adder KS_1819(s1819, c1819, in1819_1, in1819_2);
    wire[3:0] s1820, in1820_1, in1820_2;
    wire c1820;
    assign in1820_1 = {c1748,s1775[1],s86[2],s89[1]};
    assign in1820_2 = {c1749,s1776[1],s88[0],s90[1]};
    CLA_4 KS_1820(s1820, c1820, in1820_1, in1820_2);
    wire[0:0] s1821, in1821_1, in1821_2;
    wire c1821;
    assign in1821_1 = {c1750};
    assign in1821_2 = {c1751};
    Half_Adder KS_1821(s1821, c1821, in1821_1, in1821_2);
    wire[1:0] s1822, in1822_1, in1822_2;
    wire c1822;
    assign in1822_1 = {c1752,s1777[1]};
    assign in1822_2 = {c1753,s1778[1]};
    CLA_2 KS_1822(s1822, c1822, in1822_1, in1822_2);
    wire[0:0] s1823, in1823_1, in1823_2;
    wire c1823;
    assign in1823_1 = {c1754};
    assign in1823_2 = {c1755};
    Half_Adder KS_1823(s1823, c1823, in1823_1, in1823_2);
    wire[2:0] s1824, in1824_1, in1824_2;
    wire c1824;
    assign in1824_1 = {c1756,s1779[1],s89[0]};
    assign in1824_2 = {c1757,s1780[1],s90[0]};
    CLA_3 KS_1824(s1824, c1824, in1824_1, in1824_2);
    wire[0:0] s1825, in1825_1, in1825_2;
    wire c1825;
    assign in1825_1 = {c1758};
    assign in1825_2 = {c1759};
    Half_Adder KS_1825(s1825, c1825, in1825_1, in1825_2);
    wire[1:0] s1826, in1826_1, in1826_2;
    wire c1826;
    assign in1826_1 = {c1760,s1781[1]};
    assign in1826_2 = {c1761,s1782[1]};
    CLA_2 KS_1826(s1826, c1826, in1826_1, in1826_2);
    wire[0:0] s1827, in1827_1, in1827_2;
    wire c1827;
    assign in1827_1 = {c1765};
    assign in1827_2 = {c1769};
    Half_Adder KS_1827(s1827, c1827, in1827_1, in1827_2);
    wire[3:0] s1828, in1828_1, in1828_2;
    wire c1828;
    assign in1828_1 = {s1773[0],s1783[1],s91[0],s91[1]};
    assign in1828_2 = {s1774[0],s1784[1],s92[0],s92[1]};
    CLA_4 KS_1828(s1828, c1828, in1828_1, in1828_2);
    wire[0:0] s1829, in1829_1, in1829_2;
    wire c1829;
    assign in1829_1 = {s1775[0]};
    assign in1829_2 = {s1776[0]};
    Half_Adder KS_1829(s1829, c1829, in1829_1, in1829_2);
    wire[1:0] s1830, in1830_1, in1830_2;
    wire c1830;
    assign in1830_1 = {s1777[0],s1785[1]};
    assign in1830_2 = {s1778[0],s1786[1]};
    CLA_2 KS_1830(s1830, c1830, in1830_1, in1830_2);
    wire[0:0] s1831, in1831_1, in1831_2;
    wire c1831;
    assign in1831_1 = {s1779[0]};
    assign in1831_2 = {s1780[0]};
    Half_Adder KS_1831(s1831, c1831, in1831_1, in1831_2);
    wire[2:0] s1832, in1832_1, in1832_2;
    wire c1832;
    assign in1832_1 = {s1781[0],s1787[1],s1773[2]};
    assign in1832_2 = {s1782[0],s1788[1],s1774[2]};
    CLA_3 KS_1832(s1832, c1832, in1832_1, in1832_2);
    wire[0:0] s1833, in1833_1, in1833_2;
    wire c1833;
    assign in1833_1 = {s1783[0]};
    assign in1833_2 = {s1784[0]};
    Half_Adder KS_1833(s1833, c1833, in1833_1, in1833_2);
    wire[1:0] s1834, in1834_1, in1834_2;
    wire c1834;
    assign in1834_1 = {s1785[0],s1789[1]};
    assign in1834_2 = {s1786[0],s1790[1]};
    CLA_2 KS_1834(s1834, c1834, in1834_1, in1834_2);
    wire[0:0] s1835, in1835_1, in1835_2;
    wire c1835;
    assign in1835_1 = {s1787[0]};
    assign in1835_2 = {s1788[0]};
    Half_Adder KS_1835(s1835, c1835, in1835_1, in1835_2);
    wire[3:0] s1836, in1836_1, in1836_2;
    wire c1836;
    assign in1836_1 = {s1790[0],s1791[1],s1775[2],s93[0]};
    assign in1836_2 = {s1791[0],s1792[1],s1776[2],s94[0]};
    CLA_4_c KS_1836(s1836, c1836, in1836_1, in1836_2, s1789[0]);
    wire[3:0] s1837, in1837_1, in1837_2;
    wire c1837;
    assign in1837_1 = {pp83[17],pp68[33],pp63[39],pp67[36]};
    assign in1837_2 = {pp84[16],pp69[32],pp64[38],pp68[35]};
    CLA_4 KS_1837(s1837, c1837, in1837_1, in1837_2);
    wire[3:0] s1838, in1838_1, in1838_2;
    wire c1838;
    assign in1838_1 = {pp85[15],pp70[31],pp65[37],pp69[34]};
    assign in1838_2 = {pp86[14],pp71[30],pp66[36],pp70[33]};
    CLA_4 KS_1838(s1838, c1838, in1838_1, in1838_2);
    wire[3:0] s1839, in1839_1, in1839_2;
    wire c1839;
    assign in1839_1 = {pp87[13],pp72[29],pp67[35],pp71[32]};
    assign in1839_2 = {pp88[12],pp73[28],pp68[34],pp72[31]};
    CLA_4 KS_1839(s1839, c1839, in1839_1, in1839_2);
    wire[3:0] s1840, in1840_1, in1840_2;
    wire c1840;
    assign in1840_1 = {pp89[11],pp74[27],pp69[33],pp73[30]};
    assign in1840_2 = {pp90[10],pp75[26],pp70[32],pp74[29]};
    CLA_4 KS_1840(s1840, c1840, in1840_1, in1840_2);
    wire[3:0] s1841, in1841_1, in1841_2;
    wire c1841;
    assign in1841_1 = {pp91[9],pp76[25],pp71[31],pp75[28]};
    assign in1841_2 = {pp92[8],pp77[24],pp72[30],pp76[27]};
    CLA_4 KS_1841(s1841, c1841, in1841_1, in1841_2);
    wire[3:0] s1842, in1842_1, in1842_2;
    wire c1842;
    assign in1842_1 = {pp93[7],pp78[23],pp73[29],pp77[26]};
    assign in1842_2 = {pp94[6],pp79[22],pp74[28],pp78[25]};
    CLA_4 KS_1842(s1842, c1842, in1842_1, in1842_2);
    wire[3:0] s1843, in1843_1, in1843_2;
    wire c1843;
    assign in1843_1 = {pp95[5],pp80[21],pp75[27],pp79[24]};
    assign in1843_2 = {pp96[4],pp81[20],pp76[26],pp80[23]};
    CLA_4 KS_1843(s1843, c1843, in1843_1, in1843_2);
    wire[3:0] s1844, in1844_1, in1844_2;
    wire c1844;
    assign in1844_1 = {pp97[3],pp82[19],pp77[25],pp81[22]};
    assign in1844_2 = {pp98[2],pp83[18],pp78[24],pp82[21]};
    CLA_4 KS_1844(s1844, c1844, in1844_1, in1844_2);
    wire[3:0] s1845, in1845_1, in1845_2;
    wire c1845;
    assign in1845_1 = {pp99[1],pp84[17],pp79[23],pp83[20]};
    assign in1845_2 = {pp100[0],pp85[16],pp80[22],pp84[19]};
    CLA_4 KS_1845(s1845, c1845, in1845_1, in1845_2);
    wire[3:0] s1846, in1846_1, in1846_2;
    wire c1846;
    assign in1846_1 = {c67,pp86[15],pp81[21],pp85[18]};
    assign in1846_2 = {c68,pp87[14],pp82[20],pp86[17]};
    CLA_4 KS_1846(s1846, c1846, in1846_1, in1846_2);
    wire[3:0] s1847, in1847_1, in1847_2;
    wire c1847;
    assign in1847_1 = {c69,pp88[13],pp83[19],pp87[16]};
    assign in1847_2 = {c70,pp89[12],pp84[18],pp88[15]};
    CLA_4 KS_1847(s1847, c1847, in1847_1, in1847_2);
    wire[3:0] s1848, in1848_1, in1848_2;
    wire c1848;
    assign in1848_1 = {c71,pp90[11],pp85[17],pp89[14]};
    assign in1848_2 = {c72,pp91[10],pp86[16],pp90[13]};
    CLA_4 KS_1848(s1848, c1848, in1848_1, in1848_2);
    wire[3:0] s1849, in1849_1, in1849_2;
    wire c1849;
    assign in1849_1 = {c73,pp92[9],pp87[15],pp91[12]};
    assign in1849_2 = {c74,pp93[8],pp88[14],pp92[11]};
    CLA_4 KS_1849(s1849, c1849, in1849_1, in1849_2);
    wire[3:0] s1850, in1850_1, in1850_2;
    wire c1850;
    assign in1850_1 = {c75,pp94[7],pp89[13],pp93[10]};
    assign in1850_2 = {c76,pp95[6],pp90[12],pp94[9]};
    CLA_4 KS_1850(s1850, c1850, in1850_1, in1850_2);
    wire[3:0] s1851, in1851_1, in1851_2;
    wire c1851;
    assign in1851_1 = {c77,pp96[5],pp91[11],pp95[8]};
    assign in1851_2 = {c78,pp97[4],pp92[10],pp96[7]};
    CLA_4 KS_1851(s1851, c1851, in1851_1, in1851_2);
    wire[3:0] s1852, in1852_1, in1852_2;
    wire c1852;
    assign in1852_1 = {c79,pp98[3],pp93[9],pp97[6]};
    assign in1852_2 = {c80,pp99[2],pp94[8],pp98[5]};
    CLA_4 KS_1852(s1852, c1852, in1852_1, in1852_2);
    wire[3:0] s1853, in1853_1, in1853_2;
    wire c1853;
    assign in1853_1 = {c82,pp100[1],pp95[7],pp99[4]};
    assign in1853_2 = {c84,pp101[0],pp96[6],pp100[3]};
    CLA_4 KS_1853(s1853, c1853, in1853_1, in1853_2);
    wire[3:0] s1854, in1854_1, in1854_2;
    wire c1854;
    assign in1854_1 = {c86,s88[3],pp97[5],pp101[2]};
    assign in1854_2 = {s88[2],s89[3],pp98[4],pp102[1]};
    CLA_4 KS_1854(s1854, c1854, in1854_1, in1854_2);
    wire[3:0] s1855, in1855_1, in1855_2;
    wire c1855;
    assign in1855_1 = {s89[2],s90[3],pp99[3],pp103[0]};
    assign in1855_2 = {s90[2],s91[3],pp100[2],c93};
    CLA_4 KS_1855(s1855, c1855, in1855_1, in1855_2);
    wire[3:0] s1856, in1856_1, in1856_2;
    wire c1856;
    assign in1856_1 = {s91[2],s92[3],pp101[1],c94};
    assign in1856_2 = {s92[2],s93[2],pp102[0],c95};
    CLA_4 KS_1856(s1856, c1856, in1856_1, in1856_2);
    wire[3:0] s1857, in1857_1, in1857_2;
    wire c1857;
    assign in1857_1 = {s93[1],s94[2],c88,c96};
    assign in1857_2 = {s94[1],s95[2],c89,c97};
    CLA_4 KS_1857(s1857, c1857, in1857_1, in1857_2);
    wire[3:0] s1858, in1858_1, in1858_2;
    wire c1858;
    assign in1858_1 = {s95[1],s96[2],c90,c98};
    assign in1858_2 = {s96[1],s97[2],c91,s99[3]};
    CLA_4 KS_1858(s1858, c1858, in1858_1, in1858_2);
    wire[3:0] s1859, in1859_1, in1859_2;
    wire c1859;
    assign in1859_1 = {s97[1],s98[2],c92,s100[3]};
    assign in1859_2 = {s98[1],s99[1],s93[3],s101[3]};
    CLA_4 KS_1859(s1859, c1859, in1859_1, in1859_2);
    wire[3:0] s1860, in1860_1, in1860_2;
    wire c1860;
    assign in1860_1 = {s99[0],s100[1],s94[3],s102[3]};
    assign in1860_2 = {s100[0],s101[1],s95[3],s103[3]};
    CLA_4 KS_1860(s1860, c1860, in1860_1, in1860_2);
    wire[3:0] s1861, in1861_1, in1861_2;
    wire c1861;
    assign in1861_1 = {s101[0],s102[1],s96[3],s104[3]};
    assign in1861_2 = {s102[0],s103[1],s97[3],s105[3]};
    CLA_4 KS_1861(s1861, c1861, in1861_1, in1861_2);
    wire[3:0] s1862, in1862_1, in1862_2;
    wire c1862;
    assign in1862_1 = {s103[0],s104[1],s98[3],s106[3]};
    assign in1862_2 = {s104[0],s105[1],s99[2],s107[3]};
    CLA_4 KS_1862(s1862, c1862, in1862_1, in1862_2);
    wire[3:0] s1863, in1863_1, in1863_2;
    wire c1863;
    assign in1863_1 = {s105[0],s106[1],s100[2],s108[3]};
    assign in1863_2 = {s106[0],s107[1],s101[2],s109[3]};
    CLA_4 KS_1863(s1863, c1863, in1863_1, in1863_2);
    wire[3:0] s1864, in1864_1, in1864_2;
    wire c1864;
    assign in1864_1 = {s107[0],s108[1],s102[2],s110[3]};
    assign in1864_2 = {s108[0],s109[1],s103[2],s111[3]};
    CLA_4 KS_1864(s1864, c1864, in1864_1, in1864_2);
    wire[3:0] s1865, in1865_1, in1865_2;
    wire c1865;
    assign in1865_1 = {s109[0],s110[1],s104[2],s112[3]};
    assign in1865_2 = {s110[0],s111[1],s105[2],s113[3]};
    CLA_4 KS_1865(s1865, c1865, in1865_1, in1865_2);
    wire[3:0] s1866, in1866_1, in1866_2;
    wire c1866;
    assign in1866_1 = {s111[0],s112[1],s106[2],s114[3]};
    assign in1866_2 = {s112[0],s113[1],s107[2],s116[3]};
    CLA_4 KS_1866(s1866, c1866, in1866_1, in1866_2);
    wire[3:0] s1867, in1867_1, in1867_2;
    wire c1867;
    assign in1867_1 = {s113[0],s114[1],s108[2],s118[3]};
    assign in1867_2 = {s114[0],c115,s109[2],s120[3]};
    CLA_4 KS_1867(s1867, c1867, in1867_1, in1867_2);
    wire[0:0] s1868, in1868_1, in1868_2;
    wire c1868;
    assign in1868_1 = {s115[0]};
    assign in1868_2 = {s116[0]};
    Half_Adder KS_1868(s1868, c1868, in1868_1, in1868_2);
    wire[3:0] s1869, in1869_1, in1869_2;
    wire c1869;
    assign in1869_1 = {s117[0],s116[1],s110[2],s122[3]};
    assign in1869_2 = {s118[0],c117,s111[2],s124[3]};
    CLA_4 KS_1869(s1869, c1869, in1869_1, in1869_2);
    wire[0:0] s1870, in1870_1, in1870_2;
    wire c1870;
    assign in1870_1 = {s119[0]};
    assign in1870_2 = {s120[0]};
    Half_Adder KS_1870(s1870, c1870, in1870_1, in1870_2);
    wire[1:0] s1871, in1871_1, in1871_2;
    wire c1871;
    assign in1871_1 = {s121[0],s118[1]};
    assign in1871_2 = {s122[0],c119};
    CLA_2 KS_1871(s1871, c1871, in1871_1, in1871_2);
    wire[0:0] s1872, in1872_1, in1872_2;
    wire c1872;
    assign in1872_1 = {s123[0]};
    assign in1872_2 = {s124[0]};
    Half_Adder KS_1872(s1872, c1872, in1872_1, in1872_2);
    wire[2:0] s1873, in1873_1, in1873_2;
    wire c1873;
    assign in1873_1 = {s125[0],s120[1],s112[2]};
    assign in1873_2 = {s126[0],c121,s113[2]};
    CLA_3 KS_1873(s1873, c1873, in1873_1, in1873_2);
    wire[0:0] s1874, in1874_1, in1874_2;
    wire c1874;
    assign in1874_1 = {s127[0]};
    assign in1874_2 = {s128[0]};
    Half_Adder KS_1874(s1874, c1874, in1874_1, in1874_2);
    wire[1:0] s1875, in1875_1, in1875_2;
    wire c1875;
    assign in1875_1 = {c1773,s122[1]};
    assign in1875_2 = {c1774,c123};
    CLA_2 KS_1875(s1875, c1875, in1875_1, in1875_2);
    wire[0:0] s1876, in1876_1, in1876_2;
    wire c1876;
    assign in1876_1 = {c1775};
    assign in1876_2 = {c1776};
    Half_Adder KS_1876(s1876, c1876, in1876_1, in1876_2);
    wire[3:0] s1877, in1877_1, in1877_2;
    wire c1877;
    assign in1877_1 = {c1777,s124[1],s114[2],s126[3]};
    assign in1877_2 = {c1778,c125,s116[2],s128[3]};
    CLA_4 KS_1877(s1877, c1877, in1877_1, in1877_2);
    wire[0:0] s1878, in1878_1, in1878_2;
    wire c1878;
    assign in1878_1 = {c1779};
    assign in1878_2 = {c1780};
    Half_Adder KS_1878(s1878, c1878, in1878_1, in1878_2);
    wire[1:0] s1879, in1879_1, in1879_2;
    wire c1879;
    assign in1879_1 = {c1781,s126[1]};
    assign in1879_2 = {c1782,c127};
    CLA_2 KS_1879(s1879, c1879, in1879_1, in1879_2);
    wire[0:0] s1880, in1880_1, in1880_2;
    wire c1880;
    assign in1880_1 = {c1783};
    assign in1880_2 = {c1784};
    Half_Adder KS_1880(s1880, c1880, in1880_1, in1880_2);
    wire[2:0] s1881, in1881_1, in1881_2;
    wire c1881;
    assign in1881_1 = {c1785,s128[1],s118[2]};
    assign in1881_2 = {c1786,s1837[1],s120[2]};
    CLA_3 KS_1881(s1881, c1881, in1881_1, in1881_2);
    wire[0:0] s1882, in1882_1, in1882_2;
    wire c1882;
    assign in1882_1 = {c1787};
    assign in1882_2 = {c1788};
    Half_Adder KS_1882(s1882, c1882, in1882_1, in1882_2);
    wire[1:0] s1883, in1883_1, in1883_2;
    wire c1883;
    assign in1883_1 = {c1789,s1838[1]};
    assign in1883_2 = {c1790,s1839[1]};
    CLA_2 KS_1883(s1883, c1883, in1883_1, in1883_2);
    wire[0:0] s1884, in1884_1, in1884_2;
    wire c1884;
    assign in1884_1 = {c1791};
    assign in1884_2 = {c1792};
    Half_Adder KS_1884(s1884, c1884, in1884_1, in1884_2);
    wire[3:0] s1885, in1885_1, in1885_2;
    wire c1885;
    assign in1885_1 = {c1793,s1840[1],s122[2],s129[1]};
    assign in1885_2 = {c1794,s1841[1],s124[2],s130[1]};
    CLA_4 KS_1885(s1885, c1885, in1885_1, in1885_2);
    wire[0:0] s1886, in1886_1, in1886_2;
    wire c1886;
    assign in1886_1 = {c1795};
    assign in1886_2 = {c1796};
    Half_Adder KS_1886(s1886, c1886, in1886_1, in1886_2);
    wire[1:0] s1887, in1887_1, in1887_2;
    wire c1887;
    assign in1887_1 = {c1797,s1842[1]};
    assign in1887_2 = {c1798,s1843[1]};
    CLA_2 KS_1887(s1887, c1887, in1887_1, in1887_2);
    wire[0:0] s1888, in1888_1, in1888_2;
    wire c1888;
    assign in1888_1 = {c1799};
    assign in1888_2 = {c1800};
    Half_Adder KS_1888(s1888, c1888, in1888_1, in1888_2);
    wire[2:0] s1889, in1889_1, in1889_2;
    wire c1889;
    assign in1889_1 = {c1801,s1844[1],s126[2]};
    assign in1889_2 = {c1802,s1845[1],s128[2]};
    CLA_3 KS_1889(s1889, c1889, in1889_1, in1889_2);
    wire[0:0] s1890, in1890_1, in1890_2;
    wire c1890;
    assign in1890_1 = {c1803};
    assign in1890_2 = {c1804};
    Half_Adder KS_1890(s1890, c1890, in1890_1, in1890_2);
    wire[1:0] s1891, in1891_1, in1891_2;
    wire c1891;
    assign in1891_1 = {c1812,s1846[1]};
    assign in1891_2 = {c1820,s1847[1]};
    CLA_2 KS_1891(s1891, c1891, in1891_1, in1891_2);
    wire[0:0] s1892, in1892_1, in1892_2;
    wire c1892;
    assign in1892_1 = {c1828};
    assign in1892_2 = {c1836};
    Half_Adder KS_1892(s1892, c1892, in1892_1, in1892_2);
    wire[3:0] s1893, in1893_1, in1893_2;
    wire c1893;
    assign in1893_1 = {s1837[0],s1848[1],s129[0],s131[0]};
    assign in1893_2 = {s1838[0],s1849[1],s130[0],s132[0]};
    CLA_4 KS_1893(s1893, c1893, in1893_1, in1893_2);
    wire[0:0] s1894, in1894_1, in1894_2;
    wire c1894;
    assign in1894_1 = {s1839[0]};
    assign in1894_2 = {s1840[0]};
    Half_Adder KS_1894(s1894, c1894, in1894_1, in1894_2);
    wire[1:0] s1895, in1895_1, in1895_2;
    wire c1895;
    assign in1895_1 = {s1841[0],s1850[1]};
    assign in1895_2 = {s1842[0],s1851[1]};
    CLA_2 KS_1895(s1895, c1895, in1895_1, in1895_2);
    wire[0:0] s1896, in1896_1, in1896_2;
    wire c1896;
    assign in1896_1 = {s1843[0]};
    assign in1896_2 = {s1844[0]};
    Half_Adder KS_1896(s1896, c1896, in1896_1, in1896_2);
    wire[2:0] s1897, in1897_1, in1897_2;
    wire c1897;
    assign in1897_1 = {s1845[0],s1852[1],s1837[2]};
    assign in1897_2 = {s1846[0],s1853[1],s1838[2]};
    CLA_3 KS_1897(s1897, c1897, in1897_1, in1897_2);
    wire[0:0] s1898, in1898_1, in1898_2;
    wire c1898;
    assign in1898_1 = {s1847[0]};
    assign in1898_2 = {s1848[0]};
    Half_Adder KS_1898(s1898, c1898, in1898_1, in1898_2);
    wire[1:0] s1899, in1899_1, in1899_2;
    wire c1899;
    assign in1899_1 = {s1849[0],s1854[1]};
    assign in1899_2 = {s1850[0],s1855[1]};
    CLA_2 KS_1899(s1899, c1899, in1899_1, in1899_2);
    wire[0:0] s1900, in1900_1, in1900_2;
    wire c1900;
    assign in1900_1 = {s1851[0]};
    assign in1900_2 = {s1852[0]};
    Half_Adder KS_1900(s1900, c1900, in1900_1, in1900_2);
    wire[3:0] s1901, in1901_1, in1901_2;
    wire c1901;
    assign in1901_1 = {s1853[0],s1856[1],s1839[2],s133[0]};
    assign in1901_2 = {s1854[0],s1857[1],s1840[2],s134[0]};
    CLA_4 KS_1901(s1901, c1901, in1901_1, in1901_2);
    wire[0:0] s1902, in1902_1, in1902_2;
    wire c1902;
    assign in1902_1 = {s1856[0]};
    assign in1902_2 = {s1857[0]};
    Full_Adder KS_1902(s1902, c1902, in1902_1, in1902_2, s1855[0]);
    wire[3:0] s1903, in1903_1, in1903_2;
    wire c1903;
    assign in1903_1 = {pp103[1],pp82[23],pp72[34],pp79[28]};
    assign in1903_2 = {pp104[0],pp83[22],pp73[33],pp80[27]};
    CLA_4 KS_1903(s1903, c1903, in1903_1, in1903_2);
    wire[3:0] s1904, in1904_1, in1904_2;
    wire c1904;
    assign in1904_1 = {c99,pp84[21],pp74[32],pp81[26]};
    assign in1904_2 = {c100,pp85[20],pp75[31],pp82[25]};
    CLA_4 KS_1904(s1904, c1904, in1904_1, in1904_2);
    wire[3:0] s1905, in1905_1, in1905_2;
    wire c1905;
    assign in1905_1 = {c101,pp86[19],pp76[30],pp83[24]};
    assign in1905_2 = {c102,pp87[18],pp77[29],pp84[23]};
    CLA_4 KS_1905(s1905, c1905, in1905_1, in1905_2);
    wire[3:0] s1906, in1906_1, in1906_2;
    wire c1906;
    assign in1906_1 = {c103,pp88[17],pp78[28],pp85[22]};
    assign in1906_2 = {c104,pp89[16],pp79[27],pp86[21]};
    CLA_4 KS_1906(s1906, c1906, in1906_1, in1906_2);
    wire[3:0] s1907, in1907_1, in1907_2;
    wire c1907;
    assign in1907_1 = {c105,pp90[15],pp80[26],pp87[20]};
    assign in1907_2 = {c106,pp91[14],pp81[25],pp88[19]};
    CLA_4 KS_1907(s1907, c1907, in1907_1, in1907_2);
    wire[3:0] s1908, in1908_1, in1908_2;
    wire c1908;
    assign in1908_1 = {c107,pp92[13],pp82[24],pp89[18]};
    assign in1908_2 = {c108,pp93[12],pp83[23],pp90[17]};
    CLA_4 KS_1908(s1908, c1908, in1908_1, in1908_2);
    wire[3:0] s1909, in1909_1, in1909_2;
    wire c1909;
    assign in1909_1 = {c109,pp94[11],pp84[22],pp91[16]};
    assign in1909_2 = {c110,pp95[10],pp85[21],pp92[15]};
    CLA_4 KS_1909(s1909, c1909, in1909_1, in1909_2);
    wire[3:0] s1910, in1910_1, in1910_2;
    wire c1910;
    assign in1910_1 = {c111,pp96[9],pp86[20],pp93[14]};
    assign in1910_2 = {c112,pp97[8],pp87[19],pp94[13]};
    CLA_4 KS_1910(s1910, c1910, in1910_1, in1910_2);
    wire[3:0] s1911, in1911_1, in1911_2;
    wire c1911;
    assign in1911_1 = {c113,pp98[7],pp88[18],pp95[12]};
    assign in1911_2 = {c114,pp99[6],pp89[17],pp96[11]};
    CLA_4 KS_1911(s1911, c1911, in1911_1, in1911_2);
    wire[3:0] s1912, in1912_1, in1912_2;
    wire c1912;
    assign in1912_1 = {c116,pp100[5],pp90[16],pp97[10]};
    assign in1912_2 = {c118,pp101[4],pp91[15],pp98[9]};
    CLA_4 KS_1912(s1912, c1912, in1912_1, in1912_2);
    wire[3:0] s1913, in1913_1, in1913_2;
    wire c1913;
    assign in1913_1 = {c120,pp102[3],pp92[14],pp99[8]};
    assign in1913_2 = {c122,pp103[2],pp93[13],pp100[7]};
    CLA_4 KS_1913(s1913, c1913, in1913_1, in1913_2);
    wire[3:0] s1914, in1914_1, in1914_2;
    wire c1914;
    assign in1914_1 = {c124,pp104[1],pp94[12],pp101[6]};
    assign in1914_2 = {c126,pp105[0],pp95[11],pp102[5]};
    CLA_4 KS_1914(s1914, c1914, in1914_1, in1914_2);
    wire[3:0] s1915, in1915_1, in1915_2;
    wire c1915;
    assign in1915_1 = {c128,s129[3],pp96[10],pp103[4]};
    assign in1915_2 = {s129[2],s130[3],pp97[9],pp104[3]};
    CLA_4 KS_1915(s1915, c1915, in1915_1, in1915_2);
    wire[3:0] s1916, in1916_1, in1916_2;
    wire c1916;
    assign in1916_1 = {s130[2],s131[2],pp98[8],pp105[2]};
    assign in1916_2 = {s131[1],s132[2],pp99[7],pp106[1]};
    CLA_4 KS_1916(s1916, c1916, in1916_1, in1916_2);
    wire[3:0] s1917, in1917_1, in1917_2;
    wire c1917;
    assign in1917_1 = {s132[1],s133[2],pp100[6],pp107[0]};
    assign in1917_2 = {s133[1],s134[2],pp101[5],c131};
    CLA_4 KS_1917(s1917, c1917, in1917_1, in1917_2);
    wire[3:0] s1918, in1918_1, in1918_2;
    wire c1918;
    assign in1918_1 = {s134[1],s135[2],pp102[4],c132};
    assign in1918_2 = {s135[1],s136[2],pp103[3],c133};
    CLA_4 KS_1918(s1918, c1918, in1918_1, in1918_2);
    wire[3:0] s1919, in1919_1, in1919_2;
    wire c1919;
    assign in1919_1 = {s136[1],s137[2],pp104[2],c134};
    assign in1919_2 = {s137[1],s138[2],pp105[1],c135};
    CLA_4 KS_1919(s1919, c1919, in1919_1, in1919_2);
    wire[3:0] s1920, in1920_1, in1920_2;
    wire c1920;
    assign in1920_1 = {s138[1],s139[1],pp106[0],c136};
    assign in1920_2 = {s139[0],s140[1],c129,c137};
    CLA_4 KS_1920(s1920, c1920, in1920_1, in1920_2);
    wire[3:0] s1921, in1921_1, in1921_2;
    wire c1921;
    assign in1921_1 = {s140[0],s141[1],c130,c138};
    assign in1921_2 = {s141[0],s142[1],s131[3],s139[3]};
    CLA_4 KS_1921(s1921, c1921, in1921_1, in1921_2);
    wire[3:0] s1922, in1922_1, in1922_2;
    wire c1922;
    assign in1922_1 = {s142[0],s143[1],s132[3],s140[3]};
    assign in1922_2 = {s143[0],s144[1],s133[3],s141[3]};
    CLA_4 KS_1922(s1922, c1922, in1922_1, in1922_2);
    wire[3:0] s1923, in1923_1, in1923_2;
    wire c1923;
    assign in1923_1 = {s144[0],s145[1],s134[3],s142[3]};
    assign in1923_2 = {s145[0],s146[1],s135[3],s143[3]};
    CLA_4 KS_1923(s1923, c1923, in1923_1, in1923_2);
    wire[3:0] s1924, in1924_1, in1924_2;
    wire c1924;
    assign in1924_1 = {s146[0],s147[1],s136[3],s144[3]};
    assign in1924_2 = {s147[0],s148[1],s137[3],s145[3]};
    CLA_4 KS_1924(s1924, c1924, in1924_1, in1924_2);
    wire[3:0] s1925, in1925_1, in1925_2;
    wire c1925;
    assign in1925_1 = {s148[0],s149[1],s138[3],s146[3]};
    assign in1925_2 = {s149[0],s150[1],s139[2],s147[3]};
    CLA_4 KS_1925(s1925, c1925, in1925_1, in1925_2);
    wire[3:0] s1926, in1926_1, in1926_2;
    wire c1926;
    assign in1926_1 = {s150[0],s151[1],s140[2],s148[3]};
    assign in1926_2 = {s151[0],s152[1],s141[2],s149[3]};
    CLA_4 KS_1926(s1926, c1926, in1926_1, in1926_2);
    wire[3:0] s1927, in1927_1, in1927_2;
    wire c1927;
    assign in1927_1 = {s152[0],s153[1],s142[2],s150[3]};
    assign in1927_2 = {s153[0],s154[1],s143[2],s151[3]};
    CLA_4 KS_1927(s1927, c1927, in1927_1, in1927_2);
    wire[3:0] s1928, in1928_1, in1928_2;
    wire c1928;
    assign in1928_1 = {s154[0],s155[1],s144[2],s152[3]};
    assign in1928_2 = {s155[0],s156[1],s145[2],s153[3]};
    CLA_4 KS_1928(s1928, c1928, in1928_1, in1928_2);
    wire[3:0] s1929, in1929_1, in1929_2;
    wire c1929;
    assign in1929_1 = {s156[0],s157[1],s146[2],s154[3]};
    assign in1929_2 = {s157[0],s158[1],s147[2],s155[3]};
    CLA_4 KS_1929(s1929, c1929, in1929_1, in1929_2);
    wire[3:0] s1930, in1930_1, in1930_2;
    wire c1930;
    assign in1930_1 = {s158[0],s159[1],s148[2],s156[3]};
    assign in1930_2 = {s159[0],c160,s149[2],s157[3]};
    CLA_4 KS_1930(s1930, c1930, in1930_1, in1930_2);
    wire[3:0] s1931, in1931_1, in1931_2;
    wire c1931;
    assign in1931_1 = {s160[0],s161[1],s150[2],s158[3]};
    assign in1931_2 = {s161[0],c162,s151[2],s159[3]};
    CLA_4 KS_1931(s1931, c1931, in1931_1, in1931_2);
    wire[3:0] s1932, in1932_1, in1932_2;
    wire c1932;
    assign in1932_1 = {s162[0],s163[1],s152[2],s161[3]};
    assign in1932_2 = {s163[0],c164,s153[2],s163[3]};
    CLA_4 KS_1932(s1932, c1932, in1932_1, in1932_2);
    wire[3:0] s1933, in1933_1, in1933_2;
    wire c1933;
    assign in1933_1 = {s164[0],s165[1],s154[2],s165[3]};
    assign in1933_2 = {s165[0],c166,s155[2],s167[3]};
    CLA_4 KS_1933(s1933, c1933, in1933_1, in1933_2);
    wire[0:0] s1934, in1934_1, in1934_2;
    wire c1934;
    assign in1934_1 = {s166[0]};
    assign in1934_2 = {s167[0]};
    Half_Adder KS_1934(s1934, c1934, in1934_1, in1934_2);
    wire[3:0] s1935, in1935_1, in1935_2;
    wire c1935;
    assign in1935_1 = {s168[0],s167[1],s156[2],s169[3]};
    assign in1935_2 = {s169[0],c168,s157[2],s173[3]};
    CLA_4 KS_1935(s1935, c1935, in1935_1, in1935_2);
    wire[0:0] s1936, in1936_1, in1936_2;
    wire c1936;
    assign in1936_1 = {s170[0]};
    assign in1936_2 = {s171[0]};
    Half_Adder KS_1936(s1936, c1936, in1936_1, in1936_2);
    wire[1:0] s1937, in1937_1, in1937_2;
    wire c1937;
    assign in1937_1 = {s172[0],s169[1]};
    assign in1937_2 = {s173[0],c170};
    CLA_2 KS_1937(s1937, c1937, in1937_1, in1937_2);
    wire[0:0] s1938, in1938_1, in1938_2;
    wire c1938;
    assign in1938_1 = {s174[0]};
    assign in1938_2 = {s175[0]};
    Half_Adder KS_1938(s1938, c1938, in1938_1, in1938_2);
    wire[2:0] s1939, in1939_1, in1939_2;
    wire c1939;
    assign in1939_1 = {s176[0],s171[1],s158[2]};
    assign in1939_2 = {s177[0],c172,s159[2]};
    CLA_3 KS_1939(s1939, c1939, in1939_1, in1939_2);
    wire[0:0] s1940, in1940_1, in1940_2;
    wire c1940;
    assign in1940_1 = {s178[0]};
    assign in1940_2 = {s179[0]};
    Half_Adder KS_1940(s1940, c1940, in1940_1, in1940_2);
    wire[1:0] s1941, in1941_1, in1941_2;
    wire c1941;
    assign in1941_1 = {c1837,s173[1]};
    assign in1941_2 = {c1838,c174};
    CLA_2 KS_1941(s1941, c1941, in1941_1, in1941_2);
    wire[0:0] s1942, in1942_1, in1942_2;
    wire c1942;
    assign in1942_1 = {c1839};
    assign in1942_2 = {c1840};
    Half_Adder KS_1942(s1942, c1942, in1942_1, in1942_2);
    wire[3:0] s1943, in1943_1, in1943_2;
    wire c1943;
    assign in1943_1 = {c1841,s175[1],s161[2],s177[3]};
    assign in1943_2 = {c1842,c176,s163[2],s180[0]};
    CLA_4 KS_1943(s1943, c1943, in1943_1, in1943_2);
    wire[0:0] s1944, in1944_1, in1944_2;
    wire c1944;
    assign in1944_1 = {c1843};
    assign in1944_2 = {c1844};
    Half_Adder KS_1944(s1944, c1944, in1944_1, in1944_2);
    wire[1:0] s1945, in1945_1, in1945_2;
    wire c1945;
    assign in1945_1 = {c1845,s177[1]};
    assign in1945_2 = {c1846,c178};
    CLA_2 KS_1945(s1945, c1945, in1945_1, in1945_2);
    wire[0:0] s1946, in1946_1, in1946_2;
    wire c1946;
    assign in1946_1 = {c1847};
    assign in1946_2 = {c1848};
    Half_Adder KS_1946(s1946, c1946, in1946_1, in1946_2);
    wire[2:0] s1947, in1947_1, in1947_2;
    wire c1947;
    assign in1947_1 = {c1849,s179[1],s165[2]};
    assign in1947_2 = {c1850,s1903[1],s167[2]};
    CLA_3 KS_1947(s1947, c1947, in1947_1, in1947_2);
    wire[0:0] s1948, in1948_1, in1948_2;
    wire c1948;
    assign in1948_1 = {c1851};
    assign in1948_2 = {c1852};
    Half_Adder KS_1948(s1948, c1948, in1948_1, in1948_2);
    wire[1:0] s1949, in1949_1, in1949_2;
    wire c1949;
    assign in1949_1 = {c1853,s1904[1]};
    assign in1949_2 = {c1854,s1905[1]};
    CLA_2 KS_1949(s1949, c1949, in1949_1, in1949_2);
    wire[0:0] s1950, in1950_1, in1950_2;
    wire c1950;
    assign in1950_1 = {c1855};
    assign in1950_2 = {c1856};
    Half_Adder KS_1950(s1950, c1950, in1950_1, in1950_2);
    wire[3:0] s1951, in1951_1, in1951_2;
    wire c1951;
    assign in1951_1 = {c1857,s1906[1],s169[2],s181[0]};
    assign in1951_2 = {c1858,s1907[1],c171,s182[0]};
    CLA_4 KS_1951(s1951, c1951, in1951_1, in1951_2);
    wire[0:0] s1952, in1952_1, in1952_2;
    wire c1952;
    assign in1952_1 = {c1859};
    assign in1952_2 = {c1860};
    Half_Adder KS_1952(s1952, c1952, in1952_1, in1952_2);
    wire[1:0] s1953, in1953_1, in1953_2;
    wire c1953;
    assign in1953_1 = {c1861,s1908[1]};
    assign in1953_2 = {c1862,s1909[1]};
    CLA_2 KS_1953(s1953, c1953, in1953_1, in1953_2);
    wire[0:0] s1954, in1954_1, in1954_2;
    wire c1954;
    assign in1954_1 = {c1863};
    assign in1954_2 = {c1864};
    Half_Adder KS_1954(s1954, c1954, in1954_1, in1954_2);
    wire[2:0] s1955, in1955_1, in1955_2;
    wire c1955;
    assign in1955_1 = {c1865,s1910[1],s173[2]};
    assign in1955_2 = {c1866,s1911[1],c175};
    CLA_3 KS_1955(s1955, c1955, in1955_1, in1955_2);
    wire[0:0] s1956, in1956_1, in1956_2;
    wire c1956;
    assign in1956_1 = {c1867};
    assign in1956_2 = {c1869};
    Half_Adder KS_1956(s1956, c1956, in1956_1, in1956_2);
    wire[1:0] s1957, in1957_1, in1957_2;
    wire c1957;
    assign in1957_1 = {c1877,s1912[1]};
    assign in1957_2 = {c1885,s1913[1]};
    CLA_2 KS_1957(s1957, c1957, in1957_1, in1957_2);
    wire[0:0] s1958, in1958_1, in1958_2;
    wire c1958;
    assign in1958_1 = {c1893};
    assign in1958_2 = {c1901};
    Half_Adder KS_1958(s1958, c1958, in1958_1, in1958_2);
    wire[3:0] s1959, in1959_1, in1959_2;
    wire c1959;
    assign in1959_1 = {s1903[0],s1914[1],s177[2],s183[0]};
    assign in1959_2 = {s1904[0],s1915[1],c179,s184[0]};
    CLA_4 KS_1959(s1959, c1959, in1959_1, in1959_2);
    wire[0:0] s1960, in1960_1, in1960_2;
    wire c1960;
    assign in1960_1 = {s1905[0]};
    assign in1960_2 = {s1906[0]};
    Half_Adder KS_1960(s1960, c1960, in1960_1, in1960_2);
    wire[1:0] s1961, in1961_1, in1961_2;
    wire c1961;
    assign in1961_1 = {s1907[0],s1916[1]};
    assign in1961_2 = {s1908[0],s1917[1]};
    CLA_2 KS_1961(s1961, c1961, in1961_1, in1961_2);
    wire[0:0] s1962, in1962_1, in1962_2;
    wire c1962;
    assign in1962_1 = {s1909[0]};
    assign in1962_2 = {s1910[0]};
    Half_Adder KS_1962(s1962, c1962, in1962_1, in1962_2);
    wire[2:0] s1963, in1963_1, in1963_2;
    wire c1963;
    assign in1963_1 = {s1911[0],s1918[1],s1903[2]};
    assign in1963_2 = {s1912[0],s1919[1],s1904[2]};
    CLA_3 KS_1963(s1963, c1963, in1963_1, in1963_2);
    wire[0:0] s1964, in1964_1, in1964_2;
    wire c1964;
    assign in1964_1 = {s1913[0]};
    assign in1964_2 = {s1914[0]};
    Half_Adder KS_1964(s1964, c1964, in1964_1, in1964_2);
    wire[1:0] s1965, in1965_1, in1965_2;
    wire c1965;
    assign in1965_1 = {s1915[0],s1920[1]};
    assign in1965_2 = {s1916[0],s1921[1]};
    CLA_2 KS_1965(s1965, c1965, in1965_1, in1965_2);
    wire[0:0] s1966, in1966_1, in1966_2;
    wire c1966;
    assign in1966_1 = {s1917[0]};
    assign in1966_2 = {s1918[0]};
    Half_Adder KS_1966(s1966, c1966, in1966_1, in1966_2);
    wire[3:0] s1967, in1967_1, in1967_2;
    wire c1967;
    assign in1967_1 = {s1919[0],s1922[1],s1905[2],s185[0]};
    assign in1967_2 = {s1920[0],s1923[1],s1906[2],s186[0]};
    CLA_4 KS_1967(s1967, c1967, in1967_1, in1967_2);
    wire[0:0] s1968, in1968_1, in1968_2;
    wire c1968;
    assign in1968_1 = {s1922[0]};
    assign in1968_2 = {s1923[0]};
    Full_Adder KS_1968(s1968, c1968, in1968_1, in1968_2, s1921[0]);
    wire[3:0] s1969, in1969_1, in1969_2;
    wire c1969;
    assign in1969_1 = {c151,pp94[15],pp82[28],pp93[18]};
    assign in1969_2 = {c152,pp95[14],pp83[27],pp94[17]};
    CLA_4 KS_1969(s1969, c1969, in1969_1, in1969_2);
    wire[3:0] s1970, in1970_1, in1970_2;
    wire c1970;
    assign in1970_1 = {c153,pp96[13],pp84[26],pp95[16]};
    assign in1970_2 = {c154,pp97[12],pp85[25],pp96[15]};
    CLA_4 KS_1970(s1970, c1970, in1970_1, in1970_2);
    wire[3:0] s1971, in1971_1, in1971_2;
    wire c1971;
    assign in1971_1 = {c155,pp98[11],pp86[24],pp97[14]};
    assign in1971_2 = {c156,pp99[10],pp87[23],pp98[13]};
    CLA_4 KS_1971(s1971, c1971, in1971_1, in1971_2);
    wire[3:0] s1972, in1972_1, in1972_2;
    wire c1972;
    assign in1972_1 = {c157,pp100[9],pp88[22],pp99[12]};
    assign in1972_2 = {c158,pp101[8],pp89[21],pp100[11]};
    CLA_4 KS_1972(s1972, c1972, in1972_1, in1972_2);
    wire[3:0] s1973, in1973_1, in1973_2;
    wire c1973;
    assign in1973_1 = {c159,pp102[7],pp90[20],pp101[10]};
    assign in1973_2 = {c161,pp103[6],pp91[19],pp102[9]};
    CLA_4 KS_1973(s1973, c1973, in1973_1, in1973_2);
    wire[3:0] s1974, in1974_1, in1974_2;
    wire c1974;
    assign in1974_1 = {c163,pp104[5],pp92[18],pp103[8]};
    assign in1974_2 = {c165,pp105[4],pp93[17],pp104[7]};
    CLA_4 KS_1974(s1974, c1974, in1974_1, in1974_2);
    wire[3:0] s1975, in1975_1, in1975_2;
    wire c1975;
    assign in1975_1 = {c167,pp106[3],pp94[16],pp105[6]};
    assign in1975_2 = {c169,pp107[2],pp95[15],pp106[5]};
    CLA_4 KS_1975(s1975, c1975, in1975_1, in1975_2);
    wire[3:0] s1976, in1976_1, in1976_2;
    wire c1976;
    assign in1976_1 = {c173,pp108[1],pp96[14],pp107[4]};
    assign in1976_2 = {c177,pp109[0],pp97[13],pp108[3]};
    CLA_4 KS_1976(s1976, c1976, in1976_1, in1976_2);
    wire[3:0] s1977, in1977_1, in1977_2;
    wire c1977;
    assign in1977_1 = {s180[1],s180[2],pp98[12],pp109[2]};
    assign in1977_2 = {s181[1],s181[2],pp99[11],pp110[1]};
    CLA_4 KS_1977(s1977, c1977, in1977_1, in1977_2);
    wire[3:0] s1978, in1978_1, in1978_2;
    wire c1978;
    assign in1978_1 = {s182[1],s182[2],pp100[10],pp111[0]};
    assign in1978_2 = {s183[1],s183[2],pp101[9],c180};
    CLA_4 KS_1978(s1978, c1978, in1978_1, in1978_2);
    wire[3:0] s1979, in1979_1, in1979_2;
    wire c1979;
    assign in1979_1 = {s184[1],s184[2],pp102[8],c181};
    assign in1979_2 = {s185[1],s185[2],pp103[7],c182};
    CLA_4 KS_1979(s1979, c1979, in1979_1, in1979_2);
    wire[3:0] s1980, in1980_1, in1980_2;
    wire c1980;
    assign in1980_1 = {s186[1],s186[2],pp104[6],c183};
    assign in1980_2 = {s187[1],s187[2],pp105[5],c184};
    CLA_4 KS_1980(s1980, c1980, in1980_1, in1980_2);
    wire[3:0] s1981, in1981_1, in1981_2;
    wire c1981;
    assign in1981_1 = {s188[1],s188[2],pp106[4],c185};
    assign in1981_2 = {s189[1],s189[2],pp107[3],c186};
    CLA_4 KS_1981(s1981, c1981, in1981_1, in1981_2);
    wire[3:0] s1982, in1982_1, in1982_2;
    wire c1982;
    assign in1982_1 = {s190[1],s190[2],pp108[2],c187};
    assign in1982_2 = {s191[0],s191[1],pp109[1],c188};
    CLA_4 KS_1982(s1982, c1982, in1982_1, in1982_2);
    wire[3:0] s1983, in1983_1, in1983_2;
    wire c1983;
    assign in1983_1 = {s192[0],s192[1],pp110[0],c189};
    assign in1983_2 = {s193[0],s193[1],s180[3],c190};
    CLA_4 KS_1983(s1983, c1983, in1983_1, in1983_2);
    wire[3:0] s1984, in1984_1, in1984_2;
    wire c1984;
    assign in1984_1 = {s194[0],s194[1],s181[3],s191[3]};
    assign in1984_2 = {s195[0],s195[1],s182[3],s192[3]};
    CLA_4 KS_1984(s1984, c1984, in1984_1, in1984_2);
    wire[3:0] s1985, in1985_1, in1985_2;
    wire c1985;
    assign in1985_1 = {s196[0],s196[1],s183[3],s193[3]};
    assign in1985_2 = {s197[0],s197[1],s184[3],s194[3]};
    CLA_4 KS_1985(s1985, c1985, in1985_1, in1985_2);
    wire[3:0] s1986, in1986_1, in1986_2;
    wire c1986;
    assign in1986_1 = {s198[0],s198[1],s185[3],s195[3]};
    assign in1986_2 = {s199[0],s199[1],s186[3],s196[3]};
    CLA_4 KS_1986(s1986, c1986, in1986_1, in1986_2);
    wire[3:0] s1987, in1987_1, in1987_2;
    wire c1987;
    assign in1987_1 = {s200[0],s200[1],s187[3],s197[3]};
    assign in1987_2 = {s201[0],s201[1],s188[3],s198[3]};
    CLA_4 KS_1987(s1987, c1987, in1987_1, in1987_2);
    wire[3:0] s1988, in1988_1, in1988_2;
    wire c1988;
    assign in1988_1 = {s202[0],s202[1],s189[3],s199[3]};
    assign in1988_2 = {s203[0],s203[1],s190[3],s200[3]};
    CLA_4 KS_1988(s1988, c1988, in1988_1, in1988_2);
    wire[3:0] s1989, in1989_1, in1989_2;
    wire c1989;
    assign in1989_1 = {s204[0],s204[1],s191[2],s201[3]};
    assign in1989_2 = {s205[0],s205[1],s192[2],s202[3]};
    CLA_4 KS_1989(s1989, c1989, in1989_1, in1989_2);
    wire[3:0] s1990, in1990_1, in1990_2;
    wire c1990;
    assign in1990_1 = {s206[0],s206[1],s193[2],s203[3]};
    assign in1990_2 = {s207[0],s207[1],s194[2],s204[3]};
    CLA_4 KS_1990(s1990, c1990, in1990_1, in1990_2);
    wire[3:0] s1991, in1991_1, in1991_2;
    wire c1991;
    assign in1991_1 = {s208[0],s208[1],s195[2],s205[3]};
    assign in1991_2 = {s209[0],s209[1],s196[2],s206[3]};
    CLA_4 KS_1991(s1991, c1991, in1991_1, in1991_2);
    wire[3:0] s1992, in1992_1, in1992_2;
    wire c1992;
    assign in1992_1 = {s210[0],s210[1],s197[2],s207[3]};
    assign in1992_2 = {s211[0],s211[1],s198[2],s208[3]};
    CLA_4 KS_1992(s1992, c1992, in1992_1, in1992_2);
    wire[3:0] s1993, in1993_1, in1993_2;
    wire c1993;
    assign in1993_1 = {s212[0],s212[1],s199[2],s209[3]};
    assign in1993_2 = {s213[0],s213[1],s200[2],s210[3]};
    CLA_4 KS_1993(s1993, c1993, in1993_1, in1993_2);
    wire[3:0] s1994, in1994_1, in1994_2;
    wire c1994;
    assign in1994_1 = {s214[0],s214[1],s201[2],s211[3]};
    assign in1994_2 = {s215[0],c215,s202[2],s212[3]};
    CLA_4 KS_1994(s1994, c1994, in1994_1, in1994_2);
    wire[3:0] s1995, in1995_1, in1995_2;
    wire c1995;
    assign in1995_1 = {s216[0],s216[1],s203[2],s213[3]};
    assign in1995_2 = {s217[0],c217,s204[2],s214[3]};
    CLA_4 KS_1995(s1995, c1995, in1995_1, in1995_2);
    wire[3:0] s1996, in1996_1, in1996_2;
    wire c1996;
    assign in1996_1 = {s218[0],s218[1],s205[2],s216[3]};
    assign in1996_2 = {s219[0],c219,s206[2],s220[3]};
    CLA_4 KS_1996(s1996, c1996, in1996_1, in1996_2);
    wire[3:0] s1997, in1997_1, in1997_2;
    wire c1997;
    assign in1997_1 = {s220[0],s220[1],s207[2],s224[3]};
    assign in1997_2 = {s221[0],c221,s208[2],s228[3]};
    CLA_4 KS_1997(s1997, c1997, in1997_1, in1997_2);
    wire[3:0] s1998, in1998_1, in1998_2;
    wire c1998;
    assign in1998_1 = {s222[0],s222[1],s209[2],s232[3]};
    assign in1998_2 = {s223[0],c223,s210[2],s236[3]};
    CLA_4 KS_1998(s1998, c1998, in1998_1, in1998_2);
    wire[3:0] s1999, in1999_1, in1999_2;
    wire c1999;
    assign in1999_1 = {s224[0],s224[1],s211[2],s240[0]};
    assign in1999_2 = {s225[0],c225,s212[2],s241[0]};
    CLA_4 KS_1999(s1999, c1999, in1999_1, in1999_2);
    wire[3:0] s2000, in2000_1, in2000_2;
    wire c2000;
    assign in2000_1 = {s226[0],s226[1],s213[2],s242[0]};
    assign in2000_2 = {s227[0],c227,s214[2],s243[0]};
    CLA_4 KS_2000(s2000, c2000, in2000_1, in2000_2);
    wire[0:0] s2001, in2001_1, in2001_2;
    wire c2001;
    assign in2001_1 = {s228[0]};
    assign in2001_2 = {s229[0]};
    Half_Adder KS_2001(s2001, c2001, in2001_1, in2001_2);
    wire[1:0] s2002, in2002_1, in2002_2;
    wire c2002;
    assign in2002_1 = {s230[0],s228[1]};
    assign in2002_2 = {s231[0],c229};
    CLA_2 KS_2002(s2002, c2002, in2002_1, in2002_2);
    wire[0:0] s2003, in2003_1, in2003_2;
    wire c2003;
    assign in2003_1 = {s232[0]};
    assign in2003_2 = {s233[0]};
    Half_Adder KS_2003(s2003, c2003, in2003_1, in2003_2);
    wire[2:0] s2004, in2004_1, in2004_2;
    wire c2004;
    assign in2004_1 = {s234[0],s230[1],s216[2]};
    assign in2004_2 = {s235[0],c231,c218};
    CLA_3 KS_2004(s2004, c2004, in2004_1, in2004_2);
    wire[0:0] s2005, in2005_1, in2005_2;
    wire c2005;
    assign in2005_1 = {s236[0]};
    assign in2005_2 = {s237[0]};
    Half_Adder KS_2005(s2005, c2005, in2005_1, in2005_2);
    wire[1:0] s2006, in2006_1, in2006_2;
    wire c2006;
    assign in2006_1 = {s238[0],s232[1]};
    assign in2006_2 = {s239[0],c233};
    CLA_2 KS_2006(s2006, c2006, in2006_1, in2006_2);
    wire[0:0] s2007, in2007_1, in2007_2;
    wire c2007;
    assign in2007_1 = {c1903};
    assign in2007_2 = {c1904};
    Half_Adder KS_2007(s2007, c2007, in2007_1, in2007_2);
    wire[3:0] s2008, in2008_1, in2008_2;
    wire c2008;
    assign in2008_1 = {c1905,s234[1],s220[2],s244[0]};
    assign in2008_2 = {c1906,c235,c222,s245[0]};
    CLA_4 KS_2008(s2008, c2008, in2008_1, in2008_2);
    wire[0:0] s2009, in2009_1, in2009_2;
    wire c2009;
    assign in2009_1 = {c1907};
    assign in2009_2 = {c1908};
    Half_Adder KS_2009(s2009, c2009, in2009_1, in2009_2);
    wire[1:0] s2010, in2010_1, in2010_2;
    wire c2010;
    assign in2010_1 = {c1909,s236[1]};
    assign in2010_2 = {c1910,c237};
    CLA_2 KS_2010(s2010, c2010, in2010_1, in2010_2);
    wire[0:0] s2011, in2011_1, in2011_2;
    wire c2011;
    assign in2011_1 = {c1911};
    assign in2011_2 = {c1912};
    Half_Adder KS_2011(s2011, c2011, in2011_1, in2011_2);
    wire[2:0] s2012, in2012_1, in2012_2;
    wire c2012;
    assign in2012_1 = {c1913,s238[1],s224[2]};
    assign in2012_2 = {c1914,c239,c226};
    CLA_3 KS_2012(s2012, c2012, in2012_1, in2012_2);
    wire[0:0] s2013, in2013_1, in2013_2;
    wire c2013;
    assign in2013_1 = {c1915};
    assign in2013_2 = {c1916};
    Half_Adder KS_2013(s2013, c2013, in2013_1, in2013_2);
    wire[1:0] s2014, in2014_1, in2014_2;
    wire c2014;
    assign in2014_1 = {c1917,s1969[1]};
    assign in2014_2 = {c1918,s1970[1]};
    CLA_2 KS_2014(s2014, c2014, in2014_1, in2014_2);
    wire[0:0] s2015, in2015_1, in2015_2;
    wire c2015;
    assign in2015_1 = {c1919};
    assign in2015_2 = {c1920};
    Half_Adder KS_2015(s2015, c2015, in2015_1, in2015_2);
    wire[3:0] s2016, in2016_1, in2016_2;
    wire c2016;
    assign in2016_1 = {c1921,s1971[1],s228[2],s246[0]};
    assign in2016_2 = {c1922,s1972[1],c230,s247[0]};
    CLA_4 KS_2016(s2016, c2016, in2016_1, in2016_2);
    wire[0:0] s2017, in2017_1, in2017_2;
    wire c2017;
    assign in2017_1 = {c1923};
    assign in2017_2 = {c1924};
    Half_Adder KS_2017(s2017, c2017, in2017_1, in2017_2);
    wire[1:0] s2018, in2018_1, in2018_2;
    wire c2018;
    assign in2018_1 = {c1925,s1973[1]};
    assign in2018_2 = {c1926,s1974[1]};
    CLA_2 KS_2018(s2018, c2018, in2018_1, in2018_2);
    wire[0:0] s2019, in2019_1, in2019_2;
    wire c2019;
    assign in2019_1 = {c1927};
    assign in2019_2 = {c1928};
    Half_Adder KS_2019(s2019, c2019, in2019_1, in2019_2);
    wire[2:0] s2020, in2020_1, in2020_2;
    wire c2020;
    assign in2020_1 = {c1929,s1975[1],s232[2]};
    assign in2020_2 = {c1930,s1976[1],c234};
    CLA_3 KS_2020(s2020, c2020, in2020_1, in2020_2);
    wire[0:0] s2021, in2021_1, in2021_2;
    wire c2021;
    assign in2021_1 = {c1931};
    assign in2021_2 = {c1932};
    Half_Adder KS_2021(s2021, c2021, in2021_1, in2021_2);
    wire[1:0] s2022, in2022_1, in2022_2;
    wire c2022;
    assign in2022_1 = {c1933,s1977[1]};
    assign in2022_2 = {c1935,s1978[1]};
    CLA_2 KS_2022(s2022, c2022, in2022_1, in2022_2);
    wire[0:0] s2023, in2023_1, in2023_2;
    wire c2023;
    assign in2023_1 = {c1943};
    assign in2023_2 = {c1951};
    Half_Adder KS_2023(s2023, c2023, in2023_1, in2023_2);
    wire[3:0] s2024, in2024_1, in2024_2;
    wire c2024;
    assign in2024_1 = {c1959,s1979[1],s236[2],s248[0]};
    assign in2024_2 = {c1967,s1980[1],c238,s249[0]};
    CLA_4 KS_2024(s2024, c2024, in2024_1, in2024_2);
    wire[0:0] s2025, in2025_1, in2025_2;
    wire c2025;
    assign in2025_1 = {s1969[0]};
    assign in2025_2 = {s1970[0]};
    Half_Adder KS_2025(s2025, c2025, in2025_1, in2025_2);
    wire[1:0] s2026, in2026_1, in2026_2;
    wire c2026;
    assign in2026_1 = {s1971[0],s1981[1]};
    assign in2026_2 = {s1972[0],s1982[1]};
    CLA_2 KS_2026(s2026, c2026, in2026_1, in2026_2);
    wire[0:0] s2027, in2027_1, in2027_2;
    wire c2027;
    assign in2027_1 = {s1973[0]};
    assign in2027_2 = {s1974[0]};
    Half_Adder KS_2027(s2027, c2027, in2027_1, in2027_2);
    wire[2:0] s2028, in2028_1, in2028_2;
    wire c2028;
    assign in2028_1 = {s1975[0],s1983[1],s1969[2]};
    assign in2028_2 = {s1976[0],s1984[1],s1970[2]};
    CLA_3 KS_2028(s2028, c2028, in2028_1, in2028_2);
    wire[0:0] s2029, in2029_1, in2029_2;
    wire c2029;
    assign in2029_1 = {s1977[0]};
    assign in2029_2 = {s1978[0]};
    Half_Adder KS_2029(s2029, c2029, in2029_1, in2029_2);
    wire[1:0] s2030, in2030_1, in2030_2;
    wire c2030;
    assign in2030_1 = {s1979[0],s1985[1]};
    assign in2030_2 = {s1980[0],s1986[1]};
    CLA_2 KS_2030(s2030, c2030, in2030_1, in2030_2);
    wire[0:0] s2031, in2031_1, in2031_2;
    wire c2031;
    assign in2031_1 = {s1981[0]};
    assign in2031_2 = {s1982[0]};
    Half_Adder KS_2031(s2031, c2031, in2031_1, in2031_2);
    wire[3:0] s2032, in2032_1, in2032_2;
    wire c2032;
    assign in2032_1 = {s1983[0],s1987[1],s1971[2],s250[0]};
    assign in2032_2 = {s1984[0],s1988[1],s1972[2],s251[0]};
    CLA_4 KS_2032(s2032, c2032, in2032_1, in2032_2);
    wire[0:0] s2033, in2033_1, in2033_2;
    wire c2033;
    assign in2033_1 = {s1985[0]};
    assign in2033_2 = {s1986[0]};
    Half_Adder KS_2033(s2033, c2033, in2033_1, in2033_2);
    wire[1:0] s2034, in2034_1, in2034_2;
    wire c2034;
    assign in2034_1 = {s1988[0],s1989[1]};
    assign in2034_2 = {s1989[0],s1990[1]};
    CLA_2_c KS_2034(s2034, c2034, in2034_1, in2034_2, s1987[0]);
    wire[3:0] s2035, in2035_1, in2035_2;
    wire c2035;
    assign in2035_1 = {c211,pp104[9],pp92[22],pp111[4]};
    assign in2035_2 = {c212,pp105[8],pp93[21],pp112[3]};
    CLA_4 KS_2035(s2035, c2035, in2035_1, in2035_2);
    wire[3:0] s2036, in2036_1, in2036_2;
    wire c2036;
    assign in2036_1 = {c213,pp106[7],pp94[20],pp113[2]};
    assign in2036_2 = {c214,pp107[6],pp95[19],pp114[1]};
    CLA_4 KS_2036(s2036, c2036, in2036_1, in2036_2);
    wire[3:0] s2037, in2037_1, in2037_2;
    wire c2037;
    assign in2037_1 = {c216,pp108[5],pp96[18],pp115[0]};
    assign in2037_2 = {c220,pp109[4],pp97[17],c240};
    CLA_4 KS_2037(s2037, c2037, in2037_1, in2037_2);
    wire[3:0] s2038, in2038_1, in2038_2;
    wire c2038;
    assign in2038_1 = {c224,pp110[3],pp98[16],c241};
    assign in2038_2 = {c228,pp111[2],pp99[15],c242};
    CLA_4 KS_2038(s2038, c2038, in2038_1, in2038_2);
    wire[3:0] s2039, in2039_1, in2039_2;
    wire c2039;
    assign in2039_1 = {c232,pp112[1],pp100[14],c243};
    assign in2039_2 = {c236,pp113[0],pp101[13],c244};
    CLA_4 KS_2039(s2039, c2039, in2039_1, in2039_2);
    wire[3:0] s2040, in2040_1, in2040_2;
    wire c2040;
    assign in2040_1 = {s240[1],s240[2],pp102[12],c245};
    assign in2040_2 = {s241[1],s241[2],pp103[11],c246};
    CLA_4 KS_2040(s2040, c2040, in2040_1, in2040_2);
    wire[3:0] s2041, in2041_1, in2041_2;
    wire c2041;
    assign in2041_1 = {s242[1],s242[2],pp104[10],c247};
    assign in2041_2 = {s243[1],s243[2],pp105[9],c248};
    CLA_4 KS_2041(s2041, c2041, in2041_1, in2041_2);
    wire[3:0] s2042, in2042_1, in2042_2;
    wire c2042;
    assign in2042_1 = {s244[1],s244[2],pp106[8],c249};
    assign in2042_2 = {s245[1],s245[2],pp107[7],c250};
    CLA_4 KS_2042(s2042, c2042, in2042_1, in2042_2);
    wire[3:0] s2043, in2043_1, in2043_2;
    wire c2043;
    assign in2043_1 = {s246[1],s246[2],pp108[6],c251};
    assign in2043_2 = {s247[1],s247[2],pp109[5],c252};
    CLA_4 KS_2043(s2043, c2043, in2043_1, in2043_2);
    wire[3:0] s2044, in2044_1, in2044_2;
    wire c2044;
    assign in2044_1 = {s248[1],s248[2],pp110[4],c253};
    assign in2044_2 = {s249[1],s249[2],pp111[3],c254};
    CLA_4 KS_2044(s2044, c2044, in2044_1, in2044_2);
    wire[3:0] s2045, in2045_1, in2045_2;
    wire c2045;
    assign in2045_1 = {s250[1],s250[2],pp112[2],c255};
    assign in2045_2 = {s251[1],s251[2],pp113[1],s256[3]};
    CLA_4 KS_2045(s2045, c2045, in2045_1, in2045_2);
    wire[3:0] s2046, in2046_1, in2046_2;
    wire c2046;
    assign in2046_1 = {s252[1],s252[2],pp114[0],s257[3]};
    assign in2046_2 = {s253[1],s253[2],s240[3],s258[3]};
    CLA_4 KS_2046(s2046, c2046, in2046_1, in2046_2);
    wire[3:0] s2047, in2047_1, in2047_2;
    wire c2047;
    assign in2047_1 = {s254[1],s254[2],s241[3],s259[3]};
    assign in2047_2 = {s255[1],s255[2],s242[3],s260[3]};
    CLA_4 KS_2047(s2047, c2047, in2047_1, in2047_2);
    wire[3:0] s2048, in2048_1, in2048_2;
    wire c2048;
    assign in2048_1 = {s256[0],s256[1],s243[3],s261[3]};
    assign in2048_2 = {s257[0],s257[1],s244[3],s262[3]};
    CLA_4 KS_2048(s2048, c2048, in2048_1, in2048_2);
    wire[3:0] s2049, in2049_1, in2049_2;
    wire c2049;
    assign in2049_1 = {s258[0],s258[1],s245[3],s263[3]};
    assign in2049_2 = {s259[0],s259[1],s246[3],s264[3]};
    CLA_4 KS_2049(s2049, c2049, in2049_1, in2049_2);
    wire[3:0] s2050, in2050_1, in2050_2;
    wire c2050;
    assign in2050_1 = {s260[0],s260[1],s247[3],s265[3]};
    assign in2050_2 = {s261[0],s261[1],s248[3],s266[3]};
    CLA_4 KS_2050(s2050, c2050, in2050_1, in2050_2);
    wire[3:0] s2051, in2051_1, in2051_2;
    wire c2051;
    assign in2051_1 = {s262[0],s262[1],s249[3],s267[3]};
    assign in2051_2 = {s263[0],s263[1],s250[3],s268[3]};
    CLA_4 KS_2051(s2051, c2051, in2051_1, in2051_2);
    wire[3:0] s2052, in2052_1, in2052_2;
    wire c2052;
    assign in2052_1 = {s264[0],s264[1],s251[3],s269[3]};
    assign in2052_2 = {s265[0],s265[1],s252[3],s270[3]};
    CLA_4 KS_2052(s2052, c2052, in2052_1, in2052_2);
    wire[3:0] s2053, in2053_1, in2053_2;
    wire c2053;
    assign in2053_1 = {s266[0],s266[1],s253[3],s271[3]};
    assign in2053_2 = {s267[0],s267[1],s254[3],s272[3]};
    CLA_4 KS_2053(s2053, c2053, in2053_1, in2053_2);
    wire[3:0] s2054, in2054_1, in2054_2;
    wire c2054;
    assign in2054_1 = {s268[0],s268[1],s255[3],s273[3]};
    assign in2054_2 = {s269[0],s269[1],s256[2],s274[3]};
    CLA_4 KS_2054(s2054, c2054, in2054_1, in2054_2);
    wire[3:0] s2055, in2055_1, in2055_2;
    wire c2055;
    assign in2055_1 = {s270[0],s270[1],s257[2],s275[3]};
    assign in2055_2 = {s271[0],s271[1],s258[2],s276[3]};
    CLA_4 KS_2055(s2055, c2055, in2055_1, in2055_2);
    wire[3:0] s2056, in2056_1, in2056_2;
    wire c2056;
    assign in2056_1 = {s272[0],s272[1],s259[2],s277[3]};
    assign in2056_2 = {s273[0],s273[1],s260[2],s278[3]};
    CLA_4 KS_2056(s2056, c2056, in2056_1, in2056_2);
    wire[3:0] s2057, in2057_1, in2057_2;
    wire c2057;
    assign in2057_1 = {s274[0],s274[1],s261[2],s280[3]};
    assign in2057_2 = {s275[0],s275[1],s262[2],s284[3]};
    CLA_4 KS_2057(s2057, c2057, in2057_1, in2057_2);
    wire[3:0] s2058, in2058_1, in2058_2;
    wire c2058;
    assign in2058_1 = {s276[0],s276[1],s263[2],s288[3]};
    assign in2058_2 = {s277[0],s277[1],s264[2],s292[3]};
    CLA_4 KS_2058(s2058, c2058, in2058_1, in2058_2);
    wire[3:0] s2059, in2059_1, in2059_2;
    wire c2059;
    assign in2059_1 = {s278[0],s278[1],s265[2],s296[3]};
    assign in2059_2 = {s279[0],c279,s266[2],s300[3]};
    CLA_4 KS_2059(s2059, c2059, in2059_1, in2059_2);
    wire[3:0] s2060, in2060_1, in2060_2;
    wire c2060;
    assign in2060_1 = {s280[0],s280[1],s267[2],s304[3]};
    assign in2060_2 = {s281[0],c281,s268[2],s306[0]};
    CLA_4 KS_2060(s2060, c2060, in2060_1, in2060_2);
    wire[3:0] s2061, in2061_1, in2061_2;
    wire c2061;
    assign in2061_1 = {s282[0],s282[1],s269[2],s307[0]};
    assign in2061_2 = {s283[0],c283,s270[2],s308[0]};
    CLA_4 KS_2061(s2061, c2061, in2061_1, in2061_2);
    wire[3:0] s2062, in2062_1, in2062_2;
    wire c2062;
    assign in2062_1 = {s284[0],s284[1],s271[2],s309[0]};
    assign in2062_2 = {s285[0],c285,s272[2],s310[0]};
    CLA_4 KS_2062(s2062, c2062, in2062_1, in2062_2);
    wire[3:0] s2063, in2063_1, in2063_2;
    wire c2063;
    assign in2063_1 = {s286[0],s286[1],s273[2],s311[0]};
    assign in2063_2 = {s287[0],c287,s274[2],s312[0]};
    CLA_4 KS_2063(s2063, c2063, in2063_1, in2063_2);
    wire[3:0] s2064, in2064_1, in2064_2;
    wire c2064;
    assign in2064_1 = {s288[0],s288[1],s275[2],s313[0]};
    assign in2064_2 = {s289[0],c289,s276[2],s314[0]};
    CLA_4 KS_2064(s2064, c2064, in2064_1, in2064_2);
    wire[3:0] s2065, in2065_1, in2065_2;
    wire c2065;
    assign in2065_1 = {s290[0],s290[1],s277[2],s315[0]};
    assign in2065_2 = {s291[0],c291,s278[2],s316[0]};
    CLA_4 KS_2065(s2065, c2065, in2065_1, in2065_2);
    wire[1:0] s2066, in2066_1, in2066_2;
    wire c2066;
    assign in2066_1 = {s292[0],s292[1]};
    assign in2066_2 = {s293[0],c293};
    CLA_2 KS_2066(s2066, c2066, in2066_1, in2066_2);
    wire[0:0] s2067, in2067_1, in2067_2;
    wire c2067;
    assign in2067_1 = {s294[0]};
    assign in2067_2 = {s295[0]};
    Half_Adder KS_2067(s2067, c2067, in2067_1, in2067_2);
    wire[3:0] s2068, in2068_1, in2068_2;
    wire c2068;
    assign in2068_1 = {s296[0],s294[1],s280[2],s317[0]};
    assign in2068_2 = {s297[0],c295,c282,s318[0]};
    CLA_4 KS_2068(s2068, c2068, in2068_1, in2068_2);
    wire[0:0] s2069, in2069_1, in2069_2;
    wire c2069;
    assign in2069_1 = {s298[0]};
    assign in2069_2 = {s299[0]};
    Half_Adder KS_2069(s2069, c2069, in2069_1, in2069_2);
    wire[1:0] s2070, in2070_1, in2070_2;
    wire c2070;
    assign in2070_1 = {s300[0],s296[1]};
    assign in2070_2 = {s301[0],c297};
    CLA_2 KS_2070(s2070, c2070, in2070_1, in2070_2);
    wire[0:0] s2071, in2071_1, in2071_2;
    wire c2071;
    assign in2071_1 = {s302[0]};
    assign in2071_2 = {s303[0]};
    Half_Adder KS_2071(s2071, c2071, in2071_1, in2071_2);
    wire[2:0] s2072, in2072_1, in2072_2;
    wire c2072;
    assign in2072_1 = {s304[0],s298[1],s284[2]};
    assign in2072_2 = {s305[0],c299,c286};
    CLA_3 KS_2072(s2072, c2072, in2072_1, in2072_2);
    wire[0:0] s2073, in2073_1, in2073_2;
    wire c2073;
    assign in2073_1 = {c1969};
    assign in2073_2 = {c1970};
    Half_Adder KS_2073(s2073, c2073, in2073_1, in2073_2);
    wire[1:0] s2074, in2074_1, in2074_2;
    wire c2074;
    assign in2074_1 = {c1971,s300[1]};
    assign in2074_2 = {c1972,c301};
    CLA_2 KS_2074(s2074, c2074, in2074_1, in2074_2);
    wire[0:0] s2075, in2075_1, in2075_2;
    wire c2075;
    assign in2075_1 = {c1973};
    assign in2075_2 = {c1974};
    Half_Adder KS_2075(s2075, c2075, in2075_1, in2075_2);
    wire[3:0] s2076, in2076_1, in2076_2;
    wire c2076;
    assign in2076_1 = {c1975,s302[1],s288[2],s319[0]};
    assign in2076_2 = {c1976,c303,c290,s320[0]};
    CLA_4 KS_2076(s2076, c2076, in2076_1, in2076_2);
    wire[0:0] s2077, in2077_1, in2077_2;
    wire c2077;
    assign in2077_1 = {c1977};
    assign in2077_2 = {c1978};
    Half_Adder KS_2077(s2077, c2077, in2077_1, in2077_2);
    wire[1:0] s2078, in2078_1, in2078_2;
    wire c2078;
    assign in2078_1 = {c1979,s304[1]};
    assign in2078_2 = {c1980,c305};
    CLA_2 KS_2078(s2078, c2078, in2078_1, in2078_2);
    wire[0:0] s2079, in2079_1, in2079_2;
    wire c2079;
    assign in2079_1 = {c1981};
    assign in2079_2 = {c1982};
    Half_Adder KS_2079(s2079, c2079, in2079_1, in2079_2);
    wire[2:0] s2080, in2080_1, in2080_2;
    wire c2080;
    assign in2080_1 = {c1983,s2035[1],s292[2]};
    assign in2080_2 = {c1984,s2036[1],c294};
    CLA_3 KS_2080(s2080, c2080, in2080_1, in2080_2);
    wire[0:0] s2081, in2081_1, in2081_2;
    wire c2081;
    assign in2081_1 = {c1985};
    assign in2081_2 = {c1986};
    Half_Adder KS_2081(s2081, c2081, in2081_1, in2081_2);
    wire[1:0] s2082, in2082_1, in2082_2;
    wire c2082;
    assign in2082_1 = {c1987,s2037[1]};
    assign in2082_2 = {c1988,s2038[1]};
    CLA_2 KS_2082(s2082, c2082, in2082_1, in2082_2);
    wire[0:0] s2083, in2083_1, in2083_2;
    wire c2083;
    assign in2083_1 = {c1989};
    assign in2083_2 = {c1990};
    Half_Adder KS_2083(s2083, c2083, in2083_1, in2083_2);
    wire[3:0] s2084, in2084_1, in2084_2;
    wire c2084;
    assign in2084_1 = {c1991,s2039[1],s296[2],s321[0]};
    assign in2084_2 = {c1992,s2040[1],c298,s322[0]};
    CLA_4 KS_2084(s2084, c2084, in2084_1, in2084_2);
    wire[0:0] s2085, in2085_1, in2085_2;
    wire c2085;
    assign in2085_1 = {c1993};
    assign in2085_2 = {c1994};
    Half_Adder KS_2085(s2085, c2085, in2085_1, in2085_2);
    wire[1:0] s2086, in2086_1, in2086_2;
    wire c2086;
    assign in2086_1 = {c1995,s2041[1]};
    assign in2086_2 = {c1996,s2042[1]};
    CLA_2 KS_2086(s2086, c2086, in2086_1, in2086_2);
    wire[0:0] s2087, in2087_1, in2087_2;
    wire c2087;
    assign in2087_1 = {c1997};
    assign in2087_2 = {c1998};
    Half_Adder KS_2087(s2087, c2087, in2087_1, in2087_2);
    wire[2:0] s2088, in2088_1, in2088_2;
    wire c2088;
    assign in2088_1 = {c1999,s2043[1],s300[2]};
    assign in2088_2 = {c2000,s2044[1],c302};
    CLA_3 KS_2088(s2088, c2088, in2088_1, in2088_2);
    wire[0:0] s2089, in2089_1, in2089_2;
    wire c2089;
    assign in2089_1 = {c2008};
    assign in2089_2 = {c2016};
    Half_Adder KS_2089(s2089, c2089, in2089_1, in2089_2);
    wire[1:0] s2090, in2090_1, in2090_2;
    wire c2090;
    assign in2090_1 = {c2024,s2045[1]};
    assign in2090_2 = {c2032,s2046[1]};
    CLA_2 KS_2090(s2090, c2090, in2090_1, in2090_2);
    wire[0:0] s2091, in2091_1, in2091_2;
    wire c2091;
    assign in2091_1 = {s2035[0]};
    assign in2091_2 = {s2036[0]};
    Half_Adder KS_2091(s2091, c2091, in2091_1, in2091_2);
    wire[3:0] s2092, in2092_1, in2092_2;
    wire c2092;
    assign in2092_1 = {s2037[0],s2047[1],s304[2],s323[0]};
    assign in2092_2 = {s2038[0],s2048[1],s2035[2],s324[0]};
    CLA_4 KS_2092(s2092, c2092, in2092_1, in2092_2);
    wire[0:0] s2093, in2093_1, in2093_2;
    wire c2093;
    assign in2093_1 = {s2039[0]};
    assign in2093_2 = {s2040[0]};
    Half_Adder KS_2093(s2093, c2093, in2093_1, in2093_2);
    wire[1:0] s2094, in2094_1, in2094_2;
    wire c2094;
    assign in2094_1 = {s2041[0],s2049[1]};
    assign in2094_2 = {s2042[0],s2050[1]};
    CLA_2 KS_2094(s2094, c2094, in2094_1, in2094_2);
    wire[0:0] s2095, in2095_1, in2095_2;
    wire c2095;
    assign in2095_1 = {s2043[0]};
    assign in2095_2 = {s2044[0]};
    Half_Adder KS_2095(s2095, c2095, in2095_1, in2095_2);
    wire[2:0] s2096, in2096_1, in2096_2;
    wire c2096;
    assign in2096_1 = {s2045[0],s2051[1],s2036[2]};
    assign in2096_2 = {s2046[0],s2052[1],s2037[2]};
    CLA_3 KS_2096(s2096, c2096, in2096_1, in2096_2);
    wire[0:0] s2097, in2097_1, in2097_2;
    wire c2097;
    assign in2097_1 = {s2047[0]};
    assign in2097_2 = {s2048[0]};
    Half_Adder KS_2097(s2097, c2097, in2097_1, in2097_2);
    wire[1:0] s2098, in2098_1, in2098_2;
    wire c2098;
    assign in2098_1 = {s2049[0],s2053[1]};
    assign in2098_2 = {s2050[0],s2054[1]};
    CLA_2 KS_2098(s2098, c2098, in2098_1, in2098_2);
    wire[0:0] s2099, in2099_1, in2099_2;
    wire c2099;
    assign in2099_1 = {s2051[0]};
    assign in2099_2 = {s2052[0]};
    Half_Adder KS_2099(s2099, c2099, in2099_1, in2099_2);
    wire[3:0] s2100, in2100_1, in2100_2;
    wire c2100;
    assign in2100_1 = {s2054[0],s2055[1],s2038[2],s325[0]};
    assign in2100_2 = {s2055[0],s2056[1],s2039[2],s326[0]};
    CLA_4_c KS_2100(s2100, c2100, in2100_1, in2100_2, s2053[0]);
    wire[3:0] s2101, in2101_1, in2101_2;
    wire c2101;
    assign in2101_1 = {c284,pp112[5],pp100[18],c323};
    assign in2101_2 = {c288,pp113[4],pp101[17],c324};
    CLA_4 KS_2101(s2101, c2101, in2101_1, in2101_2);
    wire[3:0] s2102, in2102_1, in2102_2;
    wire c2102;
    assign in2102_1 = {c292,pp114[3],pp102[16],c325};
    assign in2102_2 = {c296,pp115[2],pp103[15],c326};
    CLA_4 KS_2102(s2102, c2102, in2102_1, in2102_2);
    wire[3:0] s2103, in2103_1, in2103_2;
    wire c2103;
    assign in2103_1 = {c300,pp116[1],pp104[14],c327};
    assign in2103_2 = {c304,pp117[0],pp105[13],c328};
    CLA_4 KS_2103(s2103, c2103, in2103_1, in2103_2);
    wire[3:0] s2104, in2104_1, in2104_2;
    wire c2104;
    assign in2104_1 = {s306[1],s306[2],pp106[12],c329};
    assign in2104_2 = {s307[1],s307[2],pp107[11],c330};
    CLA_4 KS_2104(s2104, c2104, in2104_1, in2104_2);
    wire[3:0] s2105, in2105_1, in2105_2;
    wire c2105;
    assign in2105_1 = {s308[1],s308[2],pp108[10],s331[3]};
    assign in2105_2 = {s309[1],s309[2],pp109[9],s332[3]};
    CLA_4 KS_2105(s2105, c2105, in2105_1, in2105_2);
    wire[3:0] s2106, in2106_1, in2106_2;
    wire c2106;
    assign in2106_1 = {s310[1],s310[2],pp110[8],s333[3]};
    assign in2106_2 = {s311[1],s311[2],pp111[7],s334[3]};
    CLA_4 KS_2106(s2106, c2106, in2106_1, in2106_2);
    wire[3:0] s2107, in2107_1, in2107_2;
    wire c2107;
    assign in2107_1 = {s312[1],s312[2],pp112[6],s335[3]};
    assign in2107_2 = {s313[1],s313[2],pp113[5],s336[3]};
    CLA_4 KS_2107(s2107, c2107, in2107_1, in2107_2);
    wire[3:0] s2108, in2108_1, in2108_2;
    wire c2108;
    assign in2108_1 = {s314[1],s314[2],pp114[4],s337[3]};
    assign in2108_2 = {s315[1],s315[2],pp115[3],s338[3]};
    CLA_4 KS_2108(s2108, c2108, in2108_1, in2108_2);
    wire[3:0] s2109, in2109_1, in2109_2;
    wire c2109;
    assign in2109_1 = {s316[1],s316[2],pp116[2],s339[3]};
    assign in2109_2 = {s317[1],s317[2],pp117[1],s340[3]};
    CLA_4 KS_2109(s2109, c2109, in2109_1, in2109_2);
    wire[3:0] s2110, in2110_1, in2110_2;
    wire c2110;
    assign in2110_1 = {s318[1],s318[2],pp118[0],s341[3]};
    assign in2110_2 = {s319[1],s319[2],s306[3],s342[3]};
    CLA_4 KS_2110(s2110, c2110, in2110_1, in2110_2);
    wire[3:0] s2111, in2111_1, in2111_2;
    wire c2111;
    assign in2111_1 = {s320[1],s320[2],s307[3],s343[3]};
    assign in2111_2 = {s321[1],s321[2],s308[3],s344[3]};
    CLA_4 KS_2111(s2111, c2111, in2111_1, in2111_2);
    wire[3:0] s2112, in2112_1, in2112_2;
    wire c2112;
    assign in2112_1 = {s322[1],s322[2],s309[3],s345[3]};
    assign in2112_2 = {s323[1],s323[2],s310[3],s346[3]};
    CLA_4 KS_2112(s2112, c2112, in2112_1, in2112_2);
    wire[3:0] s2113, in2113_1, in2113_2;
    wire c2113;
    assign in2113_1 = {s324[1],s324[2],s311[3],s347[3]};
    assign in2113_2 = {s325[1],s325[2],s312[3],s348[3]};
    CLA_4 KS_2113(s2113, c2113, in2113_1, in2113_2);
    wire[3:0] s2114, in2114_1, in2114_2;
    wire c2114;
    assign in2114_1 = {s326[1],s326[2],s313[3],s350[3]};
    assign in2114_2 = {s327[1],s327[2],s314[3],s354[3]};
    CLA_4 KS_2114(s2114, c2114, in2114_1, in2114_2);
    wire[3:0] s2115, in2115_1, in2115_2;
    wire c2115;
    assign in2115_1 = {s328[1],s328[2],s315[3],s358[3]};
    assign in2115_2 = {s329[1],s329[2],s316[3],s362[3]};
    CLA_4 KS_2115(s2115, c2115, in2115_1, in2115_2);
    wire[3:0] s2116, in2116_1, in2116_2;
    wire c2116;
    assign in2116_1 = {s330[1],s330[2],s317[3],s366[3]};
    assign in2116_2 = {s331[0],s331[1],s318[3],s370[3]};
    CLA_4 KS_2116(s2116, c2116, in2116_1, in2116_2);
    wire[3:0] s2117, in2117_1, in2117_2;
    wire c2117;
    assign in2117_1 = {s332[0],s332[1],s319[3],s374[3]};
    assign in2117_2 = {s333[0],s333[1],s320[3],s376[0]};
    CLA_4 KS_2117(s2117, c2117, in2117_1, in2117_2);
    wire[3:0] s2118, in2118_1, in2118_2;
    wire c2118;
    assign in2118_1 = {s334[0],s334[1],s321[3],s377[0]};
    assign in2118_2 = {s335[0],s335[1],s322[3],s378[0]};
    CLA_4 KS_2118(s2118, c2118, in2118_1, in2118_2);
    wire[3:0] s2119, in2119_1, in2119_2;
    wire c2119;
    assign in2119_1 = {s336[0],s336[1],s323[3],s379[0]};
    assign in2119_2 = {s337[0],s337[1],s324[3],s380[0]};
    CLA_4 KS_2119(s2119, c2119, in2119_1, in2119_2);
    wire[3:0] s2120, in2120_1, in2120_2;
    wire c2120;
    assign in2120_1 = {s338[0],s338[1],s325[3],s381[0]};
    assign in2120_2 = {s339[0],s339[1],s326[3],s382[0]};
    CLA_4 KS_2120(s2120, c2120, in2120_1, in2120_2);
    wire[3:0] s2121, in2121_1, in2121_2;
    wire c2121;
    assign in2121_1 = {s340[0],s340[1],s327[3],s383[0]};
    assign in2121_2 = {s341[0],s341[1],s328[3],s384[0]};
    CLA_4 KS_2121(s2121, c2121, in2121_1, in2121_2);
    wire[3:0] s2122, in2122_1, in2122_2;
    wire c2122;
    assign in2122_1 = {s342[0],s342[1],s329[3],s385[0]};
    assign in2122_2 = {s343[0],s343[1],s330[3],s386[0]};
    CLA_4 KS_2122(s2122, c2122, in2122_1, in2122_2);
    wire[3:0] s2123, in2123_1, in2123_2;
    wire c2123;
    assign in2123_1 = {s344[0],s344[1],s331[2],s387[0]};
    assign in2123_2 = {s345[0],s345[1],s332[2],s388[0]};
    CLA_4 KS_2123(s2123, c2123, in2123_1, in2123_2);
    wire[3:0] s2124, in2124_1, in2124_2;
    wire c2124;
    assign in2124_1 = {s346[0],s346[1],s333[2],s389[0]};
    assign in2124_2 = {s347[0],s347[1],s334[2],s390[0]};
    CLA_4 KS_2124(s2124, c2124, in2124_1, in2124_2);
    wire[3:0] s2125, in2125_1, in2125_2;
    wire c2125;
    assign in2125_1 = {s348[0],s348[1],s335[2],s391[0]};
    assign in2125_2 = {s349[0],c349,s336[2],s392[0]};
    CLA_4 KS_2125(s2125, c2125, in2125_1, in2125_2);
    wire[3:0] s2126, in2126_1, in2126_2;
    wire c2126;
    assign in2126_1 = {s350[0],s350[1],s337[2],s393[0]};
    assign in2126_2 = {s351[0],c351,s338[2],s394[0]};
    CLA_4 KS_2126(s2126, c2126, in2126_1, in2126_2);
    wire[3:0] s2127, in2127_1, in2127_2;
    wire c2127;
    assign in2127_1 = {s352[0],s352[1],s339[2],s395[0]};
    assign in2127_2 = {s353[0],c353,s340[2],s396[0]};
    CLA_4 KS_2127(s2127, c2127, in2127_1, in2127_2);
    wire[3:0] s2128, in2128_1, in2128_2;
    wire c2128;
    assign in2128_1 = {s354[0],s354[1],s341[2],s397[0]};
    assign in2128_2 = {s355[0],c355,s342[2],s398[0]};
    CLA_4 KS_2128(s2128, c2128, in2128_1, in2128_2);
    wire[3:0] s2129, in2129_1, in2129_2;
    wire c2129;
    assign in2129_1 = {s356[0],s356[1],s343[2],s399[0]};
    assign in2129_2 = {s357[0],c357,s344[2],s400[0]};
    CLA_4 KS_2129(s2129, c2129, in2129_1, in2129_2);
    wire[3:0] s2130, in2130_1, in2130_2;
    wire c2130;
    assign in2130_1 = {s358[0],s358[1],s345[2],s401[0]};
    assign in2130_2 = {s359[0],c359,s346[2],s402[0]};
    CLA_4 KS_2130(s2130, c2130, in2130_1, in2130_2);
    wire[3:0] s2131, in2131_1, in2131_2;
    wire c2131;
    assign in2131_1 = {s360[0],s360[1],s347[2],s403[0]};
    assign in2131_2 = {s361[0],c361,s348[2],s404[0]};
    CLA_4 KS_2131(s2131, c2131, in2131_1, in2131_2);
    wire[1:0] s2132, in2132_1, in2132_2;
    wire c2132;
    assign in2132_1 = {s362[0],s362[1]};
    assign in2132_2 = {s363[0],c363};
    CLA_2 KS_2132(s2132, c2132, in2132_1, in2132_2);
    wire[0:0] s2133, in2133_1, in2133_2;
    wire c2133;
    assign in2133_1 = {s364[0]};
    assign in2133_2 = {s365[0]};
    Half_Adder KS_2133(s2133, c2133, in2133_1, in2133_2);
    wire[3:0] s2134, in2134_1, in2134_2;
    wire c2134;
    assign in2134_1 = {s366[0],s364[1],s350[2],s405[0]};
    assign in2134_2 = {s367[0],c365,c352,s406[0]};
    CLA_4 KS_2134(s2134, c2134, in2134_1, in2134_2);
    wire[0:0] s2135, in2135_1, in2135_2;
    wire c2135;
    assign in2135_1 = {s368[0]};
    assign in2135_2 = {s369[0]};
    Half_Adder KS_2135(s2135, c2135, in2135_1, in2135_2);
    wire[1:0] s2136, in2136_1, in2136_2;
    wire c2136;
    assign in2136_1 = {s370[0],s366[1]};
    assign in2136_2 = {s371[0],c367};
    CLA_2 KS_2136(s2136, c2136, in2136_1, in2136_2);
    wire[0:0] s2137, in2137_1, in2137_2;
    wire c2137;
    assign in2137_1 = {s372[0]};
    assign in2137_2 = {s373[0]};
    Half_Adder KS_2137(s2137, c2137, in2137_1, in2137_2);
    wire[2:0] s2138, in2138_1, in2138_2;
    wire c2138;
    assign in2138_1 = {s374[0],s368[1],s354[2]};
    assign in2138_2 = {s375[0],c369,c356};
    CLA_3 KS_2138(s2138, c2138, in2138_1, in2138_2);
    wire[0:0] s2139, in2139_1, in2139_2;
    wire c2139;
    assign in2139_1 = {c2035};
    assign in2139_2 = {c2036};
    Half_Adder KS_2139(s2139, c2139, in2139_1, in2139_2);
    wire[1:0] s2140, in2140_1, in2140_2;
    wire c2140;
    assign in2140_1 = {c2037,s370[1]};
    assign in2140_2 = {c2038,c371};
    CLA_2 KS_2140(s2140, c2140, in2140_1, in2140_2);
    wire[0:0] s2141, in2141_1, in2141_2;
    wire c2141;
    assign in2141_1 = {c2039};
    assign in2141_2 = {c2040};
    Half_Adder KS_2141(s2141, c2141, in2141_1, in2141_2);
    wire[3:0] s2142, in2142_1, in2142_2;
    wire c2142;
    assign in2142_1 = {c2041,s372[1],s358[2],s407[0]};
    assign in2142_2 = {c2042,c373,c360,s408[0]};
    CLA_4 KS_2142(s2142, c2142, in2142_1, in2142_2);
    wire[0:0] s2143, in2143_1, in2143_2;
    wire c2143;
    assign in2143_1 = {c2043};
    assign in2143_2 = {c2044};
    Half_Adder KS_2143(s2143, c2143, in2143_1, in2143_2);
    wire[1:0] s2144, in2144_1, in2144_2;
    wire c2144;
    assign in2144_1 = {c2045,s374[1]};
    assign in2144_2 = {c2046,c375};
    CLA_2 KS_2144(s2144, c2144, in2144_1, in2144_2);
    wire[0:0] s2145, in2145_1, in2145_2;
    wire c2145;
    assign in2145_1 = {c2047};
    assign in2145_2 = {c2048};
    Half_Adder KS_2145(s2145, c2145, in2145_1, in2145_2);
    wire[2:0] s2146, in2146_1, in2146_2;
    wire c2146;
    assign in2146_1 = {c2049,s2101[1],s362[2]};
    assign in2146_2 = {c2050,s2102[1],c364};
    CLA_3 KS_2146(s2146, c2146, in2146_1, in2146_2);
    wire[0:0] s2147, in2147_1, in2147_2;
    wire c2147;
    assign in2147_1 = {c2051};
    assign in2147_2 = {c2052};
    Half_Adder KS_2147(s2147, c2147, in2147_1, in2147_2);
    wire[1:0] s2148, in2148_1, in2148_2;
    wire c2148;
    assign in2148_1 = {c2053,s2103[1]};
    assign in2148_2 = {c2054,s2104[1]};
    CLA_2 KS_2148(s2148, c2148, in2148_1, in2148_2);
    wire[0:0] s2149, in2149_1, in2149_2;
    wire c2149;
    assign in2149_1 = {c2055};
    assign in2149_2 = {c2056};
    Half_Adder KS_2149(s2149, c2149, in2149_1, in2149_2);
    wire[3:0] s2150, in2150_1, in2150_2;
    wire c2150;
    assign in2150_1 = {c2057,s2105[1],s366[2],s409[0]};
    assign in2150_2 = {c2058,s2106[1],c368,s410[0]};
    CLA_4 KS_2150(s2150, c2150, in2150_1, in2150_2);
    wire[0:0] s2151, in2151_1, in2151_2;
    wire c2151;
    assign in2151_1 = {c2059};
    assign in2151_2 = {c2060};
    Half_Adder KS_2151(s2151, c2151, in2151_1, in2151_2);
    wire[1:0] s2152, in2152_1, in2152_2;
    wire c2152;
    assign in2152_1 = {c2061,s2107[1]};
    assign in2152_2 = {c2062,s2108[1]};
    CLA_2 KS_2152(s2152, c2152, in2152_1, in2152_2);
    wire[0:0] s2153, in2153_1, in2153_2;
    wire c2153;
    assign in2153_1 = {c2063};
    assign in2153_2 = {c2064};
    Half_Adder KS_2153(s2153, c2153, in2153_1, in2153_2);
    wire[2:0] s2154, in2154_1, in2154_2;
    wire c2154;
    assign in2154_1 = {c2065,s2109[1],s370[2]};
    assign in2154_2 = {c2068,s2110[1],c372};
    CLA_3 KS_2154(s2154, c2154, in2154_1, in2154_2);
    wire[0:0] s2155, in2155_1, in2155_2;
    wire c2155;
    assign in2155_1 = {c2076};
    assign in2155_2 = {c2084};
    Half_Adder KS_2155(s2155, c2155, in2155_1, in2155_2);
    wire[1:0] s2156, in2156_1, in2156_2;
    wire c2156;
    assign in2156_1 = {c2092,s2111[1]};
    assign in2156_2 = {c2100,s2112[1]};
    CLA_2 KS_2156(s2156, c2156, in2156_1, in2156_2);
    wire[0:0] s2157, in2157_1, in2157_2;
    wire c2157;
    assign in2157_1 = {s2101[0]};
    assign in2157_2 = {s2102[0]};
    Half_Adder KS_2157(s2157, c2157, in2157_1, in2157_2);
    wire[3:0] s2158, in2158_1, in2158_2;
    wire c2158;
    assign in2158_1 = {s2103[0],s2113[1],s374[2],s411[0]};
    assign in2158_2 = {s2104[0],s2114[1],s2101[2],s412[0]};
    CLA_4 KS_2158(s2158, c2158, in2158_1, in2158_2);
    wire[0:0] s2159, in2159_1, in2159_2;
    wire c2159;
    assign in2159_1 = {s2105[0]};
    assign in2159_2 = {s2106[0]};
    Half_Adder KS_2159(s2159, c2159, in2159_1, in2159_2);
    wire[1:0] s2160, in2160_1, in2160_2;
    wire c2160;
    assign in2160_1 = {s2107[0],s2115[1]};
    assign in2160_2 = {s2108[0],s2116[1]};
    CLA_2 KS_2160(s2160, c2160, in2160_1, in2160_2);
    wire[0:0] s2161, in2161_1, in2161_2;
    wire c2161;
    assign in2161_1 = {s2109[0]};
    assign in2161_2 = {s2110[0]};
    Half_Adder KS_2161(s2161, c2161, in2161_1, in2161_2);
    wire[2:0] s2162, in2162_1, in2162_2;
    wire c2162;
    assign in2162_1 = {s2111[0],s2117[1],s2102[2]};
    assign in2162_2 = {s2112[0],s2118[1],s2103[2]};
    CLA_3 KS_2162(s2162, c2162, in2162_1, in2162_2);
    wire[0:0] s2163, in2163_1, in2163_2;
    wire c2163;
    assign in2163_1 = {s2113[0]};
    assign in2163_2 = {s2114[0]};
    Half_Adder KS_2163(s2163, c2163, in2163_1, in2163_2);
    wire[1:0] s2164, in2164_1, in2164_2;
    wire c2164;
    assign in2164_1 = {s2115[0],s2119[1]};
    assign in2164_2 = {s2116[0],s2120[1]};
    CLA_2 KS_2164(s2164, c2164, in2164_1, in2164_2);
    wire[0:0] s2165, in2165_1, in2165_2;
    wire c2165;
    assign in2165_1 = {s2117[0]};
    assign in2165_2 = {s2118[0]};
    Half_Adder KS_2165(s2165, c2165, in2165_1, in2165_2);
    wire[3:0] s2166, in2166_1, in2166_2;
    wire c2166;
    assign in2166_1 = {s2120[0],s2121[1],s2104[2],s413[0]};
    assign in2166_2 = {s2121[0],s2122[1],s2105[2],s414[0]};
    CLA_4_c KS_2166(s2166, c2166, in2166_1, in2166_2, s2119[0]);
    wire[3:0] s2167, in2167_1, in2167_2;
    wire c2167;
    assign in2167_1 = {c350,pp116[5],pp106[16],s449[0]};
    assign in2167_2 = {c354,pp117[4],pp107[15],s450[0]};
    CLA_4 KS_2167(s2167, c2167, in2167_1, in2167_2);
    wire[3:0] s2168, in2168_1, in2168_2;
    wire c2168;
    assign in2168_1 = {c358,pp118[3],pp108[14],s451[0]};
    assign in2168_2 = {c362,pp119[2],pp109[13],s452[0]};
    CLA_4 KS_2168(s2168, c2168, in2168_1, in2168_2);
    wire[3:0] s2169, in2169_1, in2169_2;
    wire c2169;
    assign in2169_1 = {c366,pp120[1],pp110[12],s453[0]};
    assign in2169_2 = {c370,pp121[0],pp111[11],s454[0]};
    CLA_4 KS_2169(s2169, c2169, in2169_1, in2169_2);
    wire[3:0] s2170, in2170_1, in2170_2;
    wire c2170;
    assign in2170_1 = {c374,s376[2],pp112[10],s455[0]};
    assign in2170_2 = {s376[1],s377[2],pp113[9],s456[0]};
    CLA_4 KS_2170(s2170, c2170, in2170_1, in2170_2);
    wire[3:0] s2171, in2171_1, in2171_2;
    wire c2171;
    assign in2171_1 = {s377[1],s378[2],pp114[8],s457[0]};
    assign in2171_2 = {s378[1],s379[2],pp115[7],s458[0]};
    CLA_4 KS_2171(s2171, c2171, in2171_1, in2171_2);
    wire[3:0] s2172, in2172_1, in2172_2;
    wire c2172;
    assign in2172_1 = {s379[1],s380[2],pp116[6],s459[0]};
    assign in2172_2 = {s380[1],s381[2],pp117[5],s460[0]};
    CLA_4 KS_2172(s2172, c2172, in2172_1, in2172_2);
    wire[3:0] s2173, in2173_1, in2173_2;
    wire c2173;
    assign in2173_1 = {s381[1],s382[2],pp118[4],s461[0]};
    assign in2173_2 = {s382[1],s383[2],pp119[3],s462[0]};
    CLA_4 KS_2173(s2173, c2173, in2173_1, in2173_2);
    wire[3:0] s2174, in2174_1, in2174_2;
    wire c2174;
    assign in2174_1 = {s383[1],s384[2],pp120[2],s463[0]};
    assign in2174_2 = {s384[1],s385[2],pp121[1],s464[0]};
    CLA_4 KS_2174(s2174, c2174, in2174_1, in2174_2);
    wire[3:0] s2175, in2175_1, in2175_2;
    wire c2175;
    assign in2175_1 = {s385[1],s386[2],pp122[0],s465[0]};
    assign in2175_2 = {s386[1],s387[2],s376[3],s466[0]};
    CLA_4 KS_2175(s2175, c2175, in2175_1, in2175_2);
    wire[3:0] s2176, in2176_1, in2176_2;
    wire c2176;
    assign in2176_1 = {s387[1],s388[2],s377[3],s467[0]};
    assign in2176_2 = {s388[1],s389[2],s378[3],s468[0]};
    CLA_4 KS_2176(s2176, c2176, in2176_1, in2176_2);
    wire[3:0] s2177, in2177_1, in2177_2;
    wire c2177;
    assign in2177_1 = {s389[1],s390[2],s379[3],s469[0]};
    assign in2177_2 = {s390[1],s391[2],s380[3],s470[0]};
    CLA_4 KS_2177(s2177, c2177, in2177_1, in2177_2);
    wire[3:0] s2178, in2178_1, in2178_2;
    wire c2178;
    assign in2178_1 = {s391[1],s392[2],s381[3],s471[0]};
    assign in2178_2 = {s392[1],s393[2],s382[3],s472[0]};
    CLA_4 KS_2178(s2178, c2178, in2178_1, in2178_2);
    wire[3:0] s2179, in2179_1, in2179_2;
    wire c2179;
    assign in2179_1 = {s393[1],s394[2],s383[3],s473[0]};
    assign in2179_2 = {s394[1],s395[2],s384[3],s474[0]};
    CLA_4 KS_2179(s2179, c2179, in2179_1, in2179_2);
    wire[3:0] s2180, in2180_1, in2180_2;
    wire c2180;
    assign in2180_1 = {s395[1],s396[2],s385[3],s475[0]};
    assign in2180_2 = {s396[1],s397[2],s386[3],s476[0]};
    CLA_4 KS_2180(s2180, c2180, in2180_1, in2180_2);
    wire[3:0] s2181, in2181_1, in2181_2;
    wire c2181;
    assign in2181_1 = {s397[1],s398[2],s387[3],s477[0]};
    assign in2181_2 = {s398[1],s399[2],s388[3],s478[0]};
    CLA_4 KS_2181(s2181, c2181, in2181_1, in2181_2);
    wire[3:0] s2182, in2182_1, in2182_2;
    wire c2182;
    assign in2182_1 = {s399[1],s400[2],s389[3],s479[0]};
    assign in2182_2 = {s400[1],s401[2],s390[3],s480[0]};
    CLA_4 KS_2182(s2182, c2182, in2182_1, in2182_2);
    wire[3:0] s2183, in2183_1, in2183_2;
    wire c2183;
    assign in2183_1 = {s401[1],s402[2],s391[3],s481[0]};
    assign in2183_2 = {s402[1],s403[2],s392[3],s482[0]};
    CLA_4 KS_2183(s2183, c2183, in2183_1, in2183_2);
    wire[3:0] s2184, in2184_1, in2184_2;
    wire c2184;
    assign in2184_1 = {s403[1],s404[2],s393[3],s483[0]};
    assign in2184_2 = {s404[1],s405[2],s394[3],s484[0]};
    CLA_4 KS_2184(s2184, c2184, in2184_1, in2184_2);
    wire[3:0] s2185, in2185_1, in2185_2;
    wire c2185;
    assign in2185_1 = {s405[1],s406[2],s395[3],s485[0]};
    assign in2185_2 = {s406[1],s407[2],s396[3],s486[0]};
    CLA_4 KS_2185(s2185, c2185, in2185_1, in2185_2);
    wire[3:0] s2186, in2186_1, in2186_2;
    wire c2186;
    assign in2186_1 = {s407[1],s408[2],s397[3],s487[0]};
    assign in2186_2 = {s408[1],s409[2],s398[3],s488[0]};
    CLA_4 KS_2186(s2186, c2186, in2186_1, in2186_2);
    wire[3:0] s2187, in2187_1, in2187_2;
    wire c2187;
    assign in2187_1 = {s409[1],s410[2],s399[3],s489[0]};
    assign in2187_2 = {s410[1],s411[2],s400[3],s490[0]};
    CLA_4 KS_2187(s2187, c2187, in2187_1, in2187_2);
    wire[3:0] s2188, in2188_1, in2188_2;
    wire c2188;
    assign in2188_1 = {s411[1],s412[2],s401[3],s491[0]};
    assign in2188_2 = {s412[1],s413[2],s402[3],s492[0]};
    CLA_4 KS_2188(s2188, c2188, in2188_1, in2188_2);
    wire[3:0] s2189, in2189_1, in2189_2;
    wire c2189;
    assign in2189_1 = {s413[1],s414[2],s403[3],s493[0]};
    assign in2189_2 = {s414[1],s415[2],s404[3],s494[0]};
    CLA_4 KS_2189(s2189, c2189, in2189_1, in2189_2);
    wire[3:0] s2190, in2190_1, in2190_2;
    wire c2190;
    assign in2190_1 = {s415[1],s416[2],s405[3],s495[0]};
    assign in2190_2 = {s416[1],s417[2],s406[3],s496[0]};
    CLA_4 KS_2190(s2190, c2190, in2190_1, in2190_2);
    wire[3:0] s2191, in2191_1, in2191_2;
    wire c2191;
    assign in2191_1 = {s417[1],s418[2],s407[3],s497[0]};
    assign in2191_2 = {s418[1],s419[1],s408[3],s498[0]};
    CLA_4 KS_2191(s2191, c2191, in2191_1, in2191_2);
    wire[3:0] s2192, in2192_1, in2192_2;
    wire c2192;
    assign in2192_1 = {s419[0],s420[1],s409[3],s499[0]};
    assign in2192_2 = {s420[0],s421[1],s410[3],s500[0]};
    CLA_4 KS_2192(s2192, c2192, in2192_1, in2192_2);
    wire[3:0] s2193, in2193_1, in2193_2;
    wire c2193;
    assign in2193_1 = {s421[0],s422[1],s411[3],s501[0]};
    assign in2193_2 = {s422[0],c423,s412[3],s502[0]};
    CLA_4 KS_2193(s2193, c2193, in2193_1, in2193_2);
    wire[3:0] s2194, in2194_1, in2194_2;
    wire c2194;
    assign in2194_1 = {s423[0],s424[1],s413[3],s503[0]};
    assign in2194_2 = {s424[0],c425,s414[3],s504[0]};
    CLA_4 KS_2194(s2194, c2194, in2194_1, in2194_2);
    wire[3:0] s2195, in2195_1, in2195_2;
    wire c2195;
    assign in2195_1 = {s425[0],s426[1],s415[3],s505[0]};
    assign in2195_2 = {s426[0],c427,s416[3],s506[0]};
    CLA_4 KS_2195(s2195, c2195, in2195_1, in2195_2);
    wire[3:0] s2196, in2196_1, in2196_2;
    wire c2196;
    assign in2196_1 = {s427[0],s428[1],s417[3],s507[0]};
    assign in2196_2 = {s428[0],c429,s418[3],s508[0]};
    CLA_4 KS_2196(s2196, c2196, in2196_1, in2196_2);
    wire[3:0] s2197, in2197_1, in2197_2;
    wire c2197;
    assign in2197_1 = {s429[0],s430[1],s419[2],s509[0]};
    assign in2197_2 = {s430[0],c431,s420[2],s510[0]};
    CLA_4 KS_2197(s2197, c2197, in2197_1, in2197_2);
    wire[0:0] s2198, in2198_1, in2198_2;
    wire c2198;
    assign in2198_1 = {s431[0]};
    assign in2198_2 = {s432[0]};
    Half_Adder KS_2198(s2198, c2198, in2198_1, in2198_2);
    wire[1:0] s2199, in2199_1, in2199_2;
    wire c2199;
    assign in2199_1 = {s433[0],s432[1]};
    assign in2199_2 = {s434[0],c433};
    CLA_2 KS_2199(s2199, c2199, in2199_1, in2199_2);
    wire[0:0] s2200, in2200_1, in2200_2;
    wire c2200;
    assign in2200_1 = {s435[0]};
    assign in2200_2 = {s436[0]};
    Half_Adder KS_2200(s2200, c2200, in2200_1, in2200_2);
    wire[3:0] s2201, in2201_1, in2201_2;
    wire c2201;
    assign in2201_1 = {s437[0],s434[1],s421[2],s511[0]};
    assign in2201_2 = {s438[0],c435,s422[2],s512[0]};
    CLA_4 KS_2201(s2201, c2201, in2201_1, in2201_2);
    wire[0:0] s2202, in2202_1, in2202_2;
    wire c2202;
    assign in2202_1 = {s439[0]};
    assign in2202_2 = {s440[0]};
    Half_Adder KS_2202(s2202, c2202, in2202_1, in2202_2);
    wire[1:0] s2203, in2203_1, in2203_2;
    wire c2203;
    assign in2203_1 = {s441[0],s436[1]};
    assign in2203_2 = {s442[0],c437};
    CLA_2 KS_2203(s2203, c2203, in2203_1, in2203_2);
    wire[0:0] s2204, in2204_1, in2204_2;
    wire c2204;
    assign in2204_1 = {s443[0]};
    assign in2204_2 = {s444[0]};
    Half_Adder KS_2204(s2204, c2204, in2204_1, in2204_2);
    wire[2:0] s2205, in2205_1, in2205_2;
    wire c2205;
    assign in2205_1 = {c2101,s438[1],s424[2]};
    assign in2205_2 = {c2102,c439,c426};
    CLA_3 KS_2205(s2205, c2205, in2205_1, in2205_2);
    wire[0:0] s2206, in2206_1, in2206_2;
    wire c2206;
    assign in2206_1 = {c2103};
    assign in2206_2 = {c2104};
    Half_Adder KS_2206(s2206, c2206, in2206_1, in2206_2);
    wire[1:0] s2207, in2207_1, in2207_2;
    wire c2207;
    assign in2207_1 = {c2105,s440[1]};
    assign in2207_2 = {c2106,c441};
    CLA_2 KS_2207(s2207, c2207, in2207_1, in2207_2);
    wire[0:0] s2208, in2208_1, in2208_2;
    wire c2208;
    assign in2208_1 = {c2107};
    assign in2208_2 = {c2108};
    Half_Adder KS_2208(s2208, c2208, in2208_1, in2208_2);
    wire[3:0] s2209, in2209_1, in2209_2;
    wire c2209;
    assign in2209_1 = {c2109,s442[1],s428[2],s513[0]};
    assign in2209_2 = {c2110,c443,c430,s514[0]};
    CLA_4 KS_2209(s2209, c2209, in2209_1, in2209_2);
    wire[0:0] s2210, in2210_1, in2210_2;
    wire c2210;
    assign in2210_1 = {c2111};
    assign in2210_2 = {c2112};
    Half_Adder KS_2210(s2210, c2210, in2210_1, in2210_2);
    wire[1:0] s2211, in2211_1, in2211_2;
    wire c2211;
    assign in2211_1 = {c2113,s444[1]};
    assign in2211_2 = {c2114,s2167[1]};
    CLA_2 KS_2211(s2211, c2211, in2211_1, in2211_2);
    wire[0:0] s2212, in2212_1, in2212_2;
    wire c2212;
    assign in2212_1 = {c2115};
    assign in2212_2 = {c2116};
    Half_Adder KS_2212(s2212, c2212, in2212_1, in2212_2);
    wire[2:0] s2213, in2213_1, in2213_2;
    wire c2213;
    assign in2213_1 = {c2117,s2168[1],s432[2]};
    assign in2213_2 = {c2118,s2169[1],c434};
    CLA_3 KS_2213(s2213, c2213, in2213_1, in2213_2);
    wire[0:0] s2214, in2214_1, in2214_2;
    wire c2214;
    assign in2214_1 = {c2119};
    assign in2214_2 = {c2120};
    Half_Adder KS_2214(s2214, c2214, in2214_1, in2214_2);
    wire[1:0] s2215, in2215_1, in2215_2;
    wire c2215;
    assign in2215_1 = {c2121,s2170[1]};
    assign in2215_2 = {c2122,s2171[1]};
    CLA_2 KS_2215(s2215, c2215, in2215_1, in2215_2);
    wire[0:0] s2216, in2216_1, in2216_2;
    wire c2216;
    assign in2216_1 = {c2123};
    assign in2216_2 = {c2124};
    Half_Adder KS_2216(s2216, c2216, in2216_1, in2216_2);
    wire[3:0] s2217, in2217_1, in2217_2;
    wire c2217;
    assign in2217_1 = {c2125,s2172[1],s436[2],s515[0]};
    assign in2217_2 = {c2126,s2173[1],c438,s516[0]};
    CLA_4 KS_2217(s2217, c2217, in2217_1, in2217_2);
    wire[0:0] s2218, in2218_1, in2218_2;
    wire c2218;
    assign in2218_1 = {c2127};
    assign in2218_2 = {c2128};
    Half_Adder KS_2218(s2218, c2218, in2218_1, in2218_2);
    wire[1:0] s2219, in2219_1, in2219_2;
    wire c2219;
    assign in2219_1 = {c2129,s2174[1]};
    assign in2219_2 = {c2130,s2175[1]};
    CLA_2 KS_2219(s2219, c2219, in2219_1, in2219_2);
    wire[0:0] s2220, in2220_1, in2220_2;
    wire c2220;
    assign in2220_1 = {c2131};
    assign in2220_2 = {c2134};
    Half_Adder KS_2220(s2220, c2220, in2220_1, in2220_2);
    wire[2:0] s2221, in2221_1, in2221_2;
    wire c2221;
    assign in2221_1 = {c2142,s2176[1],s440[2]};
    assign in2221_2 = {c2150,s2177[1],c442};
    CLA_3 KS_2221(s2221, c2221, in2221_1, in2221_2);
    wire[0:0] s2222, in2222_1, in2222_2;
    wire c2222;
    assign in2222_1 = {c2158};
    assign in2222_2 = {c2166};
    Half_Adder KS_2222(s2222, c2222, in2222_1, in2222_2);
    wire[1:0] s2223, in2223_1, in2223_2;
    wire c2223;
    assign in2223_1 = {s2167[0],s2178[1]};
    assign in2223_2 = {s2168[0],s2179[1]};
    CLA_2 KS_2223(s2223, c2223, in2223_1, in2223_2);
    wire[0:0] s2224, in2224_1, in2224_2;
    wire c2224;
    assign in2224_1 = {s2169[0]};
    assign in2224_2 = {s2170[0]};
    Half_Adder KS_2224(s2224, c2224, in2224_1, in2224_2);
    wire[3:0] s2225, in2225_1, in2225_2;
    wire c2225;
    assign in2225_1 = {s2171[0],s2180[1],s444[2],s517[0]};
    assign in2225_2 = {s2172[0],s2181[1],s2167[2],s518[0]};
    CLA_4 KS_2225(s2225, c2225, in2225_1, in2225_2);
    wire[0:0] s2226, in2226_1, in2226_2;
    wire c2226;
    assign in2226_1 = {s2173[0]};
    assign in2226_2 = {s2174[0]};
    Half_Adder KS_2226(s2226, c2226, in2226_1, in2226_2);
    wire[1:0] s2227, in2227_1, in2227_2;
    wire c2227;
    assign in2227_1 = {s2175[0],s2182[1]};
    assign in2227_2 = {s2176[0],s2183[1]};
    CLA_2 KS_2227(s2227, c2227, in2227_1, in2227_2);
    wire[0:0] s2228, in2228_1, in2228_2;
    wire c2228;
    assign in2228_1 = {s2177[0]};
    assign in2228_2 = {s2178[0]};
    Half_Adder KS_2228(s2228, c2228, in2228_1, in2228_2);
    wire[2:0] s2229, in2229_1, in2229_2;
    wire c2229;
    assign in2229_1 = {s2179[0],s2184[1],s2168[2]};
    assign in2229_2 = {s2180[0],s2185[1],s2169[2]};
    CLA_3 KS_2229(s2229, c2229, in2229_1, in2229_2);
    wire[0:0] s2230, in2230_1, in2230_2;
    wire c2230;
    assign in2230_1 = {s2181[0]};
    assign in2230_2 = {s2182[0]};
    Half_Adder KS_2230(s2230, c2230, in2230_1, in2230_2);
    wire[1:0] s2231, in2231_1, in2231_2;
    wire c2231;
    assign in2231_1 = {s2183[0],s2186[1]};
    assign in2231_2 = {s2184[0],s2187[1]};
    CLA_2 KS_2231(s2231, c2231, in2231_1, in2231_2);
    wire[0:0] s2232, in2232_1, in2232_2;
    wire c2232;
    assign in2232_1 = {s2186[0]};
    assign in2232_2 = {s2187[0]};
    Full_Adder KS_2232(s2232, c2232, in2232_1, in2232_2, s2185[0]);
    wire[3:0] s2233, in2233_1, in2233_2;
    wire c2233;
    assign in2233_1 = {s450[1],pp120[5],pp112[14],s556[0]};
    assign in2233_2 = {s451[1],pp121[4],pp113[13],s557[0]};
    CLA_4 KS_2233(s2233, c2233, in2233_1, in2233_2);
    wire[3:0] s2234, in2234_1, in2234_2;
    wire c2234;
    assign in2234_1 = {s452[1],pp122[3],pp114[12],s558[0]};
    assign in2234_2 = {s453[1],pp123[2],pp115[11],s559[0]};
    CLA_4 KS_2234(s2234, c2234, in2234_1, in2234_2);
    wire[3:0] s2235, in2235_1, in2235_2;
    wire c2235;
    assign in2235_1 = {s454[1],pp124[1],pp116[10],s560[0]};
    assign in2235_2 = {s455[1],pp125[0],pp117[9],s561[0]};
    CLA_4 KS_2235(s2235, c2235, in2235_1, in2235_2);
    wire[3:0] s2236, in2236_1, in2236_2;
    wire c2236;
    assign in2236_1 = {s456[1],s445[2],pp118[8],s562[0]};
    assign in2236_2 = {s457[1],s446[2],pp119[7],s563[0]};
    CLA_4 KS_2236(s2236, c2236, in2236_1, in2236_2);
    wire[3:0] s2237, in2237_1, in2237_2;
    wire c2237;
    assign in2237_1 = {s458[1],s447[2],pp120[6],s564[0]};
    assign in2237_2 = {s459[1],s448[2],pp121[5],s565[0]};
    CLA_4 KS_2237(s2237, c2237, in2237_1, in2237_2);
    wire[3:0] s2238, in2238_1, in2238_2;
    wire c2238;
    assign in2238_1 = {s460[1],s449[2],pp122[4],s566[0]};
    assign in2238_2 = {s461[1],s450[2],pp123[3],s567[0]};
    CLA_4 KS_2238(s2238, c2238, in2238_1, in2238_2);
    wire[3:0] s2239, in2239_1, in2239_2;
    wire c2239;
    assign in2239_1 = {s462[1],s451[2],pp124[2],s568[0]};
    assign in2239_2 = {s463[1],s452[2],pp125[1],s569[0]};
    CLA_4 KS_2239(s2239, c2239, in2239_1, in2239_2);
    wire[3:0] s2240, in2240_1, in2240_2;
    wire c2240;
    assign in2240_1 = {s464[1],s453[2],pp126[0],s570[0]};
    assign in2240_2 = {s465[1],s454[2],s445[3],s571[0]};
    CLA_4 KS_2240(s2240, c2240, in2240_1, in2240_2);
    wire[3:0] s2241, in2241_1, in2241_2;
    wire c2241;
    assign in2241_1 = {s466[1],s455[2],s446[3],s572[0]};
    assign in2241_2 = {s467[1],s456[2],s447[3],s573[0]};
    CLA_4 KS_2241(s2241, c2241, in2241_1, in2241_2);
    wire[3:0] s2242, in2242_1, in2242_2;
    wire c2242;
    assign in2242_1 = {s468[1],s457[2],s448[3],s574[0]};
    assign in2242_2 = {s469[1],s458[2],s449[3],s575[0]};
    CLA_4 KS_2242(s2242, c2242, in2242_1, in2242_2);
    wire[3:0] s2243, in2243_1, in2243_2;
    wire c2243;
    assign in2243_1 = {s470[1],s459[2],s450[3],s576[0]};
    assign in2243_2 = {s471[1],s460[2],s451[3],s577[0]};
    CLA_4 KS_2243(s2243, c2243, in2243_1, in2243_2);
    wire[3:0] s2244, in2244_1, in2244_2;
    wire c2244;
    assign in2244_1 = {s472[1],s461[2],s452[3],s578[0]};
    assign in2244_2 = {s473[1],s462[2],s453[3],s579[0]};
    CLA_4 KS_2244(s2244, c2244, in2244_1, in2244_2);
    wire[3:0] s2245, in2245_1, in2245_2;
    wire c2245;
    assign in2245_1 = {s474[1],s463[2],s454[3],s580[0]};
    assign in2245_2 = {s475[1],s464[2],s455[3],s581[0]};
    CLA_4 KS_2245(s2245, c2245, in2245_1, in2245_2);
    wire[3:0] s2246, in2246_1, in2246_2;
    wire c2246;
    assign in2246_1 = {s476[1],s465[2],s456[3],s582[0]};
    assign in2246_2 = {s477[1],s466[2],s457[3],s583[0]};
    CLA_4 KS_2246(s2246, c2246, in2246_1, in2246_2);
    wire[3:0] s2247, in2247_1, in2247_2;
    wire c2247;
    assign in2247_1 = {s478[1],s467[2],s458[3],s584[0]};
    assign in2247_2 = {s479[1],s468[2],s459[3],s585[0]};
    CLA_4 KS_2247(s2247, c2247, in2247_1, in2247_2);
    wire[3:0] s2248, in2248_1, in2248_2;
    wire c2248;
    assign in2248_1 = {s480[1],s469[2],s460[3],s586[0]};
    assign in2248_2 = {s481[1],s470[2],s461[3],s587[0]};
    CLA_4 KS_2248(s2248, c2248, in2248_1, in2248_2);
    wire[3:0] s2249, in2249_1, in2249_2;
    wire c2249;
    assign in2249_1 = {s482[1],s471[2],s462[3],s588[0]};
    assign in2249_2 = {s483[1],s472[2],s463[3],s589[0]};
    CLA_4 KS_2249(s2249, c2249, in2249_1, in2249_2);
    wire[3:0] s2250, in2250_1, in2250_2;
    wire c2250;
    assign in2250_1 = {s484[1],s473[2],s464[3],s590[0]};
    assign in2250_2 = {s485[1],s474[2],s465[3],s591[0]};
    CLA_4 KS_2250(s2250, c2250, in2250_1, in2250_2);
    wire[3:0] s2251, in2251_1, in2251_2;
    wire c2251;
    assign in2251_1 = {s486[1],s475[2],s466[3],s592[0]};
    assign in2251_2 = {s487[1],s476[2],s467[3],s593[0]};
    CLA_4 KS_2251(s2251, c2251, in2251_1, in2251_2);
    wire[3:0] s2252, in2252_1, in2252_2;
    wire c2252;
    assign in2252_1 = {s488[1],s477[2],s468[3],s594[0]};
    assign in2252_2 = {s489[1],s478[2],s469[3],s595[0]};
    CLA_4 KS_2252(s2252, c2252, in2252_1, in2252_2);
    wire[3:0] s2253, in2253_1, in2253_2;
    wire c2253;
    assign in2253_1 = {s490[1],s479[2],s470[3],s596[0]};
    assign in2253_2 = {s491[1],s480[2],s471[3],s597[0]};
    CLA_4 KS_2253(s2253, c2253, in2253_1, in2253_2);
    wire[3:0] s2254, in2254_1, in2254_2;
    wire c2254;
    assign in2254_1 = {s492[1],s481[2],s472[3],s598[0]};
    assign in2254_2 = {s493[1],s482[2],s473[3],s599[0]};
    CLA_4 KS_2254(s2254, c2254, in2254_1, in2254_2);
    wire[3:0] s2255, in2255_1, in2255_2;
    wire c2255;
    assign in2255_1 = {s494[1],s483[2],s474[3],s600[0]};
    assign in2255_2 = {s495[1],s484[2],s475[3],s601[0]};
    CLA_4 KS_2255(s2255, c2255, in2255_1, in2255_2);
    wire[3:0] s2256, in2256_1, in2256_2;
    wire c2256;
    assign in2256_1 = {s496[1],s485[2],s476[3],s602[0]};
    assign in2256_2 = {s497[1],s486[2],s477[3],s603[0]};
    CLA_4 KS_2256(s2256, c2256, in2256_1, in2256_2);
    wire[3:0] s2257, in2257_1, in2257_2;
    wire c2257;
    assign in2257_1 = {s498[1],s487[2],s478[3],s604[0]};
    assign in2257_2 = {s499[1],s488[2],s479[3],s605[0]};
    CLA_4 KS_2257(s2257, c2257, in2257_1, in2257_2);
    wire[3:0] s2258, in2258_1, in2258_2;
    wire c2258;
    assign in2258_1 = {s500[1],s489[2],s480[3],s606[0]};
    assign in2258_2 = {s501[1],s490[2],s481[3],s607[0]};
    CLA_4 KS_2258(s2258, c2258, in2258_1, in2258_2);
    wire[3:0] s2259, in2259_1, in2259_2;
    wire c2259;
    assign in2259_1 = {s502[1],s491[2],s482[3],s608[0]};
    assign in2259_2 = {s503[1],s492[2],s483[3],s609[0]};
    CLA_4 KS_2259(s2259, c2259, in2259_1, in2259_2);
    wire[3:0] s2260, in2260_1, in2260_2;
    wire c2260;
    assign in2260_1 = {s504[1],s493[2],s484[3],s610[0]};
    assign in2260_2 = {c505,s494[2],s485[3],s611[0]};
    CLA_4 KS_2260(s2260, c2260, in2260_1, in2260_2);
    wire[3:0] s2261, in2261_1, in2261_2;
    wire c2261;
    assign in2261_1 = {s506[1],s495[2],s486[3],s612[0]};
    assign in2261_2 = {c507,c496,s487[3],s613[0]};
    CLA_4 KS_2261(s2261, c2261, in2261_1, in2261_2);
    wire[3:0] s2262, in2262_1, in2262_2;
    wire c2262;
    assign in2262_1 = {s508[1],s497[2],s488[3],s614[0]};
    assign in2262_2 = {c509,c498,s489[3],s615[0]};
    CLA_4 KS_2262(s2262, c2262, in2262_1, in2262_2);
    wire[3:0] s2263, in2263_1, in2263_2;
    wire c2263;
    assign in2263_1 = {s510[1],s499[2],s490[3],s616[0]};
    assign in2263_2 = {c511,c500,s491[3],s617[0]};
    CLA_4 KS_2263(s2263, c2263, in2263_1, in2263_2);
    wire[1:0] s2264, in2264_1, in2264_2;
    wire c2264;
    assign in2264_1 = {s512[1],s501[2]};
    assign in2264_2 = {c513,c502};
    CLA_2 KS_2264(s2264, c2264, in2264_1, in2264_2);
    wire[0:0] s2265, in2265_1, in2265_2;
    wire c2265;
    assign in2265_1 = {s514[1]};
    assign in2265_2 = {c515};
    Half_Adder KS_2265(s2265, c2265, in2265_1, in2265_2);
    wire[3:0] s2266, in2266_1, in2266_2;
    wire c2266;
    assign in2266_1 = {s516[1],s503[2],s492[3],s618[0]};
    assign in2266_2 = {c517,c504,s493[3],s619[0]};
    CLA_4 KS_2266(s2266, c2266, in2266_1, in2266_2);
    wire[0:0] s2267, in2267_1, in2267_2;
    wire c2267;
    assign in2267_1 = {s518[1]};
    assign in2267_2 = {c519};
    Half_Adder KS_2267(s2267, c2267, in2267_1, in2267_2);
    wire[1:0] s2268, in2268_1, in2268_2;
    wire c2268;
    assign in2268_1 = {s520[1],s506[2]};
    assign in2268_2 = {c521,c508};
    CLA_2 KS_2268(s2268, c2268, in2268_1, in2268_2);
    wire[0:0] s2269, in2269_1, in2269_2;
    wire c2269;
    assign in2269_1 = {s522[1]};
    assign in2269_2 = {c523};
    Half_Adder KS_2269(s2269, c2269, in2269_1, in2269_2);
    wire[2:0] s2270, in2270_1, in2270_2;
    wire c2270;
    assign in2270_1 = {s524[1],s510[2],s494[3]};
    assign in2270_2 = {c2167,c512,s495[3]};
    CLA_3 KS_2270(s2270, c2270, in2270_1, in2270_2);
    wire[0:0] s2271, in2271_1, in2271_2;
    wire c2271;
    assign in2271_1 = {c2168};
    assign in2271_2 = {c2169};
    Half_Adder KS_2271(s2271, c2271, in2271_1, in2271_2);
    wire[1:0] s2272, in2272_1, in2272_2;
    wire c2272;
    assign in2272_1 = {c2170,s514[2]};
    assign in2272_2 = {c2171,c516};
    CLA_2 KS_2272(s2272, c2272, in2272_1, in2272_2);
    wire[0:0] s2273, in2273_1, in2273_2;
    wire c2273;
    assign in2273_1 = {c2172};
    assign in2273_2 = {c2173};
    Half_Adder KS_2273(s2273, c2273, in2273_1, in2273_2);
    wire[3:0] s2274, in2274_1, in2274_2;
    wire c2274;
    assign in2274_1 = {c2174,s518[2],s497[3],s620[0]};
    assign in2274_2 = {c2175,c520,c499,s621[0]};
    CLA_4 KS_2274(s2274, c2274, in2274_1, in2274_2);
    wire[0:0] s2275, in2275_1, in2275_2;
    wire c2275;
    assign in2275_1 = {c2176};
    assign in2275_2 = {c2177};
    Half_Adder KS_2275(s2275, c2275, in2275_1, in2275_2);
    wire[1:0] s2276, in2276_1, in2276_2;
    wire c2276;
    assign in2276_1 = {c2178,s522[2]};
    assign in2276_2 = {c2179,c524};
    CLA_2 KS_2276(s2276, c2276, in2276_1, in2276_2);
    wire[0:0] s2277, in2277_1, in2277_2;
    wire c2277;
    assign in2277_1 = {c2180};
    assign in2277_2 = {c2181};
    Half_Adder KS_2277(s2277, c2277, in2277_1, in2277_2);
    wire[2:0] s2278, in2278_1, in2278_2;
    wire c2278;
    assign in2278_1 = {c2182,s2233[1],s501[3]};
    assign in2278_2 = {c2183,s2234[1],c503};
    CLA_3 KS_2278(s2278, c2278, in2278_1, in2278_2);
    wire[0:0] s2279, in2279_1, in2279_2;
    wire c2279;
    assign in2279_1 = {c2184};
    assign in2279_2 = {c2185};
    Half_Adder KS_2279(s2279, c2279, in2279_1, in2279_2);
    wire[1:0] s2280, in2280_1, in2280_2;
    wire c2280;
    assign in2280_1 = {c2186,s2235[1]};
    assign in2280_2 = {c2187,s2236[1]};
    CLA_2 KS_2280(s2280, c2280, in2280_1, in2280_2);
    wire[0:0] s2281, in2281_1, in2281_2;
    wire c2281;
    assign in2281_1 = {c2188};
    assign in2281_2 = {c2189};
    Half_Adder KS_2281(s2281, c2281, in2281_1, in2281_2);
    wire[3:0] s2282, in2282_1, in2282_2;
    wire c2282;
    assign in2282_1 = {c2190,s2237[1],s506[3],s622[0]};
    assign in2282_2 = {c2191,s2238[1],c510,s623[0]};
    CLA_4 KS_2282(s2282, c2282, in2282_1, in2282_2);
    wire[0:0] s2283, in2283_1, in2283_2;
    wire c2283;
    assign in2283_1 = {c2192};
    assign in2283_2 = {c2193};
    Half_Adder KS_2283(s2283, c2283, in2283_1, in2283_2);
    wire[1:0] s2284, in2284_1, in2284_2;
    wire c2284;
    assign in2284_1 = {c2194,s2239[1]};
    assign in2284_2 = {c2195,s2240[1]};
    CLA_2 KS_2284(s2284, c2284, in2284_1, in2284_2);
    wire[0:0] s2285, in2285_1, in2285_2;
    wire c2285;
    assign in2285_1 = {c2196};
    assign in2285_2 = {c2197};
    Half_Adder KS_2285(s2285, c2285, in2285_1, in2285_2);
    wire[2:0] s2286, in2286_1, in2286_2;
    wire c2286;
    assign in2286_1 = {c2201,s2241[1],s514[3]};
    assign in2286_2 = {c2209,s2242[1],c518};
    CLA_3 KS_2286(s2286, c2286, in2286_1, in2286_2);
    wire[0:0] s2287, in2287_1, in2287_2;
    wire c2287;
    assign in2287_1 = {c2217};
    assign in2287_2 = {c2225};
    Half_Adder KS_2287(s2287, c2287, in2287_1, in2287_2);
    wire[1:0] s2288, in2288_1, in2288_2;
    wire c2288;
    assign in2288_1 = {s2233[0],s2243[1]};
    assign in2288_2 = {s2234[0],s2244[1]};
    CLA_2 KS_2288(s2288, c2288, in2288_1, in2288_2);
    wire[0:0] s2289, in2289_1, in2289_2;
    wire c2289;
    assign in2289_1 = {s2235[0]};
    assign in2289_2 = {s2236[0]};
    Half_Adder KS_2289(s2289, c2289, in2289_1, in2289_2);
    wire[3:0] s2290, in2290_1, in2290_2;
    wire c2290;
    assign in2290_1 = {s2237[0],s2245[1],s522[3],s624[0]};
    assign in2290_2 = {s2238[0],s2246[1],s2233[2],s625[0]};
    CLA_4 KS_2290(s2290, c2290, in2290_1, in2290_2);
    wire[0:0] s2291, in2291_1, in2291_2;
    wire c2291;
    assign in2291_1 = {s2239[0]};
    assign in2291_2 = {s2240[0]};
    Half_Adder KS_2291(s2291, c2291, in2291_1, in2291_2);
    wire[1:0] s2292, in2292_1, in2292_2;
    wire c2292;
    assign in2292_1 = {s2241[0],s2247[1]};
    assign in2292_2 = {s2242[0],s2248[1]};
    CLA_2 KS_2292(s2292, c2292, in2292_1, in2292_2);
    wire[0:0] s2293, in2293_1, in2293_2;
    wire c2293;
    assign in2293_1 = {s2243[0]};
    assign in2293_2 = {s2244[0]};
    Half_Adder KS_2293(s2293, c2293, in2293_1, in2293_2);
    wire[2:0] s2294, in2294_1, in2294_2;
    wire c2294;
    assign in2294_1 = {s2245[0],s2249[1],s2234[2]};
    assign in2294_2 = {s2246[0],s2250[1],s2235[2]};
    CLA_3 KS_2294(s2294, c2294, in2294_1, in2294_2);
    wire[0:0] s2295, in2295_1, in2295_2;
    wire c2295;
    assign in2295_1 = {s2247[0]};
    assign in2295_2 = {s2248[0]};
    Half_Adder KS_2295(s2295, c2295, in2295_1, in2295_2);
    wire[1:0] s2296, in2296_1, in2296_2;
    wire c2296;
    assign in2296_1 = {s2250[0],s2251[1]};
    assign in2296_2 = {s2251[0],s2252[1]};
    CLA_2_c KS_2296(s2296, c2296, in2296_1, in2296_2, s2249[0]);
    wire[3:0] s2297, in2297_1, in2297_2;
    wire c2297;
    assign in2297_1 = {s557[1],s529[2],pp117[13],s660[0]};
    assign in2297_2 = {s558[1],s530[2],pp118[12],s661[0]};
    CLA_4 KS_2297(s2297, c2297, in2297_1, in2297_2);
    wire[3:0] s2298, in2298_1, in2298_2;
    wire c2298;
    assign in2298_1 = {s559[1],s531[2],pp119[11],s662[0]};
    assign in2298_2 = {s560[1],s532[2],pp120[10],s663[0]};
    CLA_4 KS_2298(s2298, c2298, in2298_1, in2298_2);
    wire[3:0] s2299, in2299_1, in2299_2;
    wire c2299;
    assign in2299_1 = {s561[1],s533[2],pp121[9],s664[0]};
    assign in2299_2 = {s562[1],s534[2],pp122[8],s665[0]};
    CLA_4 KS_2299(s2299, c2299, in2299_1, in2299_2);
    wire[3:0] s2300, in2300_1, in2300_2;
    wire c2300;
    assign in2300_1 = {s563[1],s535[2],pp123[7],s666[0]};
    assign in2300_2 = {s564[1],s536[2],pp124[6],s667[0]};
    CLA_4 KS_2300(s2300, c2300, in2300_1, in2300_2);
    wire[3:0] s2301, in2301_1, in2301_2;
    wire c2301;
    assign in2301_1 = {s565[1],s537[2],pp125[5],s668[0]};
    assign in2301_2 = {s566[1],s538[2],pp126[4],s669[0]};
    CLA_4 KS_2301(s2301, c2301, in2301_1, in2301_2);
    wire[3:0] s2302, in2302_1, in2302_2;
    wire c2302;
    assign in2302_1 = {s567[1],s539[2],pp127[3],s670[0]};
    assign in2302_2 = {s568[1],s540[2],s525[3],s671[0]};
    CLA_4 KS_2302(s2302, c2302, in2302_1, in2302_2);
    wire[3:0] s2303, in2303_1, in2303_2;
    wire c2303;
    assign in2303_1 = {s569[1],s541[2],s526[3],s672[0]};
    assign in2303_2 = {s570[1],s542[2],s527[3],s673[0]};
    CLA_4 KS_2303(s2303, c2303, in2303_1, in2303_2);
    wire[3:0] s2304, in2304_1, in2304_2;
    wire c2304;
    assign in2304_1 = {s571[1],s543[2],s528[3],s674[0]};
    assign in2304_2 = {s572[1],s544[2],s529[3],s675[0]};
    CLA_4 KS_2304(s2304, c2304, in2304_1, in2304_2);
    wire[3:0] s2305, in2305_1, in2305_2;
    wire c2305;
    assign in2305_1 = {s573[1],s545[2],s530[3],s676[0]};
    assign in2305_2 = {s574[1],s546[2],s531[3],s677[0]};
    CLA_4 KS_2305(s2305, c2305, in2305_1, in2305_2);
    wire[3:0] s2306, in2306_1, in2306_2;
    wire c2306;
    assign in2306_1 = {s575[1],s547[2],s532[3],s678[0]};
    assign in2306_2 = {s576[1],s548[2],s533[3],s679[0]};
    CLA_4 KS_2306(s2306, c2306, in2306_1, in2306_2);
    wire[3:0] s2307, in2307_1, in2307_2;
    wire c2307;
    assign in2307_1 = {s577[1],s549[2],s534[3],s680[0]};
    assign in2307_2 = {c578,s550[2],s535[3],s681[0]};
    CLA_4 KS_2307(s2307, c2307, in2307_1, in2307_2);
    wire[3:0] s2308, in2308_1, in2308_2;
    wire c2308;
    assign in2308_1 = {s579[1],s551[2],s536[3],s682[0]};
    assign in2308_2 = {c580,s552[2],s537[3],s683[0]};
    CLA_4 KS_2308(s2308, c2308, in2308_1, in2308_2);
    wire[3:0] s2309, in2309_1, in2309_2;
    wire c2309;
    assign in2309_1 = {s581[1],s553[2],s538[3],s684[0]};
    assign in2309_2 = {c582,s554[2],s539[3],s685[0]};
    CLA_4 KS_2309(s2309, c2309, in2309_1, in2309_2);
    wire[3:0] s2310, in2310_1, in2310_2;
    wire c2310;
    assign in2310_1 = {s583[1],s555[2],s540[3],s686[0]};
    assign in2310_2 = {c584,s556[2],s541[3],s687[0]};
    CLA_4 KS_2310(s2310, c2310, in2310_1, in2310_2);
    wire[3:0] s2311, in2311_1, in2311_2;
    wire c2311;
    assign in2311_1 = {s585[1],s557[2],s542[3],s688[0]};
    assign in2311_2 = {c586,s558[2],s543[3],s689[0]};
    CLA_4 KS_2311(s2311, c2311, in2311_1, in2311_2);
    wire[3:0] s2312, in2312_1, in2312_2;
    wire c2312;
    assign in2312_1 = {s587[1],s559[2],s544[3],s690[0]};
    assign in2312_2 = {c588,s560[2],s545[3],s691[0]};
    CLA_4 KS_2312(s2312, c2312, in2312_1, in2312_2);
    wire[3:0] s2313, in2313_1, in2313_2;
    wire c2313;
    assign in2313_1 = {s589[1],s561[2],s546[3],s692[0]};
    assign in2313_2 = {c590,s562[2],s547[3],s693[0]};
    CLA_4 KS_2313(s2313, c2313, in2313_1, in2313_2);
    wire[3:0] s2314, in2314_1, in2314_2;
    wire c2314;
    assign in2314_1 = {s591[1],s563[2],s548[3],s694[0]};
    assign in2314_2 = {c592,s564[2],s549[3],s695[0]};
    CLA_4 KS_2314(s2314, c2314, in2314_1, in2314_2);
    wire[3:0] s2315, in2315_1, in2315_2;
    wire c2315;
    assign in2315_1 = {s593[1],s565[2],s550[3],s696[0]};
    assign in2315_2 = {c594,s566[2],s551[3],s697[0]};
    CLA_4 KS_2315(s2315, c2315, in2315_1, in2315_2);
    wire[3:0] s2316, in2316_1, in2316_2;
    wire c2316;
    assign in2316_1 = {s595[1],s567[2],s552[3],s698[0]};
    assign in2316_2 = {c596,s568[2],s553[3],s699[0]};
    CLA_4 KS_2316(s2316, c2316, in2316_1, in2316_2);
    wire[3:0] s2317, in2317_1, in2317_2;
    wire c2317;
    assign in2317_1 = {s597[1],s569[2],s554[3],s700[0]};
    assign in2317_2 = {c598,s570[2],s555[3],s701[0]};
    CLA_4 KS_2317(s2317, c2317, in2317_1, in2317_2);
    wire[3:0] s2318, in2318_1, in2318_2;
    wire c2318;
    assign in2318_1 = {s599[1],s571[2],s556[3],s702[0]};
    assign in2318_2 = {c600,s572[2],s557[3],s703[0]};
    CLA_4 KS_2318(s2318, c2318, in2318_1, in2318_2);
    wire[3:0] s2319, in2319_1, in2319_2;
    wire c2319;
    assign in2319_1 = {s601[1],s573[2],s558[3],s704[0]};
    assign in2319_2 = {c602,s574[2],s559[3],s705[0]};
    CLA_4 KS_2319(s2319, c2319, in2319_1, in2319_2);
    wire[3:0] s2320, in2320_1, in2320_2;
    wire c2320;
    assign in2320_1 = {s603[1],s575[2],s560[3],s706[0]};
    assign in2320_2 = {c604,c576,s561[3],s707[0]};
    CLA_4 KS_2320(s2320, c2320, in2320_1, in2320_2);
    wire[3:0] s2321, in2321_1, in2321_2;
    wire c2321;
    assign in2321_1 = {s605[1],s577[2],s562[3],s708[0]};
    assign in2321_2 = {c606,c579,s563[3],s709[0]};
    CLA_4 KS_2321(s2321, c2321, in2321_1, in2321_2);
    wire[3:0] s2322, in2322_1, in2322_2;
    wire c2322;
    assign in2322_1 = {s607[1],s581[2],s564[3],s710[0]};
    assign in2322_2 = {c608,c583,s565[3],s711[0]};
    CLA_4 KS_2322(s2322, c2322, in2322_1, in2322_2);
    wire[3:0] s2323, in2323_1, in2323_2;
    wire c2323;
    assign in2323_1 = {s609[1],s585[2],s566[3],s712[0]};
    assign in2323_2 = {c610,c587,s567[3],s713[0]};
    CLA_4 KS_2323(s2323, c2323, in2323_1, in2323_2);
    wire[3:0] s2324, in2324_1, in2324_2;
    wire c2324;
    assign in2324_1 = {s611[1],s589[2],s568[3],s714[0]};
    assign in2324_2 = {c612,c591,s569[3],s715[0]};
    CLA_4 KS_2324(s2324, c2324, in2324_1, in2324_2);
    wire[3:0] s2325, in2325_1, in2325_2;
    wire c2325;
    assign in2325_1 = {s613[1],s593[2],s570[3],s716[0]};
    assign in2325_2 = {c614,c595,s571[3],s717[0]};
    CLA_4 KS_2325(s2325, c2325, in2325_1, in2325_2);
    wire[3:0] s2326, in2326_1, in2326_2;
    wire c2326;
    assign in2326_1 = {s615[1],s597[2],s572[3],s718[0]};
    assign in2326_2 = {c616,c599,s573[3],s719[0]};
    CLA_4 KS_2326(s2326, c2326, in2326_1, in2326_2);
    wire[3:0] s2327, in2327_1, in2327_2;
    wire c2327;
    assign in2327_1 = {s617[1],s601[2],s574[3],s720[0]};
    assign in2327_2 = {c618,c603,c575,s721[0]};
    CLA_4 KS_2327(s2327, c2327, in2327_1, in2327_2);
    wire[3:0] s2328, in2328_1, in2328_2;
    wire c2328;
    assign in2328_1 = {s619[1],s605[2],s577[3],s722[0]};
    assign in2328_2 = {c620,c607,c581,s723[0]};
    CLA_4 KS_2328(s2328, c2328, in2328_1, in2328_2);
    wire[0:0] s2329, in2329_1, in2329_2;
    wire c2329;
    assign in2329_1 = {s621[1]};
    assign in2329_2 = {c622};
    Half_Adder KS_2329(s2329, c2329, in2329_1, in2329_2);
    wire[1:0] s2330, in2330_1, in2330_2;
    wire c2330;
    assign in2330_1 = {s623[1],s609[2]};
    assign in2330_2 = {c624,c611};
    CLA_2 KS_2330(s2330, c2330, in2330_1, in2330_2);
    wire[0:0] s2331, in2331_1, in2331_2;
    wire c2331;
    assign in2331_1 = {s625[1]};
    assign in2331_2 = {c626};
    Half_Adder KS_2331(s2331, c2331, in2331_1, in2331_2);
    wire[2:0] s2332, in2332_1, in2332_2;
    wire c2332;
    assign in2332_1 = {s627[1],s613[2],s585[3]};
    assign in2332_2 = {c628,c615,c589};
    CLA_3 KS_2332(s2332, c2332, in2332_1, in2332_2);
    wire[0:0] s2333, in2333_1, in2333_2;
    wire c2333;
    assign in2333_1 = {s629[1]};
    assign in2333_2 = {c630};
    Half_Adder KS_2333(s2333, c2333, in2333_1, in2333_2);
    wire[1:0] s2334, in2334_1, in2334_2;
    wire c2334;
    assign in2334_1 = {s631[1],s617[2]};
    assign in2334_2 = {c2233,c619};
    CLA_2 KS_2334(s2334, c2334, in2334_1, in2334_2);
    wire[0:0] s2335, in2335_1, in2335_2;
    wire c2335;
    assign in2335_1 = {c2234};
    assign in2335_2 = {c2235};
    Half_Adder KS_2335(s2335, c2335, in2335_1, in2335_2);
    wire[3:0] s2336, in2336_1, in2336_2;
    wire c2336;
    assign in2336_1 = {c2236,s621[2],s593[3],s724[0]};
    assign in2336_2 = {c2237,c623,c597,s725[0]};
    CLA_4 KS_2336(s2336, c2336, in2336_1, in2336_2);
    wire[0:0] s2337, in2337_1, in2337_2;
    wire c2337;
    assign in2337_1 = {c2238};
    assign in2337_2 = {c2239};
    Half_Adder KS_2337(s2337, c2337, in2337_1, in2337_2);
    wire[1:0] s2338, in2338_1, in2338_2;
    wire c2338;
    assign in2338_1 = {c2240,s625[2]};
    assign in2338_2 = {c2241,c627};
    CLA_2 KS_2338(s2338, c2338, in2338_1, in2338_2);
    wire[0:0] s2339, in2339_1, in2339_2;
    wire c2339;
    assign in2339_1 = {c2242};
    assign in2339_2 = {c2243};
    Half_Adder KS_2339(s2339, c2339, in2339_1, in2339_2);
    wire[2:0] s2340, in2340_1, in2340_2;
    wire c2340;
    assign in2340_1 = {c2244,s629[2],s601[3]};
    assign in2340_2 = {c2245,c631,c605};
    CLA_3 KS_2340(s2340, c2340, in2340_1, in2340_2);
    wire[0:0] s2341, in2341_1, in2341_2;
    wire c2341;
    assign in2341_1 = {c2246};
    assign in2341_2 = {c2247};
    Half_Adder KS_2341(s2341, c2341, in2341_1, in2341_2);
    wire[1:0] s2342, in2342_1, in2342_2;
    wire c2342;
    assign in2342_1 = {c2248,s2297[1]};
    assign in2342_2 = {c2249,s2298[1]};
    CLA_2 KS_2342(s2342, c2342, in2342_1, in2342_2);
    wire[0:0] s2343, in2343_1, in2343_2;
    wire c2343;
    assign in2343_1 = {c2250};
    assign in2343_2 = {c2251};
    Half_Adder KS_2343(s2343, c2343, in2343_1, in2343_2);
    wire[3:0] s2344, in2344_1, in2344_2;
    wire c2344;
    assign in2344_1 = {c2252,s2299[1],s609[3],s726[0]};
    assign in2344_2 = {c2253,s2300[1],c613,s727[0]};
    CLA_4 KS_2344(s2344, c2344, in2344_1, in2344_2);
    wire[0:0] s2345, in2345_1, in2345_2;
    wire c2345;
    assign in2345_1 = {c2254};
    assign in2345_2 = {c2255};
    Half_Adder KS_2345(s2345, c2345, in2345_1, in2345_2);
    wire[1:0] s2346, in2346_1, in2346_2;
    wire c2346;
    assign in2346_1 = {c2256,s2301[1]};
    assign in2346_2 = {c2257,s2302[1]};
    CLA_2 KS_2346(s2346, c2346, in2346_1, in2346_2);
    wire[0:0] s2347, in2347_1, in2347_2;
    wire c2347;
    assign in2347_1 = {c2258};
    assign in2347_2 = {c2259};
    Half_Adder KS_2347(s2347, c2347, in2347_1, in2347_2);
    wire[2:0] s2348, in2348_1, in2348_2;
    wire c2348;
    assign in2348_1 = {c2260,s2303[1],s617[3]};
    assign in2348_2 = {c2261,s2304[1],c621};
    CLA_3 KS_2348(s2348, c2348, in2348_1, in2348_2);
    wire[0:0] s2349, in2349_1, in2349_2;
    wire c2349;
    assign in2349_1 = {c2262};
    assign in2349_2 = {c2263};
    Half_Adder KS_2349(s2349, c2349, in2349_1, in2349_2);
    wire[1:0] s2350, in2350_1, in2350_2;
    wire c2350;
    assign in2350_1 = {c2266,s2305[1]};
    assign in2350_2 = {c2274,s2306[1]};
    CLA_2 KS_2350(s2350, c2350, in2350_1, in2350_2);
    wire[0:0] s2351, in2351_1, in2351_2;
    wire c2351;
    assign in2351_1 = {c2282};
    assign in2351_2 = {c2290};
    Half_Adder KS_2351(s2351, c2351, in2351_1, in2351_2);
    wire[3:0] s2352, in2352_1, in2352_2;
    wire c2352;
    assign in2352_1 = {s2297[0],s2307[1],s625[3],s728[0]};
    assign in2352_2 = {s2298[0],s2308[1],c629,s729[0]};
    CLA_4 KS_2352(s2352, c2352, in2352_1, in2352_2);
    wire[0:0] s2353, in2353_1, in2353_2;
    wire c2353;
    assign in2353_1 = {s2299[0]};
    assign in2353_2 = {s2300[0]};
    Half_Adder KS_2353(s2353, c2353, in2353_1, in2353_2);
    wire[1:0] s2354, in2354_1, in2354_2;
    wire c2354;
    assign in2354_1 = {s2301[0],s2309[1]};
    assign in2354_2 = {s2302[0],s2310[1]};
    CLA_2 KS_2354(s2354, c2354, in2354_1, in2354_2);
    wire[0:0] s2355, in2355_1, in2355_2;
    wire c2355;
    assign in2355_1 = {s2303[0]};
    assign in2355_2 = {s2304[0]};
    Half_Adder KS_2355(s2355, c2355, in2355_1, in2355_2);
    wire[2:0] s2356, in2356_1, in2356_2;
    wire c2356;
    assign in2356_1 = {s2305[0],s2311[1],s2297[2]};
    assign in2356_2 = {s2306[0],s2312[1],s2298[2]};
    CLA_3 KS_2356(s2356, c2356, in2356_1, in2356_2);
    wire[0:0] s2357, in2357_1, in2357_2;
    wire c2357;
    assign in2357_1 = {s2307[0]};
    assign in2357_2 = {s2308[0]};
    Half_Adder KS_2357(s2357, c2357, in2357_1, in2357_2);
    wire[1:0] s2358, in2358_1, in2358_2;
    wire c2358;
    assign in2358_1 = {s2309[0],s2313[1]};
    assign in2358_2 = {s2310[0],s2314[1]};
    CLA_2 KS_2358(s2358, c2358, in2358_1, in2358_2);
    wire[0:0] s2359, in2359_1, in2359_2;
    wire c2359;
    assign in2359_1 = {s2311[0]};
    assign in2359_2 = {s2312[0]};
    Half_Adder KS_2359(s2359, c2359, in2359_1, in2359_2);
    wire[3:0] s2360, in2360_1, in2360_2;
    wire c2360;
    assign in2360_1 = {s2314[0],s2315[1],s2299[2],s730[0]};
    assign in2360_2 = {s2315[0],s2316[1],s2300[2],s731[0]};
    CLA_4_c KS_2360(s2360, c2360, in2360_1, in2360_2, s2313[0]);
    wire[3:0] s2361, in2361_1, in2361_2;
    wire c2361;
    assign in2361_1 = {s661[1],s632[2],pp113[21],s756[0]};
    assign in2361_2 = {s662[1],s633[2],pp114[20],s757[0]};
    CLA_4 KS_2361(s2361, c2361, in2361_1, in2361_2);
    wire[3:0] s2362, in2362_1, in2362_2;
    wire c2362;
    assign in2362_1 = {s663[1],s634[2],pp115[19],s758[0]};
    assign in2362_2 = {s664[1],s635[2],pp116[18],s759[0]};
    CLA_4 KS_2362(s2362, c2362, in2362_1, in2362_2);
    wire[3:0] s2363, in2363_1, in2363_2;
    wire c2363;
    assign in2363_1 = {s665[1],s636[2],pp117[17],s760[0]};
    assign in2363_2 = {s666[1],s637[2],pp118[16],s761[0]};
    CLA_4 KS_2363(s2363, c2363, in2363_1, in2363_2);
    wire[3:0] s2364, in2364_1, in2364_2;
    wire c2364;
    assign in2364_1 = {s667[1],s638[2],pp119[15],s762[0]};
    assign in2364_2 = {s668[1],s639[2],pp120[14],s763[0]};
    CLA_4 KS_2364(s2364, c2364, in2364_1, in2364_2);
    wire[3:0] s2365, in2365_1, in2365_2;
    wire c2365;
    assign in2365_1 = {s669[1],s640[2],pp121[13],s764[0]};
    assign in2365_2 = {s670[1],s641[2],pp122[12],s765[0]};
    CLA_4 KS_2365(s2365, c2365, in2365_1, in2365_2);
    wire[3:0] s2366, in2366_1, in2366_2;
    wire c2366;
    assign in2366_1 = {s671[1],s642[2],pp123[11],s766[0]};
    assign in2366_2 = {s672[1],s643[2],pp124[10],s767[0]};
    CLA_4 KS_2366(s2366, c2366, in2366_1, in2366_2);
    wire[3:0] s2367, in2367_1, in2367_2;
    wire c2367;
    assign in2367_1 = {s673[1],s644[2],pp125[9],s768[0]};
    assign in2367_2 = {s674[1],s645[2],pp126[8],s769[0]};
    CLA_4 KS_2367(s2367, c2367, in2367_1, in2367_2);
    wire[3:0] s2368, in2368_1, in2368_2;
    wire c2368;
    assign in2368_1 = {s675[1],s646[2],pp127[7],s770[0]};
    assign in2368_2 = {s676[1],s647[2],s632[3],s771[0]};
    CLA_4 KS_2368(s2368, c2368, in2368_1, in2368_2);
    wire[3:0] s2369, in2369_1, in2369_2;
    wire c2369;
    assign in2369_1 = {s677[1],s648[2],s633[3],s772[0]};
    assign in2369_2 = {s678[1],s649[2],s634[3],s773[0]};
    CLA_4 KS_2369(s2369, c2369, in2369_1, in2369_2);
    wire[3:0] s2370, in2370_1, in2370_2;
    wire c2370;
    assign in2370_1 = {s679[1],s650[2],s635[3],s774[0]};
    assign in2370_2 = {c680,s651[2],s636[3],s775[0]};
    CLA_4 KS_2370(s2370, c2370, in2370_1, in2370_2);
    wire[3:0] s2371, in2371_1, in2371_2;
    wire c2371;
    assign in2371_1 = {s681[1],s652[2],s637[3],s776[0]};
    assign in2371_2 = {c682,s653[2],s638[3],s777[0]};
    CLA_4 KS_2371(s2371, c2371, in2371_1, in2371_2);
    wire[3:0] s2372, in2372_1, in2372_2;
    wire c2372;
    assign in2372_1 = {s683[1],s654[2],s639[3],s778[0]};
    assign in2372_2 = {c684,s655[2],s640[3],s779[0]};
    CLA_4 KS_2372(s2372, c2372, in2372_1, in2372_2);
    wire[3:0] s2373, in2373_1, in2373_2;
    wire c2373;
    assign in2373_1 = {s685[1],s656[2],s641[3],s780[0]};
    assign in2373_2 = {c686,s657[2],s642[3],s781[0]};
    CLA_4 KS_2373(s2373, c2373, in2373_1, in2373_2);
    wire[3:0] s2374, in2374_1, in2374_2;
    wire c2374;
    assign in2374_1 = {s687[1],s658[2],s643[3],s782[0]};
    assign in2374_2 = {c688,s659[2],s644[3],s783[0]};
    CLA_4 KS_2374(s2374, c2374, in2374_1, in2374_2);
    wire[3:0] s2375, in2375_1, in2375_2;
    wire c2375;
    assign in2375_1 = {s689[1],s660[2],s645[3],s784[0]};
    assign in2375_2 = {c690,s661[2],s646[3],s785[0]};
    CLA_4 KS_2375(s2375, c2375, in2375_1, in2375_2);
    wire[3:0] s2376, in2376_1, in2376_2;
    wire c2376;
    assign in2376_1 = {s691[1],s662[2],s647[3],s786[0]};
    assign in2376_2 = {c692,s663[2],s648[3],s787[0]};
    CLA_4 KS_2376(s2376, c2376, in2376_1, in2376_2);
    wire[3:0] s2377, in2377_1, in2377_2;
    wire c2377;
    assign in2377_1 = {s693[1],s664[2],s649[3],s788[0]};
    assign in2377_2 = {c694,s665[2],s650[3],s789[0]};
    CLA_4 KS_2377(s2377, c2377, in2377_1, in2377_2);
    wire[3:0] s2378, in2378_1, in2378_2;
    wire c2378;
    assign in2378_1 = {s695[1],s666[2],s651[3],s790[0]};
    assign in2378_2 = {c696,s667[2],s652[3],s791[0]};
    CLA_4 KS_2378(s2378, c2378, in2378_1, in2378_2);
    wire[3:0] s2379, in2379_1, in2379_2;
    wire c2379;
    assign in2379_1 = {s697[1],s668[2],s653[3],s792[0]};
    assign in2379_2 = {c698,s669[2],s654[3],s793[0]};
    CLA_4 KS_2379(s2379, c2379, in2379_1, in2379_2);
    wire[3:0] s2380, in2380_1, in2380_2;
    wire c2380;
    assign in2380_1 = {s699[1],s670[2],s655[3],s794[0]};
    assign in2380_2 = {c700,s671[2],s656[3],s795[0]};
    CLA_4 KS_2380(s2380, c2380, in2380_1, in2380_2);
    wire[3:0] s2381, in2381_1, in2381_2;
    wire c2381;
    assign in2381_1 = {s701[1],s672[2],s657[3],s796[0]};
    assign in2381_2 = {c702,s673[2],s658[3],s797[0]};
    CLA_4 KS_2381(s2381, c2381, in2381_1, in2381_2);
    wire[3:0] s2382, in2382_1, in2382_2;
    wire c2382;
    assign in2382_1 = {s703[1],s674[2],s659[3],s798[0]};
    assign in2382_2 = {c704,s675[2],s660[3],s799[0]};
    CLA_4 KS_2382(s2382, c2382, in2382_1, in2382_2);
    wire[3:0] s2383, in2383_1, in2383_2;
    wire c2383;
    assign in2383_1 = {s705[1],s676[2],s661[3],s800[0]};
    assign in2383_2 = {c706,s677[2],s662[3],s801[0]};
    CLA_4 KS_2383(s2383, c2383, in2383_1, in2383_2);
    wire[3:0] s2384, in2384_1, in2384_2;
    wire c2384;
    assign in2384_1 = {s707[1],s678[2],s663[3],s802[0]};
    assign in2384_2 = {c708,c679,s664[3],s803[0]};
    CLA_4 KS_2384(s2384, c2384, in2384_1, in2384_2);
    wire[3:0] s2385, in2385_1, in2385_2;
    wire c2385;
    assign in2385_1 = {s709[1],s681[2],s665[3],s804[0]};
    assign in2385_2 = {c710,c683,s666[3],s805[0]};
    CLA_4 KS_2385(s2385, c2385, in2385_1, in2385_2);
    wire[3:0] s2386, in2386_1, in2386_2;
    wire c2386;
    assign in2386_1 = {s711[1],s685[2],s667[3],s806[0]};
    assign in2386_2 = {c712,c687,s668[3],s807[0]};
    CLA_4 KS_2386(s2386, c2386, in2386_1, in2386_2);
    wire[3:0] s2387, in2387_1, in2387_2;
    wire c2387;
    assign in2387_1 = {s713[1],s689[2],s669[3],s808[0]};
    assign in2387_2 = {c714,c691,s670[3],s809[0]};
    CLA_4 KS_2387(s2387, c2387, in2387_1, in2387_2);
    wire[3:0] s2388, in2388_1, in2388_2;
    wire c2388;
    assign in2388_1 = {s715[1],s693[2],s671[3],s810[0]};
    assign in2388_2 = {c716,c695,s672[3],s811[0]};
    CLA_4 KS_2388(s2388, c2388, in2388_1, in2388_2);
    wire[3:0] s2389, in2389_1, in2389_2;
    wire c2389;
    assign in2389_1 = {s717[1],s697[2],s673[3],s812[0]};
    assign in2389_2 = {c718,c699,s674[3],s813[0]};
    CLA_4 KS_2389(s2389, c2389, in2389_1, in2389_2);
    wire[3:0] s2390, in2390_1, in2390_2;
    wire c2390;
    assign in2390_1 = {s719[1],s701[2],s675[3],s814[0]};
    assign in2390_2 = {c720,c703,s676[3],s815[0]};
    CLA_4 KS_2390(s2390, c2390, in2390_1, in2390_2);
    wire[3:0] s2391, in2391_1, in2391_2;
    wire c2391;
    assign in2391_1 = {s721[1],s705[2],s677[3],s816[0]};
    assign in2391_2 = {c722,c707,c678,s817[0]};
    CLA_4 KS_2391(s2391, c2391, in2391_1, in2391_2);
    wire[3:0] s2392, in2392_1, in2392_2;
    wire c2392;
    assign in2392_1 = {s723[1],s709[2],s681[3],s818[0]};
    assign in2392_2 = {c724,c711,c685,s819[0]};
    CLA_4 KS_2392(s2392, c2392, in2392_1, in2392_2);
    wire[0:0] s2393, in2393_1, in2393_2;
    wire c2393;
    assign in2393_1 = {s725[1]};
    assign in2393_2 = {c726};
    Half_Adder KS_2393(s2393, c2393, in2393_1, in2393_2);
    wire[1:0] s2394, in2394_1, in2394_2;
    wire c2394;
    assign in2394_1 = {s727[1],s713[2]};
    assign in2394_2 = {c728,c715};
    CLA_2 KS_2394(s2394, c2394, in2394_1, in2394_2);
    wire[0:0] s2395, in2395_1, in2395_2;
    wire c2395;
    assign in2395_1 = {s729[1]};
    assign in2395_2 = {c730};
    Half_Adder KS_2395(s2395, c2395, in2395_1, in2395_2);
    wire[2:0] s2396, in2396_1, in2396_2;
    wire c2396;
    assign in2396_1 = {s731[1],s717[2],s689[3]};
    assign in2396_2 = {c732,c719,c693};
    CLA_3 KS_2396(s2396, c2396, in2396_1, in2396_2);
    wire[0:0] s2397, in2397_1, in2397_2;
    wire c2397;
    assign in2397_1 = {s733[1]};
    assign in2397_2 = {c734};
    Half_Adder KS_2397(s2397, c2397, in2397_1, in2397_2);
    wire[1:0] s2398, in2398_1, in2398_2;
    wire c2398;
    assign in2398_1 = {s735[1],s721[2]};
    assign in2398_2 = {c2297,c723};
    CLA_2 KS_2398(s2398, c2398, in2398_1, in2398_2);
    wire[0:0] s2399, in2399_1, in2399_2;
    wire c2399;
    assign in2399_1 = {c2298};
    assign in2399_2 = {c2299};
    Half_Adder KS_2399(s2399, c2399, in2399_1, in2399_2);
    wire[3:0] s2400, in2400_1, in2400_2;
    wire c2400;
    assign in2400_1 = {c2300,s725[2],s697[3],s820[0]};
    assign in2400_2 = {c2301,c727,c701,s821[0]};
    CLA_4 KS_2400(s2400, c2400, in2400_1, in2400_2);
    wire[0:0] s2401, in2401_1, in2401_2;
    wire c2401;
    assign in2401_1 = {c2302};
    assign in2401_2 = {c2303};
    Half_Adder KS_2401(s2401, c2401, in2401_1, in2401_2);
    wire[1:0] s2402, in2402_1, in2402_2;
    wire c2402;
    assign in2402_1 = {c2304,s729[2]};
    assign in2402_2 = {c2305,c731};
    CLA_2 KS_2402(s2402, c2402, in2402_1, in2402_2);
    wire[0:0] s2403, in2403_1, in2403_2;
    wire c2403;
    assign in2403_1 = {c2306};
    assign in2403_2 = {c2307};
    Half_Adder KS_2403(s2403, c2403, in2403_1, in2403_2);
    wire[2:0] s2404, in2404_1, in2404_2;
    wire c2404;
    assign in2404_1 = {c2308,s733[2],s705[3]};
    assign in2404_2 = {c2309,c735,c709};
    CLA_3 KS_2404(s2404, c2404, in2404_1, in2404_2);
    wire[0:0] s2405, in2405_1, in2405_2;
    wire c2405;
    assign in2405_1 = {c2310};
    assign in2405_2 = {c2311};
    Half_Adder KS_2405(s2405, c2405, in2405_1, in2405_2);
    wire[1:0] s2406, in2406_1, in2406_2;
    wire c2406;
    assign in2406_1 = {c2312,s2361[1]};
    assign in2406_2 = {c2313,s2362[1]};
    CLA_2 KS_2406(s2406, c2406, in2406_1, in2406_2);
    wire[0:0] s2407, in2407_1, in2407_2;
    wire c2407;
    assign in2407_1 = {c2314};
    assign in2407_2 = {c2315};
    Half_Adder KS_2407(s2407, c2407, in2407_1, in2407_2);
    wire[3:0] s2408, in2408_1, in2408_2;
    wire c2408;
    assign in2408_1 = {c2316,s2363[1],s713[3],s822[0]};
    assign in2408_2 = {c2317,s2364[1],c717,s823[0]};
    CLA_4 KS_2408(s2408, c2408, in2408_1, in2408_2);
    wire[0:0] s2409, in2409_1, in2409_2;
    wire c2409;
    assign in2409_1 = {c2318};
    assign in2409_2 = {c2319};
    Half_Adder KS_2409(s2409, c2409, in2409_1, in2409_2);
    wire[1:0] s2410, in2410_1, in2410_2;
    wire c2410;
    assign in2410_1 = {c2320,s2365[1]};
    assign in2410_2 = {c2321,s2366[1]};
    CLA_2 KS_2410(s2410, c2410, in2410_1, in2410_2);
    wire[0:0] s2411, in2411_1, in2411_2;
    wire c2411;
    assign in2411_1 = {c2322};
    assign in2411_2 = {c2323};
    Half_Adder KS_2411(s2411, c2411, in2411_1, in2411_2);
    wire[2:0] s2412, in2412_1, in2412_2;
    wire c2412;
    assign in2412_1 = {c2324,s2367[1],s721[3]};
    assign in2412_2 = {c2325,s2368[1],c725};
    CLA_3 KS_2412(s2412, c2412, in2412_1, in2412_2);
    wire[0:0] s2413, in2413_1, in2413_2;
    wire c2413;
    assign in2413_1 = {c2326};
    assign in2413_2 = {c2327};
    Half_Adder KS_2413(s2413, c2413, in2413_1, in2413_2);
    wire[1:0] s2414, in2414_1, in2414_2;
    wire c2414;
    assign in2414_1 = {c2328,s2369[1]};
    assign in2414_2 = {c2336,s2370[1]};
    CLA_2 KS_2414(s2414, c2414, in2414_1, in2414_2);
    wire[0:0] s2415, in2415_1, in2415_2;
    wire c2415;
    assign in2415_1 = {c2344};
    assign in2415_2 = {c2352};
    Half_Adder KS_2415(s2415, c2415, in2415_1, in2415_2);
    wire[3:0] s2416, in2416_1, in2416_2;
    wire c2416;
    assign in2416_1 = {c2360,s2371[1],s729[3],s824[0]};
    assign in2416_2 = {s2361[0],s2372[1],c733,s825[0]};
    CLA_4 KS_2416(s2416, c2416, in2416_1, in2416_2);
    wire[0:0] s2417, in2417_1, in2417_2;
    wire c2417;
    assign in2417_1 = {s2362[0]};
    assign in2417_2 = {s2363[0]};
    Half_Adder KS_2417(s2417, c2417, in2417_1, in2417_2);
    wire[1:0] s2418, in2418_1, in2418_2;
    wire c2418;
    assign in2418_1 = {s2364[0],s2373[1]};
    assign in2418_2 = {s2365[0],s2374[1]};
    CLA_2 KS_2418(s2418, c2418, in2418_1, in2418_2);
    wire[0:0] s2419, in2419_1, in2419_2;
    wire c2419;
    assign in2419_1 = {s2366[0]};
    assign in2419_2 = {s2367[0]};
    Half_Adder KS_2419(s2419, c2419, in2419_1, in2419_2);
    wire[2:0] s2420, in2420_1, in2420_2;
    wire c2420;
    assign in2420_1 = {s2368[0],s2375[1],s2361[2]};
    assign in2420_2 = {s2369[0],s2376[1],s2362[2]};
    CLA_3 KS_2420(s2420, c2420, in2420_1, in2420_2);
    wire[0:0] s2421, in2421_1, in2421_2;
    wire c2421;
    assign in2421_1 = {s2370[0]};
    assign in2421_2 = {s2371[0]};
    Half_Adder KS_2421(s2421, c2421, in2421_1, in2421_2);
    wire[1:0] s2422, in2422_1, in2422_2;
    wire c2422;
    assign in2422_1 = {s2372[0],s2377[1]};
    assign in2422_2 = {s2373[0],s2378[1]};
    CLA_2 KS_2422(s2422, c2422, in2422_1, in2422_2);
    wire[0:0] s2423, in2423_1, in2423_2;
    wire c2423;
    assign in2423_1 = {s2374[0]};
    assign in2423_2 = {s2375[0]};
    Half_Adder KS_2423(s2423, c2423, in2423_1, in2423_2);
    wire[3:0] s2424, in2424_1, in2424_2;
    wire c2424;
    assign in2424_1 = {s2376[0],s2379[1],s2363[2],s826[0]};
    assign in2424_2 = {s2377[0],s2380[1],s2364[2],s827[0]};
    CLA_4 KS_2424(s2424, c2424, in2424_1, in2424_2);
    wire[0:0] s2425, in2425_1, in2425_2;
    wire c2425;
    assign in2425_1 = {s2379[0]};
    assign in2425_2 = {s2380[0]};
    Full_Adder KS_2425(s2425, c2425, in2425_1, in2425_2, s2378[0]);
    wire[3:0] s2426, in2426_1, in2426_2;
    wire c2426;
    assign in2426_1 = {s757[1],pp122[15],pp109[29],s844[0]};
    assign in2426_2 = {s758[1],pp123[14],pp110[28],s845[0]};
    CLA_4 KS_2426(s2426, c2426, in2426_1, in2426_2);
    wire[3:0] s2427, in2427_1, in2427_2;
    wire c2427;
    assign in2427_1 = {s759[1],pp124[13],pp111[27],s846[0]};
    assign in2427_2 = {s760[1],pp125[12],pp112[26],s847[0]};
    CLA_4 KS_2427(s2427, c2427, in2427_1, in2427_2);
    wire[3:0] s2428, in2428_1, in2428_2;
    wire c2428;
    assign in2428_1 = {s761[1],pp126[11],pp113[25],s848[0]};
    assign in2428_2 = {s762[1],pp127[10],pp114[24],s849[0]};
    CLA_4 KS_2428(s2428, c2428, in2428_1, in2428_2);
    wire[3:0] s2429, in2429_1, in2429_2;
    wire c2429;
    assign in2429_1 = {s763[1],s736[2],pp115[23],s850[0]};
    assign in2429_2 = {s764[1],s737[2],pp116[22],s851[0]};
    CLA_4 KS_2429(s2429, c2429, in2429_1, in2429_2);
    wire[3:0] s2430, in2430_1, in2430_2;
    wire c2430;
    assign in2430_1 = {s765[1],s738[2],pp117[21],s852[0]};
    assign in2430_2 = {s766[1],s739[2],pp118[20],s853[0]};
    CLA_4 KS_2430(s2430, c2430, in2430_1, in2430_2);
    wire[3:0] s2431, in2431_1, in2431_2;
    wire c2431;
    assign in2431_1 = {s767[1],s740[2],pp119[19],s854[0]};
    assign in2431_2 = {s768[1],s741[2],pp120[18],s855[0]};
    CLA_4 KS_2431(s2431, c2431, in2431_1, in2431_2);
    wire[3:0] s2432, in2432_1, in2432_2;
    wire c2432;
    assign in2432_1 = {s769[1],s742[2],pp121[17],s856[0]};
    assign in2432_2 = {s770[1],s743[2],pp122[16],s857[0]};
    CLA_4 KS_2432(s2432, c2432, in2432_1, in2432_2);
    wire[3:0] s2433, in2433_1, in2433_2;
    wire c2433;
    assign in2433_1 = {s771[1],s744[2],pp123[15],s858[0]};
    assign in2433_2 = {s772[1],s745[2],pp124[14],s859[0]};
    CLA_4 KS_2433(s2433, c2433, in2433_1, in2433_2);
    wire[3:0] s2434, in2434_1, in2434_2;
    wire c2434;
    assign in2434_1 = {s773[1],s746[2],pp125[13],s860[0]};
    assign in2434_2 = {s774[1],s747[2],pp126[12],s861[0]};
    CLA_4 KS_2434(s2434, c2434, in2434_1, in2434_2);
    wire[3:0] s2435, in2435_1, in2435_2;
    wire c2435;
    assign in2435_1 = {s775[1],s748[2],pp127[11],s862[0]};
    assign in2435_2 = {s776[1],s749[2],s736[3],s863[0]};
    CLA_4 KS_2435(s2435, c2435, in2435_1, in2435_2);
    wire[3:0] s2436, in2436_1, in2436_2;
    wire c2436;
    assign in2436_1 = {s777[1],s750[2],s737[3],s864[0]};
    assign in2436_2 = {s778[1],s751[2],s738[3],s865[0]};
    CLA_4 KS_2436(s2436, c2436, in2436_1, in2436_2);
    wire[3:0] s2437, in2437_1, in2437_2;
    wire c2437;
    assign in2437_1 = {s779[1],s752[2],s739[3],s866[0]};
    assign in2437_2 = {c780,s753[2],s740[3],s867[0]};
    CLA_4 KS_2437(s2437, c2437, in2437_1, in2437_2);
    wire[3:0] s2438, in2438_1, in2438_2;
    wire c2438;
    assign in2438_1 = {s781[1],s754[2],s741[3],s868[0]};
    assign in2438_2 = {c782,s755[2],s742[3],s869[0]};
    CLA_4 KS_2438(s2438, c2438, in2438_1, in2438_2);
    wire[3:0] s2439, in2439_1, in2439_2;
    wire c2439;
    assign in2439_1 = {s783[1],s756[2],s743[3],s870[0]};
    assign in2439_2 = {c784,s757[2],s744[3],s871[0]};
    CLA_4 KS_2439(s2439, c2439, in2439_1, in2439_2);
    wire[3:0] s2440, in2440_1, in2440_2;
    wire c2440;
    assign in2440_1 = {s785[1],s758[2],s745[3],s872[0]};
    assign in2440_2 = {c786,s759[2],s746[3],s873[0]};
    CLA_4 KS_2440(s2440, c2440, in2440_1, in2440_2);
    wire[3:0] s2441, in2441_1, in2441_2;
    wire c2441;
    assign in2441_1 = {s787[1],s760[2],s747[3],s874[0]};
    assign in2441_2 = {c788,s761[2],s748[3],s875[0]};
    CLA_4 KS_2441(s2441, c2441, in2441_1, in2441_2);
    wire[3:0] s2442, in2442_1, in2442_2;
    wire c2442;
    assign in2442_1 = {s789[1],s762[2],s749[3],s876[0]};
    assign in2442_2 = {c790,s763[2],s750[3],s877[0]};
    CLA_4 KS_2442(s2442, c2442, in2442_1, in2442_2);
    wire[3:0] s2443, in2443_1, in2443_2;
    wire c2443;
    assign in2443_1 = {s791[1],s764[2],s751[3],s878[0]};
    assign in2443_2 = {c792,s765[2],s752[3],s879[0]};
    CLA_4 KS_2443(s2443, c2443, in2443_1, in2443_2);
    wire[3:0] s2444, in2444_1, in2444_2;
    wire c2444;
    assign in2444_1 = {s793[1],s766[2],s753[3],s880[0]};
    assign in2444_2 = {c794,s767[2],s754[3],s881[0]};
    CLA_4 KS_2444(s2444, c2444, in2444_1, in2444_2);
    wire[3:0] s2445, in2445_1, in2445_2;
    wire c2445;
    assign in2445_1 = {s795[1],s768[2],s755[3],s882[0]};
    assign in2445_2 = {c796,s769[2],s756[3],s883[0]};
    CLA_4 KS_2445(s2445, c2445, in2445_1, in2445_2);
    wire[3:0] s2446, in2446_1, in2446_2;
    wire c2446;
    assign in2446_1 = {s797[1],s770[2],s757[3],s884[0]};
    assign in2446_2 = {c798,s771[2],s758[3],s885[0]};
    CLA_4 KS_2446(s2446, c2446, in2446_1, in2446_2);
    wire[3:0] s2447, in2447_1, in2447_2;
    wire c2447;
    assign in2447_1 = {s799[1],s772[2],s759[3],s886[0]};
    assign in2447_2 = {c800,s773[2],s760[3],s887[0]};
    CLA_4 KS_2447(s2447, c2447, in2447_1, in2447_2);
    wire[3:0] s2448, in2448_1, in2448_2;
    wire c2448;
    assign in2448_1 = {s801[1],s774[2],s761[3],s888[0]};
    assign in2448_2 = {c802,s775[2],s762[3],s889[0]};
    CLA_4 KS_2448(s2448, c2448, in2448_1, in2448_2);
    wire[3:0] s2449, in2449_1, in2449_2;
    wire c2449;
    assign in2449_1 = {s803[1],s776[2],s763[3],s890[0]};
    assign in2449_2 = {c804,s777[2],s764[3],s891[0]};
    CLA_4 KS_2449(s2449, c2449, in2449_1, in2449_2);
    wire[3:0] s2450, in2450_1, in2450_2;
    wire c2450;
    assign in2450_1 = {s805[1],s778[2],s765[3],s892[0]};
    assign in2450_2 = {c806,c779,s766[3],s893[0]};
    CLA_4 KS_2450(s2450, c2450, in2450_1, in2450_2);
    wire[3:0] s2451, in2451_1, in2451_2;
    wire c2451;
    assign in2451_1 = {s807[1],s781[2],s767[3],s894[0]};
    assign in2451_2 = {c808,c783,s768[3],s895[0]};
    CLA_4 KS_2451(s2451, c2451, in2451_1, in2451_2);
    wire[3:0] s2452, in2452_1, in2452_2;
    wire c2452;
    assign in2452_1 = {s809[1],s785[2],s769[3],s896[0]};
    assign in2452_2 = {c810,c787,s770[3],s897[0]};
    CLA_4 KS_2452(s2452, c2452, in2452_1, in2452_2);
    wire[3:0] s2453, in2453_1, in2453_2;
    wire c2453;
    assign in2453_1 = {s811[1],s789[2],s771[3],s898[0]};
    assign in2453_2 = {c812,c791,s772[3],s899[0]};
    CLA_4 KS_2453(s2453, c2453, in2453_1, in2453_2);
    wire[3:0] s2454, in2454_1, in2454_2;
    wire c2454;
    assign in2454_1 = {s813[1],s793[2],s773[3],s900[0]};
    assign in2454_2 = {c814,c795,s774[3],s901[0]};
    CLA_4 KS_2454(s2454, c2454, in2454_1, in2454_2);
    wire[3:0] s2455, in2455_1, in2455_2;
    wire c2455;
    assign in2455_1 = {s815[1],s797[2],s775[3],s902[0]};
    assign in2455_2 = {c816,c799,s776[3],s903[0]};
    CLA_4 KS_2455(s2455, c2455, in2455_1, in2455_2);
    wire[3:0] s2456, in2456_1, in2456_2;
    wire c2456;
    assign in2456_1 = {s817[1],s801[2],s777[3],s904[0]};
    assign in2456_2 = {c818,c803,c778,s905[0]};
    CLA_4 KS_2456(s2456, c2456, in2456_1, in2456_2);
    wire[1:0] s2457, in2457_1, in2457_2;
    wire c2457;
    assign in2457_1 = {s819[1],s805[2]};
    assign in2457_2 = {c820,c807};
    CLA_2 KS_2457(s2457, c2457, in2457_1, in2457_2);
    wire[0:0] s2458, in2458_1, in2458_2;
    wire c2458;
    assign in2458_1 = {s821[1]};
    assign in2458_2 = {c822};
    Half_Adder KS_2458(s2458, c2458, in2458_1, in2458_2);
    wire[3:0] s2459, in2459_1, in2459_2;
    wire c2459;
    assign in2459_1 = {s823[1],s809[2],s781[3],s906[0]};
    assign in2459_2 = {c824,c811,c785,s907[0]};
    CLA_4 KS_2459(s2459, c2459, in2459_1, in2459_2);
    wire[0:0] s2460, in2460_1, in2460_2;
    wire c2460;
    assign in2460_1 = {s825[1]};
    assign in2460_2 = {c826};
    Half_Adder KS_2460(s2460, c2460, in2460_1, in2460_2);
    wire[1:0] s2461, in2461_1, in2461_2;
    wire c2461;
    assign in2461_1 = {s827[1],s813[2]};
    assign in2461_2 = {c828,c815};
    CLA_2 KS_2461(s2461, c2461, in2461_1, in2461_2);
    wire[0:0] s2462, in2462_1, in2462_2;
    wire c2462;
    assign in2462_1 = {s829[1]};
    assign in2462_2 = {c830};
    Half_Adder KS_2462(s2462, c2462, in2462_1, in2462_2);
    wire[2:0] s2463, in2463_1, in2463_2;
    wire c2463;
    assign in2463_1 = {s831[1],s817[2],s789[3]};
    assign in2463_2 = {c2361,c819,c793};
    CLA_3 KS_2463(s2463, c2463, in2463_1, in2463_2);
    wire[0:0] s2464, in2464_1, in2464_2;
    wire c2464;
    assign in2464_1 = {c2362};
    assign in2464_2 = {c2363};
    Half_Adder KS_2464(s2464, c2464, in2464_1, in2464_2);
    wire[1:0] s2465, in2465_1, in2465_2;
    wire c2465;
    assign in2465_1 = {c2364,s821[2]};
    assign in2465_2 = {c2365,c823};
    CLA_2 KS_2465(s2465, c2465, in2465_1, in2465_2);
    wire[0:0] s2466, in2466_1, in2466_2;
    wire c2466;
    assign in2466_1 = {c2366};
    assign in2466_2 = {c2367};
    Half_Adder KS_2466(s2466, c2466, in2466_1, in2466_2);
    wire[3:0] s2467, in2467_1, in2467_2;
    wire c2467;
    assign in2467_1 = {c2368,s825[2],s797[3],s908[0]};
    assign in2467_2 = {c2369,c827,c801,s909[0]};
    CLA_4 KS_2467(s2467, c2467, in2467_1, in2467_2);
    wire[0:0] s2468, in2468_1, in2468_2;
    wire c2468;
    assign in2468_1 = {c2370};
    assign in2468_2 = {c2371};
    Half_Adder KS_2468(s2468, c2468, in2468_1, in2468_2);
    wire[1:0] s2469, in2469_1, in2469_2;
    wire c2469;
    assign in2469_1 = {c2372,s829[2]};
    assign in2469_2 = {c2373,c831};
    CLA_2 KS_2469(s2469, c2469, in2469_1, in2469_2);
    wire[0:0] s2470, in2470_1, in2470_2;
    wire c2470;
    assign in2470_1 = {c2374};
    assign in2470_2 = {c2375};
    Half_Adder KS_2470(s2470, c2470, in2470_1, in2470_2);
    wire[2:0] s2471, in2471_1, in2471_2;
    wire c2471;
    assign in2471_1 = {c2376,s2426[1],s805[3]};
    assign in2471_2 = {c2377,s2427[1],c809};
    CLA_3 KS_2471(s2471, c2471, in2471_1, in2471_2);
    wire[0:0] s2472, in2472_1, in2472_2;
    wire c2472;
    assign in2472_1 = {c2378};
    assign in2472_2 = {c2379};
    Half_Adder KS_2472(s2472, c2472, in2472_1, in2472_2);
    wire[1:0] s2473, in2473_1, in2473_2;
    wire c2473;
    assign in2473_1 = {c2380,s2428[1]};
    assign in2473_2 = {c2381,s2429[1]};
    CLA_2 KS_2473(s2473, c2473, in2473_1, in2473_2);
    wire[0:0] s2474, in2474_1, in2474_2;
    wire c2474;
    assign in2474_1 = {c2382};
    assign in2474_2 = {c2383};
    Half_Adder KS_2474(s2474, c2474, in2474_1, in2474_2);
    wire[3:0] s2475, in2475_1, in2475_2;
    wire c2475;
    assign in2475_1 = {c2384,s2430[1],s813[3],s910[0]};
    assign in2475_2 = {c2385,s2431[1],c817,s911[0]};
    CLA_4 KS_2475(s2475, c2475, in2475_1, in2475_2);
    wire[0:0] s2476, in2476_1, in2476_2;
    wire c2476;
    assign in2476_1 = {c2386};
    assign in2476_2 = {c2387};
    Half_Adder KS_2476(s2476, c2476, in2476_1, in2476_2);
    wire[1:0] s2477, in2477_1, in2477_2;
    wire c2477;
    assign in2477_1 = {c2388,s2432[1]};
    assign in2477_2 = {c2389,s2433[1]};
    CLA_2 KS_2477(s2477, c2477, in2477_1, in2477_2);
    wire[0:0] s2478, in2478_1, in2478_2;
    wire c2478;
    assign in2478_1 = {c2390};
    assign in2478_2 = {c2391};
    Half_Adder KS_2478(s2478, c2478, in2478_1, in2478_2);
    wire[2:0] s2479, in2479_1, in2479_2;
    wire c2479;
    assign in2479_1 = {c2392,s2434[1],s821[3]};
    assign in2479_2 = {c2400,s2435[1],c825};
    CLA_3 KS_2479(s2479, c2479, in2479_1, in2479_2);
    wire[0:0] s2480, in2480_1, in2480_2;
    wire c2480;
    assign in2480_1 = {c2408};
    assign in2480_2 = {c2416};
    Half_Adder KS_2480(s2480, c2480, in2480_1, in2480_2);
    wire[1:0] s2481, in2481_1, in2481_2;
    wire c2481;
    assign in2481_1 = {c2424,s2436[1]};
    assign in2481_2 = {s2426[0],s2437[1]};
    CLA_2 KS_2481(s2481, c2481, in2481_1, in2481_2);
    wire[0:0] s2482, in2482_1, in2482_2;
    wire c2482;
    assign in2482_1 = {s2427[0]};
    assign in2482_2 = {s2428[0]};
    Half_Adder KS_2482(s2482, c2482, in2482_1, in2482_2);
    wire[3:0] s2483, in2483_1, in2483_2;
    wire c2483;
    assign in2483_1 = {s2429[0],s2438[1],s829[3],s912[0]};
    assign in2483_2 = {s2430[0],s2439[1],s2426[2],s913[0]};
    CLA_4 KS_2483(s2483, c2483, in2483_1, in2483_2);
    wire[0:0] s2484, in2484_1, in2484_2;
    wire c2484;
    assign in2484_1 = {s2431[0]};
    assign in2484_2 = {s2432[0]};
    Half_Adder KS_2484(s2484, c2484, in2484_1, in2484_2);
    wire[1:0] s2485, in2485_1, in2485_2;
    wire c2485;
    assign in2485_1 = {s2433[0],s2440[1]};
    assign in2485_2 = {s2434[0],s2441[1]};
    CLA_2 KS_2485(s2485, c2485, in2485_1, in2485_2);
    wire[0:0] s2486, in2486_1, in2486_2;
    wire c2486;
    assign in2486_1 = {s2435[0]};
    assign in2486_2 = {s2436[0]};
    Half_Adder KS_2486(s2486, c2486, in2486_1, in2486_2);
    wire[2:0] s2487, in2487_1, in2487_2;
    wire c2487;
    assign in2487_1 = {s2437[0],s2442[1],s2427[2]};
    assign in2487_2 = {s2438[0],s2443[1],s2428[2]};
    CLA_3 KS_2487(s2487, c2487, in2487_1, in2487_2);
    wire[0:0] s2488, in2488_1, in2488_2;
    wire c2488;
    assign in2488_1 = {s2439[0]};
    assign in2488_2 = {s2440[0]};
    Half_Adder KS_2488(s2488, c2488, in2488_1, in2488_2);
    wire[1:0] s2489, in2489_1, in2489_2;
    wire c2489;
    assign in2489_1 = {s2441[0],s2444[1]};
    assign in2489_2 = {s2442[0],s2445[1]};
    CLA_2 KS_2489(s2489, c2489, in2489_1, in2489_2);
    wire[0:0] s2490, in2490_1, in2490_2;
    wire c2490;
    assign in2490_1 = {s2444[0]};
    assign in2490_2 = {s2445[0]};
    Full_Adder KS_2490(s2490, c2490, in2490_1, in2490_2, s2443[0]);
    wire[3:0] s2491, in2491_1, in2491_2;
    wire c2491;
    assign in2491_1 = {s845[1],pp116[25],pp103[39],s923[0]};
    assign in2491_2 = {s846[1],pp117[24],pp104[38],s924[0]};
    CLA_4 KS_2491(s2491, c2491, in2491_1, in2491_2);
    wire[3:0] s2492, in2492_1, in2492_2;
    wire c2492;
    assign in2492_1 = {s847[1],pp118[23],pp105[37],s925[0]};
    assign in2492_2 = {s848[1],pp119[22],pp106[36],s926[0]};
    CLA_4 KS_2492(s2492, c2492, in2492_1, in2492_2);
    wire[3:0] s2493, in2493_1, in2493_2;
    wire c2493;
    assign in2493_1 = {s849[1],pp120[21],pp107[35],s927[0]};
    assign in2493_2 = {s850[1],pp121[20],pp108[34],s928[0]};
    CLA_4 KS_2493(s2493, c2493, in2493_1, in2493_2);
    wire[3:0] s2494, in2494_1, in2494_2;
    wire c2494;
    assign in2494_1 = {s851[1],pp122[19],pp109[33],s929[0]};
    assign in2494_2 = {s852[1],pp123[18],pp110[32],s930[0]};
    CLA_4 KS_2494(s2494, c2494, in2494_1, in2494_2);
    wire[3:0] s2495, in2495_1, in2495_2;
    wire c2495;
    assign in2495_1 = {s853[1],pp124[17],pp111[31],s931[0]};
    assign in2495_2 = {s854[1],pp125[16],pp112[30],s932[0]};
    CLA_4 KS_2495(s2495, c2495, in2495_1, in2495_2);
    wire[3:0] s2496, in2496_1, in2496_2;
    wire c2496;
    assign in2496_1 = {s855[1],pp126[15],pp113[29],s933[0]};
    assign in2496_2 = {s856[1],pp127[14],pp114[28],s934[0]};
    CLA_4 KS_2496(s2496, c2496, in2496_1, in2496_2);
    wire[3:0] s2497, in2497_1, in2497_2;
    wire c2497;
    assign in2497_1 = {s857[1],s832[2],pp115[27],s935[0]};
    assign in2497_2 = {s858[1],s833[2],pp116[26],s936[0]};
    CLA_4 KS_2497(s2497, c2497, in2497_1, in2497_2);
    wire[3:0] s2498, in2498_1, in2498_2;
    wire c2498;
    assign in2498_1 = {s859[1],s834[2],pp117[25],s937[0]};
    assign in2498_2 = {s860[1],s835[2],pp118[24],s938[0]};
    CLA_4 KS_2498(s2498, c2498, in2498_1, in2498_2);
    wire[3:0] s2499, in2499_1, in2499_2;
    wire c2499;
    assign in2499_1 = {s861[1],s836[2],pp119[23],s939[0]};
    assign in2499_2 = {s862[1],s837[2],pp120[22],s940[0]};
    CLA_4 KS_2499(s2499, c2499, in2499_1, in2499_2);
    wire[3:0] s2500, in2500_1, in2500_2;
    wire c2500;
    assign in2500_1 = {s863[1],s838[2],pp121[21],s941[0]};
    assign in2500_2 = {s864[1],s839[2],pp122[20],s942[0]};
    CLA_4 KS_2500(s2500, c2500, in2500_1, in2500_2);
    wire[3:0] s2501, in2501_1, in2501_2;
    wire c2501;
    assign in2501_1 = {s865[1],s840[2],pp123[19],s943[0]};
    assign in2501_2 = {s866[1],s841[2],pp124[18],s944[0]};
    CLA_4 KS_2501(s2501, c2501, in2501_1, in2501_2);
    wire[3:0] s2502, in2502_1, in2502_2;
    wire c2502;
    assign in2502_1 = {s867[1],s842[2],pp125[17],s945[0]};
    assign in2502_2 = {s868[1],s843[2],pp126[16],s946[0]};
    CLA_4 KS_2502(s2502, c2502, in2502_1, in2502_2);
    wire[3:0] s2503, in2503_1, in2503_2;
    wire c2503;
    assign in2503_1 = {s869[1],s844[2],pp127[15],s947[0]};
    assign in2503_2 = {s870[1],s845[2],s832[3],s948[0]};
    CLA_4 KS_2503(s2503, c2503, in2503_1, in2503_2);
    wire[3:0] s2504, in2504_1, in2504_2;
    wire c2504;
    assign in2504_1 = {s871[1],s846[2],s833[3],s949[0]};
    assign in2504_2 = {c872,s847[2],s834[3],s950[0]};
    CLA_4 KS_2504(s2504, c2504, in2504_1, in2504_2);
    wire[3:0] s2505, in2505_1, in2505_2;
    wire c2505;
    assign in2505_1 = {s873[1],s848[2],s835[3],s951[0]};
    assign in2505_2 = {c874,s849[2],s836[3],s952[0]};
    CLA_4 KS_2505(s2505, c2505, in2505_1, in2505_2);
    wire[3:0] s2506, in2506_1, in2506_2;
    wire c2506;
    assign in2506_1 = {s875[1],s850[2],s837[3],s953[0]};
    assign in2506_2 = {c876,s851[2],s838[3],s954[0]};
    CLA_4 KS_2506(s2506, c2506, in2506_1, in2506_2);
    wire[3:0] s2507, in2507_1, in2507_2;
    wire c2507;
    assign in2507_1 = {s877[1],s852[2],s839[3],s955[0]};
    assign in2507_2 = {c878,s853[2],s840[3],s956[0]};
    CLA_4 KS_2507(s2507, c2507, in2507_1, in2507_2);
    wire[3:0] s2508, in2508_1, in2508_2;
    wire c2508;
    assign in2508_1 = {s879[1],s854[2],s841[3],s957[0]};
    assign in2508_2 = {c880,s855[2],s842[3],s958[0]};
    CLA_4 KS_2508(s2508, c2508, in2508_1, in2508_2);
    wire[3:0] s2509, in2509_1, in2509_2;
    wire c2509;
    assign in2509_1 = {s881[1],s856[2],s843[3],s959[0]};
    assign in2509_2 = {c882,s857[2],s844[3],s960[0]};
    CLA_4 KS_2509(s2509, c2509, in2509_1, in2509_2);
    wire[3:0] s2510, in2510_1, in2510_2;
    wire c2510;
    assign in2510_1 = {s883[1],s858[2],s845[3],s961[0]};
    assign in2510_2 = {c884,s859[2],s846[3],s962[0]};
    CLA_4 KS_2510(s2510, c2510, in2510_1, in2510_2);
    wire[3:0] s2511, in2511_1, in2511_2;
    wire c2511;
    assign in2511_1 = {s885[1],s860[2],s847[3],s963[0]};
    assign in2511_2 = {c886,s861[2],s848[3],s964[0]};
    CLA_4 KS_2511(s2511, c2511, in2511_1, in2511_2);
    wire[3:0] s2512, in2512_1, in2512_2;
    wire c2512;
    assign in2512_1 = {s887[1],s862[2],s849[3],s965[0]};
    assign in2512_2 = {c888,s863[2],s850[3],s966[0]};
    CLA_4 KS_2512(s2512, c2512, in2512_1, in2512_2);
    wire[3:0] s2513, in2513_1, in2513_2;
    wire c2513;
    assign in2513_1 = {s889[1],s864[2],s851[3],s967[0]};
    assign in2513_2 = {c890,s865[2],s852[3],s968[0]};
    CLA_4 KS_2513(s2513, c2513, in2513_1, in2513_2);
    wire[3:0] s2514, in2514_1, in2514_2;
    wire c2514;
    assign in2514_1 = {s891[1],s866[2],s853[3],s969[0]};
    assign in2514_2 = {c892,s867[2],s854[3],s970[0]};
    CLA_4 KS_2514(s2514, c2514, in2514_1, in2514_2);
    wire[3:0] s2515, in2515_1, in2515_2;
    wire c2515;
    assign in2515_1 = {s893[1],s868[2],s855[3],s971[0]};
    assign in2515_2 = {c894,s869[2],s856[3],s972[0]};
    CLA_4 KS_2515(s2515, c2515, in2515_1, in2515_2);
    wire[3:0] s2516, in2516_1, in2516_2;
    wire c2516;
    assign in2516_1 = {s895[1],s870[2],s857[3],s973[0]};
    assign in2516_2 = {c896,c871,s858[3],s974[0]};
    CLA_4 KS_2516(s2516, c2516, in2516_1, in2516_2);
    wire[3:0] s2517, in2517_1, in2517_2;
    wire c2517;
    assign in2517_1 = {s897[1],s873[2],s859[3],s975[0]};
    assign in2517_2 = {c898,c875,s860[3],s976[0]};
    CLA_4 KS_2517(s2517, c2517, in2517_1, in2517_2);
    wire[3:0] s2518, in2518_1, in2518_2;
    wire c2518;
    assign in2518_1 = {s899[1],s877[2],s861[3],s977[0]};
    assign in2518_2 = {c900,c879,s862[3],s978[0]};
    CLA_4 KS_2518(s2518, c2518, in2518_1, in2518_2);
    wire[3:0] s2519, in2519_1, in2519_2;
    wire c2519;
    assign in2519_1 = {s901[1],s881[2],s863[3],s979[0]};
    assign in2519_2 = {c902,c883,s864[3],s980[0]};
    CLA_4 KS_2519(s2519, c2519, in2519_1, in2519_2);
    wire[3:0] s2520, in2520_1, in2520_2;
    wire c2520;
    assign in2520_1 = {s903[1],s885[2],s865[3],s981[0]};
    assign in2520_2 = {c904,c887,s866[3],s982[0]};
    CLA_4 KS_2520(s2520, c2520, in2520_1, in2520_2);
    wire[3:0] s2521, in2521_1, in2521_2;
    wire c2521;
    assign in2521_1 = {s905[1],s889[2],s867[3],s983[0]};
    assign in2521_2 = {c906,c891,s868[3],s984[0]};
    CLA_4 KS_2521(s2521, c2521, in2521_1, in2521_2);
    wire[3:0] s2522, in2522_1, in2522_2;
    wire c2522;
    assign in2522_1 = {s907[1],s893[2],s869[3],s985[0]};
    assign in2522_2 = {c908,c895,c870,s986[0]};
    CLA_4 KS_2522(s2522, c2522, in2522_1, in2522_2);
    wire[0:0] s2523, in2523_1, in2523_2;
    wire c2523;
    assign in2523_1 = {s909[1]};
    assign in2523_2 = {c910};
    Half_Adder KS_2523(s2523, c2523, in2523_1, in2523_2);
    wire[1:0] s2524, in2524_1, in2524_2;
    wire c2524;
    assign in2524_1 = {s911[1],s897[2]};
    assign in2524_2 = {c912,c899};
    CLA_2 KS_2524(s2524, c2524, in2524_1, in2524_2);
    wire[0:0] s2525, in2525_1, in2525_2;
    wire c2525;
    assign in2525_1 = {s913[1]};
    assign in2525_2 = {c914};
    Half_Adder KS_2525(s2525, c2525, in2525_1, in2525_2);
    wire[2:0] s2526, in2526_1, in2526_2;
    wire c2526;
    assign in2526_1 = {s915[1],s901[2],s873[3]};
    assign in2526_2 = {c916,c903,c877};
    CLA_3 KS_2526(s2526, c2526, in2526_1, in2526_2);
    wire[0:0] s2527, in2527_1, in2527_2;
    wire c2527;
    assign in2527_1 = {s917[1]};
    assign in2527_2 = {c918};
    Half_Adder KS_2527(s2527, c2527, in2527_1, in2527_2);
    wire[1:0] s2528, in2528_1, in2528_2;
    wire c2528;
    assign in2528_1 = {s919[1],s905[2]};
    assign in2528_2 = {c2426,c907};
    CLA_2 KS_2528(s2528, c2528, in2528_1, in2528_2);
    wire[0:0] s2529, in2529_1, in2529_2;
    wire c2529;
    assign in2529_1 = {c2427};
    assign in2529_2 = {c2428};
    Half_Adder KS_2529(s2529, c2529, in2529_1, in2529_2);
    wire[3:0] s2530, in2530_1, in2530_2;
    wire c2530;
    assign in2530_1 = {c2429,s909[2],s881[3],s987[0]};
    assign in2530_2 = {c2430,c911,c885,s988[0]};
    CLA_4 KS_2530(s2530, c2530, in2530_1, in2530_2);
    wire[0:0] s2531, in2531_1, in2531_2;
    wire c2531;
    assign in2531_1 = {c2431};
    assign in2531_2 = {c2432};
    Half_Adder KS_2531(s2531, c2531, in2531_1, in2531_2);
    wire[1:0] s2532, in2532_1, in2532_2;
    wire c2532;
    assign in2532_1 = {c2433,s913[2]};
    assign in2532_2 = {c2434,c915};
    CLA_2 KS_2532(s2532, c2532, in2532_1, in2532_2);
    wire[0:0] s2533, in2533_1, in2533_2;
    wire c2533;
    assign in2533_1 = {c2435};
    assign in2533_2 = {c2436};
    Half_Adder KS_2533(s2533, c2533, in2533_1, in2533_2);
    wire[2:0] s2534, in2534_1, in2534_2;
    wire c2534;
    assign in2534_1 = {c2437,s917[2],s889[3]};
    assign in2534_2 = {c2438,c919,c893};
    CLA_3 KS_2534(s2534, c2534, in2534_1, in2534_2);
    wire[0:0] s2535, in2535_1, in2535_2;
    wire c2535;
    assign in2535_1 = {c2439};
    assign in2535_2 = {c2440};
    Half_Adder KS_2535(s2535, c2535, in2535_1, in2535_2);
    wire[1:0] s2536, in2536_1, in2536_2;
    wire c2536;
    assign in2536_1 = {c2441,s2491[1]};
    assign in2536_2 = {c2442,s2492[1]};
    CLA_2 KS_2536(s2536, c2536, in2536_1, in2536_2);
    wire[0:0] s2537, in2537_1, in2537_2;
    wire c2537;
    assign in2537_1 = {c2443};
    assign in2537_2 = {c2444};
    Half_Adder KS_2537(s2537, c2537, in2537_1, in2537_2);
    wire[3:0] s2538, in2538_1, in2538_2;
    wire c2538;
    assign in2538_1 = {c2445,s2493[1],s897[3],s989[0]};
    assign in2538_2 = {c2446,s2494[1],c901,s990[0]};
    CLA_4 KS_2538(s2538, c2538, in2538_1, in2538_2);
    wire[0:0] s2539, in2539_1, in2539_2;
    wire c2539;
    assign in2539_1 = {c2447};
    assign in2539_2 = {c2448};
    Half_Adder KS_2539(s2539, c2539, in2539_1, in2539_2);
    wire[1:0] s2540, in2540_1, in2540_2;
    wire c2540;
    assign in2540_1 = {c2449,s2495[1]};
    assign in2540_2 = {c2450,s2496[1]};
    CLA_2 KS_2540(s2540, c2540, in2540_1, in2540_2);
    wire[0:0] s2541, in2541_1, in2541_2;
    wire c2541;
    assign in2541_1 = {c2451};
    assign in2541_2 = {c2452};
    Half_Adder KS_2541(s2541, c2541, in2541_1, in2541_2);
    wire[2:0] s2542, in2542_1, in2542_2;
    wire c2542;
    assign in2542_1 = {c2453,s2497[1],s905[3]};
    assign in2542_2 = {c2454,s2498[1],c909};
    CLA_3 KS_2542(s2542, c2542, in2542_1, in2542_2);
    wire[0:0] s2543, in2543_1, in2543_2;
    wire c2543;
    assign in2543_1 = {c2455};
    assign in2543_2 = {c2456};
    Half_Adder KS_2543(s2543, c2543, in2543_1, in2543_2);
    wire[1:0] s2544, in2544_1, in2544_2;
    wire c2544;
    assign in2544_1 = {c2459,s2499[1]};
    assign in2544_2 = {c2467,s2500[1]};
    CLA_2 KS_2544(s2544, c2544, in2544_1, in2544_2);
    wire[0:0] s2545, in2545_1, in2545_2;
    wire c2545;
    assign in2545_1 = {c2475};
    assign in2545_2 = {c2483};
    Half_Adder KS_2545(s2545, c2545, in2545_1, in2545_2);
    wire[3:0] s2546, in2546_1, in2546_2;
    wire c2546;
    assign in2546_1 = {s2491[0],s2501[1],s913[3],s991[0]};
    assign in2546_2 = {s2492[0],s2502[1],c917,s992[0]};
    CLA_4 KS_2546(s2546, c2546, in2546_1, in2546_2);
    wire[0:0] s2547, in2547_1, in2547_2;
    wire c2547;
    assign in2547_1 = {s2493[0]};
    assign in2547_2 = {s2494[0]};
    Half_Adder KS_2547(s2547, c2547, in2547_1, in2547_2);
    wire[1:0] s2548, in2548_1, in2548_2;
    wire c2548;
    assign in2548_1 = {s2495[0],s2503[1]};
    assign in2548_2 = {s2496[0],s2504[1]};
    CLA_2 KS_2548(s2548, c2548, in2548_1, in2548_2);
    wire[0:0] s2549, in2549_1, in2549_2;
    wire c2549;
    assign in2549_1 = {s2497[0]};
    assign in2549_2 = {s2498[0]};
    Half_Adder KS_2549(s2549, c2549, in2549_1, in2549_2);
    wire[2:0] s2550, in2550_1, in2550_2;
    wire c2550;
    assign in2550_1 = {s2499[0],s2505[1],s2491[2]};
    assign in2550_2 = {s2500[0],s2506[1],s2492[2]};
    CLA_3 KS_2550(s2550, c2550, in2550_1, in2550_2);
    wire[0:0] s2551, in2551_1, in2551_2;
    wire c2551;
    assign in2551_1 = {s2501[0]};
    assign in2551_2 = {s2502[0]};
    Half_Adder KS_2551(s2551, c2551, in2551_1, in2551_2);
    wire[1:0] s2552, in2552_1, in2552_2;
    wire c2552;
    assign in2552_1 = {s2503[0],s2507[1]};
    assign in2552_2 = {s2504[0],s2508[1]};
    CLA_2 KS_2552(s2552, c2552, in2552_1, in2552_2);
    wire[0:0] s2553, in2553_1, in2553_2;
    wire c2553;
    assign in2553_1 = {s2505[0]};
    assign in2553_2 = {s2506[0]};
    Half_Adder KS_2553(s2553, c2553, in2553_1, in2553_2);
    wire[3:0] s2554, in2554_1, in2554_2;
    wire c2554;
    assign in2554_1 = {s2508[0],s2509[1],s2493[2],s993[0]};
    assign in2554_2 = {s2509[0],s2510[1],s2494[2],s994[0]};
    CLA_4_c KS_2554(s2554, c2554, in2554_1, in2554_2, s2507[0]);
    wire[3:0] s2555, in2555_1, in2555_2;
    wire c2555;
    assign in2555_1 = {s923[1],pp110[35],pp99[47],c965};
    assign in2555_2 = {s924[1],pp111[34],pp100[46],c973};
    CLA_4 KS_2555(s2555, c2555, in2555_1, in2555_2);
    wire[3:0] s2556, in2556_1, in2556_2;
    wire c2556;
    assign in2556_1 = {s925[1],pp112[33],pp101[45],c981};
    assign in2556_2 = {s926[1],pp113[32],pp102[44],c989};
    CLA_4 KS_2556(s2556, c2556, in2556_1, in2556_2);
    wire[3:0] s2557, in2557_1, in2557_2;
    wire c2557;
    assign in2557_1 = {s927[1],pp114[31],pp103[43],c997};
    assign in2557_2 = {s928[1],pp115[30],pp104[42],s999[0]};
    CLA_4 KS_2557(s2557, c2557, in2557_1, in2557_2);
    wire[3:0] s2558, in2558_1, in2558_2;
    wire c2558;
    assign in2558_1 = {s929[1],pp116[29],pp105[41],s1000[0]};
    assign in2558_2 = {s930[1],pp117[28],pp106[40],s1001[0]};
    CLA_4 KS_2558(s2558, c2558, in2558_1, in2558_2);
    wire[3:0] s2559, in2559_1, in2559_2;
    wire c2559;
    assign in2559_1 = {s931[1],pp118[27],pp107[39],s1002[0]};
    assign in2559_2 = {s932[1],pp119[26],pp108[38],s1003[0]};
    CLA_4 KS_2559(s2559, c2559, in2559_1, in2559_2);
    wire[3:0] s2560, in2560_1, in2560_2;
    wire c2560;
    assign in2560_1 = {s933[1],pp120[25],pp109[37],s1004[0]};
    assign in2560_2 = {s934[1],pp121[24],pp110[36],s1005[0]};
    CLA_4 KS_2560(s2560, c2560, in2560_1, in2560_2);
    wire[3:0] s2561, in2561_1, in2561_2;
    wire c2561;
    assign in2561_1 = {s935[1],pp122[23],pp111[35],s1006[0]};
    assign in2561_2 = {s936[1],pp123[22],pp112[34],s1007[0]};
    CLA_4 KS_2561(s2561, c2561, in2561_1, in2561_2);
    wire[3:0] s2562, in2562_1, in2562_2;
    wire c2562;
    assign in2562_1 = {s937[1],pp124[21],pp113[33],s1008[0]};
    assign in2562_2 = {s938[1],pp125[20],pp114[32],s1009[0]};
    CLA_4 KS_2562(s2562, c2562, in2562_1, in2562_2);
    wire[3:0] s2563, in2563_1, in2563_2;
    wire c2563;
    assign in2563_1 = {s939[1],pp126[19],pp115[31],s1010[0]};
    assign in2563_2 = {s940[1],pp127[18],pp116[30],s1011[0]};
    CLA_4 KS_2563(s2563, c2563, in2563_1, in2563_2);
    wire[3:0] s2564, in2564_1, in2564_2;
    wire c2564;
    assign in2564_1 = {s941[1],s920[2],pp117[29],s1012[0]};
    assign in2564_2 = {s942[1],s921[2],pp118[28],s1013[0]};
    CLA_4 KS_2564(s2564, c2564, in2564_1, in2564_2);
    wire[3:0] s2565, in2565_1, in2565_2;
    wire c2565;
    assign in2565_1 = {s943[1],s922[2],pp119[27],s1014[0]};
    assign in2565_2 = {s944[1],s923[2],pp120[26],s1015[0]};
    CLA_4 KS_2565(s2565, c2565, in2565_1, in2565_2);
    wire[3:0] s2566, in2566_1, in2566_2;
    wire c2566;
    assign in2566_1 = {s945[1],s924[2],pp121[25],s1016[0]};
    assign in2566_2 = {s946[1],s925[2],pp122[24],s1017[0]};
    CLA_4 KS_2566(s2566, c2566, in2566_1, in2566_2);
    wire[3:0] s2567, in2567_1, in2567_2;
    wire c2567;
    assign in2567_1 = {s947[1],s926[2],pp123[23],s1018[0]};
    assign in2567_2 = {s948[1],s927[2],pp124[22],s1019[0]};
    CLA_4 KS_2567(s2567, c2567, in2567_1, in2567_2);
    wire[3:0] s2568, in2568_1, in2568_2;
    wire c2568;
    assign in2568_1 = {s949[1],s928[2],pp125[21],s1020[0]};
    assign in2568_2 = {s950[1],s929[2],pp126[20],s1021[0]};
    CLA_4 KS_2568(s2568, c2568, in2568_1, in2568_2);
    wire[3:0] s2569, in2569_1, in2569_2;
    wire c2569;
    assign in2569_1 = {s951[1],s930[2],pp127[19],s1022[0]};
    assign in2569_2 = {s952[1],s931[2],s920[3],s1023[0]};
    CLA_4 KS_2569(s2569, c2569, in2569_1, in2569_2);
    wire[3:0] s2570, in2570_1, in2570_2;
    wire c2570;
    assign in2570_1 = {s953[1],s932[2],s921[3],s1024[0]};
    assign in2570_2 = {s954[1],s933[2],s922[3],s1025[0]};
    CLA_4 KS_2570(s2570, c2570, in2570_1, in2570_2);
    wire[3:0] s2571, in2571_1, in2571_2;
    wire c2571;
    assign in2571_1 = {s955[1],s934[2],s923[3],s1026[0]};
    assign in2571_2 = {c956,s935[2],s924[3],s1027[0]};
    CLA_4 KS_2571(s2571, c2571, in2571_1, in2571_2);
    wire[3:0] s2572, in2572_1, in2572_2;
    wire c2572;
    assign in2572_1 = {s957[1],s936[2],s925[3],s1028[0]};
    assign in2572_2 = {c958,s937[2],s926[3],s1029[0]};
    CLA_4 KS_2572(s2572, c2572, in2572_1, in2572_2);
    wire[3:0] s2573, in2573_1, in2573_2;
    wire c2573;
    assign in2573_1 = {s959[1],s938[2],s927[3],s1030[0]};
    assign in2573_2 = {c960,s939[2],s928[3],s1031[0]};
    CLA_4 KS_2573(s2573, c2573, in2573_1, in2573_2);
    wire[3:0] s2574, in2574_1, in2574_2;
    wire c2574;
    assign in2574_1 = {s961[1],s940[2],s929[3],s1032[0]};
    assign in2574_2 = {c962,s941[2],s930[3],s1033[0]};
    CLA_4 KS_2574(s2574, c2574, in2574_1, in2574_2);
    wire[3:0] s2575, in2575_1, in2575_2;
    wire c2575;
    assign in2575_1 = {s963[1],s942[2],s931[3],s1034[0]};
    assign in2575_2 = {c964,s943[2],s932[3],s1035[0]};
    CLA_4 KS_2575(s2575, c2575, in2575_1, in2575_2);
    wire[3:0] s2576, in2576_1, in2576_2;
    wire c2576;
    assign in2576_1 = {s965[1],s944[2],s933[3],s1036[0]};
    assign in2576_2 = {c966,s945[2],s934[3],s1037[0]};
    CLA_4 KS_2576(s2576, c2576, in2576_1, in2576_2);
    wire[3:0] s2577, in2577_1, in2577_2;
    wire c2577;
    assign in2577_1 = {s967[1],s946[2],s935[3],s1038[0]};
    assign in2577_2 = {c968,s947[2],s936[3],s1039[0]};
    CLA_4 KS_2577(s2577, c2577, in2577_1, in2577_2);
    wire[3:0] s2578, in2578_1, in2578_2;
    wire c2578;
    assign in2578_1 = {s969[1],s948[2],s937[3],s1040[0]};
    assign in2578_2 = {c970,s949[2],s938[3],s1041[0]};
    CLA_4 KS_2578(s2578, c2578, in2578_1, in2578_2);
    wire[3:0] s2579, in2579_1, in2579_2;
    wire c2579;
    assign in2579_1 = {s971[1],s950[2],s939[3],s1042[0]};
    assign in2579_2 = {c972,s951[2],s940[3],s1043[0]};
    CLA_4 KS_2579(s2579, c2579, in2579_1, in2579_2);
    wire[3:0] s2580, in2580_1, in2580_2;
    wire c2580;
    assign in2580_1 = {s973[1],s952[2],s941[3],s1044[0]};
    assign in2580_2 = {c974,s953[2],s942[3],s1045[0]};
    CLA_4 KS_2580(s2580, c2580, in2580_1, in2580_2);
    wire[3:0] s2581, in2581_1, in2581_2;
    wire c2581;
    assign in2581_1 = {s975[1],s954[2],s943[3],s1046[0]};
    assign in2581_2 = {c976,c955,s944[3],s1047[0]};
    CLA_4 KS_2581(s2581, c2581, in2581_1, in2581_2);
    wire[3:0] s2582, in2582_1, in2582_2;
    wire c2582;
    assign in2582_1 = {s977[1],s957[2],s945[3],s1048[0]};
    assign in2582_2 = {c978,c959,s946[3],s1049[0]};
    CLA_4 KS_2582(s2582, c2582, in2582_1, in2582_2);
    wire[3:0] s2583, in2583_1, in2583_2;
    wire c2583;
    assign in2583_1 = {s979[1],s961[2],s947[3],s1050[0]};
    assign in2583_2 = {c980,c963,s948[3],s1051[0]};
    CLA_4 KS_2583(s2583, c2583, in2583_1, in2583_2);
    wire[3:0] s2584, in2584_1, in2584_2;
    wire c2584;
    assign in2584_1 = {s981[1],s965[2],s949[3],s1052[0]};
    assign in2584_2 = {c982,c967,s950[3],s1053[0]};
    CLA_4 KS_2584(s2584, c2584, in2584_1, in2584_2);
    wire[3:0] s2585, in2585_1, in2585_2;
    wire c2585;
    assign in2585_1 = {s983[1],s969[2],s951[3],s1054[0]};
    assign in2585_2 = {c984,c971,s952[3],s1055[0]};
    CLA_4 KS_2585(s2585, c2585, in2585_1, in2585_2);
    wire[0:0] s2586, in2586_1, in2586_2;
    wire c2586;
    assign in2586_1 = {s985[1]};
    assign in2586_2 = {c986};
    Half_Adder KS_2586(s2586, c2586, in2586_1, in2586_2);
    wire[1:0] s2587, in2587_1, in2587_2;
    wire c2587;
    assign in2587_1 = {s987[1],s973[2]};
    assign in2587_2 = {c988,c975};
    CLA_2 KS_2587(s2587, c2587, in2587_1, in2587_2);
    wire[0:0] s2588, in2588_1, in2588_2;
    wire c2588;
    assign in2588_1 = {s989[1]};
    assign in2588_2 = {c990};
    Half_Adder KS_2588(s2588, c2588, in2588_1, in2588_2);
    wire[3:0] s2589, in2589_1, in2589_2;
    wire c2589;
    assign in2589_1 = {s991[1],s977[2],s953[3],s1056[0]};
    assign in2589_2 = {c992,c979,c954,s1057[0]};
    CLA_4 KS_2589(s2589, c2589, in2589_1, in2589_2);
    wire[0:0] s2590, in2590_1, in2590_2;
    wire c2590;
    assign in2590_1 = {s993[1]};
    assign in2590_2 = {c994};
    Half_Adder KS_2590(s2590, c2590, in2590_1, in2590_2);
    wire[1:0] s2591, in2591_1, in2591_2;
    wire c2591;
    assign in2591_1 = {s995[1],s981[2]};
    assign in2591_2 = {c996,c983};
    CLA_2 KS_2591(s2591, c2591, in2591_1, in2591_2);
    wire[0:0] s2592, in2592_1, in2592_2;
    wire c2592;
    assign in2592_1 = {s997[1]};
    assign in2592_2 = {c998};
    Half_Adder KS_2592(s2592, c2592, in2592_1, in2592_2);
    wire[2:0] s2593, in2593_1, in2593_2;
    wire c2593;
    assign in2593_1 = {c2491,s985[2],s957[3]};
    assign in2593_2 = {c2492,c987,c961};
    CLA_3 KS_2593(s2593, c2593, in2593_1, in2593_2);
    wire[0:0] s2594, in2594_1, in2594_2;
    wire c2594;
    assign in2594_1 = {c2493};
    assign in2594_2 = {c2494};
    Half_Adder KS_2594(s2594, c2594, in2594_1, in2594_2);
    wire[1:0] s2595, in2595_1, in2595_2;
    wire c2595;
    assign in2595_1 = {c2495,s989[2]};
    assign in2595_2 = {c2496,c991};
    CLA_2 KS_2595(s2595, c2595, in2595_1, in2595_2);
    wire[0:0] s2596, in2596_1, in2596_2;
    wire c2596;
    assign in2596_1 = {c2497};
    assign in2596_2 = {c2498};
    Half_Adder KS_2596(s2596, c2596, in2596_1, in2596_2);
    wire[3:0] s2597, in2597_1, in2597_2;
    wire c2597;
    assign in2597_1 = {c2499,s993[2],s965[3],s1058[0]};
    assign in2597_2 = {c2500,c995,c969,s1059[0]};
    CLA_4 KS_2597(s2597, c2597, in2597_1, in2597_2);
    wire[0:0] s2598, in2598_1, in2598_2;
    wire c2598;
    assign in2598_1 = {c2501};
    assign in2598_2 = {c2502};
    Half_Adder KS_2598(s2598, c2598, in2598_1, in2598_2);
    wire[1:0] s2599, in2599_1, in2599_2;
    wire c2599;
    assign in2599_1 = {c2503,s997[2]};
    assign in2599_2 = {c2504,s2555[1]};
    CLA_2 KS_2599(s2599, c2599, in2599_1, in2599_2);
    wire[0:0] s2600, in2600_1, in2600_2;
    wire c2600;
    assign in2600_1 = {c2505};
    assign in2600_2 = {c2506};
    Half_Adder KS_2600(s2600, c2600, in2600_1, in2600_2);
    wire[2:0] s2601, in2601_1, in2601_2;
    wire c2601;
    assign in2601_1 = {c2507,s2556[1],s973[3]};
    assign in2601_2 = {c2508,s2557[1],c977};
    CLA_3 KS_2601(s2601, c2601, in2601_1, in2601_2);
    wire[0:0] s2602, in2602_1, in2602_2;
    wire c2602;
    assign in2602_1 = {c2509};
    assign in2602_2 = {c2510};
    Half_Adder KS_2602(s2602, c2602, in2602_1, in2602_2);
    wire[1:0] s2603, in2603_1, in2603_2;
    wire c2603;
    assign in2603_1 = {c2511,s2558[1]};
    assign in2603_2 = {c2512,s2559[1]};
    CLA_2 KS_2603(s2603, c2603, in2603_1, in2603_2);
    wire[0:0] s2604, in2604_1, in2604_2;
    wire c2604;
    assign in2604_1 = {c2513};
    assign in2604_2 = {c2514};
    Half_Adder KS_2604(s2604, c2604, in2604_1, in2604_2);
    wire[3:0] s2605, in2605_1, in2605_2;
    wire c2605;
    assign in2605_1 = {c2515,s2560[1],s981[3],s1060[0]};
    assign in2605_2 = {c2516,s2561[1],c985,s1061[0]};
    CLA_4 KS_2605(s2605, c2605, in2605_1, in2605_2);
    wire[0:0] s2606, in2606_1, in2606_2;
    wire c2606;
    assign in2606_1 = {c2517};
    assign in2606_2 = {c2518};
    Half_Adder KS_2606(s2606, c2606, in2606_1, in2606_2);
    wire[1:0] s2607, in2607_1, in2607_2;
    wire c2607;
    assign in2607_1 = {c2519,s2562[1]};
    assign in2607_2 = {c2520,s2563[1]};
    CLA_2 KS_2607(s2607, c2607, in2607_1, in2607_2);
    wire[0:0] s2608, in2608_1, in2608_2;
    wire c2608;
    assign in2608_1 = {c2521};
    assign in2608_2 = {c2522};
    Half_Adder KS_2608(s2608, c2608, in2608_1, in2608_2);
    wire[2:0] s2609, in2609_1, in2609_2;
    wire c2609;
    assign in2609_1 = {c2530,s2564[1],s989[3]};
    assign in2609_2 = {c2538,s2565[1],c993};
    CLA_3 KS_2609(s2609, c2609, in2609_1, in2609_2);
    wire[0:0] s2610, in2610_1, in2610_2;
    wire c2610;
    assign in2610_1 = {c2546};
    assign in2610_2 = {c2554};
    Half_Adder KS_2610(s2610, c2610, in2610_1, in2610_2);
    wire[1:0] s2611, in2611_1, in2611_2;
    wire c2611;
    assign in2611_1 = {s2555[0],s2566[1]};
    assign in2611_2 = {s2556[0],s2567[1]};
    CLA_2 KS_2611(s2611, c2611, in2611_1, in2611_2);
    wire[0:0] s2612, in2612_1, in2612_2;
    wire c2612;
    assign in2612_1 = {s2557[0]};
    assign in2612_2 = {s2558[0]};
    Half_Adder KS_2612(s2612, c2612, in2612_1, in2612_2);
    wire[3:0] s2613, in2613_1, in2613_2;
    wire c2613;
    assign in2613_1 = {s2559[0],s2568[1],s997[3],s1062[0]};
    assign in2613_2 = {s2560[0],s2569[1],s2555[2],s1063[0]};
    CLA_4 KS_2613(s2613, c2613, in2613_1, in2613_2);
    wire[0:0] s2614, in2614_1, in2614_2;
    wire c2614;
    assign in2614_1 = {s2561[0]};
    assign in2614_2 = {s2562[0]};
    Half_Adder KS_2614(s2614, c2614, in2614_1, in2614_2);
    wire[1:0] s2615, in2615_1, in2615_2;
    wire c2615;
    assign in2615_1 = {s2563[0],s2570[1]};
    assign in2615_2 = {s2564[0],s2571[1]};
    CLA_2 KS_2615(s2615, c2615, in2615_1, in2615_2);
    wire[0:0] s2616, in2616_1, in2616_2;
    wire c2616;
    assign in2616_1 = {s2565[0]};
    assign in2616_2 = {s2566[0]};
    Half_Adder KS_2616(s2616, c2616, in2616_1, in2616_2);
    wire[2:0] s2617, in2617_1, in2617_2;
    wire c2617;
    assign in2617_1 = {s2567[0],s2572[1],s2556[2]};
    assign in2617_2 = {s2568[0],s2573[1],s2557[2]};
    CLA_3 KS_2617(s2617, c2617, in2617_1, in2617_2);
    wire[0:0] s2618, in2618_1, in2618_2;
    wire c2618;
    assign in2618_1 = {s2569[0]};
    assign in2618_2 = {s2570[0]};
    Half_Adder KS_2618(s2618, c2618, in2618_1, in2618_2);
    wire[1:0] s2619, in2619_1, in2619_2;
    wire c2619;
    assign in2619_1 = {s2571[0],s2574[1]};
    assign in2619_2 = {s2572[0],s2575[1]};
    CLA_2 KS_2619(s2619, c2619, in2619_1, in2619_2);
    wire[0:0] s2620, in2620_1, in2620_2;
    wire c2620;
    assign in2620_1 = {s2574[0]};
    assign in2620_2 = {s2575[0]};
    Full_Adder KS_2620(s2620, c2620, in2620_1, in2620_2, s2573[0]);
    wire[3:0] s2621, in2621_1, in2621_2;
    wire c2621;
    assign in2621_1 = {pp123[25],pp104[45],pp93[57],c1020};
    assign in2621_2 = {pp124[24],pp105[44],pp94[56],c1021};
    CLA_4 KS_2621(s2621, c2621, in2621_1, in2621_2);
    wire[3:0] s2622, in2622_1, in2622_2;
    wire c2622;
    assign in2622_1 = {pp125[23],pp106[43],pp95[55],c1022};
    assign in2622_2 = {pp126[22],pp107[42],pp96[54],c1023};
    CLA_4 KS_2622(s2622, c2622, in2622_1, in2622_2);
    wire[3:0] s2623, in2623_1, in2623_2;
    wire c2623;
    assign in2623_1 = {pp127[21],pp108[41],pp97[53],c1024};
    assign in2623_2 = {s999[1],pp109[40],pp98[52],c1025};
    CLA_4 KS_2623(s2623, c2623, in2623_1, in2623_2);
    wire[3:0] s2624, in2624_1, in2624_2;
    wire c2624;
    assign in2624_1 = {s1000[1],pp110[39],pp99[51],c1026};
    assign in2624_2 = {s1001[1],pp111[38],pp100[50],c1027};
    CLA_4 KS_2624(s2624, c2624, in2624_1, in2624_2);
    wire[3:0] s2625, in2625_1, in2625_2;
    wire c2625;
    assign in2625_1 = {s1002[1],pp112[37],pp101[49],c1028};
    assign in2625_2 = {s1003[1],pp113[36],pp102[48],c1032};
    CLA_4 KS_2625(s2625, c2625, in2625_1, in2625_2);
    wire[3:0] s2626, in2626_1, in2626_2;
    wire c2626;
    assign in2626_1 = {s1004[1],pp114[35],pp103[47],c1040};
    assign in2626_2 = {s1005[1],pp115[34],pp104[46],c1048};
    CLA_4 KS_2626(s2626, c2626, in2626_1, in2626_2);
    wire[3:0] s2627, in2627_1, in2627_2;
    wire c2627;
    assign in2627_1 = {s1006[1],pp116[33],pp105[45],c1056};
    assign in2627_2 = {s1007[1],pp117[32],pp106[44],c1064};
    CLA_4 KS_2627(s2627, c2627, in2627_1, in2627_2);
    wire[3:0] s2628, in2628_1, in2628_2;
    wire c2628;
    assign in2628_1 = {s1008[1],pp118[31],pp107[43],s1070[0]};
    assign in2628_2 = {s1009[1],pp119[30],pp108[42],s1071[0]};
    CLA_4 KS_2628(s2628, c2628, in2628_1, in2628_2);
    wire[3:0] s2629, in2629_1, in2629_2;
    wire c2629;
    assign in2629_1 = {s1010[1],pp120[29],pp109[41],s1072[0]};
    assign in2629_2 = {s1011[1],pp121[28],pp110[40],s1073[0]};
    CLA_4 KS_2629(s2629, c2629, in2629_1, in2629_2);
    wire[3:0] s2630, in2630_1, in2630_2;
    wire c2630;
    assign in2630_1 = {s1012[1],pp122[27],pp111[39],s1074[0]};
    assign in2630_2 = {s1013[1],pp123[26],pp112[38],s1075[0]};
    CLA_4 KS_2630(s2630, c2630, in2630_1, in2630_2);
    wire[3:0] s2631, in2631_1, in2631_2;
    wire c2631;
    assign in2631_1 = {s1014[1],pp124[25],pp113[37],s1076[0]};
    assign in2631_2 = {s1015[1],pp125[24],pp114[36],s1077[0]};
    CLA_4 KS_2631(s2631, c2631, in2631_1, in2631_2);
    wire[3:0] s2632, in2632_1, in2632_2;
    wire c2632;
    assign in2632_1 = {s1016[1],pp126[23],pp115[35],s1078[0]};
    assign in2632_2 = {s1017[1],pp127[22],pp116[34],s1079[0]};
    CLA_4 KS_2632(s2632, c2632, in2632_1, in2632_2);
    wire[3:0] s2633, in2633_1, in2633_2;
    wire c2633;
    assign in2633_1 = {s1018[1],s999[2],pp117[33],s1080[0]};
    assign in2633_2 = {s1019[1],s1000[2],pp118[32],s1081[0]};
    CLA_4 KS_2633(s2633, c2633, in2633_1, in2633_2);
    wire[3:0] s2634, in2634_1, in2634_2;
    wire c2634;
    assign in2634_1 = {s1020[1],s1001[2],pp119[31],s1082[0]};
    assign in2634_2 = {s1021[1],s1002[2],pp120[30],s1083[0]};
    CLA_4 KS_2634(s2634, c2634, in2634_1, in2634_2);
    wire[3:0] s2635, in2635_1, in2635_2;
    wire c2635;
    assign in2635_1 = {s1022[1],s1003[2],pp121[29],s1084[0]};
    assign in2635_2 = {s1023[1],s1004[2],pp122[28],s1085[0]};
    CLA_4 KS_2635(s2635, c2635, in2635_1, in2635_2);
    wire[3:0] s2636, in2636_1, in2636_2;
    wire c2636;
    assign in2636_1 = {s1024[1],s1005[2],pp123[27],s1086[0]};
    assign in2636_2 = {s1025[1],s1006[2],pp124[26],s1087[0]};
    CLA_4 KS_2636(s2636, c2636, in2636_1, in2636_2);
    wire[3:0] s2637, in2637_1, in2637_2;
    wire c2637;
    assign in2637_1 = {s1026[1],s1007[2],pp125[25],s1088[0]};
    assign in2637_2 = {s1027[1],s1008[2],pp126[24],s1089[0]};
    CLA_4 KS_2637(s2637, c2637, in2637_1, in2637_2);
    wire[3:0] s2638, in2638_1, in2638_2;
    wire c2638;
    assign in2638_1 = {s1028[1],s1009[2],pp127[23],s1090[0]};
    assign in2638_2 = {s1029[1],s1010[2],s999[3],s1091[0]};
    CLA_4 KS_2638(s2638, c2638, in2638_1, in2638_2);
    wire[3:0] s2639, in2639_1, in2639_2;
    wire c2639;
    assign in2639_1 = {s1030[1],s1011[2],s1000[3],s1092[0]};
    assign in2639_2 = {c1031,s1012[2],s1001[3],s1093[0]};
    CLA_4 KS_2639(s2639, c2639, in2639_1, in2639_2);
    wire[3:0] s2640, in2640_1, in2640_2;
    wire c2640;
    assign in2640_1 = {s1032[1],s1013[2],s1002[3],s1094[0]};
    assign in2640_2 = {c1033,s1014[2],s1003[3],s1095[0]};
    CLA_4 KS_2640(s2640, c2640, in2640_1, in2640_2);
    wire[3:0] s2641, in2641_1, in2641_2;
    wire c2641;
    assign in2641_1 = {s1034[1],s1015[2],s1004[3],s1096[0]};
    assign in2641_2 = {c1035,s1016[2],s1005[3],s1097[0]};
    CLA_4 KS_2641(s2641, c2641, in2641_1, in2641_2);
    wire[3:0] s2642, in2642_1, in2642_2;
    wire c2642;
    assign in2642_1 = {s1036[1],s1017[2],s1006[3],s1098[0]};
    assign in2642_2 = {c1037,s1018[2],s1007[3],s1099[0]};
    CLA_4 KS_2642(s2642, c2642, in2642_1, in2642_2);
    wire[3:0] s2643, in2643_1, in2643_2;
    wire c2643;
    assign in2643_1 = {s1038[1],s1019[2],s1008[3],s1100[0]};
    assign in2643_2 = {c1039,s1020[2],s1009[3],s1101[0]};
    CLA_4 KS_2643(s2643, c2643, in2643_1, in2643_2);
    wire[3:0] s2644, in2644_1, in2644_2;
    wire c2644;
    assign in2644_1 = {s1040[1],s1021[2],s1010[3],s1102[0]};
    assign in2644_2 = {c1041,s1022[2],s1011[3],s1103[0]};
    CLA_4 KS_2644(s2644, c2644, in2644_1, in2644_2);
    wire[3:0] s2645, in2645_1, in2645_2;
    wire c2645;
    assign in2645_1 = {s1042[1],s1023[2],s1012[3],s1104[0]};
    assign in2645_2 = {c1043,s1024[2],s1013[3],s1105[0]};
    CLA_4 KS_2645(s2645, c2645, in2645_1, in2645_2);
    wire[3:0] s2646, in2646_1, in2646_2;
    wire c2646;
    assign in2646_1 = {s1044[1],s1025[2],s1014[3],s1106[0]};
    assign in2646_2 = {c1045,s1026[2],s1015[3],s1107[0]};
    CLA_4 KS_2646(s2646, c2646, in2646_1, in2646_2);
    wire[3:0] s2647, in2647_1, in2647_2;
    wire c2647;
    assign in2647_1 = {s1046[1],s1027[2],s1016[3],s1108[0]};
    assign in2647_2 = {c1047,s1028[2],s1017[3],s1109[0]};
    CLA_4 KS_2647(s2647, c2647, in2647_1, in2647_2);
    wire[3:0] s2648, in2648_1, in2648_2;
    wire c2648;
    assign in2648_1 = {s1048[1],s1029[2],s1018[3],s1110[0]};
    assign in2648_2 = {c1049,c1030,s1019[3],s1111[0]};
    CLA_4 KS_2648(s2648, c2648, in2648_1, in2648_2);
    wire[3:0] s2649, in2649_1, in2649_2;
    wire c2649;
    assign in2649_1 = {s1050[1],s1032[2],s1020[3],s1112[0]};
    assign in2649_2 = {c1051,c1034,s1021[3],s1113[0]};
    CLA_4 KS_2649(s2649, c2649, in2649_1, in2649_2);
    wire[3:0] s2650, in2650_1, in2650_2;
    wire c2650;
    assign in2650_1 = {s1052[1],s1036[2],s1022[3],s1114[0]};
    assign in2650_2 = {c1053,c1038,s1023[3],s1115[0]};
    CLA_4 KS_2650(s2650, c2650, in2650_1, in2650_2);
    wire[3:0] s2651, in2651_1, in2651_2;
    wire c2651;
    assign in2651_1 = {s1054[1],s1040[2],s1024[3],s1116[0]};
    assign in2651_2 = {c1055,c1042,s1025[3],s1117[0]};
    CLA_4 KS_2651(s2651, c2651, in2651_1, in2651_2);
    wire[0:0] s2652, in2652_1, in2652_2;
    wire c2652;
    assign in2652_1 = {s1056[1]};
    assign in2652_2 = {c1057};
    Half_Adder KS_2652(s2652, c2652, in2652_1, in2652_2);
    wire[3:0] s2653, in2653_1, in2653_2;
    wire c2653;
    assign in2653_1 = {s1058[1],s1044[2],s1026[3],s1118[0]};
    assign in2653_2 = {c1059,c1046,s1027[3],s1119[0]};
    CLA_4 KS_2653(s2653, c2653, in2653_1, in2653_2);
    wire[0:0] s2654, in2654_1, in2654_2;
    wire c2654;
    assign in2654_1 = {s1060[1]};
    assign in2654_2 = {c1061};
    Half_Adder KS_2654(s2654, c2654, in2654_1, in2654_2);
    wire[1:0] s2655, in2655_1, in2655_2;
    wire c2655;
    assign in2655_1 = {s1062[1],s1048[2]};
    assign in2655_2 = {c1063,c1050};
    CLA_2 KS_2655(s2655, c2655, in2655_1, in2655_2);
    wire[0:0] s2656, in2656_1, in2656_2;
    wire c2656;
    assign in2656_1 = {s1064[1]};
    assign in2656_2 = {c1065};
    Half_Adder KS_2656(s2656, c2656, in2656_1, in2656_2);
    wire[2:0] s2657, in2657_1, in2657_2;
    wire c2657;
    assign in2657_1 = {s1066[1],s1052[2],s1028[3]};
    assign in2657_2 = {c1067,c1054,c1029};
    CLA_3 KS_2657(s2657, c2657, in2657_1, in2657_2);
    wire[0:0] s2658, in2658_1, in2658_2;
    wire c2658;
    assign in2658_1 = {s1068[1]};
    assign in2658_2 = {c1069};
    Half_Adder KS_2658(s2658, c2658, in2658_1, in2658_2);
    wire[1:0] s2659, in2659_1, in2659_2;
    wire c2659;
    assign in2659_1 = {c2555,s1056[2]};
    assign in2659_2 = {c2556,c1058};
    CLA_2 KS_2659(s2659, c2659, in2659_1, in2659_2);
    wire[0:0] s2660, in2660_1, in2660_2;
    wire c2660;
    assign in2660_1 = {c2557};
    assign in2660_2 = {c2558};
    Half_Adder KS_2660(s2660, c2660, in2660_1, in2660_2);
    wire[3:0] s2661, in2661_1, in2661_2;
    wire c2661;
    assign in2661_1 = {c2559,s1060[2],s1032[3],s1120[0]};
    assign in2661_2 = {c2560,c1062,c1036,s1121[0]};
    CLA_4 KS_2661(s2661, c2661, in2661_1, in2661_2);
    wire[0:0] s2662, in2662_1, in2662_2;
    wire c2662;
    assign in2662_1 = {c2561};
    assign in2662_2 = {c2562};
    Half_Adder KS_2662(s2662, c2662, in2662_1, in2662_2);
    wire[1:0] s2663, in2663_1, in2663_2;
    wire c2663;
    assign in2663_1 = {c2563,s1064[2]};
    assign in2663_2 = {c2564,c1066};
    CLA_2 KS_2663(s2663, c2663, in2663_1, in2663_2);
    wire[0:0] s2664, in2664_1, in2664_2;
    wire c2664;
    assign in2664_1 = {c2565};
    assign in2664_2 = {c2566};
    Half_Adder KS_2664(s2664, c2664, in2664_1, in2664_2);
    wire[2:0] s2665, in2665_1, in2665_2;
    wire c2665;
    assign in2665_1 = {c2567,s1068[2],s1040[3]};
    assign in2665_2 = {c2568,s2621[1],c1044};
    CLA_3 KS_2665(s2665, c2665, in2665_1, in2665_2);
    wire[0:0] s2666, in2666_1, in2666_2;
    wire c2666;
    assign in2666_1 = {c2569};
    assign in2666_2 = {c2570};
    Half_Adder KS_2666(s2666, c2666, in2666_1, in2666_2);
    wire[1:0] s2667, in2667_1, in2667_2;
    wire c2667;
    assign in2667_1 = {c2571,s2622[1]};
    assign in2667_2 = {c2572,s2623[1]};
    CLA_2 KS_2667(s2667, c2667, in2667_1, in2667_2);
    wire[0:0] s2668, in2668_1, in2668_2;
    wire c2668;
    assign in2668_1 = {c2573};
    assign in2668_2 = {c2574};
    Half_Adder KS_2668(s2668, c2668, in2668_1, in2668_2);
    wire[3:0] s2669, in2669_1, in2669_2;
    wire c2669;
    assign in2669_1 = {c2575,s2624[1],s1048[3],s1122[0]};
    assign in2669_2 = {c2576,s2625[1],c1052,s1123[0]};
    CLA_4 KS_2669(s2669, c2669, in2669_1, in2669_2);
    wire[0:0] s2670, in2670_1, in2670_2;
    wire c2670;
    assign in2670_1 = {c2577};
    assign in2670_2 = {c2578};
    Half_Adder KS_2670(s2670, c2670, in2670_1, in2670_2);
    wire[1:0] s2671, in2671_1, in2671_2;
    wire c2671;
    assign in2671_1 = {c2579,s2626[1]};
    assign in2671_2 = {c2580,s2627[1]};
    CLA_2 KS_2671(s2671, c2671, in2671_1, in2671_2);
    wire[0:0] s2672, in2672_1, in2672_2;
    wire c2672;
    assign in2672_1 = {c2581};
    assign in2672_2 = {c2582};
    Half_Adder KS_2672(s2672, c2672, in2672_1, in2672_2);
    wire[2:0] s2673, in2673_1, in2673_2;
    wire c2673;
    assign in2673_1 = {c2583,s2628[1],s1056[3]};
    assign in2673_2 = {c2584,s2629[1],c1060};
    CLA_3 KS_2673(s2673, c2673, in2673_1, in2673_2);
    wire[0:0] s2674, in2674_1, in2674_2;
    wire c2674;
    assign in2674_1 = {c2585};
    assign in2674_2 = {c2589};
    Half_Adder KS_2674(s2674, c2674, in2674_1, in2674_2);
    wire[1:0] s2675, in2675_1, in2675_2;
    wire c2675;
    assign in2675_1 = {c2597,s2630[1]};
    assign in2675_2 = {c2605,s2631[1]};
    CLA_2 KS_2675(s2675, c2675, in2675_1, in2675_2);
    wire[0:0] s2676, in2676_1, in2676_2;
    wire c2676;
    assign in2676_1 = {c2613};
    assign in2676_2 = {s2621[0]};
    Half_Adder KS_2676(s2676, c2676, in2676_1, in2676_2);
    wire[3:0] s2677, in2677_1, in2677_2;
    wire c2677;
    assign in2677_1 = {s2622[0],s2632[1],s1064[3],s1124[0]};
    assign in2677_2 = {s2623[0],s2633[1],c1068,s1125[0]};
    CLA_4 KS_2677(s2677, c2677, in2677_1, in2677_2);
    wire[0:0] s2678, in2678_1, in2678_2;
    wire c2678;
    assign in2678_1 = {s2624[0]};
    assign in2678_2 = {s2625[0]};
    Half_Adder KS_2678(s2678, c2678, in2678_1, in2678_2);
    wire[1:0] s2679, in2679_1, in2679_2;
    wire c2679;
    assign in2679_1 = {s2626[0],s2634[1]};
    assign in2679_2 = {s2627[0],s2635[1]};
    CLA_2 KS_2679(s2679, c2679, in2679_1, in2679_2);
    wire[0:0] s2680, in2680_1, in2680_2;
    wire c2680;
    assign in2680_1 = {s2628[0]};
    assign in2680_2 = {s2629[0]};
    Half_Adder KS_2680(s2680, c2680, in2680_1, in2680_2);
    wire[2:0] s2681, in2681_1, in2681_2;
    wire c2681;
    assign in2681_1 = {s2630[0],s2636[1],s2621[2]};
    assign in2681_2 = {s2631[0],s2637[1],s2622[2]};
    CLA_3 KS_2681(s2681, c2681, in2681_1, in2681_2);
    wire[0:0] s2682, in2682_1, in2682_2;
    wire c2682;
    assign in2682_1 = {s2632[0]};
    assign in2682_2 = {s2633[0]};
    Half_Adder KS_2682(s2682, c2682, in2682_1, in2682_2);
    wire[1:0] s2683, in2683_1, in2683_2;
    wire c2683;
    assign in2683_1 = {s2634[0],s2638[1]};
    assign in2683_2 = {s2635[0],s2639[1]};
    CLA_2 KS_2683(s2683, c2683, in2683_1, in2683_2);
    wire[0:0] s2684, in2684_1, in2684_2;
    wire c2684;
    assign in2684_1 = {s2636[0]};
    assign in2684_2 = {s2637[0]};
    Half_Adder KS_2684(s2684, c2684, in2684_1, in2684_2);
    wire[3:0] s2685, in2685_1, in2685_2;
    wire c2685;
    assign in2685_1 = {s2639[0],s2640[1],s2623[2],s1126[0]};
    assign in2685_2 = {s2640[0],s2641[1],s2624[2],s1127[0]};
    CLA_4_c KS_2685(s2685, c2685, in2685_1, in2685_2, s2638[0]);
    wire[3:0] s2686, in2686_1, in2686_2;
    wire c2686;
    assign in2686_1 = {pp115[37],pp98[55],pp89[65],c1079};
    assign in2686_2 = {pp116[36],pp99[54],pp90[64],c1080};
    CLA_4 KS_2686(s2686, c2686, in2686_1, in2686_2);
    wire[3:0] s2687, in2687_1, in2687_2;
    wire c2687;
    assign in2687_1 = {pp117[35],pp100[53],pp91[63],c1081};
    assign in2687_2 = {pp118[34],pp101[52],pp92[62],c1082};
    CLA_4 KS_2687(s2687, c2687, in2687_1, in2687_2);
    wire[3:0] s2688, in2688_1, in2688_2;
    wire c2688;
    assign in2688_1 = {pp119[33],pp102[51],pp93[61],c1083};
    assign in2688_2 = {pp120[32],pp103[50],pp94[60],c1084};
    CLA_4 KS_2688(s2688, c2688, in2688_1, in2688_2);
    wire[3:0] s2689, in2689_1, in2689_2;
    wire c2689;
    assign in2689_1 = {pp121[31],pp104[49],pp95[59],c1085};
    assign in2689_2 = {pp122[30],pp105[48],pp96[58],c1086};
    CLA_4 KS_2689(s2689, c2689, in2689_1, in2689_2);
    wire[3:0] s2690, in2690_1, in2690_2;
    wire c2690;
    assign in2690_1 = {pp123[29],pp106[47],pp97[57],c1087};
    assign in2690_2 = {pp124[28],pp107[46],pp98[56],c1088};
    CLA_4 KS_2690(s2690, c2690, in2690_1, in2690_2);
    wire[3:0] s2691, in2691_1, in2691_2;
    wire c2691;
    assign in2691_1 = {pp125[27],pp108[45],pp99[55],c1089};
    assign in2691_2 = {pp126[26],pp109[44],pp100[54],c1090};
    CLA_4 KS_2691(s2691, c2691, in2691_1, in2691_2);
    wire[3:0] s2692, in2692_1, in2692_2;
    wire c2692;
    assign in2692_1 = {pp127[25],pp110[43],pp101[53],c1091};
    assign in2692_2 = {s1070[1],pp111[42],pp102[52],c1092};
    CLA_4 KS_2692(s2692, c2692, in2692_1, in2692_2);
    wire[3:0] s2693, in2693_1, in2693_2;
    wire c2693;
    assign in2693_1 = {s1071[1],pp112[41],pp103[51],c1093};
    assign in2693_2 = {s1072[1],pp113[40],pp104[50],c1094};
    CLA_4 KS_2693(s2693, c2693, in2693_1, in2693_2);
    wire[3:0] s2694, in2694_1, in2694_2;
    wire c2694;
    assign in2694_1 = {s1073[1],pp114[39],pp105[49],c1095};
    assign in2694_2 = {s1074[1],pp115[38],pp106[48],c1099};
    CLA_4 KS_2694(s2694, c2694, in2694_1, in2694_2);
    wire[3:0] s2695, in2695_1, in2695_2;
    wire c2695;
    assign in2695_1 = {s1075[1],pp116[37],pp107[47],c1107};
    assign in2695_2 = {s1076[1],pp117[36],pp108[46],c1115};
    CLA_4 KS_2695(s2695, c2695, in2695_1, in2695_2);
    wire[3:0] s2696, in2696_1, in2696_2;
    wire c2696;
    assign in2696_1 = {s1077[1],pp118[35],pp109[45],c1123};
    assign in2696_2 = {s1078[1],pp119[34],pp110[44],c1131};
    CLA_4 KS_2696(s2696, c2696, in2696_1, in2696_2);
    wire[3:0] s2697, in2697_1, in2697_2;
    wire c2697;
    assign in2697_1 = {s1079[1],pp120[33],pp111[43],s1132[0]};
    assign in2697_2 = {s1080[1],pp121[32],pp112[42],s1133[0]};
    CLA_4 KS_2697(s2697, c2697, in2697_1, in2697_2);
    wire[3:0] s2698, in2698_1, in2698_2;
    wire c2698;
    assign in2698_1 = {s1081[1],pp122[31],pp113[41],s1134[0]};
    assign in2698_2 = {s1082[1],pp123[30],pp114[40],s1135[0]};
    CLA_4 KS_2698(s2698, c2698, in2698_1, in2698_2);
    wire[3:0] s2699, in2699_1, in2699_2;
    wire c2699;
    assign in2699_1 = {s1083[1],pp124[29],pp115[39],s1136[0]};
    assign in2699_2 = {s1084[1],pp125[28],pp116[38],s1137[0]};
    CLA_4 KS_2699(s2699, c2699, in2699_1, in2699_2);
    wire[3:0] s2700, in2700_1, in2700_2;
    wire c2700;
    assign in2700_1 = {s1085[1],pp126[27],pp117[37],s1138[0]};
    assign in2700_2 = {s1086[1],pp127[26],pp118[36],s1139[0]};
    CLA_4 KS_2700(s2700, c2700, in2700_1, in2700_2);
    wire[3:0] s2701, in2701_1, in2701_2;
    wire c2701;
    assign in2701_1 = {s1087[1],s1070[2],pp119[35],s1140[0]};
    assign in2701_2 = {s1088[1],s1071[2],pp120[34],s1141[0]};
    CLA_4 KS_2701(s2701, c2701, in2701_1, in2701_2);
    wire[3:0] s2702, in2702_1, in2702_2;
    wire c2702;
    assign in2702_1 = {s1089[1],s1072[2],pp121[33],s1142[0]};
    assign in2702_2 = {s1090[1],s1073[2],pp122[32],s1143[0]};
    CLA_4 KS_2702(s2702, c2702, in2702_1, in2702_2);
    wire[3:0] s2703, in2703_1, in2703_2;
    wire c2703;
    assign in2703_1 = {s1091[1],s1074[2],pp123[31],s1144[0]};
    assign in2703_2 = {s1092[1],s1075[2],pp124[30],s1145[0]};
    CLA_4 KS_2703(s2703, c2703, in2703_1, in2703_2);
    wire[3:0] s2704, in2704_1, in2704_2;
    wire c2704;
    assign in2704_1 = {s1093[1],s1076[2],pp125[29],s1146[0]};
    assign in2704_2 = {s1094[1],s1077[2],pp126[28],s1147[0]};
    CLA_4 KS_2704(s2704, c2704, in2704_1, in2704_2);
    wire[3:0] s2705, in2705_1, in2705_2;
    wire c2705;
    assign in2705_1 = {s1095[1],s1078[2],pp127[27],s1148[0]};
    assign in2705_2 = {s1096[1],s1079[2],s1070[3],s1149[0]};
    CLA_4 KS_2705(s2705, c2705, in2705_1, in2705_2);
    wire[3:0] s2706, in2706_1, in2706_2;
    wire c2706;
    assign in2706_1 = {s1097[1],s1080[2],s1071[3],s1150[0]};
    assign in2706_2 = {c1098,s1081[2],s1072[3],s1151[0]};
    CLA_4 KS_2706(s2706, c2706, in2706_1, in2706_2);
    wire[3:0] s2707, in2707_1, in2707_2;
    wire c2707;
    assign in2707_1 = {s1099[1],s1082[2],s1073[3],s1152[0]};
    assign in2707_2 = {c1100,s1083[2],s1074[3],s1153[0]};
    CLA_4 KS_2707(s2707, c2707, in2707_1, in2707_2);
    wire[3:0] s2708, in2708_1, in2708_2;
    wire c2708;
    assign in2708_1 = {s1101[1],s1084[2],s1075[3],s1154[0]};
    assign in2708_2 = {c1102,s1085[2],s1076[3],s1155[0]};
    CLA_4 KS_2708(s2708, c2708, in2708_1, in2708_2);
    wire[3:0] s2709, in2709_1, in2709_2;
    wire c2709;
    assign in2709_1 = {s1103[1],s1086[2],s1077[3],s1156[0]};
    assign in2709_2 = {c1104,s1087[2],s1078[3],s1157[0]};
    CLA_4 KS_2709(s2709, c2709, in2709_1, in2709_2);
    wire[3:0] s2710, in2710_1, in2710_2;
    wire c2710;
    assign in2710_1 = {s1105[1],s1088[2],s1079[3],s1158[0]};
    assign in2710_2 = {c1106,s1089[2],s1080[3],s1159[0]};
    CLA_4 KS_2710(s2710, c2710, in2710_1, in2710_2);
    wire[3:0] s2711, in2711_1, in2711_2;
    wire c2711;
    assign in2711_1 = {s1107[1],s1090[2],s1081[3],s1160[0]};
    assign in2711_2 = {c1108,s1091[2],s1082[3],s1161[0]};
    CLA_4 KS_2711(s2711, c2711, in2711_1, in2711_2);
    wire[3:0] s2712, in2712_1, in2712_2;
    wire c2712;
    assign in2712_1 = {s1109[1],s1092[2],s1083[3],s1162[0]};
    assign in2712_2 = {c1110,s1093[2],s1084[3],s1163[0]};
    CLA_4 KS_2712(s2712, c2712, in2712_1, in2712_2);
    wire[3:0] s2713, in2713_1, in2713_2;
    wire c2713;
    assign in2713_1 = {s1111[1],s1094[2],s1085[3],s1164[0]};
    assign in2713_2 = {c1112,s1095[2],s1086[3],s1165[0]};
    CLA_4 KS_2713(s2713, c2713, in2713_1, in2713_2);
    wire[3:0] s2714, in2714_1, in2714_2;
    wire c2714;
    assign in2714_1 = {s1113[1],s1096[2],s1087[3],s1166[0]};
    assign in2714_2 = {c1114,c1097,s1088[3],s1167[0]};
    CLA_4 KS_2714(s2714, c2714, in2714_1, in2714_2);
    wire[3:0] s2715, in2715_1, in2715_2;
    wire c2715;
    assign in2715_1 = {s1115[1],s1099[2],s1089[3],s1168[0]};
    assign in2715_2 = {c1116,c1101,s1090[3],s1169[0]};
    CLA_4 KS_2715(s2715, c2715, in2715_1, in2715_2);
    wire[3:0] s2716, in2716_1, in2716_2;
    wire c2716;
    assign in2716_1 = {s1117[1],s1103[2],s1091[3],s1170[0]};
    assign in2716_2 = {c1118,c1105,s1092[3],s1171[0]};
    CLA_4 KS_2716(s2716, c2716, in2716_1, in2716_2);
    wire[0:0] s2717, in2717_1, in2717_2;
    wire c2717;
    assign in2717_1 = {s1119[1]};
    assign in2717_2 = {c1120};
    Half_Adder KS_2717(s2717, c2717, in2717_1, in2717_2);
    wire[1:0] s2718, in2718_1, in2718_2;
    wire c2718;
    assign in2718_1 = {s1121[1],s1107[2]};
    assign in2718_2 = {c1122,c1109};
    CLA_2 KS_2718(s2718, c2718, in2718_1, in2718_2);
    wire[0:0] s2719, in2719_1, in2719_2;
    wire c2719;
    assign in2719_1 = {s1123[1]};
    assign in2719_2 = {c1124};
    Half_Adder KS_2719(s2719, c2719, in2719_1, in2719_2);
    wire[3:0] s2720, in2720_1, in2720_2;
    wire c2720;
    assign in2720_1 = {s1125[1],s1111[2],s1093[3],s1172[0]};
    assign in2720_2 = {c1126,c1113,s1094[3],s1173[0]};
    CLA_4 KS_2720(s2720, c2720, in2720_1, in2720_2);
    wire[0:0] s2721, in2721_1, in2721_2;
    wire c2721;
    assign in2721_1 = {s1127[1]};
    assign in2721_2 = {c1128};
    Half_Adder KS_2721(s2721, c2721, in2721_1, in2721_2);
    wire[1:0] s2722, in2722_1, in2722_2;
    wire c2722;
    assign in2722_1 = {s1129[1],s1115[2]};
    assign in2722_2 = {c1130,c1117};
    CLA_2 KS_2722(s2722, c2722, in2722_1, in2722_2);
    wire[0:0] s2723, in2723_1, in2723_2;
    wire c2723;
    assign in2723_1 = {s1131[1]};
    assign in2723_2 = {c2621};
    Half_Adder KS_2723(s2723, c2723, in2723_1, in2723_2);
    wire[2:0] s2724, in2724_1, in2724_2;
    wire c2724;
    assign in2724_1 = {c2622,s1119[2],s1095[3]};
    assign in2724_2 = {c2623,c1121,c1096};
    CLA_3 KS_2724(s2724, c2724, in2724_1, in2724_2);
    wire[0:0] s2725, in2725_1, in2725_2;
    wire c2725;
    assign in2725_1 = {c2624};
    assign in2725_2 = {c2625};
    Half_Adder KS_2725(s2725, c2725, in2725_1, in2725_2);
    wire[1:0] s2726, in2726_1, in2726_2;
    wire c2726;
    assign in2726_1 = {c2626,s1123[2]};
    assign in2726_2 = {c2627,c1125};
    CLA_2 KS_2726(s2726, c2726, in2726_1, in2726_2);
    wire[0:0] s2727, in2727_1, in2727_2;
    wire c2727;
    assign in2727_1 = {c2628};
    assign in2727_2 = {c2629};
    Half_Adder KS_2727(s2727, c2727, in2727_1, in2727_2);
    wire[3:0] s2728, in2728_1, in2728_2;
    wire c2728;
    assign in2728_1 = {c2630,s1127[2],s1099[3],s1174[0]};
    assign in2728_2 = {c2631,c1129,c1103,s1175[0]};
    CLA_4 KS_2728(s2728, c2728, in2728_1, in2728_2);
    wire[0:0] s2729, in2729_1, in2729_2;
    wire c2729;
    assign in2729_1 = {c2632};
    assign in2729_2 = {c2633};
    Half_Adder KS_2729(s2729, c2729, in2729_1, in2729_2);
    wire[1:0] s2730, in2730_1, in2730_2;
    wire c2730;
    assign in2730_1 = {c2634,s1131[2]};
    assign in2730_2 = {c2635,s2686[1]};
    CLA_2 KS_2730(s2730, c2730, in2730_1, in2730_2);
    wire[0:0] s2731, in2731_1, in2731_2;
    wire c2731;
    assign in2731_1 = {c2636};
    assign in2731_2 = {c2637};
    Half_Adder KS_2731(s2731, c2731, in2731_1, in2731_2);
    wire[2:0] s2732, in2732_1, in2732_2;
    wire c2732;
    assign in2732_1 = {c2638,s2687[1],s1107[3]};
    assign in2732_2 = {c2639,s2688[1],c1111};
    CLA_3 KS_2732(s2732, c2732, in2732_1, in2732_2);
    wire[0:0] s2733, in2733_1, in2733_2;
    wire c2733;
    assign in2733_1 = {c2640};
    assign in2733_2 = {c2641};
    Half_Adder KS_2733(s2733, c2733, in2733_1, in2733_2);
    wire[1:0] s2734, in2734_1, in2734_2;
    wire c2734;
    assign in2734_1 = {c2642,s2689[1]};
    assign in2734_2 = {c2643,s2690[1]};
    CLA_2 KS_2734(s2734, c2734, in2734_1, in2734_2);
    wire[0:0] s2735, in2735_1, in2735_2;
    wire c2735;
    assign in2735_1 = {c2644};
    assign in2735_2 = {c2645};
    Half_Adder KS_2735(s2735, c2735, in2735_1, in2735_2);
    wire[3:0] s2736, in2736_1, in2736_2;
    wire c2736;
    assign in2736_1 = {c2646,s2691[1],s1115[3],s1176[0]};
    assign in2736_2 = {c2647,s2692[1],c1119,s1177[0]};
    CLA_4 KS_2736(s2736, c2736, in2736_1, in2736_2);
    wire[0:0] s2737, in2737_1, in2737_2;
    wire c2737;
    assign in2737_1 = {c2648};
    assign in2737_2 = {c2649};
    Half_Adder KS_2737(s2737, c2737, in2737_1, in2737_2);
    wire[1:0] s2738, in2738_1, in2738_2;
    wire c2738;
    assign in2738_1 = {c2650,s2693[1]};
    assign in2738_2 = {c2651,s2694[1]};
    CLA_2 KS_2738(s2738, c2738, in2738_1, in2738_2);
    wire[0:0] s2739, in2739_1, in2739_2;
    wire c2739;
    assign in2739_1 = {c2653};
    assign in2739_2 = {c2661};
    Half_Adder KS_2739(s2739, c2739, in2739_1, in2739_2);
    wire[2:0] s2740, in2740_1, in2740_2;
    wire c2740;
    assign in2740_1 = {c2669,s2695[1],s1123[3]};
    assign in2740_2 = {c2677,s2696[1],c1127};
    CLA_3 KS_2740(s2740, c2740, in2740_1, in2740_2);
    wire[0:0] s2741, in2741_1, in2741_2;
    wire c2741;
    assign in2741_1 = {c2685};
    assign in2741_2 = {s2686[0]};
    Half_Adder KS_2741(s2741, c2741, in2741_1, in2741_2);
    wire[1:0] s2742, in2742_1, in2742_2;
    wire c2742;
    assign in2742_1 = {s2687[0],s2697[1]};
    assign in2742_2 = {s2688[0],s2698[1]};
    CLA_2 KS_2742(s2742, c2742, in2742_1, in2742_2);
    wire[0:0] s2743, in2743_1, in2743_2;
    wire c2743;
    assign in2743_1 = {s2689[0]};
    assign in2743_2 = {s2690[0]};
    Half_Adder KS_2743(s2743, c2743, in2743_1, in2743_2);
    wire[3:0] s2744, in2744_1, in2744_2;
    wire c2744;
    assign in2744_1 = {s2691[0],s2699[1],s1131[3],s1178[0]};
    assign in2744_2 = {s2692[0],s2700[1],s2686[2],s1179[0]};
    CLA_4 KS_2744(s2744, c2744, in2744_1, in2744_2);
    wire[0:0] s2745, in2745_1, in2745_2;
    wire c2745;
    assign in2745_1 = {s2693[0]};
    assign in2745_2 = {s2694[0]};
    Half_Adder KS_2745(s2745, c2745, in2745_1, in2745_2);
    wire[1:0] s2746, in2746_1, in2746_2;
    wire c2746;
    assign in2746_1 = {s2695[0],s2701[1]};
    assign in2746_2 = {s2696[0],s2702[1]};
    CLA_2 KS_2746(s2746, c2746, in2746_1, in2746_2);
    wire[0:0] s2747, in2747_1, in2747_2;
    wire c2747;
    assign in2747_1 = {s2697[0]};
    assign in2747_2 = {s2698[0]};
    Half_Adder KS_2747(s2747, c2747, in2747_1, in2747_2);
    wire[2:0] s2748, in2748_1, in2748_2;
    wire c2748;
    assign in2748_1 = {s2699[0],s2703[1],s2687[2]};
    assign in2748_2 = {s2700[0],s2704[1],s2688[2]};
    CLA_3 KS_2748(s2748, c2748, in2748_1, in2748_2);
    wire[0:0] s2749, in2749_1, in2749_2;
    wire c2749;
    assign in2749_1 = {s2701[0]};
    assign in2749_2 = {s2702[0]};
    Half_Adder KS_2749(s2749, c2749, in2749_1, in2749_2);
    wire[1:0] s2750, in2750_1, in2750_2;
    wire c2750;
    assign in2750_1 = {s2704[0],s2705[1]};
    assign in2750_2 = {s2705[0],s2706[1]};
    CLA_2_c KS_2750(s2750, c2750, in2750_1, in2750_2, s2703[0]);
    wire[3:0] s2751, in2751_1, in2751_2;
    wire c2751;
    assign in2751_1 = {pp107[49],pp92[65],pp83[75],pp123[36]};
    assign in2751_2 = {pp108[48],pp93[64],pp84[74],pp124[35]};
    CLA_4 KS_2751(s2751, c2751, in2751_1, in2751_2);
    wire[3:0] s2752, in2752_1, in2752_2;
    wire c2752;
    assign in2752_1 = {pp109[47],pp94[63],pp85[73],pp125[34]};
    assign in2752_2 = {pp110[46],pp95[62],pp86[72],pp126[33]};
    CLA_4 KS_2752(s2752, c2752, in2752_1, in2752_2);
    wire[3:0] s2753, in2753_1, in2753_2;
    wire c2753;
    assign in2753_1 = {pp111[45],pp96[61],pp87[71],pp127[32]};
    assign in2753_2 = {pp112[44],pp97[60],pp88[70],c1132};
    CLA_4 KS_2753(s2753, c2753, in2753_1, in2753_2);
    wire[3:0] s2754, in2754_1, in2754_2;
    wire c2754;
    assign in2754_1 = {pp113[43],pp98[59],pp89[69],c1133};
    assign in2754_2 = {pp114[42],pp99[58],pp90[68],c1134};
    CLA_4 KS_2754(s2754, c2754, in2754_1, in2754_2);
    wire[3:0] s2755, in2755_1, in2755_2;
    wire c2755;
    assign in2755_1 = {pp115[41],pp100[57],pp91[67],c1135};
    assign in2755_2 = {pp116[40],pp101[56],pp92[66],c1136};
    CLA_4 KS_2755(s2755, c2755, in2755_1, in2755_2);
    wire[3:0] s2756, in2756_1, in2756_2;
    wire c2756;
    assign in2756_1 = {pp117[39],pp102[55],pp93[65],c1137};
    assign in2756_2 = {pp118[38],pp103[54],pp94[64],c1138};
    CLA_4 KS_2756(s2756, c2756, in2756_1, in2756_2);
    wire[3:0] s2757, in2757_1, in2757_2;
    wire c2757;
    assign in2757_1 = {pp119[37],pp104[53],pp95[63],c1139};
    assign in2757_2 = {pp120[36],pp105[52],pp96[62],c1140};
    CLA_4 KS_2757(s2757, c2757, in2757_1, in2757_2);
    wire[3:0] s2758, in2758_1, in2758_2;
    wire c2758;
    assign in2758_1 = {pp121[35],pp106[51],pp97[61],c1141};
    assign in2758_2 = {pp122[34],pp107[50],pp98[60],c1142};
    CLA_4 KS_2758(s2758, c2758, in2758_1, in2758_2);
    wire[3:0] s2759, in2759_1, in2759_2;
    wire c2759;
    assign in2759_1 = {pp123[33],pp108[49],pp99[59],c1143};
    assign in2759_2 = {pp124[32],pp109[48],pp100[58],c1144};
    CLA_4 KS_2759(s2759, c2759, in2759_1, in2759_2);
    wire[3:0] s2760, in2760_1, in2760_2;
    wire c2760;
    assign in2760_1 = {pp125[31],pp110[47],pp101[57],c1145};
    assign in2760_2 = {pp126[30],pp111[46],pp102[56],c1146};
    CLA_4 KS_2760(s2760, c2760, in2760_1, in2760_2);
    wire[3:0] s2761, in2761_1, in2761_2;
    wire c2761;
    assign in2761_1 = {pp127[29],pp112[45],pp103[55],c1147};
    assign in2761_2 = {s1132[1],pp113[44],pp104[54],c1148};
    CLA_4 KS_2761(s2761, c2761, in2761_1, in2761_2);
    wire[3:0] s2762, in2762_1, in2762_2;
    wire c2762;
    assign in2762_1 = {s1133[1],pp114[43],pp105[53],c1149};
    assign in2762_2 = {s1134[1],pp115[42],pp106[52],c1150};
    CLA_4 KS_2762(s2762, c2762, in2762_1, in2762_2);
    wire[3:0] s2763, in2763_1, in2763_2;
    wire c2763;
    assign in2763_1 = {s1135[1],pp116[41],pp107[51],c1151};
    assign in2763_2 = {s1136[1],pp117[40],pp108[50],c1152};
    CLA_4 KS_2763(s2763, c2763, in2763_1, in2763_2);
    wire[3:0] s2764, in2764_1, in2764_2;
    wire c2764;
    assign in2764_1 = {s1137[1],pp118[39],pp109[49],c1153};
    assign in2764_2 = {s1138[1],pp119[38],pp110[48],c1157};
    CLA_4 KS_2764(s2764, c2764, in2764_1, in2764_2);
    wire[3:0] s2765, in2765_1, in2765_2;
    wire c2765;
    assign in2765_1 = {s1139[1],pp120[37],pp111[47],c1165};
    assign in2765_2 = {s1140[1],pp121[36],pp112[46],c1173};
    CLA_4 KS_2765(s2765, c2765, in2765_1, in2765_2);
    wire[3:0] s2766, in2766_1, in2766_2;
    wire c2766;
    assign in2766_1 = {s1141[1],pp122[35],pp113[45],c1181};
    assign in2766_2 = {s1142[1],pp123[34],pp114[44],s1186[0]};
    CLA_4 KS_2766(s2766, c2766, in2766_1, in2766_2);
    wire[3:0] s2767, in2767_1, in2767_2;
    wire c2767;
    assign in2767_1 = {s1143[1],pp124[33],pp115[43],s1187[0]};
    assign in2767_2 = {s1144[1],pp125[32],pp116[42],s1188[0]};
    CLA_4 KS_2767(s2767, c2767, in2767_1, in2767_2);
    wire[3:0] s2768, in2768_1, in2768_2;
    wire c2768;
    assign in2768_1 = {s1145[1],pp126[31],pp117[41],s1189[0]};
    assign in2768_2 = {s1146[1],pp127[30],pp118[40],s1190[0]};
    CLA_4 KS_2768(s2768, c2768, in2768_1, in2768_2);
    wire[3:0] s2769, in2769_1, in2769_2;
    wire c2769;
    assign in2769_1 = {s1147[1],s1132[2],pp119[39],s1191[0]};
    assign in2769_2 = {s1148[1],s1133[2],pp120[38],s1192[0]};
    CLA_4 KS_2769(s2769, c2769, in2769_1, in2769_2);
    wire[3:0] s2770, in2770_1, in2770_2;
    wire c2770;
    assign in2770_1 = {s1149[1],s1134[2],pp121[37],s1193[0]};
    assign in2770_2 = {s1150[1],s1135[2],pp122[36],s1194[0]};
    CLA_4 KS_2770(s2770, c2770, in2770_1, in2770_2);
    wire[3:0] s2771, in2771_1, in2771_2;
    wire c2771;
    assign in2771_1 = {s1151[1],s1136[2],pp123[35],s1195[0]};
    assign in2771_2 = {s1152[1],s1137[2],pp124[34],s1196[0]};
    CLA_4 KS_2771(s2771, c2771, in2771_1, in2771_2);
    wire[3:0] s2772, in2772_1, in2772_2;
    wire c2772;
    assign in2772_1 = {s1153[1],s1138[2],pp125[33],s1197[0]};
    assign in2772_2 = {s1154[1],s1139[2],pp126[32],s1198[0]};
    CLA_4 KS_2772(s2772, c2772, in2772_1, in2772_2);
    wire[3:0] s2773, in2773_1, in2773_2;
    wire c2773;
    assign in2773_1 = {s1155[1],s1140[2],pp127[31],s1199[0]};
    assign in2773_2 = {c1156,s1141[2],s1132[3],s1200[0]};
    CLA_4 KS_2773(s2773, c2773, in2773_1, in2773_2);
    wire[3:0] s2774, in2774_1, in2774_2;
    wire c2774;
    assign in2774_1 = {s1157[1],s1142[2],s1133[3],s1201[0]};
    assign in2774_2 = {c1158,s1143[2],s1134[3],s1202[0]};
    CLA_4 KS_2774(s2774, c2774, in2774_1, in2774_2);
    wire[3:0] s2775, in2775_1, in2775_2;
    wire c2775;
    assign in2775_1 = {s1159[1],s1144[2],s1135[3],s1203[0]};
    assign in2775_2 = {c1160,s1145[2],s1136[3],s1204[0]};
    CLA_4 KS_2775(s2775, c2775, in2775_1, in2775_2);
    wire[3:0] s2776, in2776_1, in2776_2;
    wire c2776;
    assign in2776_1 = {s1161[1],s1146[2],s1137[3],s1205[0]};
    assign in2776_2 = {c1162,s1147[2],s1138[3],s1206[0]};
    CLA_4 KS_2776(s2776, c2776, in2776_1, in2776_2);
    wire[3:0] s2777, in2777_1, in2777_2;
    wire c2777;
    assign in2777_1 = {s1163[1],s1148[2],s1139[3],s1207[0]};
    assign in2777_2 = {c1164,s1149[2],s1140[3],s1208[0]};
    CLA_4 KS_2777(s2777, c2777, in2777_1, in2777_2);
    wire[3:0] s2778, in2778_1, in2778_2;
    wire c2778;
    assign in2778_1 = {s1165[1],s1150[2],s1141[3],s1209[0]};
    assign in2778_2 = {c1166,s1151[2],s1142[3],s1210[0]};
    CLA_4 KS_2778(s2778, c2778, in2778_1, in2778_2);
    wire[3:0] s2779, in2779_1, in2779_2;
    wire c2779;
    assign in2779_1 = {s1167[1],s1152[2],s1143[3],s1211[0]};
    assign in2779_2 = {c1168,s1153[2],s1144[3],s1212[0]};
    CLA_4 KS_2779(s2779, c2779, in2779_1, in2779_2);
    wire[3:0] s2780, in2780_1, in2780_2;
    wire c2780;
    assign in2780_1 = {s1169[1],s1154[2],s1145[3],s1213[0]};
    assign in2780_2 = {c1170,c1155,s1146[3],s1214[0]};
    CLA_4 KS_2780(s2780, c2780, in2780_1, in2780_2);
    wire[3:0] s2781, in2781_1, in2781_2;
    wire c2781;
    assign in2781_1 = {s1171[1],s1157[2],s1147[3],s1215[0]};
    assign in2781_2 = {c1172,c1159,s1148[3],s1216[0]};
    CLA_4 KS_2781(s2781, c2781, in2781_1, in2781_2);
    wire[0:0] s2782, in2782_1, in2782_2;
    wire c2782;
    assign in2782_1 = {s1173[1]};
    assign in2782_2 = {c1174};
    Half_Adder KS_2782(s2782, c2782, in2782_1, in2782_2);
    wire[3:0] s2783, in2783_1, in2783_2;
    wire c2783;
    assign in2783_1 = {s1175[1],s1161[2],s1149[3],s1217[0]};
    assign in2783_2 = {c1176,c1163,s1150[3],s1218[0]};
    CLA_4 KS_2783(s2783, c2783, in2783_1, in2783_2);
    wire[0:0] s2784, in2784_1, in2784_2;
    wire c2784;
    assign in2784_1 = {s1177[1]};
    assign in2784_2 = {c1178};
    Half_Adder KS_2784(s2784, c2784, in2784_1, in2784_2);
    wire[1:0] s2785, in2785_1, in2785_2;
    wire c2785;
    assign in2785_1 = {s1179[1],s1165[2]};
    assign in2785_2 = {c1180,c1167};
    CLA_2 KS_2785(s2785, c2785, in2785_1, in2785_2);
    wire[0:0] s2786, in2786_1, in2786_2;
    wire c2786;
    assign in2786_1 = {s1181[1]};
    assign in2786_2 = {c1182};
    Half_Adder KS_2786(s2786, c2786, in2786_1, in2786_2);
    wire[2:0] s2787, in2787_1, in2787_2;
    wire c2787;
    assign in2787_1 = {s1183[1],s1169[2],s1151[3]};
    assign in2787_2 = {c1184,c1171,s1152[3]};
    CLA_3 KS_2787(s2787, c2787, in2787_1, in2787_2);
    wire[0:0] s2788, in2788_1, in2788_2;
    wire c2788;
    assign in2788_1 = {s1185[1]};
    assign in2788_2 = {c2686};
    Half_Adder KS_2788(s2788, c2788, in2788_1, in2788_2);
    wire[1:0] s2789, in2789_1, in2789_2;
    wire c2789;
    assign in2789_1 = {c2687,s1173[2]};
    assign in2789_2 = {c2688,c1175};
    CLA_2 KS_2789(s2789, c2789, in2789_1, in2789_2);
    wire[0:0] s2790, in2790_1, in2790_2;
    wire c2790;
    assign in2790_1 = {c2689};
    assign in2790_2 = {c2690};
    Half_Adder KS_2790(s2790, c2790, in2790_1, in2790_2);
    wire[3:0] s2791, in2791_1, in2791_2;
    wire c2791;
    assign in2791_1 = {c2691,s1177[2],s1153[3],s1219[0]};
    assign in2791_2 = {c2692,c1179,c1154,s1220[0]};
    CLA_4 KS_2791(s2791, c2791, in2791_1, in2791_2);
    wire[0:0] s2792, in2792_1, in2792_2;
    wire c2792;
    assign in2792_1 = {c2693};
    assign in2792_2 = {c2694};
    Half_Adder KS_2792(s2792, c2792, in2792_1, in2792_2);
    wire[1:0] s2793, in2793_1, in2793_2;
    wire c2793;
    assign in2793_1 = {c2695,s1181[2]};
    assign in2793_2 = {c2696,c1183};
    CLA_2 KS_2793(s2793, c2793, in2793_1, in2793_2);
    wire[0:0] s2794, in2794_1, in2794_2;
    wire c2794;
    assign in2794_1 = {c2697};
    assign in2794_2 = {c2698};
    Half_Adder KS_2794(s2794, c2794, in2794_1, in2794_2);
    wire[2:0] s2795, in2795_1, in2795_2;
    wire c2795;
    assign in2795_1 = {c2699,s1185[2],s1157[3]};
    assign in2795_2 = {c2700,s2751[1],c1161};
    CLA_3 KS_2795(s2795, c2795, in2795_1, in2795_2);
    wire[0:0] s2796, in2796_1, in2796_2;
    wire c2796;
    assign in2796_1 = {c2701};
    assign in2796_2 = {c2702};
    Half_Adder KS_2796(s2796, c2796, in2796_1, in2796_2);
    wire[1:0] s2797, in2797_1, in2797_2;
    wire c2797;
    assign in2797_1 = {c2703,s2752[1]};
    assign in2797_2 = {c2704,s2753[1]};
    CLA_2 KS_2797(s2797, c2797, in2797_1, in2797_2);
    wire[0:0] s2798, in2798_1, in2798_2;
    wire c2798;
    assign in2798_1 = {c2705};
    assign in2798_2 = {c2706};
    Half_Adder KS_2798(s2798, c2798, in2798_1, in2798_2);
    wire[3:0] s2799, in2799_1, in2799_2;
    wire c2799;
    assign in2799_1 = {c2707,s2754[1],s1165[3],s1221[0]};
    assign in2799_2 = {c2708,s2755[1],c1169,s1222[0]};
    CLA_4 KS_2799(s2799, c2799, in2799_1, in2799_2);
    wire[0:0] s2800, in2800_1, in2800_2;
    wire c2800;
    assign in2800_1 = {c2709};
    assign in2800_2 = {c2710};
    Half_Adder KS_2800(s2800, c2800, in2800_1, in2800_2);
    wire[1:0] s2801, in2801_1, in2801_2;
    wire c2801;
    assign in2801_1 = {c2711,s2756[1]};
    assign in2801_2 = {c2712,s2757[1]};
    CLA_2 KS_2801(s2801, c2801, in2801_1, in2801_2);
    wire[0:0] s2802, in2802_1, in2802_2;
    wire c2802;
    assign in2802_1 = {c2713};
    assign in2802_2 = {c2714};
    Half_Adder KS_2802(s2802, c2802, in2802_1, in2802_2);
    wire[2:0] s2803, in2803_1, in2803_2;
    wire c2803;
    assign in2803_1 = {c2715,s2758[1],s1173[3]};
    assign in2803_2 = {c2716,s2759[1],c1177};
    CLA_3 KS_2803(s2803, c2803, in2803_1, in2803_2);
    wire[0:0] s2804, in2804_1, in2804_2;
    wire c2804;
    assign in2804_1 = {c2720};
    assign in2804_2 = {c2728};
    Half_Adder KS_2804(s2804, c2804, in2804_1, in2804_2);
    wire[1:0] s2805, in2805_1, in2805_2;
    wire c2805;
    assign in2805_1 = {c2736,s2760[1]};
    assign in2805_2 = {c2744,s2761[1]};
    CLA_2 KS_2805(s2805, c2805, in2805_1, in2805_2);
    wire[0:0] s2806, in2806_1, in2806_2;
    wire c2806;
    assign in2806_1 = {s2751[0]};
    assign in2806_2 = {s2752[0]};
    Half_Adder KS_2806(s2806, c2806, in2806_1, in2806_2);
    wire[3:0] s2807, in2807_1, in2807_2;
    wire c2807;
    assign in2807_1 = {s2753[0],s2762[1],s1181[3],s1223[0]};
    assign in2807_2 = {s2754[0],s2763[1],c1185,s1224[0]};
    CLA_4 KS_2807(s2807, c2807, in2807_1, in2807_2);
    wire[0:0] s2808, in2808_1, in2808_2;
    wire c2808;
    assign in2808_1 = {s2755[0]};
    assign in2808_2 = {s2756[0]};
    Half_Adder KS_2808(s2808, c2808, in2808_1, in2808_2);
    wire[1:0] s2809, in2809_1, in2809_2;
    wire c2809;
    assign in2809_1 = {s2757[0],s2764[1]};
    assign in2809_2 = {s2758[0],s2765[1]};
    CLA_2 KS_2809(s2809, c2809, in2809_1, in2809_2);
    wire[0:0] s2810, in2810_1, in2810_2;
    wire c2810;
    assign in2810_1 = {s2759[0]};
    assign in2810_2 = {s2760[0]};
    Half_Adder KS_2810(s2810, c2810, in2810_1, in2810_2);
    wire[2:0] s2811, in2811_1, in2811_2;
    wire c2811;
    assign in2811_1 = {s2761[0],s2766[1],s2751[2]};
    assign in2811_2 = {s2762[0],s2767[1],s2752[2]};
    CLA_3 KS_2811(s2811, c2811, in2811_1, in2811_2);
    wire[0:0] s2812, in2812_1, in2812_2;
    wire c2812;
    assign in2812_1 = {s2763[0]};
    assign in2812_2 = {s2764[0]};
    Half_Adder KS_2812(s2812, c2812, in2812_1, in2812_2);
    wire[1:0] s2813, in2813_1, in2813_2;
    wire c2813;
    assign in2813_1 = {s2765[0],s2768[1]};
    assign in2813_2 = {s2766[0],s2769[1]};
    CLA_2 KS_2813(s2813, c2813, in2813_1, in2813_2);
    wire[0:0] s2814, in2814_1, in2814_2;
    wire c2814;
    assign in2814_1 = {s2768[0]};
    assign in2814_2 = {s2769[0]};
    Full_Adder KS_2814(s2814, c2814, in2814_1, in2814_2, s2767[0]);
    wire[3:0] s2815, in2815_1, in2815_2;
    wire c2815;
    assign in2815_1 = {pp97[63],pp84[77],pp77[85],pp109[54]};
    assign in2815_2 = {pp98[62],pp85[76],pp78[84],pp110[53]};
    CLA_4 KS_2815(s2815, c2815, in2815_1, in2815_2);
    wire[3:0] s2816, in2816_1, in2816_2;
    wire c2816;
    assign in2816_1 = {pp99[61],pp86[75],pp79[83],pp111[52]};
    assign in2816_2 = {pp100[60],pp87[74],pp80[82],pp112[51]};
    CLA_4 KS_2816(s2816, c2816, in2816_1, in2816_2);
    wire[3:0] s2817, in2817_1, in2817_2;
    wire c2817;
    assign in2817_1 = {pp101[59],pp88[73],pp81[81],pp113[50]};
    assign in2817_2 = {pp102[58],pp89[72],pp82[80],pp114[49]};
    CLA_4 KS_2817(s2817, c2817, in2817_1, in2817_2);
    wire[3:0] s2818, in2818_1, in2818_2;
    wire c2818;
    assign in2818_1 = {pp103[57],pp90[71],pp83[79],pp115[48]};
    assign in2818_2 = {pp104[56],pp91[70],pp84[78],pp116[47]};
    CLA_4 KS_2818(s2818, c2818, in2818_1, in2818_2);
    wire[3:0] s2819, in2819_1, in2819_2;
    wire c2819;
    assign in2819_1 = {pp105[55],pp92[69],pp85[77],pp117[46]};
    assign in2819_2 = {pp106[54],pp93[68],pp86[76],pp118[45]};
    CLA_4 KS_2819(s2819, c2819, in2819_1, in2819_2);
    wire[3:0] s2820, in2820_1, in2820_2;
    wire c2820;
    assign in2820_1 = {pp107[53],pp94[67],pp87[75],pp119[44]};
    assign in2820_2 = {pp108[52],pp95[66],pp88[74],pp120[43]};
    CLA_4 KS_2820(s2820, c2820, in2820_1, in2820_2);
    wire[3:0] s2821, in2821_1, in2821_2;
    wire c2821;
    assign in2821_1 = {pp109[51],pp96[65],pp89[73],pp121[42]};
    assign in2821_2 = {pp110[50],pp97[64],pp90[72],pp122[41]};
    CLA_4 KS_2821(s2821, c2821, in2821_1, in2821_2);
    wire[3:0] s2822, in2822_1, in2822_2;
    wire c2822;
    assign in2822_1 = {pp111[49],pp98[63],pp91[71],pp123[40]};
    assign in2822_2 = {pp112[48],pp99[62],pp92[70],pp124[39]};
    CLA_4 KS_2822(s2822, c2822, in2822_1, in2822_2);
    wire[3:0] s2823, in2823_1, in2823_2;
    wire c2823;
    assign in2823_1 = {pp113[47],pp100[61],pp93[69],pp125[38]};
    assign in2823_2 = {pp114[46],pp101[60],pp94[68],pp126[37]};
    CLA_4 KS_2823(s2823, c2823, in2823_1, in2823_2);
    wire[3:0] s2824, in2824_1, in2824_2;
    wire c2824;
    assign in2824_1 = {pp115[45],pp102[59],pp95[67],pp127[36]};
    assign in2824_2 = {pp116[44],pp103[58],pp96[66],c1186};
    CLA_4 KS_2824(s2824, c2824, in2824_1, in2824_2);
    wire[3:0] s2825, in2825_1, in2825_2;
    wire c2825;
    assign in2825_1 = {pp117[43],pp104[57],pp97[65],c1187};
    assign in2825_2 = {pp118[42],pp105[56],pp98[64],c1188};
    CLA_4 KS_2825(s2825, c2825, in2825_1, in2825_2);
    wire[3:0] s2826, in2826_1, in2826_2;
    wire c2826;
    assign in2826_1 = {pp119[41],pp106[55],pp99[63],c1189};
    assign in2826_2 = {pp120[40],pp107[54],pp100[62],c1190};
    CLA_4 KS_2826(s2826, c2826, in2826_1, in2826_2);
    wire[3:0] s2827, in2827_1, in2827_2;
    wire c2827;
    assign in2827_1 = {pp121[39],pp108[53],pp101[61],c1191};
    assign in2827_2 = {pp122[38],pp109[52],pp102[60],c1192};
    CLA_4 KS_2827(s2827, c2827, in2827_1, in2827_2);
    wire[3:0] s2828, in2828_1, in2828_2;
    wire c2828;
    assign in2828_1 = {pp123[37],pp110[51],pp103[59],c1193};
    assign in2828_2 = {pp124[36],pp111[50],pp104[58],c1194};
    CLA_4 KS_2828(s2828, c2828, in2828_1, in2828_2);
    wire[3:0] s2829, in2829_1, in2829_2;
    wire c2829;
    assign in2829_1 = {pp125[35],pp112[49],pp105[57],c1195};
    assign in2829_2 = {pp126[34],pp113[48],pp106[56],c1196};
    CLA_4 KS_2829(s2829, c2829, in2829_1, in2829_2);
    wire[3:0] s2830, in2830_1, in2830_2;
    wire c2830;
    assign in2830_1 = {pp127[33],pp114[47],pp107[55],c1197};
    assign in2830_2 = {s1186[1],pp115[46],pp108[54],c1198};
    CLA_4 KS_2830(s2830, c2830, in2830_1, in2830_2);
    wire[3:0] s2831, in2831_1, in2831_2;
    wire c2831;
    assign in2831_1 = {s1187[1],pp116[45],pp109[53],c1199};
    assign in2831_2 = {s1188[1],pp117[44],pp110[52],c1200};
    CLA_4 KS_2831(s2831, c2831, in2831_1, in2831_2);
    wire[3:0] s2832, in2832_1, in2832_2;
    wire c2832;
    assign in2832_1 = {s1189[1],pp118[43],pp111[51],c1201};
    assign in2832_2 = {s1190[1],pp119[42],pp112[50],c1202};
    CLA_4 KS_2832(s2832, c2832, in2832_1, in2832_2);
    wire[3:0] s2833, in2833_1, in2833_2;
    wire c2833;
    assign in2833_1 = {s1191[1],pp120[41],pp113[49],c1203};
    assign in2833_2 = {s1192[1],pp121[40],pp114[48],c1207};
    CLA_4 KS_2833(s2833, c2833, in2833_1, in2833_2);
    wire[3:0] s2834, in2834_1, in2834_2;
    wire c2834;
    assign in2834_1 = {s1193[1],pp122[39],pp115[47],c1215};
    assign in2834_2 = {s1194[1],pp123[38],pp116[46],c1223};
    CLA_4 KS_2834(s2834, c2834, in2834_1, in2834_2);
    wire[3:0] s2835, in2835_1, in2835_2;
    wire c2835;
    assign in2835_1 = {s1195[1],pp124[37],pp117[45],s1231[0]};
    assign in2835_2 = {s1196[1],pp125[36],pp118[44],s1232[0]};
    CLA_4 KS_2835(s2835, c2835, in2835_1, in2835_2);
    wire[3:0] s2836, in2836_1, in2836_2;
    wire c2836;
    assign in2836_1 = {s1197[1],pp126[35],pp119[43],s1233[0]};
    assign in2836_2 = {s1198[1],pp127[34],pp120[42],s1234[0]};
    CLA_4 KS_2836(s2836, c2836, in2836_1, in2836_2);
    wire[3:0] s2837, in2837_1, in2837_2;
    wire c2837;
    assign in2837_1 = {s1199[1],s1186[2],pp121[41],s1235[0]};
    assign in2837_2 = {s1200[1],s1187[2],pp122[40],s1236[0]};
    CLA_4 KS_2837(s2837, c2837, in2837_1, in2837_2);
    wire[3:0] s2838, in2838_1, in2838_2;
    wire c2838;
    assign in2838_1 = {s1201[1],s1188[2],pp123[39],s1237[0]};
    assign in2838_2 = {s1202[1],s1189[2],pp124[38],s1238[0]};
    CLA_4 KS_2838(s2838, c2838, in2838_1, in2838_2);
    wire[3:0] s2839, in2839_1, in2839_2;
    wire c2839;
    assign in2839_1 = {s1203[1],s1190[2],pp125[37],s1239[0]};
    assign in2839_2 = {s1204[1],s1191[2],pp126[36],s1240[0]};
    CLA_4 KS_2839(s2839, c2839, in2839_1, in2839_2);
    wire[3:0] s2840, in2840_1, in2840_2;
    wire c2840;
    assign in2840_1 = {s1205[1],s1192[2],pp127[35],s1241[0]};
    assign in2840_2 = {c1206,s1193[2],s1186[3],s1242[0]};
    CLA_4 KS_2840(s2840, c2840, in2840_1, in2840_2);
    wire[3:0] s2841, in2841_1, in2841_2;
    wire c2841;
    assign in2841_1 = {s1207[1],s1194[2],s1187[3],s1243[0]};
    assign in2841_2 = {c1208,s1195[2],s1188[3],s1244[0]};
    CLA_4 KS_2841(s2841, c2841, in2841_1, in2841_2);
    wire[3:0] s2842, in2842_1, in2842_2;
    wire c2842;
    assign in2842_1 = {s1209[1],s1196[2],s1189[3],s1245[0]};
    assign in2842_2 = {c1210,s1197[2],s1190[3],s1246[0]};
    CLA_4 KS_2842(s2842, c2842, in2842_1, in2842_2);
    wire[3:0] s2843, in2843_1, in2843_2;
    wire c2843;
    assign in2843_1 = {s1211[1],s1198[2],s1191[3],s1247[0]};
    assign in2843_2 = {c1212,s1199[2],s1192[3],s1248[0]};
    CLA_4 KS_2843(s2843, c2843, in2843_1, in2843_2);
    wire[3:0] s2844, in2844_1, in2844_2;
    wire c2844;
    assign in2844_1 = {s1213[1],s1200[2],s1193[3],s1249[0]};
    assign in2844_2 = {c1214,s1201[2],s1194[3],s1250[0]};
    CLA_4 KS_2844(s2844, c2844, in2844_1, in2844_2);
    wire[3:0] s2845, in2845_1, in2845_2;
    wire c2845;
    assign in2845_1 = {s1215[1],s1202[2],s1195[3],s1251[0]};
    assign in2845_2 = {c1216,s1203[2],s1196[3],s1252[0]};
    CLA_4 KS_2845(s2845, c2845, in2845_1, in2845_2);
    wire[3:0] s2846, in2846_1, in2846_2;
    wire c2846;
    assign in2846_1 = {s1217[1],s1204[2],s1197[3],s1253[0]};
    assign in2846_2 = {c1218,c1205,s1198[3],s1254[0]};
    CLA_4 KS_2846(s2846, c2846, in2846_1, in2846_2);
    wire[0:0] s2847, in2847_1, in2847_2;
    wire c2847;
    assign in2847_1 = {s1219[1]};
    assign in2847_2 = {c1220};
    Half_Adder KS_2847(s2847, c2847, in2847_1, in2847_2);
    wire[1:0] s2848, in2848_1, in2848_2;
    wire c2848;
    assign in2848_1 = {s1221[1],s1207[2]};
    assign in2848_2 = {c1222,c1209};
    CLA_2 KS_2848(s2848, c2848, in2848_1, in2848_2);
    wire[0:0] s2849, in2849_1, in2849_2;
    wire c2849;
    assign in2849_1 = {s1223[1]};
    assign in2849_2 = {c1224};
    Half_Adder KS_2849(s2849, c2849, in2849_1, in2849_2);
    wire[2:0] s2850, in2850_1, in2850_2;
    wire c2850;
    assign in2850_1 = {s1225[1],s1211[2],s1199[3]};
    assign in2850_2 = {c1226,c1213,s1200[3]};
    CLA_3 KS_2850(s2850, c2850, in2850_1, in2850_2);
    wire[0:0] s2851, in2851_1, in2851_2;
    wire c2851;
    assign in2851_1 = {s1227[1]};
    assign in2851_2 = {c1228};
    Half_Adder KS_2851(s2851, c2851, in2851_1, in2851_2);
    wire[1:0] s2852, in2852_1, in2852_2;
    wire c2852;
    assign in2852_1 = {s1229[1],s1215[2]};
    assign in2852_2 = {c1230,c1217};
    CLA_2 KS_2852(s2852, c2852, in2852_1, in2852_2);
    wire[0:0] s2853, in2853_1, in2853_2;
    wire c2853;
    assign in2853_1 = {c2751};
    assign in2853_2 = {c2752};
    Half_Adder KS_2853(s2853, c2853, in2853_1, in2853_2);
    wire[3:0] s2854, in2854_1, in2854_2;
    wire c2854;
    assign in2854_1 = {c2753,s1219[2],s1201[3],s1255[0]};
    assign in2854_2 = {c2754,c1221,s1202[3],s1256[0]};
    CLA_4 KS_2854(s2854, c2854, in2854_1, in2854_2);
    wire[0:0] s2855, in2855_1, in2855_2;
    wire c2855;
    assign in2855_1 = {c2755};
    assign in2855_2 = {c2756};
    Half_Adder KS_2855(s2855, c2855, in2855_1, in2855_2);
    wire[1:0] s2856, in2856_1, in2856_2;
    wire c2856;
    assign in2856_1 = {c2757,s1223[2]};
    assign in2856_2 = {c2758,c1225};
    CLA_2 KS_2856(s2856, c2856, in2856_1, in2856_2);
    wire[0:0] s2857, in2857_1, in2857_2;
    wire c2857;
    assign in2857_1 = {c2759};
    assign in2857_2 = {c2760};
    Half_Adder KS_2857(s2857, c2857, in2857_1, in2857_2);
    wire[2:0] s2858, in2858_1, in2858_2;
    wire c2858;
    assign in2858_1 = {c2761,s1227[2],s1203[3]};
    assign in2858_2 = {c2762,c1229,c1204};
    CLA_3 KS_2858(s2858, c2858, in2858_1, in2858_2);
    wire[0:0] s2859, in2859_1, in2859_2;
    wire c2859;
    assign in2859_1 = {c2763};
    assign in2859_2 = {c2764};
    Half_Adder KS_2859(s2859, c2859, in2859_1, in2859_2);
    wire[1:0] s2860, in2860_1, in2860_2;
    wire c2860;
    assign in2860_1 = {c2765,s2815[1]};
    assign in2860_2 = {c2766,s2816[1]};
    CLA_2 KS_2860(s2860, c2860, in2860_1, in2860_2);
    wire[0:0] s2861, in2861_1, in2861_2;
    wire c2861;
    assign in2861_1 = {c2767};
    assign in2861_2 = {c2768};
    Half_Adder KS_2861(s2861, c2861, in2861_1, in2861_2);
    wire[3:0] s2862, in2862_1, in2862_2;
    wire c2862;
    assign in2862_1 = {c2769,s2817[1],s1207[3],s1257[0]};
    assign in2862_2 = {c2770,s2818[1],c1211,s1258[0]};
    CLA_4 KS_2862(s2862, c2862, in2862_1, in2862_2);
    wire[0:0] s2863, in2863_1, in2863_2;
    wire c2863;
    assign in2863_1 = {c2771};
    assign in2863_2 = {c2772};
    Half_Adder KS_2863(s2863, c2863, in2863_1, in2863_2);
    wire[1:0] s2864, in2864_1, in2864_2;
    wire c2864;
    assign in2864_1 = {c2773,s2819[1]};
    assign in2864_2 = {c2774,s2820[1]};
    CLA_2 KS_2864(s2864, c2864, in2864_1, in2864_2);
    wire[0:0] s2865, in2865_1, in2865_2;
    wire c2865;
    assign in2865_1 = {c2775};
    assign in2865_2 = {c2776};
    Half_Adder KS_2865(s2865, c2865, in2865_1, in2865_2);
    wire[2:0] s2866, in2866_1, in2866_2;
    wire c2866;
    assign in2866_1 = {c2777,s2821[1],s1215[3]};
    assign in2866_2 = {c2778,s2822[1],c1219};
    CLA_3 KS_2866(s2866, c2866, in2866_1, in2866_2);
    wire[0:0] s2867, in2867_1, in2867_2;
    wire c2867;
    assign in2867_1 = {c2779};
    assign in2867_2 = {c2780};
    Half_Adder KS_2867(s2867, c2867, in2867_1, in2867_2);
    wire[1:0] s2868, in2868_1, in2868_2;
    wire c2868;
    assign in2868_1 = {c2781,s2823[1]};
    assign in2868_2 = {c2783,s2824[1]};
    CLA_2 KS_2868(s2868, c2868, in2868_1, in2868_2);
    wire[0:0] s2869, in2869_1, in2869_2;
    wire c2869;
    assign in2869_1 = {c2791};
    assign in2869_2 = {c2799};
    Half_Adder KS_2869(s2869, c2869, in2869_1, in2869_2);
    wire[3:0] s2870, in2870_1, in2870_2;
    wire c2870;
    assign in2870_1 = {c2807,s2825[1],s1223[3],s1259[0]};
    assign in2870_2 = {s2815[0],s2826[1],c1227,s1260[0]};
    CLA_4 KS_2870(s2870, c2870, in2870_1, in2870_2);
    wire[0:0] s2871, in2871_1, in2871_2;
    wire c2871;
    assign in2871_1 = {s2816[0]};
    assign in2871_2 = {s2817[0]};
    Half_Adder KS_2871(s2871, c2871, in2871_1, in2871_2);
    wire[1:0] s2872, in2872_1, in2872_2;
    wire c2872;
    assign in2872_1 = {s2818[0],s2827[1]};
    assign in2872_2 = {s2819[0],s2828[1]};
    CLA_2 KS_2872(s2872, c2872, in2872_1, in2872_2);
    wire[0:0] s2873, in2873_1, in2873_2;
    wire c2873;
    assign in2873_1 = {s2820[0]};
    assign in2873_2 = {s2821[0]};
    Half_Adder KS_2873(s2873, c2873, in2873_1, in2873_2);
    wire[2:0] s2874, in2874_1, in2874_2;
    wire c2874;
    assign in2874_1 = {s2822[0],s2829[1],s2815[2]};
    assign in2874_2 = {s2823[0],s2830[1],s2816[2]};
    CLA_3 KS_2874(s2874, c2874, in2874_1, in2874_2);
    wire[0:0] s2875, in2875_1, in2875_2;
    wire c2875;
    assign in2875_1 = {s2824[0]};
    assign in2875_2 = {s2825[0]};
    Half_Adder KS_2875(s2875, c2875, in2875_1, in2875_2);
    wire[1:0] s2876, in2876_1, in2876_2;
    wire c2876;
    assign in2876_1 = {s2826[0],s2831[1]};
    assign in2876_2 = {s2827[0],s2832[1]};
    CLA_2 KS_2876(s2876, c2876, in2876_1, in2876_2);
    wire[0:0] s2877, in2877_1, in2877_2;
    wire c2877;
    assign in2877_1 = {s2828[0]};
    assign in2877_2 = {s2829[0]};
    Half_Adder KS_2877(s2877, c2877, in2877_1, in2877_2);
    wire[3:0] s2878, in2878_1, in2878_2;
    wire c2878;
    assign in2878_1 = {s2830[0],s2833[1],s2817[2],s1261[0]};
    assign in2878_2 = {s2831[0],s2834[1],s2818[2],s1262[0]};
    CLA_4 KS_2878(s2878, c2878, in2878_1, in2878_2);
    wire[0:0] s2879, in2879_1, in2879_2;
    wire c2879;
    assign in2879_1 = {s2833[0]};
    assign in2879_2 = {s2834[0]};
    Full_Adder KS_2879(s2879, c2879, in2879_1, in2879_2, s2832[0]);
    wire[3:0] s2880, in2880_1, in2880_2;
    wire c2880;
    assign in2880_1 = {pp89[75],pp78[87],pp73[93],pp97[70]};
    assign in2880_2 = {pp90[74],pp79[86],pp74[92],pp98[69]};
    CLA_4 KS_2880(s2880, c2880, in2880_1, in2880_2);
    wire[3:0] s2881, in2881_1, in2881_2;
    wire c2881;
    assign in2881_1 = {pp91[73],pp80[85],pp75[91],pp99[68]};
    assign in2881_2 = {pp92[72],pp81[84],pp76[90],pp100[67]};
    CLA_4 KS_2881(s2881, c2881, in2881_1, in2881_2);
    wire[3:0] s2882, in2882_1, in2882_2;
    wire c2882;
    assign in2882_1 = {pp93[71],pp82[83],pp77[89],pp101[66]};
    assign in2882_2 = {pp94[70],pp83[82],pp78[88],pp102[65]};
    CLA_4 KS_2882(s2882, c2882, in2882_1, in2882_2);
    wire[3:0] s2883, in2883_1, in2883_2;
    wire c2883;
    assign in2883_1 = {pp95[69],pp84[81],pp79[87],pp103[64]};
    assign in2883_2 = {pp96[68],pp85[80],pp80[86],pp104[63]};
    CLA_4 KS_2883(s2883, c2883, in2883_1, in2883_2);
    wire[3:0] s2884, in2884_1, in2884_2;
    wire c2884;
    assign in2884_1 = {pp97[67],pp86[79],pp81[85],pp105[62]};
    assign in2884_2 = {pp98[66],pp87[78],pp82[84],pp106[61]};
    CLA_4 KS_2884(s2884, c2884, in2884_1, in2884_2);
    wire[3:0] s2885, in2885_1, in2885_2;
    wire c2885;
    assign in2885_1 = {pp99[65],pp88[77],pp83[83],pp107[60]};
    assign in2885_2 = {pp100[64],pp89[76],pp84[82],pp108[59]};
    CLA_4 KS_2885(s2885, c2885, in2885_1, in2885_2);
    wire[3:0] s2886, in2886_1, in2886_2;
    wire c2886;
    assign in2886_1 = {pp101[63],pp90[75],pp85[81],pp109[58]};
    assign in2886_2 = {pp102[62],pp91[74],pp86[80],pp110[57]};
    CLA_4 KS_2886(s2886, c2886, in2886_1, in2886_2);
    wire[3:0] s2887, in2887_1, in2887_2;
    wire c2887;
    assign in2887_1 = {pp103[61],pp92[73],pp87[79],pp111[56]};
    assign in2887_2 = {pp104[60],pp93[72],pp88[78],pp112[55]};
    CLA_4 KS_2887(s2887, c2887, in2887_1, in2887_2);
    wire[3:0] s2888, in2888_1, in2888_2;
    wire c2888;
    assign in2888_1 = {pp105[59],pp94[71],pp89[77],pp113[54]};
    assign in2888_2 = {pp106[58],pp95[70],pp90[76],pp114[53]};
    CLA_4 KS_2888(s2888, c2888, in2888_1, in2888_2);
    wire[3:0] s2889, in2889_1, in2889_2;
    wire c2889;
    assign in2889_1 = {pp107[57],pp96[69],pp91[75],pp115[52]};
    assign in2889_2 = {pp108[56],pp97[68],pp92[74],pp116[51]};
    CLA_4 KS_2889(s2889, c2889, in2889_1, in2889_2);
    wire[3:0] s2890, in2890_1, in2890_2;
    wire c2890;
    assign in2890_1 = {pp109[55],pp98[67],pp93[73],pp117[50]};
    assign in2890_2 = {pp110[54],pp99[66],pp94[72],pp118[49]};
    CLA_4 KS_2890(s2890, c2890, in2890_1, in2890_2);
    wire[3:0] s2891, in2891_1, in2891_2;
    wire c2891;
    assign in2891_1 = {pp111[53],pp100[65],pp95[71],pp119[48]};
    assign in2891_2 = {pp112[52],pp101[64],pp96[70],pp120[47]};
    CLA_4 KS_2891(s2891, c2891, in2891_1, in2891_2);
    wire[3:0] s2892, in2892_1, in2892_2;
    wire c2892;
    assign in2892_1 = {pp113[51],pp102[63],pp97[69],pp121[46]};
    assign in2892_2 = {pp114[50],pp103[62],pp98[68],pp122[45]};
    CLA_4 KS_2892(s2892, c2892, in2892_1, in2892_2);
    wire[3:0] s2893, in2893_1, in2893_2;
    wire c2893;
    assign in2893_1 = {pp115[49],pp104[61],pp99[67],pp123[44]};
    assign in2893_2 = {pp116[48],pp105[60],pp100[66],pp124[43]};
    CLA_4 KS_2893(s2893, c2893, in2893_1, in2893_2);
    wire[3:0] s2894, in2894_1, in2894_2;
    wire c2894;
    assign in2894_1 = {pp117[47],pp106[59],pp101[65],pp125[42]};
    assign in2894_2 = {pp118[46],pp107[58],pp102[64],pp126[41]};
    CLA_4 KS_2894(s2894, c2894, in2894_1, in2894_2);
    wire[3:0] s2895, in2895_1, in2895_2;
    wire c2895;
    assign in2895_1 = {pp119[45],pp108[57],pp103[63],pp127[40]};
    assign in2895_2 = {pp120[44],pp109[56],pp104[62],c1231};
    CLA_4 KS_2895(s2895, c2895, in2895_1, in2895_2);
    wire[3:0] s2896, in2896_1, in2896_2;
    wire c2896;
    assign in2896_1 = {pp121[43],pp110[55],pp105[61],c1232};
    assign in2896_2 = {pp122[42],pp111[54],pp106[60],c1233};
    CLA_4 KS_2896(s2896, c2896, in2896_1, in2896_2);
    wire[3:0] s2897, in2897_1, in2897_2;
    wire c2897;
    assign in2897_1 = {pp123[41],pp112[53],pp107[59],c1234};
    assign in2897_2 = {pp124[40],pp113[52],pp108[58],c1235};
    CLA_4 KS_2897(s2897, c2897, in2897_1, in2897_2);
    wire[3:0] s2898, in2898_1, in2898_2;
    wire c2898;
    assign in2898_1 = {pp125[39],pp114[51],pp109[57],c1236};
    assign in2898_2 = {pp126[38],pp115[50],pp110[56],c1237};
    CLA_4 KS_2898(s2898, c2898, in2898_1, in2898_2);
    wire[3:0] s2899, in2899_1, in2899_2;
    wire c2899;
    assign in2899_1 = {pp127[37],pp116[49],pp111[55],c1238};
    assign in2899_2 = {s1231[1],pp117[48],pp112[54],c1239};
    CLA_4 KS_2899(s2899, c2899, in2899_1, in2899_2);
    wire[3:0] s2900, in2900_1, in2900_2;
    wire c2900;
    assign in2900_1 = {s1232[1],pp118[47],pp113[53],c1240};
    assign in2900_2 = {s1233[1],pp119[46],pp114[52],c1241};
    CLA_4 KS_2900(s2900, c2900, in2900_1, in2900_2);
    wire[3:0] s2901, in2901_1, in2901_2;
    wire c2901;
    assign in2901_1 = {s1234[1],pp120[45],pp115[51],c1242};
    assign in2901_2 = {s1235[1],pp121[44],pp116[50],c1243};
    CLA_4 KS_2901(s2901, c2901, in2901_1, in2901_2);
    wire[3:0] s2902, in2902_1, in2902_2;
    wire c2902;
    assign in2902_1 = {s1236[1],pp122[43],pp117[49],c1244};
    assign in2902_2 = {s1237[1],pp123[42],pp118[48],c1248};
    CLA_4 KS_2902(s2902, c2902, in2902_1, in2902_2);
    wire[3:0] s2903, in2903_1, in2903_2;
    wire c2903;
    assign in2903_1 = {s1238[1],pp124[41],pp119[47],c1256};
    assign in2903_2 = {s1239[1],pp125[40],pp120[46],c1264};
    CLA_4 KS_2903(s2903, c2903, in2903_1, in2903_2);
    wire[3:0] s2904, in2904_1, in2904_2;
    wire c2904;
    assign in2904_1 = {s1240[1],pp126[39],pp121[45],s1267[0]};
    assign in2904_2 = {s1241[1],pp127[38],pp122[44],s1268[0]};
    CLA_4 KS_2904(s2904, c2904, in2904_1, in2904_2);
    wire[3:0] s2905, in2905_1, in2905_2;
    wire c2905;
    assign in2905_1 = {s1242[1],s1231[2],pp123[43],s1269[0]};
    assign in2905_2 = {s1243[1],s1232[2],pp124[42],s1270[0]};
    CLA_4 KS_2905(s2905, c2905, in2905_1, in2905_2);
    wire[3:0] s2906, in2906_1, in2906_2;
    wire c2906;
    assign in2906_1 = {s1244[1],s1233[2],pp125[41],s1271[0]};
    assign in2906_2 = {s1245[1],s1234[2],pp126[40],s1272[0]};
    CLA_4 KS_2906(s2906, c2906, in2906_1, in2906_2);
    wire[3:0] s2907, in2907_1, in2907_2;
    wire c2907;
    assign in2907_1 = {s1246[1],s1235[2],pp127[39],s1273[0]};
    assign in2907_2 = {c1247,s1236[2],s1231[3],s1274[0]};
    CLA_4 KS_2907(s2907, c2907, in2907_1, in2907_2);
    wire[3:0] s2908, in2908_1, in2908_2;
    wire c2908;
    assign in2908_1 = {s1248[1],s1237[2],s1232[3],s1275[0]};
    assign in2908_2 = {c1249,s1238[2],s1233[3],s1276[0]};
    CLA_4 KS_2908(s2908, c2908, in2908_1, in2908_2);
    wire[3:0] s2909, in2909_1, in2909_2;
    wire c2909;
    assign in2909_1 = {s1250[1],s1239[2],s1234[3],s1277[0]};
    assign in2909_2 = {c1251,s1240[2],s1235[3],s1278[0]};
    CLA_4 KS_2909(s2909, c2909, in2909_1, in2909_2);
    wire[3:0] s2910, in2910_1, in2910_2;
    wire c2910;
    assign in2910_1 = {s1252[1],s1241[2],s1236[3],s1279[0]};
    assign in2910_2 = {c1253,s1242[2],s1237[3],s1280[0]};
    CLA_4 KS_2910(s2910, c2910, in2910_1, in2910_2);
    wire[1:0] s2911, in2911_1, in2911_2;
    wire c2911;
    assign in2911_1 = {s1254[1],s1243[2]};
    assign in2911_2 = {c1255,s1244[2]};
    CLA_2 KS_2911(s2911, c2911, in2911_1, in2911_2);
    wire[0:0] s2912, in2912_1, in2912_2;
    wire c2912;
    assign in2912_1 = {s1256[1]};
    assign in2912_2 = {c1257};
    Half_Adder KS_2912(s2912, c2912, in2912_1, in2912_2);
    wire[3:0] s2913, in2913_1, in2913_2;
    wire c2913;
    assign in2913_1 = {s1258[1],s1245[2],s1238[3],s1281[0]};
    assign in2913_2 = {c1259,c1246,s1239[3],s1282[0]};
    CLA_4 KS_2913(s2913, c2913, in2913_1, in2913_2);
    wire[0:0] s2914, in2914_1, in2914_2;
    wire c2914;
    assign in2914_1 = {s1260[1]};
    assign in2914_2 = {c1261};
    Half_Adder KS_2914(s2914, c2914, in2914_1, in2914_2);
    wire[1:0] s2915, in2915_1, in2915_2;
    wire c2915;
    assign in2915_1 = {s1262[1],s1248[2]};
    assign in2915_2 = {c1263,c1250};
    CLA_2 KS_2915(s2915, c2915, in2915_1, in2915_2);
    wire[0:0] s2916, in2916_1, in2916_2;
    wire c2916;
    assign in2916_1 = {s1264[1]};
    assign in2916_2 = {c1265};
    Half_Adder KS_2916(s2916, c2916, in2916_1, in2916_2);
    wire[2:0] s2917, in2917_1, in2917_2;
    wire c2917;
    assign in2917_1 = {s1266[1],s1252[2],s1240[3]};
    assign in2917_2 = {c2815,c1254,s1241[3]};
    CLA_3 KS_2917(s2917, c2917, in2917_1, in2917_2);
    wire[0:0] s2918, in2918_1, in2918_2;
    wire c2918;
    assign in2918_1 = {c2816};
    assign in2918_2 = {c2817};
    Half_Adder KS_2918(s2918, c2918, in2918_1, in2918_2);
    wire[1:0] s2919, in2919_1, in2919_2;
    wire c2919;
    assign in2919_1 = {c2818,s1256[2]};
    assign in2919_2 = {c2819,c1258};
    CLA_2 KS_2919(s2919, c2919, in2919_1, in2919_2);
    wire[0:0] s2920, in2920_1, in2920_2;
    wire c2920;
    assign in2920_1 = {c2820};
    assign in2920_2 = {c2821};
    Half_Adder KS_2920(s2920, c2920, in2920_1, in2920_2);
    wire[3:0] s2921, in2921_1, in2921_2;
    wire c2921;
    assign in2921_1 = {c2822,s1260[2],s1242[3],s1283[0]};
    assign in2921_2 = {c2823,c1262,s1243[3],s1284[0]};
    CLA_4 KS_2921(s2921, c2921, in2921_1, in2921_2);
    wire[0:0] s2922, in2922_1, in2922_2;
    wire c2922;
    assign in2922_1 = {c2824};
    assign in2922_2 = {c2825};
    Half_Adder KS_2922(s2922, c2922, in2922_1, in2922_2);
    wire[1:0] s2923, in2923_1, in2923_2;
    wire c2923;
    assign in2923_1 = {c2826,s1264[2]};
    assign in2923_2 = {c2827,c1266};
    CLA_2 KS_2923(s2923, c2923, in2923_1, in2923_2);
    wire[0:0] s2924, in2924_1, in2924_2;
    wire c2924;
    assign in2924_1 = {c2828};
    assign in2924_2 = {c2829};
    Half_Adder KS_2924(s2924, c2924, in2924_1, in2924_2);
    wire[2:0] s2925, in2925_1, in2925_2;
    wire c2925;
    assign in2925_1 = {c2830,s2880[1],s1244[3]};
    assign in2925_2 = {c2831,s2881[1],c1245};
    CLA_3 KS_2925(s2925, c2925, in2925_1, in2925_2);
    wire[0:0] s2926, in2926_1, in2926_2;
    wire c2926;
    assign in2926_1 = {c2832};
    assign in2926_2 = {c2833};
    Half_Adder KS_2926(s2926, c2926, in2926_1, in2926_2);
    wire[1:0] s2927, in2927_1, in2927_2;
    wire c2927;
    assign in2927_1 = {c2834,s2882[1]};
    assign in2927_2 = {c2835,s2883[1]};
    CLA_2 KS_2927(s2927, c2927, in2927_1, in2927_2);
    wire[0:0] s2928, in2928_1, in2928_2;
    wire c2928;
    assign in2928_1 = {c2836};
    assign in2928_2 = {c2837};
    Half_Adder KS_2928(s2928, c2928, in2928_1, in2928_2);
    wire[3:0] s2929, in2929_1, in2929_2;
    wire c2929;
    assign in2929_1 = {c2838,s2884[1],s1248[3],s1285[0]};
    assign in2929_2 = {c2839,s2885[1],c1252,s1286[0]};
    CLA_4 KS_2929(s2929, c2929, in2929_1, in2929_2);
    wire[0:0] s2930, in2930_1, in2930_2;
    wire c2930;
    assign in2930_1 = {c2840};
    assign in2930_2 = {c2841};
    Half_Adder KS_2930(s2930, c2930, in2930_1, in2930_2);
    wire[1:0] s2931, in2931_1, in2931_2;
    wire c2931;
    assign in2931_1 = {c2842,s2886[1]};
    assign in2931_2 = {c2843,s2887[1]};
    CLA_2 KS_2931(s2931, c2931, in2931_1, in2931_2);
    wire[0:0] s2932, in2932_1, in2932_2;
    wire c2932;
    assign in2932_1 = {c2844};
    assign in2932_2 = {c2845};
    Half_Adder KS_2932(s2932, c2932, in2932_1, in2932_2);
    wire[2:0] s2933, in2933_1, in2933_2;
    wire c2933;
    assign in2933_1 = {c2846,s2888[1],s1256[3]};
    assign in2933_2 = {c2854,s2889[1],c1260};
    CLA_3 KS_2933(s2933, c2933, in2933_1, in2933_2);
    wire[0:0] s2934, in2934_1, in2934_2;
    wire c2934;
    assign in2934_1 = {c2862};
    assign in2934_2 = {c2870};
    Half_Adder KS_2934(s2934, c2934, in2934_1, in2934_2);
    wire[1:0] s2935, in2935_1, in2935_2;
    wire c2935;
    assign in2935_1 = {c2878,s2890[1]};
    assign in2935_2 = {s2880[0],s2891[1]};
    CLA_2 KS_2935(s2935, c2935, in2935_1, in2935_2);
    wire[0:0] s2936, in2936_1, in2936_2;
    wire c2936;
    assign in2936_1 = {s2881[0]};
    assign in2936_2 = {s2882[0]};
    Half_Adder KS_2936(s2936, c2936, in2936_1, in2936_2);
    wire[3:0] s2937, in2937_1, in2937_2;
    wire c2937;
    assign in2937_1 = {s2883[0],s2892[1],s1264[3],s1287[0]};
    assign in2937_2 = {s2884[0],s2893[1],s2880[2],s1288[0]};
    CLA_4 KS_2937(s2937, c2937, in2937_1, in2937_2);
    wire[0:0] s2938, in2938_1, in2938_2;
    wire c2938;
    assign in2938_1 = {s2885[0]};
    assign in2938_2 = {s2886[0]};
    Half_Adder KS_2938(s2938, c2938, in2938_1, in2938_2);
    wire[1:0] s2939, in2939_1, in2939_2;
    wire c2939;
    assign in2939_1 = {s2887[0],s2894[1]};
    assign in2939_2 = {s2888[0],s2895[1]};
    CLA_2 KS_2939(s2939, c2939, in2939_1, in2939_2);
    wire[0:0] s2940, in2940_1, in2940_2;
    wire c2940;
    assign in2940_1 = {s2889[0]};
    assign in2940_2 = {s2890[0]};
    Half_Adder KS_2940(s2940, c2940, in2940_1, in2940_2);
    wire[2:0] s2941, in2941_1, in2941_2;
    wire c2941;
    assign in2941_1 = {s2891[0],s2896[1],s2881[2]};
    assign in2941_2 = {s2892[0],s2897[1],s2882[2]};
    CLA_3 KS_2941(s2941, c2941, in2941_1, in2941_2);
    wire[0:0] s2942, in2942_1, in2942_2;
    wire c2942;
    assign in2942_1 = {s2893[0]};
    assign in2942_2 = {s2894[0]};
    Half_Adder KS_2942(s2942, c2942, in2942_1, in2942_2);
    wire[1:0] s2943, in2943_1, in2943_2;
    wire c2943;
    assign in2943_1 = {s2895[0],s2898[1]};
    assign in2943_2 = {s2896[0],s2899[1]};
    CLA_2 KS_2943(s2943, c2943, in2943_1, in2943_2);
    wire[0:0] s2944, in2944_1, in2944_2;
    wire c2944;
    assign in2944_1 = {s2898[0]};
    assign in2944_2 = {s2899[0]};
    Full_Adder KS_2944(s2944, c2944, in2944_1, in2944_2, s2897[0]);
    wire[3:0] s2945, in2945_1, in2945_2;
    wire c2945;
    assign in2945_1 = {pp81[87],pp72[97],pp67[103],pp83[88]};
    assign in2945_2 = {pp82[86],pp73[96],pp68[102],pp84[87]};
    CLA_4 KS_2945(s2945, c2945, in2945_1, in2945_2);
    wire[3:0] s2946, in2946_1, in2946_2;
    wire c2946;
    assign in2946_1 = {pp83[85],pp74[95],pp69[101],pp85[86]};
    assign in2946_2 = {pp84[84],pp75[94],pp70[100],pp86[85]};
    CLA_4 KS_2946(s2946, c2946, in2946_1, in2946_2);
    wire[3:0] s2947, in2947_1, in2947_2;
    wire c2947;
    assign in2947_1 = {pp85[83],pp76[93],pp71[99],pp87[84]};
    assign in2947_2 = {pp86[82],pp77[92],pp72[98],pp88[83]};
    CLA_4 KS_2947(s2947, c2947, in2947_1, in2947_2);
    wire[3:0] s2948, in2948_1, in2948_2;
    wire c2948;
    assign in2948_1 = {pp87[81],pp78[91],pp73[97],pp89[82]};
    assign in2948_2 = {pp88[80],pp79[90],pp74[96],pp90[81]};
    CLA_4 KS_2948(s2948, c2948, in2948_1, in2948_2);
    wire[3:0] s2949, in2949_1, in2949_2;
    wire c2949;
    assign in2949_1 = {pp89[79],pp80[89],pp75[95],pp91[80]};
    assign in2949_2 = {pp90[78],pp81[88],pp76[94],pp92[79]};
    CLA_4 KS_2949(s2949, c2949, in2949_1, in2949_2);
    wire[3:0] s2950, in2950_1, in2950_2;
    wire c2950;
    assign in2950_1 = {pp91[77],pp82[87],pp77[93],pp93[78]};
    assign in2950_2 = {pp92[76],pp83[86],pp78[92],pp94[77]};
    CLA_4 KS_2950(s2950, c2950, in2950_1, in2950_2);
    wire[3:0] s2951, in2951_1, in2951_2;
    wire c2951;
    assign in2951_1 = {pp93[75],pp84[85],pp79[91],pp95[76]};
    assign in2951_2 = {pp94[74],pp85[84],pp80[90],pp96[75]};
    CLA_4 KS_2951(s2951, c2951, in2951_1, in2951_2);
    wire[3:0] s2952, in2952_1, in2952_2;
    wire c2952;
    assign in2952_1 = {pp95[73],pp86[83],pp81[89],pp97[74]};
    assign in2952_2 = {pp96[72],pp87[82],pp82[88],pp98[73]};
    CLA_4 KS_2952(s2952, c2952, in2952_1, in2952_2);
    wire[3:0] s2953, in2953_1, in2953_2;
    wire c2953;
    assign in2953_1 = {pp97[71],pp88[81],pp83[87],pp99[72]};
    assign in2953_2 = {pp98[70],pp89[80],pp84[86],pp100[71]};
    CLA_4 KS_2953(s2953, c2953, in2953_1, in2953_2);
    wire[3:0] s2954, in2954_1, in2954_2;
    wire c2954;
    assign in2954_1 = {pp99[69],pp90[79],pp85[85],pp101[70]};
    assign in2954_2 = {pp100[68],pp91[78],pp86[84],pp102[69]};
    CLA_4 KS_2954(s2954, c2954, in2954_1, in2954_2);
    wire[3:0] s2955, in2955_1, in2955_2;
    wire c2955;
    assign in2955_1 = {pp101[67],pp92[77],pp87[83],pp103[68]};
    assign in2955_2 = {pp102[66],pp93[76],pp88[82],pp104[67]};
    CLA_4 KS_2955(s2955, c2955, in2955_1, in2955_2);
    wire[3:0] s2956, in2956_1, in2956_2;
    wire c2956;
    assign in2956_1 = {pp103[65],pp94[75],pp89[81],pp105[66]};
    assign in2956_2 = {pp104[64],pp95[74],pp90[80],pp106[65]};
    CLA_4 KS_2956(s2956, c2956, in2956_1, in2956_2);
    wire[3:0] s2957, in2957_1, in2957_2;
    wire c2957;
    assign in2957_1 = {pp105[63],pp96[73],pp91[79],pp107[64]};
    assign in2957_2 = {pp106[62],pp97[72],pp92[78],pp108[63]};
    CLA_4 KS_2957(s2957, c2957, in2957_1, in2957_2);
    wire[3:0] s2958, in2958_1, in2958_2;
    wire c2958;
    assign in2958_1 = {pp107[61],pp98[71],pp93[77],pp109[62]};
    assign in2958_2 = {pp108[60],pp99[70],pp94[76],pp110[61]};
    CLA_4 KS_2958(s2958, c2958, in2958_1, in2958_2);
    wire[3:0] s2959, in2959_1, in2959_2;
    wire c2959;
    assign in2959_1 = {pp109[59],pp100[69],pp95[75],pp111[60]};
    assign in2959_2 = {pp110[58],pp101[68],pp96[74],pp112[59]};
    CLA_4 KS_2959(s2959, c2959, in2959_1, in2959_2);
    wire[3:0] s2960, in2960_1, in2960_2;
    wire c2960;
    assign in2960_1 = {pp111[57],pp102[67],pp97[73],pp113[58]};
    assign in2960_2 = {pp112[56],pp103[66],pp98[72],pp114[57]};
    CLA_4 KS_2960(s2960, c2960, in2960_1, in2960_2);
    wire[3:0] s2961, in2961_1, in2961_2;
    wire c2961;
    assign in2961_1 = {pp113[55],pp104[65],pp99[71],pp115[56]};
    assign in2961_2 = {pp114[54],pp105[64],pp100[70],pp116[55]};
    CLA_4 KS_2961(s2961, c2961, in2961_1, in2961_2);
    wire[3:0] s2962, in2962_1, in2962_2;
    wire c2962;
    assign in2962_1 = {pp115[53],pp106[63],pp101[69],pp117[54]};
    assign in2962_2 = {pp116[52],pp107[62],pp102[68],pp118[53]};
    CLA_4 KS_2962(s2962, c2962, in2962_1, in2962_2);
    wire[3:0] s2963, in2963_1, in2963_2;
    wire c2963;
    assign in2963_1 = {pp117[51],pp108[61],pp103[67],pp119[52]};
    assign in2963_2 = {pp118[50],pp109[60],pp104[66],pp120[51]};
    CLA_4 KS_2963(s2963, c2963, in2963_1, in2963_2);
    wire[3:0] s2964, in2964_1, in2964_2;
    wire c2964;
    assign in2964_1 = {pp119[49],pp110[59],pp105[65],pp121[50]};
    assign in2964_2 = {pp120[48],pp111[58],pp106[64],pp122[49]};
    CLA_4 KS_2964(s2964, c2964, in2964_1, in2964_2);
    wire[3:0] s2965, in2965_1, in2965_2;
    wire c2965;
    assign in2965_1 = {pp121[47],pp112[57],pp107[63],pp123[48]};
    assign in2965_2 = {pp122[46],pp113[56],pp108[62],pp124[47]};
    CLA_4 KS_2965(s2965, c2965, in2965_1, in2965_2);
    wire[3:0] s2966, in2966_1, in2966_2;
    wire c2966;
    assign in2966_1 = {pp123[45],pp114[55],pp109[61],pp125[46]};
    assign in2966_2 = {pp124[44],pp115[54],pp110[60],pp126[45]};
    CLA_4 KS_2966(s2966, c2966, in2966_1, in2966_2);
    wire[3:0] s2967, in2967_1, in2967_2;
    wire c2967;
    assign in2967_1 = {pp125[43],pp116[53],pp111[59],pp127[44]};
    assign in2967_2 = {pp126[42],pp117[52],pp112[58],c1267};
    CLA_4 KS_2967(s2967, c2967, in2967_1, in2967_2);
    wire[3:0] s2968, in2968_1, in2968_2;
    wire c2968;
    assign in2968_1 = {pp127[41],pp118[51],pp113[57],c1268};
    assign in2968_2 = {s1267[1],pp119[50],pp114[56],c1269};
    CLA_4 KS_2968(s2968, c2968, in2968_1, in2968_2);
    wire[3:0] s2969, in2969_1, in2969_2;
    wire c2969;
    assign in2969_1 = {s1268[1],pp120[49],pp115[55],c1270};
    assign in2969_2 = {s1269[1],pp121[48],pp116[54],c1271};
    CLA_4 KS_2969(s2969, c2969, in2969_1, in2969_2);
    wire[3:0] s2970, in2970_1, in2970_2;
    wire c2970;
    assign in2970_1 = {s1270[1],pp122[47],pp117[53],c1272};
    assign in2970_2 = {s1271[1],pp123[46],pp118[52],c1273};
    CLA_4 KS_2970(s2970, c2970, in2970_1, in2970_2);
    wire[3:0] s2971, in2971_1, in2971_2;
    wire c2971;
    assign in2971_1 = {s1272[1],pp124[45],pp119[51],c1274};
    assign in2971_2 = {s1273[1],pp125[44],pp120[50],c1275};
    CLA_4 KS_2971(s2971, c2971, in2971_1, in2971_2);
    wire[3:0] s2972, in2972_1, in2972_2;
    wire c2972;
    assign in2972_1 = {s1274[1],pp126[43],pp121[49],c1276};
    assign in2972_2 = {s1275[1],pp127[42],pp122[48],c1280};
    CLA_4 KS_2972(s2972, c2972, in2972_1, in2972_2);
    wire[3:0] s2973, in2973_1, in2973_2;
    wire c2973;
    assign in2973_1 = {s1276[1],s1267[2],pp123[47],c1288};
    assign in2973_2 = {s1277[1],s1268[2],pp124[46],s1295[0]};
    CLA_4 KS_2973(s2973, c2973, in2973_1, in2973_2);
    wire[3:0] s2974, in2974_1, in2974_2;
    wire c2974;
    assign in2974_1 = {s1278[1],s1269[2],pp125[45],s1296[0]};
    assign in2974_2 = {c1279,s1270[2],pp126[44],s1297[0]};
    CLA_4 KS_2974(s2974, c2974, in2974_1, in2974_2);
    wire[3:0] s2975, in2975_1, in2975_2;
    wire c2975;
    assign in2975_1 = {s1280[1],s1271[2],pp127[43],s1298[0]};
    assign in2975_2 = {c1281,s1272[2],s1267[3],s1299[0]};
    CLA_4 KS_2975(s2975, c2975, in2975_1, in2975_2);
    wire[3:0] s2976, in2976_1, in2976_2;
    wire c2976;
    assign in2976_1 = {s1282[1],s1273[2],s1268[3],s1300[0]};
    assign in2976_2 = {c1283,s1274[2],s1269[3],s1301[0]};
    CLA_4 KS_2976(s2976, c2976, in2976_1, in2976_2);
    wire[0:0] s2977, in2977_1, in2977_2;
    wire c2977;
    assign in2977_1 = {s1284[1]};
    assign in2977_2 = {c1285};
    Half_Adder KS_2977(s2977, c2977, in2977_1, in2977_2);
    wire[1:0] s2978, in2978_1, in2978_2;
    wire c2978;
    assign in2978_1 = {s1286[1],s1275[2]};
    assign in2978_2 = {c1287,s1276[2]};
    CLA_2 KS_2978(s2978, c2978, in2978_1, in2978_2);
    wire[0:0] s2979, in2979_1, in2979_2;
    wire c2979;
    assign in2979_1 = {s1288[1]};
    assign in2979_2 = {c1289};
    Half_Adder KS_2979(s2979, c2979, in2979_1, in2979_2);
    wire[2:0] s2980, in2980_1, in2980_2;
    wire c2980;
    assign in2980_1 = {s1290[1],s1277[2],s1270[3]};
    assign in2980_2 = {c1291,c1278,s1271[3]};
    CLA_3 KS_2980(s2980, c2980, in2980_1, in2980_2);
    wire[0:0] s2981, in2981_1, in2981_2;
    wire c2981;
    assign in2981_1 = {s1292[1]};
    assign in2981_2 = {c1293};
    Half_Adder KS_2981(s2981, c2981, in2981_1, in2981_2);
    wire[1:0] s2982, in2982_1, in2982_2;
    wire c2982;
    assign in2982_1 = {s1294[1],s1280[2]};
    assign in2982_2 = {c2880,c1282};
    CLA_2 KS_2982(s2982, c2982, in2982_1, in2982_2);
    wire[0:0] s2983, in2983_1, in2983_2;
    wire c2983;
    assign in2983_1 = {c2881};
    assign in2983_2 = {c2882};
    Half_Adder KS_2983(s2983, c2983, in2983_1, in2983_2);
    wire[3:0] s2984, in2984_1, in2984_2;
    wire c2984;
    assign in2984_1 = {c2883,s1284[2],s1272[3],s1302[0]};
    assign in2984_2 = {c2884,c1286,s1273[3],s1303[0]};
    CLA_4 KS_2984(s2984, c2984, in2984_1, in2984_2);
    wire[0:0] s2985, in2985_1, in2985_2;
    wire c2985;
    assign in2985_1 = {c2885};
    assign in2985_2 = {c2886};
    Half_Adder KS_2985(s2985, c2985, in2985_1, in2985_2);
    wire[1:0] s2986, in2986_1, in2986_2;
    wire c2986;
    assign in2986_1 = {c2887,s1288[2]};
    assign in2986_2 = {c2888,c1290};
    CLA_2 KS_2986(s2986, c2986, in2986_1, in2986_2);
    wire[0:0] s2987, in2987_1, in2987_2;
    wire c2987;
    assign in2987_1 = {c2889};
    assign in2987_2 = {c2890};
    Half_Adder KS_2987(s2987, c2987, in2987_1, in2987_2);
    wire[2:0] s2988, in2988_1, in2988_2;
    wire c2988;
    assign in2988_1 = {c2891,s1292[2],s1274[3]};
    assign in2988_2 = {c2892,c1294,s1275[3]};
    CLA_3 KS_2988(s2988, c2988, in2988_1, in2988_2);
    wire[0:0] s2989, in2989_1, in2989_2;
    wire c2989;
    assign in2989_1 = {c2893};
    assign in2989_2 = {c2894};
    Half_Adder KS_2989(s2989, c2989, in2989_1, in2989_2);
    wire[1:0] s2990, in2990_1, in2990_2;
    wire c2990;
    assign in2990_1 = {c2895,s2945[1]};
    assign in2990_2 = {c2896,s2946[1]};
    CLA_2 KS_2990(s2990, c2990, in2990_1, in2990_2);
    wire[0:0] s2991, in2991_1, in2991_2;
    wire c2991;
    assign in2991_1 = {c2897};
    assign in2991_2 = {c2898};
    Half_Adder KS_2991(s2991, c2991, in2991_1, in2991_2);
    wire[3:0] s2992, in2992_1, in2992_2;
    wire c2992;
    assign in2992_1 = {c2899,s2947[1],s1276[3],s1304[0]};
    assign in2992_2 = {c2900,s2948[1],c1277,s1305[0]};
    CLA_4 KS_2992(s2992, c2992, in2992_1, in2992_2);
    wire[0:0] s2993, in2993_1, in2993_2;
    wire c2993;
    assign in2993_1 = {c2901};
    assign in2993_2 = {c2902};
    Half_Adder KS_2993(s2993, c2993, in2993_1, in2993_2);
    wire[1:0] s2994, in2994_1, in2994_2;
    wire c2994;
    assign in2994_1 = {c2903,s2949[1]};
    assign in2994_2 = {c2904,s2950[1]};
    CLA_2 KS_2994(s2994, c2994, in2994_1, in2994_2);
    wire[0:0] s2995, in2995_1, in2995_2;
    wire c2995;
    assign in2995_1 = {c2905};
    assign in2995_2 = {c2906};
    Half_Adder KS_2995(s2995, c2995, in2995_1, in2995_2);
    wire[2:0] s2996, in2996_1, in2996_2;
    wire c2996;
    assign in2996_1 = {c2907,s2951[1],s1280[3]};
    assign in2996_2 = {c2908,s2952[1],c1284};
    CLA_3 KS_2996(s2996, c2996, in2996_1, in2996_2);
    wire[0:0] s2997, in2997_1, in2997_2;
    wire c2997;
    assign in2997_1 = {c2909};
    assign in2997_2 = {c2910};
    Half_Adder KS_2997(s2997, c2997, in2997_1, in2997_2);
    wire[1:0] s2998, in2998_1, in2998_2;
    wire c2998;
    assign in2998_1 = {c2913,s2953[1]};
    assign in2998_2 = {c2921,s2954[1]};
    CLA_2 KS_2998(s2998, c2998, in2998_1, in2998_2);
    wire[0:0] s2999, in2999_1, in2999_2;
    wire c2999;
    assign in2999_1 = {c2929};
    assign in2999_2 = {c2937};
    Half_Adder KS_2999(s2999, c2999, in2999_1, in2999_2);
    wire[3:0] s3000, in3000_1, in3000_2;
    wire c3000;
    assign in3000_1 = {s2945[0],s2955[1],s1288[3],s1306[0]};
    assign in3000_2 = {s2946[0],s2956[1],c1292,s1307[0]};
    CLA_4 KS_3000(s3000, c3000, in3000_1, in3000_2);
    wire[0:0] s3001, in3001_1, in3001_2;
    wire c3001;
    assign in3001_1 = {s2947[0]};
    assign in3001_2 = {s2948[0]};
    Half_Adder KS_3001(s3001, c3001, in3001_1, in3001_2);
    wire[1:0] s3002, in3002_1, in3002_2;
    wire c3002;
    assign in3002_1 = {s2949[0],s2957[1]};
    assign in3002_2 = {s2950[0],s2958[1]};
    CLA_2 KS_3002(s3002, c3002, in3002_1, in3002_2);
    wire[0:0] s3003, in3003_1, in3003_2;
    wire c3003;
    assign in3003_1 = {s2951[0]};
    assign in3003_2 = {s2952[0]};
    Half_Adder KS_3003(s3003, c3003, in3003_1, in3003_2);
    wire[2:0] s3004, in3004_1, in3004_2;
    wire c3004;
    assign in3004_1 = {s2953[0],s2959[1],s2945[2]};
    assign in3004_2 = {s2954[0],s2960[1],s2946[2]};
    CLA_3 KS_3004(s3004, c3004, in3004_1, in3004_2);
    wire[0:0] s3005, in3005_1, in3005_2;
    wire c3005;
    assign in3005_1 = {s2955[0]};
    assign in3005_2 = {s2956[0]};
    Half_Adder KS_3005(s3005, c3005, in3005_1, in3005_2);
    wire[1:0] s3006, in3006_1, in3006_2;
    wire c3006;
    assign in3006_1 = {s2957[0],s2961[1]};
    assign in3006_2 = {s2958[0],s2962[1]};
    CLA_2 KS_3006(s3006, c3006, in3006_1, in3006_2);
    wire[0:0] s3007, in3007_1, in3007_2;
    wire c3007;
    assign in3007_1 = {s2959[0]};
    assign in3007_2 = {s2960[0]};
    Half_Adder KS_3007(s3007, c3007, in3007_1, in3007_2);
    wire[3:0] s3008, in3008_1, in3008_2;
    wire c3008;
    assign in3008_1 = {s2962[0],s2963[1],s2947[2],s1308[0]};
    assign in3008_2 = {s2963[0],s2964[1],s2948[2],s1309[0]};
    CLA_4_c KS_3008(s3008, c3008, in3008_1, in3008_2, s2961[0]);
    wire[3:0] s3009, in3009_1, in3009_2;
    wire c3009;
    assign in3009_1 = {pp71[101],pp66[107],pp63[111],pp71[104]};
    assign in3009_2 = {pp72[100],pp67[106],pp64[110],pp72[103]};
    CLA_4 KS_3009(s3009, c3009, in3009_1, in3009_2);
    wire[3:0] s3010, in3010_1, in3010_2;
    wire c3010;
    assign in3010_1 = {pp73[99],pp68[105],pp65[109],pp73[102]};
    assign in3010_2 = {pp74[98],pp69[104],pp66[108],pp74[101]};
    CLA_4 KS_3010(s3010, c3010, in3010_1, in3010_2);
    wire[3:0] s3011, in3011_1, in3011_2;
    wire c3011;
    assign in3011_1 = {pp75[97],pp70[103],pp67[107],pp75[100]};
    assign in3011_2 = {pp76[96],pp71[102],pp68[106],pp76[99]};
    CLA_4 KS_3011(s3011, c3011, in3011_1, in3011_2);
    wire[3:0] s3012, in3012_1, in3012_2;
    wire c3012;
    assign in3012_1 = {pp77[95],pp72[101],pp69[105],pp77[98]};
    assign in3012_2 = {pp78[94],pp73[100],pp70[104],pp78[97]};
    CLA_4 KS_3012(s3012, c3012, in3012_1, in3012_2);
    wire[3:0] s3013, in3013_1, in3013_2;
    wire c3013;
    assign in3013_1 = {pp79[93],pp74[99],pp71[103],pp79[96]};
    assign in3013_2 = {pp80[92],pp75[98],pp72[102],pp80[95]};
    CLA_4 KS_3013(s3013, c3013, in3013_1, in3013_2);
    wire[3:0] s3014, in3014_1, in3014_2;
    wire c3014;
    assign in3014_1 = {pp81[91],pp76[97],pp73[101],pp81[94]};
    assign in3014_2 = {pp82[90],pp77[96],pp74[100],pp82[93]};
    CLA_4 KS_3014(s3014, c3014, in3014_1, in3014_2);
    wire[3:0] s3015, in3015_1, in3015_2;
    wire c3015;
    assign in3015_1 = {pp83[89],pp78[95],pp75[99],pp83[92]};
    assign in3015_2 = {pp84[88],pp79[94],pp76[98],pp84[91]};
    CLA_4 KS_3015(s3015, c3015, in3015_1, in3015_2);
    wire[3:0] s3016, in3016_1, in3016_2;
    wire c3016;
    assign in3016_1 = {pp85[87],pp80[93],pp77[97],pp85[90]};
    assign in3016_2 = {pp86[86],pp81[92],pp78[96],pp86[89]};
    CLA_4 KS_3016(s3016, c3016, in3016_1, in3016_2);
    wire[3:0] s3017, in3017_1, in3017_2;
    wire c3017;
    assign in3017_1 = {pp87[85],pp82[91],pp79[95],pp87[88]};
    assign in3017_2 = {pp88[84],pp83[90],pp80[94],pp88[87]};
    CLA_4 KS_3017(s3017, c3017, in3017_1, in3017_2);
    wire[3:0] s3018, in3018_1, in3018_2;
    wire c3018;
    assign in3018_1 = {pp89[83],pp84[89],pp81[93],pp89[86]};
    assign in3018_2 = {pp90[82],pp85[88],pp82[92],pp90[85]};
    CLA_4 KS_3018(s3018, c3018, in3018_1, in3018_2);
    wire[3:0] s3019, in3019_1, in3019_2;
    wire c3019;
    assign in3019_1 = {pp91[81],pp86[87],pp83[91],pp91[84]};
    assign in3019_2 = {pp92[80],pp87[86],pp84[90],pp92[83]};
    CLA_4 KS_3019(s3019, c3019, in3019_1, in3019_2);
    wire[3:0] s3020, in3020_1, in3020_2;
    wire c3020;
    assign in3020_1 = {pp93[79],pp88[85],pp85[89],pp93[82]};
    assign in3020_2 = {pp94[78],pp89[84],pp86[88],pp94[81]};
    CLA_4 KS_3020(s3020, c3020, in3020_1, in3020_2);
    wire[3:0] s3021, in3021_1, in3021_2;
    wire c3021;
    assign in3021_1 = {pp95[77],pp90[83],pp87[87],pp95[80]};
    assign in3021_2 = {pp96[76],pp91[82],pp88[86],pp96[79]};
    CLA_4 KS_3021(s3021, c3021, in3021_1, in3021_2);
    wire[3:0] s3022, in3022_1, in3022_2;
    wire c3022;
    assign in3022_1 = {pp97[75],pp92[81],pp89[85],pp97[78]};
    assign in3022_2 = {pp98[74],pp93[80],pp90[84],pp98[77]};
    CLA_4 KS_3022(s3022, c3022, in3022_1, in3022_2);
    wire[3:0] s3023, in3023_1, in3023_2;
    wire c3023;
    assign in3023_1 = {pp99[73],pp94[79],pp91[83],pp99[76]};
    assign in3023_2 = {pp100[72],pp95[78],pp92[82],pp100[75]};
    CLA_4 KS_3023(s3023, c3023, in3023_1, in3023_2);
    wire[3:0] s3024, in3024_1, in3024_2;
    wire c3024;
    assign in3024_1 = {pp101[71],pp96[77],pp93[81],pp101[74]};
    assign in3024_2 = {pp102[70],pp97[76],pp94[80],pp102[73]};
    CLA_4 KS_3024(s3024, c3024, in3024_1, in3024_2);
    wire[3:0] s3025, in3025_1, in3025_2;
    wire c3025;
    assign in3025_1 = {pp103[69],pp98[75],pp95[79],pp103[72]};
    assign in3025_2 = {pp104[68],pp99[74],pp96[78],pp104[71]};
    CLA_4 KS_3025(s3025, c3025, in3025_1, in3025_2);
    wire[3:0] s3026, in3026_1, in3026_2;
    wire c3026;
    assign in3026_1 = {pp105[67],pp100[73],pp97[77],pp105[70]};
    assign in3026_2 = {pp106[66],pp101[72],pp98[76],pp106[69]};
    CLA_4 KS_3026(s3026, c3026, in3026_1, in3026_2);
    wire[3:0] s3027, in3027_1, in3027_2;
    wire c3027;
    assign in3027_1 = {pp107[65],pp102[71],pp99[75],pp107[68]};
    assign in3027_2 = {pp108[64],pp103[70],pp100[74],pp108[67]};
    CLA_4 KS_3027(s3027, c3027, in3027_1, in3027_2);
    wire[3:0] s3028, in3028_1, in3028_2;
    wire c3028;
    assign in3028_1 = {pp109[63],pp104[69],pp101[73],pp109[66]};
    assign in3028_2 = {pp110[62],pp105[68],pp102[72],pp110[65]};
    CLA_4 KS_3028(s3028, c3028, in3028_1, in3028_2);
    wire[3:0] s3029, in3029_1, in3029_2;
    wire c3029;
    assign in3029_1 = {pp111[61],pp106[67],pp103[71],pp111[64]};
    assign in3029_2 = {pp112[60],pp107[66],pp104[70],pp112[63]};
    CLA_4 KS_3029(s3029, c3029, in3029_1, in3029_2);
    wire[3:0] s3030, in3030_1, in3030_2;
    wire c3030;
    assign in3030_1 = {pp113[59],pp108[65],pp105[69],pp113[62]};
    assign in3030_2 = {pp114[58],pp109[64],pp106[68],pp114[61]};
    CLA_4 KS_3030(s3030, c3030, in3030_1, in3030_2);
    wire[3:0] s3031, in3031_1, in3031_2;
    wire c3031;
    assign in3031_1 = {pp115[57],pp110[63],pp107[67],pp115[60]};
    assign in3031_2 = {pp116[56],pp111[62],pp108[66],pp116[59]};
    CLA_4 KS_3031(s3031, c3031, in3031_1, in3031_2);
    wire[3:0] s3032, in3032_1, in3032_2;
    wire c3032;
    assign in3032_1 = {pp117[55],pp112[61],pp109[65],pp117[58]};
    assign in3032_2 = {pp118[54],pp113[60],pp110[64],pp118[57]};
    CLA_4 KS_3032(s3032, c3032, in3032_1, in3032_2);
    wire[3:0] s3033, in3033_1, in3033_2;
    wire c3033;
    assign in3033_1 = {pp119[53],pp114[59],pp111[63],pp119[56]};
    assign in3033_2 = {pp120[52],pp115[58],pp112[62],pp120[55]};
    CLA_4 KS_3033(s3033, c3033, in3033_1, in3033_2);
    wire[3:0] s3034, in3034_1, in3034_2;
    wire c3034;
    assign in3034_1 = {pp121[51],pp116[57],pp113[61],pp121[54]};
    assign in3034_2 = {pp122[50],pp117[56],pp114[60],pp122[53]};
    CLA_4 KS_3034(s3034, c3034, in3034_1, in3034_2);
    wire[3:0] s3035, in3035_1, in3035_2;
    wire c3035;
    assign in3035_1 = {pp123[49],pp118[55],pp115[59],pp123[52]};
    assign in3035_2 = {pp124[48],pp119[54],pp116[58],pp124[51]};
    CLA_4 KS_3035(s3035, c3035, in3035_1, in3035_2);
    wire[3:0] s3036, in3036_1, in3036_2;
    wire c3036;
    assign in3036_1 = {pp125[47],pp120[53],pp117[57],pp125[50]};
    assign in3036_2 = {pp126[46],pp121[52],pp118[56],pp126[49]};
    CLA_4 KS_3036(s3036, c3036, in3036_1, in3036_2);
    wire[3:0] s3037, in3037_1, in3037_2;
    wire c3037;
    assign in3037_1 = {pp127[45],pp122[51],pp119[55],pp127[48]};
    assign in3037_2 = {s1295[1],pp123[50],pp120[54],c1295};
    CLA_4 KS_3037(s3037, c3037, in3037_1, in3037_2);
    wire[3:0] s3038, in3038_1, in3038_2;
    wire c3038;
    assign in3038_1 = {s1296[1],pp124[49],pp121[53],c1296};
    assign in3038_2 = {s1297[1],pp125[48],pp122[52],c1297};
    CLA_4 KS_3038(s3038, c3038, in3038_1, in3038_2);
    wire[3:0] s3039, in3039_1, in3039_2;
    wire c3039;
    assign in3039_1 = {s1298[1],pp126[47],pp123[51],c1298};
    assign in3039_2 = {s1299[1],pp127[46],pp124[50],c1299};
    CLA_4 KS_3039(s3039, c3039, in3039_1, in3039_2);
    wire[0:0] s3040, in3040_1, in3040_2;
    wire c3040;
    assign in3040_1 = {s1300[1]};
    assign in3040_2 = {s1301[1]};
    Half_Adder KS_3040(s3040, c3040, in3040_1, in3040_2);
    wire[1:0] s3041, in3041_1, in3041_2;
    wire c3041;
    assign in3041_1 = {s1302[1],s1295[2]};
    assign in3041_2 = {c1303,s1296[2]};
    CLA_2 KS_3041(s3041, c3041, in3041_1, in3041_2);
    wire[0:0] s3042, in3042_1, in3042_2;
    wire c3042;
    assign in3042_1 = {s1304[1]};
    assign in3042_2 = {c1305};
    Half_Adder KS_3042(s3042, c3042, in3042_1, in3042_2);
    wire[3:0] s3043, in3043_1, in3043_2;
    wire c3043;
    assign in3043_1 = {s1306[1],s1297[2],pp125[49],c1300};
    assign in3043_2 = {c1307,s1298[2],pp126[48],c1304};
    CLA_4 KS_3043(s3043, c3043, in3043_1, in3043_2);
    wire[0:0] s3044, in3044_1, in3044_2;
    wire c3044;
    assign in3044_1 = {s1308[1]};
    assign in3044_2 = {c1309};
    Half_Adder KS_3044(s3044, c3044, in3044_1, in3044_2);
    wire[1:0] s3045, in3045_1, in3045_2;
    wire c3045;
    assign in3045_1 = {s1310[1],s1299[2]};
    assign in3045_2 = {c1311,s1300[2]};
    CLA_2 KS_3045(s3045, c3045, in3045_1, in3045_2);
    wire[0:0] s3046, in3046_1, in3046_2;
    wire c3046;
    assign in3046_1 = {s1312[1]};
    assign in3046_2 = {c1313};
    Half_Adder KS_3046(s3046, c3046, in3046_1, in3046_2);
    wire[2:0] s3047, in3047_1, in3047_2;
    wire c3047;
    assign in3047_1 = {c2945,s1301[2],pp127[47]};
    assign in3047_2 = {c2946,c1302,s1295[3]};
    CLA_3 KS_3047(s3047, c3047, in3047_1, in3047_2);
    wire[0:0] s3048, in3048_1, in3048_2;
    wire c3048;
    assign in3048_1 = {c2947};
    assign in3048_2 = {c2948};
    Half_Adder KS_3048(s3048, c3048, in3048_1, in3048_2);
    wire[1:0] s3049, in3049_1, in3049_2;
    wire c3049;
    assign in3049_1 = {c2949,s1304[2]};
    assign in3049_2 = {c2950,c1306};
    CLA_2 KS_3049(s3049, c3049, in3049_1, in3049_2);
    wire[0:0] s3050, in3050_1, in3050_2;
    wire c3050;
    assign in3050_1 = {c2951};
    assign in3050_2 = {c2952};
    Half_Adder KS_3050(s3050, c3050, in3050_1, in3050_2);
    wire[3:0] s3051, in3051_1, in3051_2;
    wire c3051;
    assign in3051_1 = {c2953,s1308[2],s1296[3],c1312};
    assign in3051_2 = {c2954,c1310,s1297[3],s1314[0]};
    CLA_4 KS_3051(s3051, c3051, in3051_1, in3051_2);
    wire[0:0] s3052, in3052_1, in3052_2;
    wire c3052;
    assign in3052_1 = {c2955};
    assign in3052_2 = {c2956};
    Half_Adder KS_3052(s3052, c3052, in3052_1, in3052_2);
    wire[1:0] s3053, in3053_1, in3053_2;
    wire c3053;
    assign in3053_1 = {c2957,s1312[2]};
    assign in3053_2 = {c2958,s3009[1]};
    CLA_2 KS_3053(s3053, c3053, in3053_1, in3053_2);
    wire[0:0] s3054, in3054_1, in3054_2;
    wire c3054;
    assign in3054_1 = {c2959};
    assign in3054_2 = {c2960};
    Half_Adder KS_3054(s3054, c3054, in3054_1, in3054_2);
    wire[2:0] s3055, in3055_1, in3055_2;
    wire c3055;
    assign in3055_1 = {c2961,s3010[1],s1298[3]};
    assign in3055_2 = {c2962,s3011[1],s1299[3]};
    CLA_3 KS_3055(s3055, c3055, in3055_1, in3055_2);
    wire[0:0] s3056, in3056_1, in3056_2;
    wire c3056;
    assign in3056_1 = {c2963};
    assign in3056_2 = {c2964};
    Half_Adder KS_3056(s3056, c3056, in3056_1, in3056_2);
    wire[1:0] s3057, in3057_1, in3057_2;
    wire c3057;
    assign in3057_1 = {c2965,s3012[1]};
    assign in3057_2 = {c2966,s3013[1]};
    CLA_2 KS_3057(s3057, c3057, in3057_1, in3057_2);
    wire[0:0] s3058, in3058_1, in3058_2;
    wire c3058;
    assign in3058_1 = {c2967};
    assign in3058_2 = {c2968};
    Half_Adder KS_3058(s3058, c3058, in3058_1, in3058_2);
    wire[3:0] s3059, in3059_1, in3059_2;
    wire c3059;
    assign in3059_1 = {c2969,s3014[1],s1300[3],s1315[0]};
    assign in3059_2 = {c2970,s3015[1],c1301,s1316[0]};
    CLA_4 KS_3059(s3059, c3059, in3059_1, in3059_2);
    wire[0:0] s3060, in3060_1, in3060_2;
    wire c3060;
    assign in3060_1 = {c2971};
    assign in3060_2 = {c2972};
    Half_Adder KS_3060(s3060, c3060, in3060_1, in3060_2);
    wire[1:0] s3061, in3061_1, in3061_2;
    wire c3061;
    assign in3061_1 = {c2973,s3016[1]};
    assign in3061_2 = {c2974,s3017[1]};
    CLA_2 KS_3061(s3061, c3061, in3061_1, in3061_2);
    wire[0:0] s3062, in3062_1, in3062_2;
    wire c3062;
    assign in3062_1 = {c2975};
    assign in3062_2 = {c2976};
    Half_Adder KS_3062(s3062, c3062, in3062_1, in3062_2);
    wire[2:0] s3063, in3063_1, in3063_2;
    wire c3063;
    assign in3063_1 = {c2984,s3018[1],s1304[3]};
    assign in3063_2 = {c2992,s3019[1],c1308};
    CLA_3 KS_3063(s3063, c3063, in3063_1, in3063_2);
    wire[0:0] s3064, in3064_1, in3064_2;
    wire c3064;
    assign in3064_1 = {c3000};
    assign in3064_2 = {c3008};
    Half_Adder KS_3064(s3064, c3064, in3064_1, in3064_2);
    wire[1:0] s3065, in3065_1, in3065_2;
    wire c3065;
    assign in3065_1 = {s3009[0],s3020[1]};
    assign in3065_2 = {s3010[0],s3021[1]};
    CLA_2 KS_3065(s3065, c3065, in3065_1, in3065_2);
    wire[0:0] s3066, in3066_1, in3066_2;
    wire c3066;
    assign in3066_1 = {s3011[0]};
    assign in3066_2 = {s3012[0]};
    Half_Adder KS_3066(s3066, c3066, in3066_1, in3066_2);
    wire[3:0] s3067, in3067_1, in3067_2;
    wire c3067;
    assign in3067_1 = {s3013[0],s3022[1],s1312[3],s1317[0]};
    assign in3067_2 = {s3014[0],s3023[1],s3009[2],s1318[0]};
    CLA_4 KS_3067(s3067, c3067, in3067_1, in3067_2);
    wire[0:0] s3068, in3068_1, in3068_2;
    wire c3068;
    assign in3068_1 = {s3015[0]};
    assign in3068_2 = {s3016[0]};
    Half_Adder KS_3068(s3068, c3068, in3068_1, in3068_2);
    wire[1:0] s3069, in3069_1, in3069_2;
    wire c3069;
    assign in3069_1 = {s3017[0],s3024[1]};
    assign in3069_2 = {s3018[0],s3025[1]};
    CLA_2 KS_3069(s3069, c3069, in3069_1, in3069_2);
    wire[0:0] s3070, in3070_1, in3070_2;
    wire c3070;
    assign in3070_1 = {s3019[0]};
    assign in3070_2 = {s3020[0]};
    Half_Adder KS_3070(s3070, c3070, in3070_1, in3070_2);
    wire[2:0] s3071, in3071_1, in3071_2;
    wire c3071;
    assign in3071_1 = {s3021[0],s3026[1],s3010[2]};
    assign in3071_2 = {s3022[0],s3027[1],s3011[2]};
    CLA_3 KS_3071(s3071, c3071, in3071_1, in3071_2);
    wire[0:0] s3072, in3072_1, in3072_2;
    wire c3072;
    assign in3072_1 = {s3023[0]};
    assign in3072_2 = {s3024[0]};
    Half_Adder KS_3072(s3072, c3072, in3072_1, in3072_2);
    wire[1:0] s3073, in3073_1, in3073_2;
    wire c3073;
    assign in3073_1 = {s3025[0],s3028[1]};
    assign in3073_2 = {s3026[0],s3029[1]};
    CLA_2 KS_3073(s3073, c3073, in3073_1, in3073_2);
    wire[0:0] s3074, in3074_1, in3074_2;
    wire c3074;
    assign in3074_1 = {s3028[0]};
    assign in3074_2 = {s3029[0]};
    Full_Adder KS_3074(s3074, c3074, in3074_1, in3074_2, s3027[0]);
    wire[3:0] s3075, in3075_1, in3075_2;
    wire c3075;
    assign in3075_1 = {pp63[113],pp60[117],pp57[121],pp57[122]};
    assign in3075_2 = {pp64[112],pp61[116],pp58[120],pp58[121]};
    CLA_4 KS_3075(s3075, c3075, in3075_1, in3075_2);
    wire[3:0] s3076, in3076_1, in3076_2;
    wire c3076;
    assign in3076_1 = {pp65[111],pp62[115],pp59[119],pp59[120]};
    assign in3076_2 = {pp66[110],pp63[114],pp60[118],pp60[119]};
    CLA_4 KS_3076(s3076, c3076, in3076_1, in3076_2);
    wire[3:0] s3077, in3077_1, in3077_2;
    wire c3077;
    assign in3077_1 = {pp67[109],pp64[113],pp61[117],pp61[118]};
    assign in3077_2 = {pp68[108],pp65[112],pp62[116],pp62[117]};
    CLA_4 KS_3077(s3077, c3077, in3077_1, in3077_2);
    wire[3:0] s3078, in3078_1, in3078_2;
    wire c3078;
    assign in3078_1 = {pp69[107],pp66[111],pp63[115],pp63[116]};
    assign in3078_2 = {pp70[106],pp67[110],pp64[114],pp64[115]};
    CLA_4 KS_3078(s3078, c3078, in3078_1, in3078_2);
    wire[3:0] s3079, in3079_1, in3079_2;
    wire c3079;
    assign in3079_1 = {pp71[105],pp68[109],pp65[113],pp65[114]};
    assign in3079_2 = {pp72[104],pp69[108],pp66[112],pp66[113]};
    CLA_4 KS_3079(s3079, c3079, in3079_1, in3079_2);
    wire[3:0] s3080, in3080_1, in3080_2;
    wire c3080;
    assign in3080_1 = {pp73[103],pp70[107],pp67[111],pp67[112]};
    assign in3080_2 = {pp74[102],pp71[106],pp68[110],pp68[111]};
    CLA_4 KS_3080(s3080, c3080, in3080_1, in3080_2);
    wire[3:0] s3081, in3081_1, in3081_2;
    wire c3081;
    assign in3081_1 = {pp75[101],pp72[105],pp69[109],pp69[110]};
    assign in3081_2 = {pp76[100],pp73[104],pp70[108],pp70[109]};
    CLA_4 KS_3081(s3081, c3081, in3081_1, in3081_2);
    wire[3:0] s3082, in3082_1, in3082_2;
    wire c3082;
    assign in3082_1 = {pp77[99],pp74[103],pp71[107],pp71[108]};
    assign in3082_2 = {pp78[98],pp75[102],pp72[106],pp72[107]};
    CLA_4 KS_3082(s3082, c3082, in3082_1, in3082_2);
    wire[3:0] s3083, in3083_1, in3083_2;
    wire c3083;
    assign in3083_1 = {pp79[97],pp76[101],pp73[105],pp73[106]};
    assign in3083_2 = {pp80[96],pp77[100],pp74[104],pp74[105]};
    CLA_4 KS_3083(s3083, c3083, in3083_1, in3083_2);
    wire[3:0] s3084, in3084_1, in3084_2;
    wire c3084;
    assign in3084_1 = {pp81[95],pp78[99],pp75[103],pp75[104]};
    assign in3084_2 = {pp82[94],pp79[98],pp76[102],pp76[103]};
    CLA_4 KS_3084(s3084, c3084, in3084_1, in3084_2);
    wire[3:0] s3085, in3085_1, in3085_2;
    wire c3085;
    assign in3085_1 = {pp83[93],pp80[97],pp77[101],pp77[102]};
    assign in3085_2 = {pp84[92],pp81[96],pp78[100],pp78[101]};
    CLA_4 KS_3085(s3085, c3085, in3085_1, in3085_2);
    wire[3:0] s3086, in3086_1, in3086_2;
    wire c3086;
    assign in3086_1 = {pp85[91],pp82[95],pp79[99],pp79[100]};
    assign in3086_2 = {pp86[90],pp83[94],pp80[98],pp80[99]};
    CLA_4 KS_3086(s3086, c3086, in3086_1, in3086_2);
    wire[3:0] s3087, in3087_1, in3087_2;
    wire c3087;
    assign in3087_1 = {pp87[89],pp84[93],pp81[97],pp81[98]};
    assign in3087_2 = {pp88[88],pp85[92],pp82[96],pp82[97]};
    CLA_4 KS_3087(s3087, c3087, in3087_1, in3087_2);
    wire[3:0] s3088, in3088_1, in3088_2;
    wire c3088;
    assign in3088_1 = {pp89[87],pp86[91],pp83[95],pp83[96]};
    assign in3088_2 = {pp90[86],pp87[90],pp84[94],pp84[95]};
    CLA_4 KS_3088(s3088, c3088, in3088_1, in3088_2);
    wire[3:0] s3089, in3089_1, in3089_2;
    wire c3089;
    assign in3089_1 = {pp91[85],pp88[89],pp85[93],pp85[94]};
    assign in3089_2 = {pp92[84],pp89[88],pp86[92],pp86[93]};
    CLA_4 KS_3089(s3089, c3089, in3089_1, in3089_2);
    wire[3:0] s3090, in3090_1, in3090_2;
    wire c3090;
    assign in3090_1 = {pp93[83],pp90[87],pp87[91],pp87[92]};
    assign in3090_2 = {pp94[82],pp91[86],pp88[90],pp88[91]};
    CLA_4 KS_3090(s3090, c3090, in3090_1, in3090_2);
    wire[3:0] s3091, in3091_1, in3091_2;
    wire c3091;
    assign in3091_1 = {pp95[81],pp92[85],pp89[89],pp89[90]};
    assign in3091_2 = {pp96[80],pp93[84],pp90[88],pp90[89]};
    CLA_4 KS_3091(s3091, c3091, in3091_1, in3091_2);
    wire[3:0] s3092, in3092_1, in3092_2;
    wire c3092;
    assign in3092_1 = {pp97[79],pp94[83],pp91[87],pp91[88]};
    assign in3092_2 = {pp98[78],pp95[82],pp92[86],pp92[87]};
    CLA_4 KS_3092(s3092, c3092, in3092_1, in3092_2);
    wire[3:0] s3093, in3093_1, in3093_2;
    wire c3093;
    assign in3093_1 = {pp99[77],pp96[81],pp93[85],pp93[86]};
    assign in3093_2 = {pp100[76],pp97[80],pp94[84],pp94[85]};
    CLA_4 KS_3093(s3093, c3093, in3093_1, in3093_2);
    wire[3:0] s3094, in3094_1, in3094_2;
    wire c3094;
    assign in3094_1 = {pp101[75],pp98[79],pp95[83],pp95[84]};
    assign in3094_2 = {pp102[74],pp99[78],pp96[82],pp96[83]};
    CLA_4 KS_3094(s3094, c3094, in3094_1, in3094_2);
    wire[3:0] s3095, in3095_1, in3095_2;
    wire c3095;
    assign in3095_1 = {pp103[73],pp100[77],pp97[81],pp97[82]};
    assign in3095_2 = {pp104[72],pp101[76],pp98[80],pp98[81]};
    CLA_4 KS_3095(s3095, c3095, in3095_1, in3095_2);
    wire[3:0] s3096, in3096_1, in3096_2;
    wire c3096;
    assign in3096_1 = {pp105[71],pp102[75],pp99[79],pp99[80]};
    assign in3096_2 = {pp106[70],pp103[74],pp100[78],pp100[79]};
    CLA_4 KS_3096(s3096, c3096, in3096_1, in3096_2);
    wire[3:0] s3097, in3097_1, in3097_2;
    wire c3097;
    assign in3097_1 = {pp107[69],pp104[73],pp101[77],pp101[78]};
    assign in3097_2 = {pp108[68],pp105[72],pp102[76],pp102[77]};
    CLA_4 KS_3097(s3097, c3097, in3097_1, in3097_2);
    wire[3:0] s3098, in3098_1, in3098_2;
    wire c3098;
    assign in3098_1 = {pp109[67],pp106[71],pp103[75],pp103[76]};
    assign in3098_2 = {pp110[66],pp107[70],pp104[74],pp104[75]};
    CLA_4 KS_3098(s3098, c3098, in3098_1, in3098_2);
    wire[3:0] s3099, in3099_1, in3099_2;
    wire c3099;
    assign in3099_1 = {pp111[65],pp108[69],pp105[73],pp105[74]};
    assign in3099_2 = {pp112[64],pp109[68],pp106[72],pp106[73]};
    CLA_4 KS_3099(s3099, c3099, in3099_1, in3099_2);
    wire[3:0] s3100, in3100_1, in3100_2;
    wire c3100;
    assign in3100_1 = {pp113[63],pp110[67],pp107[71],pp107[72]};
    assign in3100_2 = {pp114[62],pp111[66],pp108[70],pp108[71]};
    CLA_4 KS_3100(s3100, c3100, in3100_1, in3100_2);
    wire[3:0] s3101, in3101_1, in3101_2;
    wire c3101;
    assign in3101_1 = {pp115[61],pp112[65],pp109[69],pp109[70]};
    assign in3101_2 = {pp116[60],pp113[64],pp110[68],pp110[69]};
    CLA_4 KS_3101(s3101, c3101, in3101_1, in3101_2);
    wire[3:0] s3102, in3102_1, in3102_2;
    wire c3102;
    assign in3102_1 = {pp117[59],pp114[63],pp111[67],pp111[68]};
    assign in3102_2 = {pp118[58],pp115[62],pp112[66],pp112[67]};
    CLA_4 KS_3102(s3102, c3102, in3102_1, in3102_2);
    wire[3:0] s3103, in3103_1, in3103_2;
    wire c3103;
    assign in3103_1 = {pp119[57],pp116[61],pp113[65],pp113[66]};
    assign in3103_2 = {pp120[56],pp117[60],pp114[64],pp114[65]};
    CLA_4 KS_3103(s3103, c3103, in3103_1, in3103_2);
    wire[3:0] s3104, in3104_1, in3104_2;
    wire c3104;
    assign in3104_1 = {pp121[55],pp118[59],pp115[63],pp115[64]};
    assign in3104_2 = {pp122[54],pp119[58],pp116[62],pp116[63]};
    CLA_4 KS_3104(s3104, c3104, in3104_1, in3104_2);
    wire[3:0] s3105, in3105_1, in3105_2;
    wire c3105;
    assign in3105_1 = {pp123[53],pp120[57],pp117[61],pp117[62]};
    assign in3105_2 = {pp124[52],pp121[56],pp118[60],pp118[61]};
    CLA_4 KS_3105(s3105, c3105, in3105_1, in3105_2);
    wire[0:0] s3106, in3106_1, in3106_2;
    wire c3106;
    assign in3106_1 = {pp125[51]};
    assign in3106_2 = {pp126[50]};
    Half_Adder KS_3106(s3106, c3106, in3106_1, in3106_2);
    wire[3:0] s3107, in3107_1, in3107_2;
    wire c3107;
    assign in3107_1 = {pp127[49],pp122[55],pp119[59],pp119[60]};
    assign in3107_2 = {s1314[1],pp123[54],pp120[58],pp120[59]};
    CLA_4 KS_3107(s3107, c3107, in3107_1, in3107_2);
    wire[0:0] s3108, in3108_1, in3108_2;
    wire c3108;
    assign in3108_1 = {s1315[1]};
    assign in3108_2 = {s1316[1]};
    Half_Adder KS_3108(s3108, c3108, in3108_1, in3108_2);
    wire[1:0] s3109, in3109_1, in3109_2;
    wire c3109;
    assign in3109_1 = {s1317[1],pp124[53]};
    assign in3109_2 = {c1318,pp125[52]};
    CLA_2 KS_3109(s3109, c3109, in3109_1, in3109_2);
    wire[0:0] s3110, in3110_1, in3110_2;
    wire c3110;
    assign in3110_1 = {s1319[1]};
    assign in3110_2 = {c1320};
    Half_Adder KS_3110(s3110, c3110, in3110_1, in3110_2);
    wire[2:0] s3111, in3111_1, in3111_2;
    wire c3111;
    assign in3111_1 = {s1321[1],pp126[51],pp121[57]};
    assign in3111_2 = {c1322,pp127[50],pp122[56]};
    CLA_3 KS_3111(s3111, c3111, in3111_1, in3111_2);
    wire[0:0] s3112, in3112_1, in3112_2;
    wire c3112;
    assign in3112_1 = {s1323[1]};
    assign in3112_2 = {c1324};
    Half_Adder KS_3112(s3112, c3112, in3112_1, in3112_2);
    wire[1:0] s3113, in3113_1, in3113_2;
    wire c3113;
    assign in3113_1 = {c3009,s1314[2]};
    assign in3113_2 = {c3010,s1315[2]};
    CLA_2 KS_3113(s3113, c3113, in3113_1, in3113_2);
    wire[0:0] s3114, in3114_1, in3114_2;
    wire c3114;
    assign in3114_1 = {c3011};
    assign in3114_2 = {c3012};
    Half_Adder KS_3114(s3114, c3114, in3114_1, in3114_2);
    wire[3:0] s3115, in3115_1, in3115_2;
    wire c3115;
    assign in3115_1 = {c3013,s1316[2],pp123[55],pp121[58]};
    assign in3115_2 = {c3014,c1317,pp124[54],pp122[57]};
    CLA_4 KS_3115(s3115, c3115, in3115_1, in3115_2);
    wire[0:0] s3116, in3116_1, in3116_2;
    wire c3116;
    assign in3116_1 = {c3015};
    assign in3116_2 = {c3016};
    Half_Adder KS_3116(s3116, c3116, in3116_1, in3116_2);
    wire[1:0] s3117, in3117_1, in3117_2;
    wire c3117;
    assign in3117_1 = {c3017,s1319[2]};
    assign in3117_2 = {c3018,c1321};
    CLA_2 KS_3117(s3117, c3117, in3117_1, in3117_2);
    wire[0:0] s3118, in3118_1, in3118_2;
    wire c3118;
    assign in3118_1 = {c3019};
    assign in3118_2 = {c3020};
    Half_Adder KS_3118(s3118, c3118, in3118_1, in3118_2);
    wire[2:0] s3119, in3119_1, in3119_2;
    wire c3119;
    assign in3119_1 = {c3021,s1323[2],pp125[53]};
    assign in3119_2 = {c3022,s3075[1],pp126[52]};
    CLA_3 KS_3119(s3119, c3119, in3119_1, in3119_2);
    wire[0:0] s3120, in3120_1, in3120_2;
    wire c3120;
    assign in3120_1 = {c3023};
    assign in3120_2 = {c3024};
    Half_Adder KS_3120(s3120, c3120, in3120_1, in3120_2);
    wire[1:0] s3121, in3121_1, in3121_2;
    wire c3121;
    assign in3121_1 = {c3025,s3076[1]};
    assign in3121_2 = {c3026,s3077[1]};
    CLA_2 KS_3121(s3121, c3121, in3121_1, in3121_2);
    wire[0:0] s3122, in3122_1, in3122_2;
    wire c3122;
    assign in3122_1 = {c3027};
    assign in3122_2 = {c3028};
    Half_Adder KS_3122(s3122, c3122, in3122_1, in3122_2);
    wire[3:0] s3123, in3123_1, in3123_2;
    wire c3123;
    assign in3123_1 = {c3029,s3078[1],pp127[51],pp123[56]};
    assign in3123_2 = {c3030,s3079[1],s1314[3],pp124[55]};
    CLA_4 KS_3123(s3123, c3123, in3123_1, in3123_2);
    wire[0:0] s3124, in3124_1, in3124_2;
    wire c3124;
    assign in3124_1 = {c3031};
    assign in3124_2 = {c3032};
    Half_Adder KS_3124(s3124, c3124, in3124_1, in3124_2);
    wire[1:0] s3125, in3125_1, in3125_2;
    wire c3125;
    assign in3125_1 = {c3033,s3080[1]};
    assign in3125_2 = {c3034,s3081[1]};
    CLA_2 KS_3125(s3125, c3125, in3125_1, in3125_2);
    wire[0:0] s3126, in3126_1, in3126_2;
    wire c3126;
    assign in3126_1 = {c3035};
    assign in3126_2 = {c3036};
    Half_Adder KS_3126(s3126, c3126, in3126_1, in3126_2);
    wire[2:0] s3127, in3127_1, in3127_2;
    wire c3127;
    assign in3127_1 = {c3037,s3082[1],s1315[3]};
    assign in3127_2 = {c3038,s3083[1],c1316};
    CLA_3 KS_3127(s3127, c3127, in3127_1, in3127_2);
    wire[0:0] s3128, in3128_1, in3128_2;
    wire c3128;
    assign in3128_1 = {c3039};
    assign in3128_2 = {c3043};
    Half_Adder KS_3128(s3128, c3128, in3128_1, in3128_2);
    wire[1:0] s3129, in3129_1, in3129_2;
    wire c3129;
    assign in3129_1 = {c3051,s3084[1]};
    assign in3129_2 = {c3059,s3085[1]};
    CLA_2 KS_3129(s3129, c3129, in3129_1, in3129_2);
    wire[0:0] s3130, in3130_1, in3130_2;
    wire c3130;
    assign in3130_1 = {c3067};
    assign in3130_2 = {s3075[0]};
    Half_Adder KS_3130(s3130, c3130, in3130_1, in3130_2);
    wire[3:0] s3131, in3131_1, in3131_2;
    wire c3131;
    assign in3131_1 = {s3076[0],s3086[1],s1319[3],pp125[54]};
    assign in3131_2 = {s3077[0],s3087[1],c1323,pp126[53]};
    CLA_4 KS_3131(s3131, c3131, in3131_1, in3131_2);
    wire[0:0] s3132, in3132_1, in3132_2;
    wire c3132;
    assign in3132_1 = {s3078[0]};
    assign in3132_2 = {s3079[0]};
    Half_Adder KS_3132(s3132, c3132, in3132_1, in3132_2);
    wire[1:0] s3133, in3133_1, in3133_2;
    wire c3133;
    assign in3133_1 = {s3080[0],s3088[1]};
    assign in3133_2 = {s3081[0],s3089[1]};
    CLA_2 KS_3133(s3133, c3133, in3133_1, in3133_2);
    wire[0:0] s3134, in3134_1, in3134_2;
    wire c3134;
    assign in3134_1 = {s3082[0]};
    assign in3134_2 = {s3083[0]};
    Half_Adder KS_3134(s3134, c3134, in3134_1, in3134_2);
    wire[2:0] s3135, in3135_1, in3135_2;
    wire c3135;
    assign in3135_1 = {s3084[0],s3090[1],s3075[2]};
    assign in3135_2 = {s3085[0],s3091[1],s3076[2]};
    CLA_3 KS_3135(s3135, c3135, in3135_1, in3135_2);
    wire[0:0] s3136, in3136_1, in3136_2;
    wire c3136;
    assign in3136_1 = {s3086[0]};
    assign in3136_2 = {s3087[0]};
    Half_Adder KS_3136(s3136, c3136, in3136_1, in3136_2);
    wire[1:0] s3137, in3137_1, in3137_2;
    wire c3137;
    assign in3137_1 = {s3088[0],s3092[1]};
    assign in3137_2 = {s3089[0],s3093[1]};
    CLA_2 KS_3137(s3137, c3137, in3137_1, in3137_2);
    wire[0:0] s3138, in3138_1, in3138_2;
    wire c3138;
    assign in3138_1 = {s3090[0]};
    assign in3138_2 = {s3091[0]};
    Half_Adder KS_3138(s3138, c3138, in3138_1, in3138_2);
    wire[3:0] s3139, in3139_1, in3139_2;
    wire c3139;
    assign in3139_1 = {s3093[0],s3094[1],s3077[2],pp127[52]};
    assign in3139_2 = {s3094[0],s3095[1],s3078[2],c1314};
    CLA_4_c KS_3139(s3139, c3139, in3139_1, in3139_2, s3092[0]);
    wire[3:0] s3140, in3140_1, in3140_2;
    wire c3140;
    assign in3140_1 = {pp55[125],pp54[127],pp55[127],pp56[127]};
    assign in3140_2 = {pp56[124],pp55[126],pp56[126],pp57[126]};
    CLA_4 KS_3140(s3140, c3140, in3140_1, in3140_2);
    wire[3:0] s3141, in3141_1, in3141_2;
    wire c3141;
    assign in3141_1 = {pp57[123],pp56[125],pp57[125],pp58[125]};
    assign in3141_2 = {pp58[122],pp57[124],pp58[124],pp59[124]};
    CLA_4 KS_3141(s3141, c3141, in3141_1, in3141_2);
    wire[3:0] s3142, in3142_1, in3142_2;
    wire c3142;
    assign in3142_1 = {pp59[121],pp58[123],pp59[123],pp60[123]};
    assign in3142_2 = {pp60[120],pp59[122],pp60[122],pp61[122]};
    CLA_4 KS_3142(s3142, c3142, in3142_1, in3142_2);
    wire[3:0] s3143, in3143_1, in3143_2;
    wire c3143;
    assign in3143_1 = {pp61[119],pp60[121],pp61[121],pp62[121]};
    assign in3143_2 = {pp62[118],pp61[120],pp62[120],pp63[120]};
    CLA_4 KS_3143(s3143, c3143, in3143_1, in3143_2);
    wire[3:0] s3144, in3144_1, in3144_2;
    wire c3144;
    assign in3144_1 = {pp63[117],pp62[119],pp63[119],pp64[119]};
    assign in3144_2 = {pp64[116],pp63[118],pp64[118],pp65[118]};
    CLA_4 KS_3144(s3144, c3144, in3144_1, in3144_2);
    wire[3:0] s3145, in3145_1, in3145_2;
    wire c3145;
    assign in3145_1 = {pp65[115],pp64[117],pp65[117],pp66[117]};
    assign in3145_2 = {pp66[114],pp65[116],pp66[116],pp67[116]};
    CLA_4 KS_3145(s3145, c3145, in3145_1, in3145_2);
    wire[3:0] s3146, in3146_1, in3146_2;
    wire c3146;
    assign in3146_1 = {pp67[113],pp66[115],pp67[115],pp68[115]};
    assign in3146_2 = {pp68[112],pp67[114],pp68[114],pp69[114]};
    CLA_4 KS_3146(s3146, c3146, in3146_1, in3146_2);
    wire[3:0] s3147, in3147_1, in3147_2;
    wire c3147;
    assign in3147_1 = {pp69[111],pp68[113],pp69[113],pp70[113]};
    assign in3147_2 = {pp70[110],pp69[112],pp70[112],pp71[112]};
    CLA_4 KS_3147(s3147, c3147, in3147_1, in3147_2);
    wire[3:0] s3148, in3148_1, in3148_2;
    wire c3148;
    assign in3148_1 = {pp71[109],pp70[111],pp71[111],pp72[111]};
    assign in3148_2 = {pp72[108],pp71[110],pp72[110],pp73[110]};
    CLA_4 KS_3148(s3148, c3148, in3148_1, in3148_2);
    wire[3:0] s3149, in3149_1, in3149_2;
    wire c3149;
    assign in3149_1 = {pp73[107],pp72[109],pp73[109],pp74[109]};
    assign in3149_2 = {pp74[106],pp73[108],pp74[108],pp75[108]};
    CLA_4 KS_3149(s3149, c3149, in3149_1, in3149_2);
    wire[3:0] s3150, in3150_1, in3150_2;
    wire c3150;
    assign in3150_1 = {pp75[105],pp74[107],pp75[107],pp76[107]};
    assign in3150_2 = {pp76[104],pp75[106],pp76[106],pp77[106]};
    CLA_4 KS_3150(s3150, c3150, in3150_1, in3150_2);
    wire[3:0] s3151, in3151_1, in3151_2;
    wire c3151;
    assign in3151_1 = {pp77[103],pp76[105],pp77[105],pp78[105]};
    assign in3151_2 = {pp78[102],pp77[104],pp78[104],pp79[104]};
    CLA_4 KS_3151(s3151, c3151, in3151_1, in3151_2);
    wire[3:0] s3152, in3152_1, in3152_2;
    wire c3152;
    assign in3152_1 = {pp79[101],pp78[103],pp79[103],pp80[103]};
    assign in3152_2 = {pp80[100],pp79[102],pp80[102],pp81[102]};
    CLA_4 KS_3152(s3152, c3152, in3152_1, in3152_2);
    wire[3:0] s3153, in3153_1, in3153_2;
    wire c3153;
    assign in3153_1 = {pp81[99],pp80[101],pp81[101],pp82[101]};
    assign in3153_2 = {pp82[98],pp81[100],pp82[100],pp83[100]};
    CLA_4 KS_3153(s3153, c3153, in3153_1, in3153_2);
    wire[3:0] s3154, in3154_1, in3154_2;
    wire c3154;
    assign in3154_1 = {pp83[97],pp82[99],pp83[99],pp84[99]};
    assign in3154_2 = {pp84[96],pp83[98],pp84[98],pp85[98]};
    CLA_4 KS_3154(s3154, c3154, in3154_1, in3154_2);
    wire[3:0] s3155, in3155_1, in3155_2;
    wire c3155;
    assign in3155_1 = {pp85[95],pp84[97],pp85[97],pp86[97]};
    assign in3155_2 = {pp86[94],pp85[96],pp86[96],pp87[96]};
    CLA_4 KS_3155(s3155, c3155, in3155_1, in3155_2);
    wire[3:0] s3156, in3156_1, in3156_2;
    wire c3156;
    assign in3156_1 = {pp87[93],pp86[95],pp87[95],pp88[95]};
    assign in3156_2 = {pp88[92],pp87[94],pp88[94],pp89[94]};
    CLA_4 KS_3156(s3156, c3156, in3156_1, in3156_2);
    wire[3:0] s3157, in3157_1, in3157_2;
    wire c3157;
    assign in3157_1 = {pp89[91],pp88[93],pp89[93],pp90[93]};
    assign in3157_2 = {pp90[90],pp89[92],pp90[92],pp91[92]};
    CLA_4 KS_3157(s3157, c3157, in3157_1, in3157_2);
    wire[3:0] s3158, in3158_1, in3158_2;
    wire c3158;
    assign in3158_1 = {pp91[89],pp90[91],pp91[91],pp92[91]};
    assign in3158_2 = {pp92[88],pp91[90],pp92[90],pp93[90]};
    CLA_4 KS_3158(s3158, c3158, in3158_1, in3158_2);
    wire[3:0] s3159, in3159_1, in3159_2;
    wire c3159;
    assign in3159_1 = {pp93[87],pp92[89],pp93[89],pp94[89]};
    assign in3159_2 = {pp94[86],pp93[88],pp94[88],pp95[88]};
    CLA_4 KS_3159(s3159, c3159, in3159_1, in3159_2);
    wire[3:0] s3160, in3160_1, in3160_2;
    wire c3160;
    assign in3160_1 = {pp95[85],pp94[87],pp95[87],pp96[87]};
    assign in3160_2 = {pp96[84],pp95[86],pp96[86],pp97[86]};
    CLA_4 KS_3160(s3160, c3160, in3160_1, in3160_2);
    wire[3:0] s3161, in3161_1, in3161_2;
    wire c3161;
    assign in3161_1 = {pp97[83],pp96[85],pp97[85],pp98[85]};
    assign in3161_2 = {pp98[82],pp97[84],pp98[84],pp99[84]};
    CLA_4 KS_3161(s3161, c3161, in3161_1, in3161_2);
    wire[3:0] s3162, in3162_1, in3162_2;
    wire c3162;
    assign in3162_1 = {pp99[81],pp98[83],pp99[83],pp100[83]};
    assign in3162_2 = {pp100[80],pp99[82],pp100[82],pp101[82]};
    CLA_4 KS_3162(s3162, c3162, in3162_1, in3162_2);
    wire[3:0] s3163, in3163_1, in3163_2;
    wire c3163;
    assign in3163_1 = {pp101[79],pp100[81],pp101[81],pp102[81]};
    assign in3163_2 = {pp102[78],pp101[80],pp102[80],pp103[80]};
    CLA_4 KS_3163(s3163, c3163, in3163_1, in3163_2);
    wire[3:0] s3164, in3164_1, in3164_2;
    wire c3164;
    assign in3164_1 = {pp103[77],pp102[79],pp103[79],pp104[79]};
    assign in3164_2 = {pp104[76],pp103[78],pp104[78],pp105[78]};
    CLA_4 KS_3164(s3164, c3164, in3164_1, in3164_2);
    wire[3:0] s3165, in3165_1, in3165_2;
    wire c3165;
    assign in3165_1 = {pp105[75],pp104[77],pp105[77],pp106[77]};
    assign in3165_2 = {pp106[74],pp105[76],pp106[76],pp107[76]};
    CLA_4 KS_3165(s3165, c3165, in3165_1, in3165_2);
    wire[3:0] s3166, in3166_1, in3166_2;
    wire c3166;
    assign in3166_1 = {pp107[73],pp106[75],pp107[75],pp108[75]};
    assign in3166_2 = {pp108[72],pp107[74],pp108[74],pp109[74]};
    CLA_4 KS_3166(s3166, c3166, in3166_1, in3166_2);
    wire[3:0] s3167, in3167_1, in3167_2;
    wire c3167;
    assign in3167_1 = {pp109[71],pp108[73],pp109[73],pp110[73]};
    assign in3167_2 = {pp110[70],pp109[72],pp110[72],pp111[72]};
    CLA_4 KS_3167(s3167, c3167, in3167_1, in3167_2);
    wire[2:0] s3168, in3168_1, in3168_2;
    wire c3168;
    assign in3168_1 = {pp111[69],pp110[71],pp111[71]};
    assign in3168_2 = {pp112[68],pp111[70],pp112[70]};
    CLA_3 KS_3168(s3168, c3168, in3168_1, in3168_2);
    wire[1:0] s3169, in3169_1, in3169_2;
    wire c3169;
    assign in3169_1 = {pp113[67],pp112[69]};
    assign in3169_2 = {pp114[66],pp113[68]};
    CLA_2 KS_3169(s3169, c3169, in3169_1, in3169_2);
    wire[3:0] s3170, in3170_1, in3170_2;
    wire c3170;
    assign in3170_1 = {pp115[65],pp114[67],pp113[69],pp112[71]};
    assign in3170_2 = {pp116[64],pp115[66],pp114[68],pp113[70]};
    CLA_4 KS_3170(s3170, c3170, in3170_1, in3170_2);
    wire[0:0] s3171, in3171_1, in3171_2;
    wire c3171;
    assign in3171_1 = {pp117[63]};
    assign in3171_2 = {pp118[62]};
    Half_Adder KS_3171(s3171, c3171, in3171_1, in3171_2);
    wire[1:0] s3172, in3172_1, in3172_2;
    wire c3172;
    assign in3172_1 = {pp119[61],pp116[65]};
    assign in3172_2 = {pp120[60],pp117[64]};
    CLA_2 KS_3172(s3172, c3172, in3172_1, in3172_2);
    wire[0:0] s3173, in3173_1, in3173_2;
    wire c3173;
    assign in3173_1 = {pp121[59]};
    assign in3173_2 = {pp122[58]};
    Half_Adder KS_3173(s3173, c3173, in3173_1, in3173_2);
    wire[2:0] s3174, in3174_1, in3174_2;
    wire c3174;
    assign in3174_1 = {pp123[57],pp118[63],pp115[67]};
    assign in3174_2 = {pp124[56],pp119[62],pp116[66]};
    CLA_3 KS_3174(s3174, c3174, in3174_1, in3174_2);
    wire[0:0] s3175, in3175_1, in3175_2;
    wire c3175;
    assign in3175_1 = {pp125[55]};
    assign in3175_2 = {pp126[54]};
    Half_Adder KS_3175(s3175, c3175, in3175_1, in3175_2);
    wire[1:0] s3176, in3176_1, in3176_2;
    wire c3176;
    assign in3176_1 = {pp127[53],pp120[61]};
    assign in3176_2 = {c1325,pp121[60]};
    CLA_2 KS_3176(s3176, c3176, in3176_1, in3176_2);
    wire[0:0] s3177, in3177_1, in3177_2;
    wire c3177;
    assign in3177_1 = {s1326[1]};
    assign in3177_2 = {c3075};
    Half_Adder KS_3177(s3177, c3177, in3177_1, in3177_2);
    wire[3:0] s3178, in3178_1, in3178_2;
    wire c3178;
    assign in3178_1 = {c3076,pp122[59],pp117[65],pp114[69]};
    assign in3178_2 = {c3077,pp123[58],pp118[64],pp115[68]};
    CLA_4 KS_3178(s3178, c3178, in3178_1, in3178_2);
    wire[0:0] s3179, in3179_1, in3179_2;
    wire c3179;
    assign in3179_1 = {c3078};
    assign in3179_2 = {c3079};
    Half_Adder KS_3179(s3179, c3179, in3179_1, in3179_2);
    wire[1:0] s3180, in3180_1, in3180_2;
    wire c3180;
    assign in3180_1 = {c3080,pp124[57]};
    assign in3180_2 = {c3081,pp125[56]};
    CLA_2 KS_3180(s3180, c3180, in3180_1, in3180_2);
    wire[0:0] s3181, in3181_1, in3181_2;
    wire c3181;
    assign in3181_1 = {c3082};
    assign in3181_2 = {c3083};
    Half_Adder KS_3181(s3181, c3181, in3181_1, in3181_2);
    wire[2:0] s3182, in3182_1, in3182_2;
    wire c3182;
    assign in3182_1 = {c3084,pp126[55],pp119[63]};
    assign in3182_2 = {c3085,pp127[54],pp120[62]};
    CLA_3 KS_3182(s3182, c3182, in3182_1, in3182_2);
    wire[0:0] s3183, in3183_1, in3183_2;
    wire c3183;
    assign in3183_1 = {c3086};
    assign in3183_2 = {c3087};
    Half_Adder KS_3183(s3183, c3183, in3183_1, in3183_2);
    wire[1:0] s3184, in3184_1, in3184_2;
    wire c3184;
    assign in3184_1 = {c3088,c1326};
    assign in3184_2 = {c3089,s3140[1]};
    CLA_2 KS_3184(s3184, c3184, in3184_1, in3184_2);
    wire[0:0] s3185, in3185_1, in3185_2;
    wire c3185;
    assign in3185_1 = {c3090};
    assign in3185_2 = {c3091};
    Half_Adder KS_3185(s3185, c3185, in3185_1, in3185_2);
    wire[3:0] s3186, in3186_1, in3186_2;
    wire c3186;
    assign in3186_1 = {c3092,s3141[1],pp121[61],pp116[67]};
    assign in3186_2 = {c3093,s3142[1],pp122[60],pp117[66]};
    CLA_4 KS_3186(s3186, c3186, in3186_1, in3186_2);
    wire[0:0] s3187, in3187_1, in3187_2;
    wire c3187;
    assign in3187_1 = {c3094};
    assign in3187_2 = {c3095};
    Half_Adder KS_3187(s3187, c3187, in3187_1, in3187_2);
    wire[1:0] s3188, in3188_1, in3188_2;
    wire c3188;
    assign in3188_1 = {c3096,s3143[1]};
    assign in3188_2 = {c3097,s3144[1]};
    CLA_2 KS_3188(s3188, c3188, in3188_1, in3188_2);
    wire[0:0] s3189, in3189_1, in3189_2;
    wire c3189;
    assign in3189_1 = {c3098};
    assign in3189_2 = {c3099};
    Half_Adder KS_3189(s3189, c3189, in3189_1, in3189_2);
    wire[2:0] s3190, in3190_1, in3190_2;
    wire c3190;
    assign in3190_1 = {c3100,s3145[1],pp123[59]};
    assign in3190_2 = {c3101,s3146[1],pp124[58]};
    CLA_3 KS_3190(s3190, c3190, in3190_1, in3190_2);
    wire[0:0] s3191, in3191_1, in3191_2;
    wire c3191;
    assign in3191_1 = {c3102};
    assign in3191_2 = {c3103};
    Half_Adder KS_3191(s3191, c3191, in3191_1, in3191_2);
    wire[1:0] s3192, in3192_1, in3192_2;
    wire c3192;
    assign in3192_1 = {c3104,s3147[1]};
    assign in3192_2 = {c3105,s3148[1]};
    CLA_2 KS_3192(s3192, c3192, in3192_1, in3192_2);
    wire[0:0] s3193, in3193_1, in3193_2;
    wire c3193;
    assign in3193_1 = {c3107};
    assign in3193_2 = {c3115};
    Half_Adder KS_3193(s3193, c3193, in3193_1, in3193_2);
    wire[3:0] s3194, in3194_1, in3194_2;
    wire c3194;
    assign in3194_1 = {c3123,s3149[1],pp125[57],pp118[65]};
    assign in3194_2 = {c3131,s3150[1],pp126[56],pp119[64]};
    CLA_4 KS_3194(s3194, c3194, in3194_1, in3194_2);
    wire[0:0] s3195, in3195_1, in3195_2;
    wire c3195;
    assign in3195_1 = {c3139};
    assign in3195_2 = {s3140[0]};
    Half_Adder KS_3195(s3195, c3195, in3195_1, in3195_2);
    wire[1:0] s3196, in3196_1, in3196_2;
    wire c3196;
    assign in3196_1 = {s3141[0],s3151[1]};
    assign in3196_2 = {s3142[0],s3152[1]};
    CLA_2 KS_3196(s3196, c3196, in3196_1, in3196_2);
    wire[0:0] s3197, in3197_1, in3197_2;
    wire c3197;
    assign in3197_1 = {s3143[0]};
    assign in3197_2 = {s3144[0]};
    Half_Adder KS_3197(s3197, c3197, in3197_1, in3197_2);
    wire[2:0] s3198, in3198_1, in3198_2;
    wire c3198;
    assign in3198_1 = {s3145[0],s3153[1],pp127[55]};
    assign in3198_2 = {s3146[0],s3154[1],s3140[2]};
    CLA_3 KS_3198(s3198, c3198, in3198_1, in3198_2);
    wire[0:0] s3199, in3199_1, in3199_2;
    wire c3199;
    assign in3199_1 = {s3147[0]};
    assign in3199_2 = {s3148[0]};
    Half_Adder KS_3199(s3199, c3199, in3199_1, in3199_2);
    wire[1:0] s3200, in3200_1, in3200_2;
    wire c3200;
    assign in3200_1 = {s3149[0],s3155[1]};
    assign in3200_2 = {s3150[0],s3156[1]};
    CLA_2 KS_3200(s3200, c3200, in3200_1, in3200_2);
    wire[0:0] s3201, in3201_1, in3201_2;
    wire c3201;
    assign in3201_1 = {s3151[0]};
    assign in3201_2 = {s3152[0]};
    Half_Adder KS_3201(s3201, c3201, in3201_1, in3201_2);
    wire[3:0] s3202, in3202_1, in3202_2;
    wire c3202;
    assign in3202_1 = {s3153[0],s3157[1],s3141[2],pp120[63]};
    assign in3202_2 = {s3154[0],s3158[1],s3142[2],pp121[62]};
    CLA_4 KS_3202(s3202, c3202, in3202_1, in3202_2);
    wire[0:0] s3203, in3203_1, in3203_2;
    wire c3203;
    assign in3203_1 = {s3155[0]};
    assign in3203_2 = {s3156[0]};
    Half_Adder KS_3203(s3203, c3203, in3203_1, in3203_2);
    wire[1:0] s3204, in3204_1, in3204_2;
    wire c3204;
    assign in3204_1 = {s3158[0],s3159[1]};
    assign in3204_2 = {s3159[0],s3160[1]};
    CLA_2_c KS_3204(s3204, c3204, in3204_1, in3204_2, s3157[0]);
    wire[3:0] s3205, in3205_1, in3205_2;
    wire c3205;
    assign in3205_1 = {pp57[127],pp58[127],pp59[127],pp60[127]};
    assign in3205_2 = {pp58[126],pp59[126],pp60[126],pp61[126]};
    CLA_4 KS_3205(s3205, c3205, in3205_1, in3205_2);
    wire[3:0] s3206, in3206_1, in3206_2;
    wire c3206;
    assign in3206_1 = {pp59[125],pp60[125],pp61[125],pp62[125]};
    assign in3206_2 = {pp60[124],pp61[124],pp62[124],pp63[124]};
    CLA_4 KS_3206(s3206, c3206, in3206_1, in3206_2);
    wire[3:0] s3207, in3207_1, in3207_2;
    wire c3207;
    assign in3207_1 = {pp61[123],pp62[123],pp63[123],pp64[123]};
    assign in3207_2 = {pp62[122],pp63[122],pp64[122],pp65[122]};
    CLA_4 KS_3207(s3207, c3207, in3207_1, in3207_2);
    wire[3:0] s3208, in3208_1, in3208_2;
    wire c3208;
    assign in3208_1 = {pp63[121],pp64[121],pp65[121],pp66[121]};
    assign in3208_2 = {pp64[120],pp65[120],pp66[120],pp67[120]};
    CLA_4 KS_3208(s3208, c3208, in3208_1, in3208_2);
    wire[3:0] s3209, in3209_1, in3209_2;
    wire c3209;
    assign in3209_1 = {pp65[119],pp66[119],pp67[119],pp68[119]};
    assign in3209_2 = {pp66[118],pp67[118],pp68[118],pp69[118]};
    CLA_4 KS_3209(s3209, c3209, in3209_1, in3209_2);
    wire[3:0] s3210, in3210_1, in3210_2;
    wire c3210;
    assign in3210_1 = {pp67[117],pp68[117],pp69[117],pp70[117]};
    assign in3210_2 = {pp68[116],pp69[116],pp70[116],pp71[116]};
    CLA_4 KS_3210(s3210, c3210, in3210_1, in3210_2);
    wire[3:0] s3211, in3211_1, in3211_2;
    wire c3211;
    assign in3211_1 = {pp69[115],pp70[115],pp71[115],pp72[115]};
    assign in3211_2 = {pp70[114],pp71[114],pp72[114],pp73[114]};
    CLA_4 KS_3211(s3211, c3211, in3211_1, in3211_2);
    wire[3:0] s3212, in3212_1, in3212_2;
    wire c3212;
    assign in3212_1 = {pp71[113],pp72[113],pp73[113],pp74[113]};
    assign in3212_2 = {pp72[112],pp73[112],pp74[112],pp75[112]};
    CLA_4 KS_3212(s3212, c3212, in3212_1, in3212_2);
    wire[3:0] s3213, in3213_1, in3213_2;
    wire c3213;
    assign in3213_1 = {pp73[111],pp74[111],pp75[111],pp76[111]};
    assign in3213_2 = {pp74[110],pp75[110],pp76[110],pp77[110]};
    CLA_4 KS_3213(s3213, c3213, in3213_1, in3213_2);
    wire[3:0] s3214, in3214_1, in3214_2;
    wire c3214;
    assign in3214_1 = {pp75[109],pp76[109],pp77[109],pp78[109]};
    assign in3214_2 = {pp76[108],pp77[108],pp78[108],pp79[108]};
    CLA_4 KS_3214(s3214, c3214, in3214_1, in3214_2);
    wire[3:0] s3215, in3215_1, in3215_2;
    wire c3215;
    assign in3215_1 = {pp77[107],pp78[107],pp79[107],pp80[107]};
    assign in3215_2 = {pp78[106],pp79[106],pp80[106],pp81[106]};
    CLA_4 KS_3215(s3215, c3215, in3215_1, in3215_2);
    wire[3:0] s3216, in3216_1, in3216_2;
    wire c3216;
    assign in3216_1 = {pp79[105],pp80[105],pp81[105],pp82[105]};
    assign in3216_2 = {pp80[104],pp81[104],pp82[104],pp83[104]};
    CLA_4 KS_3216(s3216, c3216, in3216_1, in3216_2);
    wire[3:0] s3217, in3217_1, in3217_2;
    wire c3217;
    assign in3217_1 = {pp81[103],pp82[103],pp83[103],pp84[103]};
    assign in3217_2 = {pp82[102],pp83[102],pp84[102],pp85[102]};
    CLA_4 KS_3217(s3217, c3217, in3217_1, in3217_2);
    wire[3:0] s3218, in3218_1, in3218_2;
    wire c3218;
    assign in3218_1 = {pp83[101],pp84[101],pp85[101],pp86[101]};
    assign in3218_2 = {pp84[100],pp85[100],pp86[100],pp87[100]};
    CLA_4 KS_3218(s3218, c3218, in3218_1, in3218_2);
    wire[3:0] s3219, in3219_1, in3219_2;
    wire c3219;
    assign in3219_1 = {pp85[99],pp86[99],pp87[99],pp88[99]};
    assign in3219_2 = {pp86[98],pp87[98],pp88[98],pp89[98]};
    CLA_4 KS_3219(s3219, c3219, in3219_1, in3219_2);
    wire[3:0] s3220, in3220_1, in3220_2;
    wire c3220;
    assign in3220_1 = {pp87[97],pp88[97],pp89[97],pp90[97]};
    assign in3220_2 = {pp88[96],pp89[96],pp90[96],pp91[96]};
    CLA_4 KS_3220(s3220, c3220, in3220_1, in3220_2);
    wire[3:0] s3221, in3221_1, in3221_2;
    wire c3221;
    assign in3221_1 = {pp89[95],pp90[95],pp91[95],pp92[95]};
    assign in3221_2 = {pp90[94],pp91[94],pp92[94],pp93[94]};
    CLA_4 KS_3221(s3221, c3221, in3221_1, in3221_2);
    wire[3:0] s3222, in3222_1, in3222_2;
    wire c3222;
    assign in3222_1 = {pp91[93],pp92[93],pp93[93],pp94[93]};
    assign in3222_2 = {pp92[92],pp93[92],pp94[92],pp95[92]};
    CLA_4 KS_3222(s3222, c3222, in3222_1, in3222_2);
    wire[3:0] s3223, in3223_1, in3223_2;
    wire c3223;
    assign in3223_1 = {pp93[91],pp94[91],pp95[91],pp96[91]};
    assign in3223_2 = {pp94[90],pp95[90],pp96[90],pp97[90]};
    CLA_4 KS_3223(s3223, c3223, in3223_1, in3223_2);
    wire[3:0] s3224, in3224_1, in3224_2;
    wire c3224;
    assign in3224_1 = {pp95[89],pp96[89],pp97[89],pp98[89]};
    assign in3224_2 = {pp96[88],pp97[88],pp98[88],pp99[88]};
    CLA_4 KS_3224(s3224, c3224, in3224_1, in3224_2);
    wire[3:0] s3225, in3225_1, in3225_2;
    wire c3225;
    assign in3225_1 = {pp97[87],pp98[87],pp99[87],pp100[87]};
    assign in3225_2 = {pp98[86],pp99[86],pp100[86],pp101[86]};
    CLA_4 KS_3225(s3225, c3225, in3225_1, in3225_2);
    wire[3:0] s3226, in3226_1, in3226_2;
    wire c3226;
    assign in3226_1 = {pp99[85],pp100[85],pp101[85],pp102[85]};
    assign in3226_2 = {pp100[84],pp101[84],pp102[84],pp103[84]};
    CLA_4 KS_3226(s3226, c3226, in3226_1, in3226_2);
    wire[3:0] s3227, in3227_1, in3227_2;
    wire c3227;
    assign in3227_1 = {pp101[83],pp102[83],pp103[83],pp104[83]};
    assign in3227_2 = {pp102[82],pp103[82],pp104[82],pp105[82]};
    CLA_4 KS_3227(s3227, c3227, in3227_1, in3227_2);
    wire[3:0] s3228, in3228_1, in3228_2;
    wire c3228;
    assign in3228_1 = {pp103[81],pp104[81],pp105[81],pp106[81]};
    assign in3228_2 = {pp104[80],pp105[80],pp106[80],pp107[80]};
    CLA_4 KS_3228(s3228, c3228, in3228_1, in3228_2);
    wire[2:0] s3229, in3229_1, in3229_2;
    wire c3229;
    assign in3229_1 = {pp105[79],pp106[79],pp107[79]};
    assign in3229_2 = {pp106[78],pp107[78],pp108[78]};
    CLA_3 KS_3229(s3229, c3229, in3229_1, in3229_2);
    wire[1:0] s3230, in3230_1, in3230_2;
    wire c3230;
    assign in3230_1 = {pp107[77],pp108[77]};
    assign in3230_2 = {pp108[76],pp109[76]};
    CLA_2 KS_3230(s3230, c3230, in3230_1, in3230_2);
    wire[0:0] s3231, in3231_1, in3231_2;
    wire c3231;
    assign in3231_1 = {pp109[75]};
    assign in3231_2 = {pp110[74]};
    Half_Adder KS_3231(s3231, c3231, in3231_1, in3231_2);
    wire[3:0] s3232, in3232_1, in3232_2;
    wire c3232;
    assign in3232_1 = {pp111[73],pp110[75],pp109[77],pp108[79]};
    assign in3232_2 = {pp112[72],pp111[74],pp110[76],pp109[78]};
    CLA_4 KS_3232(s3232, c3232, in3232_1, in3232_2);
    wire[0:0] s3233, in3233_1, in3233_2;
    wire c3233;
    assign in3233_1 = {pp113[71]};
    assign in3233_2 = {pp114[70]};
    Half_Adder KS_3233(s3233, c3233, in3233_1, in3233_2);
    wire[1:0] s3234, in3234_1, in3234_2;
    wire c3234;
    assign in3234_1 = {pp115[69],pp112[73]};
    assign in3234_2 = {pp116[68],pp113[72]};
    CLA_2 KS_3234(s3234, c3234, in3234_1, in3234_2);
    wire[0:0] s3235, in3235_1, in3235_2;
    wire c3235;
    assign in3235_1 = {pp117[67]};
    assign in3235_2 = {pp118[66]};
    Half_Adder KS_3235(s3235, c3235, in3235_1, in3235_2);
    wire[2:0] s3236, in3236_1, in3236_2;
    wire c3236;
    assign in3236_1 = {pp119[65],pp114[71],pp111[75]};
    assign in3236_2 = {pp120[64],pp115[70],pp112[74]};
    CLA_3 KS_3236(s3236, c3236, in3236_1, in3236_2);
    wire[0:0] s3237, in3237_1, in3237_2;
    wire c3237;
    assign in3237_1 = {pp121[63]};
    assign in3237_2 = {pp122[62]};
    Half_Adder KS_3237(s3237, c3237, in3237_1, in3237_2);
    wire[1:0] s3238, in3238_1, in3238_2;
    wire c3238;
    assign in3238_1 = {pp123[61],pp116[69]};
    assign in3238_2 = {pp124[60],pp117[68]};
    CLA_2 KS_3238(s3238, c3238, in3238_1, in3238_2);
    wire[0:0] s3239, in3239_1, in3239_2;
    wire c3239;
    assign in3239_1 = {pp125[59]};
    assign in3239_2 = {pp126[58]};
    Half_Adder KS_3239(s3239, c3239, in3239_1, in3239_2);
    wire[3:0] s3240, in3240_1, in3240_2;
    wire c3240;
    assign in3240_1 = {pp127[57],pp118[67],pp113[73],pp110[77]};
    assign in3240_2 = {c3140,pp119[66],pp114[72],pp111[76]};
    CLA_4 KS_3240(s3240, c3240, in3240_1, in3240_2);
    wire[0:0] s3241, in3241_1, in3241_2;
    wire c3241;
    assign in3241_1 = {c3141};
    assign in3241_2 = {c3142};
    Half_Adder KS_3241(s3241, c3241, in3241_1, in3241_2);
    wire[1:0] s3242, in3242_1, in3242_2;
    wire c3242;
    assign in3242_1 = {c3143,pp120[65]};
    assign in3242_2 = {c3144,pp121[64]};
    CLA_2 KS_3242(s3242, c3242, in3242_1, in3242_2);
    wire[0:0] s3243, in3243_1, in3243_2;
    wire c3243;
    assign in3243_1 = {c3145};
    assign in3243_2 = {c3146};
    Half_Adder KS_3243(s3243, c3243, in3243_1, in3243_2);
    wire[2:0] s3244, in3244_1, in3244_2;
    wire c3244;
    assign in3244_1 = {c3147,pp122[63],pp115[71]};
    assign in3244_2 = {c3148,pp123[62],pp116[70]};
    CLA_3 KS_3244(s3244, c3244, in3244_1, in3244_2);
    wire[0:0] s3245, in3245_1, in3245_2;
    wire c3245;
    assign in3245_1 = {c3149};
    assign in3245_2 = {c3150};
    Half_Adder KS_3245(s3245, c3245, in3245_1, in3245_2);
    wire[1:0] s3246, in3246_1, in3246_2;
    wire c3246;
    assign in3246_1 = {c3151,pp124[61]};
    assign in3246_2 = {c3152,pp125[60]};
    CLA_2 KS_3246(s3246, c3246, in3246_1, in3246_2);
    wire[0:0] s3247, in3247_1, in3247_2;
    wire c3247;
    assign in3247_1 = {c3153};
    assign in3247_2 = {c3154};
    Half_Adder KS_3247(s3247, c3247, in3247_1, in3247_2);
    wire[3:0] s3248, in3248_1, in3248_2;
    wire c3248;
    assign in3248_1 = {c3155,pp126[59],pp117[69],pp112[75]};
    assign in3248_2 = {c3156,pp127[58],pp118[68],pp113[74]};
    CLA_4 KS_3248(s3248, c3248, in3248_1, in3248_2);
    wire[0:0] s3249, in3249_1, in3249_2;
    wire c3249;
    assign in3249_1 = {c3157};
    assign in3249_2 = {c3158};
    Half_Adder KS_3249(s3249, c3249, in3249_1, in3249_2);
    wire[1:0] s3250, in3250_1, in3250_2;
    wire c3250;
    assign in3250_1 = {c3159,s3205[1]};
    assign in3250_2 = {c3160,s3206[1]};
    CLA_2 KS_3250(s3250, c3250, in3250_1, in3250_2);
    wire[0:0] s3251, in3251_1, in3251_2;
    wire c3251;
    assign in3251_1 = {c3161};
    assign in3251_2 = {c3162};
    Half_Adder KS_3251(s3251, c3251, in3251_1, in3251_2);
    wire[2:0] s3252, in3252_1, in3252_2;
    wire c3252;
    assign in3252_1 = {c3163,s3207[1],pp119[67]};
    assign in3252_2 = {c3164,s3208[1],pp120[66]};
    CLA_3 KS_3252(s3252, c3252, in3252_1, in3252_2);
    wire[0:0] s3253, in3253_1, in3253_2;
    wire c3253;
    assign in3253_1 = {c3165};
    assign in3253_2 = {c3166};
    Half_Adder KS_3253(s3253, c3253, in3253_1, in3253_2);
    wire[1:0] s3254, in3254_1, in3254_2;
    wire c3254;
    assign in3254_1 = {c3167,s3209[1]};
    assign in3254_2 = {c3170,s3210[1]};
    CLA_2 KS_3254(s3254, c3254, in3254_1, in3254_2);
    wire[0:0] s3255, in3255_1, in3255_2;
    wire c3255;
    assign in3255_1 = {c3178};
    assign in3255_2 = {c3186};
    Half_Adder KS_3255(s3255, c3255, in3255_1, in3255_2);
    wire[3:0] s3256, in3256_1, in3256_2;
    wire c3256;
    assign in3256_1 = {c3194,s3211[1],pp121[65],pp114[73]};
    assign in3256_2 = {c3202,s3212[1],pp122[64],pp115[72]};
    CLA_4 KS_3256(s3256, c3256, in3256_1, in3256_2);
    wire[0:0] s3257, in3257_1, in3257_2;
    wire c3257;
    assign in3257_1 = {s3205[0]};
    assign in3257_2 = {s3206[0]};
    Half_Adder KS_3257(s3257, c3257, in3257_1, in3257_2);
    wire[1:0] s3258, in3258_1, in3258_2;
    wire c3258;
    assign in3258_1 = {s3207[0],s3213[1]};
    assign in3258_2 = {s3208[0],s3214[1]};
    CLA_2 KS_3258(s3258, c3258, in3258_1, in3258_2);
    wire[0:0] s3259, in3259_1, in3259_2;
    wire c3259;
    assign in3259_1 = {s3209[0]};
    assign in3259_2 = {s3210[0]};
    Half_Adder KS_3259(s3259, c3259, in3259_1, in3259_2);
    wire[2:0] s3260, in3260_1, in3260_2;
    wire c3260;
    assign in3260_1 = {s3211[0],s3215[1],pp123[63]};
    assign in3260_2 = {s3212[0],s3216[1],pp124[62]};
    CLA_3 KS_3260(s3260, c3260, in3260_1, in3260_2);
    wire[0:0] s3261, in3261_1, in3261_2;
    wire c3261;
    assign in3261_1 = {s3213[0]};
    assign in3261_2 = {s3214[0]};
    Half_Adder KS_3261(s3261, c3261, in3261_1, in3261_2);
    wire[1:0] s3262, in3262_1, in3262_2;
    wire c3262;
    assign in3262_1 = {s3216[0],s3217[1]};
    assign in3262_2 = {s3217[0],s3218[1]};
    CLA_2_c KS_3262(s3262, c3262, in3262_1, in3262_2, s3215[0]);
    wire[3:0] s3263, in3263_1, in3263_2;
    wire c3263;
    assign in3263_1 = {pp61[127],pp62[127],pp63[127],pp64[127]};
    assign in3263_2 = {pp62[126],pp63[126],pp64[126],pp65[126]};
    CLA_4 KS_3263(s3263, c3263, in3263_1, in3263_2);
    wire[3:0] s3264, in3264_1, in3264_2;
    wire c3264;
    assign in3264_1 = {pp63[125],pp64[125],pp65[125],pp66[125]};
    assign in3264_2 = {pp64[124],pp65[124],pp66[124],pp67[124]};
    CLA_4 KS_3264(s3264, c3264, in3264_1, in3264_2);
    wire[3:0] s3265, in3265_1, in3265_2;
    wire c3265;
    assign in3265_1 = {pp65[123],pp66[123],pp67[123],pp68[123]};
    assign in3265_2 = {pp66[122],pp67[122],pp68[122],pp69[122]};
    CLA_4 KS_3265(s3265, c3265, in3265_1, in3265_2);
    wire[3:0] s3266, in3266_1, in3266_2;
    wire c3266;
    assign in3266_1 = {pp67[121],pp68[121],pp69[121],pp70[121]};
    assign in3266_2 = {pp68[120],pp69[120],pp70[120],pp71[120]};
    CLA_4 KS_3266(s3266, c3266, in3266_1, in3266_2);
    wire[3:0] s3267, in3267_1, in3267_2;
    wire c3267;
    assign in3267_1 = {pp69[119],pp70[119],pp71[119],pp72[119]};
    assign in3267_2 = {pp70[118],pp71[118],pp72[118],pp73[118]};
    CLA_4 KS_3267(s3267, c3267, in3267_1, in3267_2);
    wire[3:0] s3268, in3268_1, in3268_2;
    wire c3268;
    assign in3268_1 = {pp71[117],pp72[117],pp73[117],pp74[117]};
    assign in3268_2 = {pp72[116],pp73[116],pp74[116],pp75[116]};
    CLA_4 KS_3268(s3268, c3268, in3268_1, in3268_2);
    wire[3:0] s3269, in3269_1, in3269_2;
    wire c3269;
    assign in3269_1 = {pp73[115],pp74[115],pp75[115],pp76[115]};
    assign in3269_2 = {pp74[114],pp75[114],pp76[114],pp77[114]};
    CLA_4 KS_3269(s3269, c3269, in3269_1, in3269_2);
    wire[3:0] s3270, in3270_1, in3270_2;
    wire c3270;
    assign in3270_1 = {pp75[113],pp76[113],pp77[113],pp78[113]};
    assign in3270_2 = {pp76[112],pp77[112],pp78[112],pp79[112]};
    CLA_4 KS_3270(s3270, c3270, in3270_1, in3270_2);
    wire[3:0] s3271, in3271_1, in3271_2;
    wire c3271;
    assign in3271_1 = {pp77[111],pp78[111],pp79[111],pp80[111]};
    assign in3271_2 = {pp78[110],pp79[110],pp80[110],pp81[110]};
    CLA_4 KS_3271(s3271, c3271, in3271_1, in3271_2);
    wire[3:0] s3272, in3272_1, in3272_2;
    wire c3272;
    assign in3272_1 = {pp79[109],pp80[109],pp81[109],pp82[109]};
    assign in3272_2 = {pp80[108],pp81[108],pp82[108],pp83[108]};
    CLA_4 KS_3272(s3272, c3272, in3272_1, in3272_2);
    wire[3:0] s3273, in3273_1, in3273_2;
    wire c3273;
    assign in3273_1 = {pp81[107],pp82[107],pp83[107],pp84[107]};
    assign in3273_2 = {pp82[106],pp83[106],pp84[106],pp85[106]};
    CLA_4 KS_3273(s3273, c3273, in3273_1, in3273_2);
    wire[3:0] s3274, in3274_1, in3274_2;
    wire c3274;
    assign in3274_1 = {pp83[105],pp84[105],pp85[105],pp86[105]};
    assign in3274_2 = {pp84[104],pp85[104],pp86[104],pp87[104]};
    CLA_4 KS_3274(s3274, c3274, in3274_1, in3274_2);
    wire[3:0] s3275, in3275_1, in3275_2;
    wire c3275;
    assign in3275_1 = {pp85[103],pp86[103],pp87[103],pp88[103]};
    assign in3275_2 = {pp86[102],pp87[102],pp88[102],pp89[102]};
    CLA_4 KS_3275(s3275, c3275, in3275_1, in3275_2);
    wire[3:0] s3276, in3276_1, in3276_2;
    wire c3276;
    assign in3276_1 = {pp87[101],pp88[101],pp89[101],pp90[101]};
    assign in3276_2 = {pp88[100],pp89[100],pp90[100],pp91[100]};
    CLA_4 KS_3276(s3276, c3276, in3276_1, in3276_2);
    wire[3:0] s3277, in3277_1, in3277_2;
    wire c3277;
    assign in3277_1 = {pp89[99],pp90[99],pp91[99],pp92[99]};
    assign in3277_2 = {pp90[98],pp91[98],pp92[98],pp93[98]};
    CLA_4 KS_3277(s3277, c3277, in3277_1, in3277_2);
    wire[3:0] s3278, in3278_1, in3278_2;
    wire c3278;
    assign in3278_1 = {pp91[97],pp92[97],pp93[97],pp94[97]};
    assign in3278_2 = {pp92[96],pp93[96],pp94[96],pp95[96]};
    CLA_4 KS_3278(s3278, c3278, in3278_1, in3278_2);
    wire[3:0] s3279, in3279_1, in3279_2;
    wire c3279;
    assign in3279_1 = {pp93[95],pp94[95],pp95[95],pp96[95]};
    assign in3279_2 = {pp94[94],pp95[94],pp96[94],pp97[94]};
    CLA_4 KS_3279(s3279, c3279, in3279_1, in3279_2);
    wire[3:0] s3280, in3280_1, in3280_2;
    wire c3280;
    assign in3280_1 = {pp95[93],pp96[93],pp97[93],pp98[93]};
    assign in3280_2 = {pp96[92],pp97[92],pp98[92],pp99[92]};
    CLA_4 KS_3280(s3280, c3280, in3280_1, in3280_2);
    wire[3:0] s3281, in3281_1, in3281_2;
    wire c3281;
    assign in3281_1 = {pp97[91],pp98[91],pp99[91],pp100[91]};
    assign in3281_2 = {pp98[90],pp99[90],pp100[90],pp101[90]};
    CLA_4 KS_3281(s3281, c3281, in3281_1, in3281_2);
    wire[3:0] s3282, in3282_1, in3282_2;
    wire c3282;
    assign in3282_1 = {pp99[89],pp100[89],pp101[89],pp102[89]};
    assign in3282_2 = {pp100[88],pp101[88],pp102[88],pp103[88]};
    CLA_4 KS_3282(s3282, c3282, in3282_1, in3282_2);
    wire[2:0] s3283, in3283_1, in3283_2;
    wire c3283;
    assign in3283_1 = {pp101[87],pp102[87],pp103[87]};
    assign in3283_2 = {pp102[86],pp103[86],pp104[86]};
    CLA_3 KS_3283(s3283, c3283, in3283_1, in3283_2);
    wire[1:0] s3284, in3284_1, in3284_2;
    wire c3284;
    assign in3284_1 = {pp103[85],pp104[85]};
    assign in3284_2 = {pp104[84],pp105[84]};
    CLA_2 KS_3284(s3284, c3284, in3284_1, in3284_2);
    wire[0:0] s3285, in3285_1, in3285_2;
    wire c3285;
    assign in3285_1 = {pp105[83]};
    assign in3285_2 = {pp106[82]};
    Half_Adder KS_3285(s3285, c3285, in3285_1, in3285_2);
    wire[3:0] s3286, in3286_1, in3286_2;
    wire c3286;
    assign in3286_1 = {pp107[81],pp106[83],pp105[85],pp104[87]};
    assign in3286_2 = {pp108[80],pp107[82],pp106[84],pp105[86]};
    CLA_4 KS_3286(s3286, c3286, in3286_1, in3286_2);
    wire[0:0] s3287, in3287_1, in3287_2;
    wire c3287;
    assign in3287_1 = {pp109[79]};
    assign in3287_2 = {pp110[78]};
    Half_Adder KS_3287(s3287, c3287, in3287_1, in3287_2);
    wire[1:0] s3288, in3288_1, in3288_2;
    wire c3288;
    assign in3288_1 = {pp111[77],pp108[81]};
    assign in3288_2 = {pp112[76],pp109[80]};
    CLA_2 KS_3288(s3288, c3288, in3288_1, in3288_2);
    wire[0:0] s3289, in3289_1, in3289_2;
    wire c3289;
    assign in3289_1 = {pp113[75]};
    assign in3289_2 = {pp114[74]};
    Half_Adder KS_3289(s3289, c3289, in3289_1, in3289_2);
    wire[2:0] s3290, in3290_1, in3290_2;
    wire c3290;
    assign in3290_1 = {pp115[73],pp110[79],pp107[83]};
    assign in3290_2 = {pp116[72],pp111[78],pp108[82]};
    CLA_3 KS_3290(s3290, c3290, in3290_1, in3290_2);
    wire[0:0] s3291, in3291_1, in3291_2;
    wire c3291;
    assign in3291_1 = {pp117[71]};
    assign in3291_2 = {pp118[70]};
    Half_Adder KS_3291(s3291, c3291, in3291_1, in3291_2);
    wire[1:0] s3292, in3292_1, in3292_2;
    wire c3292;
    assign in3292_1 = {pp119[69],pp112[77]};
    assign in3292_2 = {pp120[68],pp113[76]};
    CLA_2 KS_3292(s3292, c3292, in3292_1, in3292_2);
    wire[0:0] s3293, in3293_1, in3293_2;
    wire c3293;
    assign in3293_1 = {pp121[67]};
    assign in3293_2 = {pp122[66]};
    Half_Adder KS_3293(s3293, c3293, in3293_1, in3293_2);
    wire[3:0] s3294, in3294_1, in3294_2;
    wire c3294;
    assign in3294_1 = {pp123[65],pp114[75],pp109[81],pp106[85]};
    assign in3294_2 = {pp124[64],pp115[74],pp110[80],pp107[84]};
    CLA_4 KS_3294(s3294, c3294, in3294_1, in3294_2);
    wire[0:0] s3295, in3295_1, in3295_2;
    wire c3295;
    assign in3295_1 = {pp125[63]};
    assign in3295_2 = {pp126[62]};
    Half_Adder KS_3295(s3295, c3295, in3295_1, in3295_2);
    wire[1:0] s3296, in3296_1, in3296_2;
    wire c3296;
    assign in3296_1 = {pp127[61],pp116[73]};
    assign in3296_2 = {c3205,pp117[72]};
    CLA_2 KS_3296(s3296, c3296, in3296_1, in3296_2);
    wire[0:0] s3297, in3297_1, in3297_2;
    wire c3297;
    assign in3297_1 = {c3206};
    assign in3297_2 = {c3207};
    Half_Adder KS_3297(s3297, c3297, in3297_1, in3297_2);
    wire[2:0] s3298, in3298_1, in3298_2;
    wire c3298;
    assign in3298_1 = {c3208,pp118[71],pp111[79]};
    assign in3298_2 = {c3209,pp119[70],pp112[78]};
    CLA_3 KS_3298(s3298, c3298, in3298_1, in3298_2);
    wire[0:0] s3299, in3299_1, in3299_2;
    wire c3299;
    assign in3299_1 = {c3210};
    assign in3299_2 = {c3211};
    Half_Adder KS_3299(s3299, c3299, in3299_1, in3299_2);
    wire[1:0] s3300, in3300_1, in3300_2;
    wire c3300;
    assign in3300_1 = {c3212,pp120[69]};
    assign in3300_2 = {c3213,pp121[68]};
    CLA_2 KS_3300(s3300, c3300, in3300_1, in3300_2);
    wire[0:0] s3301, in3301_1, in3301_2;
    wire c3301;
    assign in3301_1 = {c3214};
    assign in3301_2 = {c3215};
    Half_Adder KS_3301(s3301, c3301, in3301_1, in3301_2);
    wire[3:0] s3302, in3302_1, in3302_2;
    wire c3302;
    assign in3302_1 = {c3216,pp122[67],pp113[77],pp108[83]};
    assign in3302_2 = {c3217,pp123[66],pp114[76],pp109[82]};
    CLA_4 KS_3302(s3302, c3302, in3302_1, in3302_2);
    wire[0:0] s3303, in3303_1, in3303_2;
    wire c3303;
    assign in3303_1 = {c3218};
    assign in3303_2 = {c3219};
    Half_Adder KS_3303(s3303, c3303, in3303_1, in3303_2);
    wire[1:0] s3304, in3304_1, in3304_2;
    wire c3304;
    assign in3304_1 = {c3220,pp124[65]};
    assign in3304_2 = {c3221,pp125[64]};
    CLA_2 KS_3304(s3304, c3304, in3304_1, in3304_2);
    wire[0:0] s3305, in3305_1, in3305_2;
    wire c3305;
    assign in3305_1 = {c3222};
    assign in3305_2 = {c3223};
    Half_Adder KS_3305(s3305, c3305, in3305_1, in3305_2);
    wire[2:0] s3306, in3306_1, in3306_2;
    wire c3306;
    assign in3306_1 = {c3224,pp126[63],pp115[75]};
    assign in3306_2 = {c3225,pp127[62],pp116[74]};
    CLA_3 KS_3306(s3306, c3306, in3306_1, in3306_2);
    wire[0:0] s3307, in3307_1, in3307_2;
    wire c3307;
    assign in3307_1 = {c3226};
    assign in3307_2 = {c3227};
    Half_Adder KS_3307(s3307, c3307, in3307_1, in3307_2);
    wire[1:0] s3308, in3308_1, in3308_2;
    wire c3308;
    assign in3308_1 = {c3228,s3263[1]};
    assign in3308_2 = {c3232,s3264[1]};
    CLA_2 KS_3308(s3308, c3308, in3308_1, in3308_2);
    wire[0:0] s3309, in3309_1, in3309_2;
    wire c3309;
    assign in3309_1 = {c3240};
    assign in3309_2 = {c3248};
    Half_Adder KS_3309(s3309, c3309, in3309_1, in3309_2);
    wire[3:0] s3310, in3310_1, in3310_2;
    wire c3310;
    assign in3310_1 = {c3256,s3265[1],pp117[73],pp110[81]};
    assign in3310_2 = {s3263[0],s3266[1],pp118[72],pp111[80]};
    CLA_4 KS_3310(s3310, c3310, in3310_1, in3310_2);
    wire[0:0] s3311, in3311_1, in3311_2;
    wire c3311;
    assign in3311_1 = {s3265[0]};
    assign in3311_2 = {s3266[0]};
    Full_Adder KS_3311(s3311, c3311, in3311_1, in3311_2, s3264[0]);
    wire[3:0] s3312, in3312_1, in3312_2;
    wire c3312;
    assign in3312_1 = {pp65[127],pp66[127],pp67[127],pp68[127]};
    assign in3312_2 = {pp66[126],pp67[126],pp68[126],pp69[126]};
    CLA_4 KS_3312(s3312, c3312, in3312_1, in3312_2);
    wire[3:0] s3313, in3313_1, in3313_2;
    wire c3313;
    assign in3313_1 = {pp67[125],pp68[125],pp69[125],pp70[125]};
    assign in3313_2 = {pp68[124],pp69[124],pp70[124],pp71[124]};
    CLA_4 KS_3313(s3313, c3313, in3313_1, in3313_2);
    wire[3:0] s3314, in3314_1, in3314_2;
    wire c3314;
    assign in3314_1 = {pp69[123],pp70[123],pp71[123],pp72[123]};
    assign in3314_2 = {pp70[122],pp71[122],pp72[122],pp73[122]};
    CLA_4 KS_3314(s3314, c3314, in3314_1, in3314_2);
    wire[3:0] s3315, in3315_1, in3315_2;
    wire c3315;
    assign in3315_1 = {pp71[121],pp72[121],pp73[121],pp74[121]};
    assign in3315_2 = {pp72[120],pp73[120],pp74[120],pp75[120]};
    CLA_4 KS_3315(s3315, c3315, in3315_1, in3315_2);
    wire[3:0] s3316, in3316_1, in3316_2;
    wire c3316;
    assign in3316_1 = {pp73[119],pp74[119],pp75[119],pp76[119]};
    assign in3316_2 = {pp74[118],pp75[118],pp76[118],pp77[118]};
    CLA_4 KS_3316(s3316, c3316, in3316_1, in3316_2);
    wire[3:0] s3317, in3317_1, in3317_2;
    wire c3317;
    assign in3317_1 = {pp75[117],pp76[117],pp77[117],pp78[117]};
    assign in3317_2 = {pp76[116],pp77[116],pp78[116],pp79[116]};
    CLA_4 KS_3317(s3317, c3317, in3317_1, in3317_2);
    wire[3:0] s3318, in3318_1, in3318_2;
    wire c3318;
    assign in3318_1 = {pp77[115],pp78[115],pp79[115],pp80[115]};
    assign in3318_2 = {pp78[114],pp79[114],pp80[114],pp81[114]};
    CLA_4 KS_3318(s3318, c3318, in3318_1, in3318_2);
    wire[3:0] s3319, in3319_1, in3319_2;
    wire c3319;
    assign in3319_1 = {pp79[113],pp80[113],pp81[113],pp82[113]};
    assign in3319_2 = {pp80[112],pp81[112],pp82[112],pp83[112]};
    CLA_4 KS_3319(s3319, c3319, in3319_1, in3319_2);
    wire[3:0] s3320, in3320_1, in3320_2;
    wire c3320;
    assign in3320_1 = {pp81[111],pp82[111],pp83[111],pp84[111]};
    assign in3320_2 = {pp82[110],pp83[110],pp84[110],pp85[110]};
    CLA_4 KS_3320(s3320, c3320, in3320_1, in3320_2);
    wire[3:0] s3321, in3321_1, in3321_2;
    wire c3321;
    assign in3321_1 = {pp83[109],pp84[109],pp85[109],pp86[109]};
    assign in3321_2 = {pp84[108],pp85[108],pp86[108],pp87[108]};
    CLA_4 KS_3321(s3321, c3321, in3321_1, in3321_2);
    wire[3:0] s3322, in3322_1, in3322_2;
    wire c3322;
    assign in3322_1 = {pp85[107],pp86[107],pp87[107],pp88[107]};
    assign in3322_2 = {pp86[106],pp87[106],pp88[106],pp89[106]};
    CLA_4 KS_3322(s3322, c3322, in3322_1, in3322_2);
    wire[3:0] s3323, in3323_1, in3323_2;
    wire c3323;
    assign in3323_1 = {pp87[105],pp88[105],pp89[105],pp90[105]};
    assign in3323_2 = {pp88[104],pp89[104],pp90[104],pp91[104]};
    CLA_4 KS_3323(s3323, c3323, in3323_1, in3323_2);
    wire[3:0] s3324, in3324_1, in3324_2;
    wire c3324;
    assign in3324_1 = {pp89[103],pp90[103],pp91[103],pp92[103]};
    assign in3324_2 = {pp90[102],pp91[102],pp92[102],pp93[102]};
    CLA_4 KS_3324(s3324, c3324, in3324_1, in3324_2);
    wire[3:0] s3325, in3325_1, in3325_2;
    wire c3325;
    assign in3325_1 = {pp91[101],pp92[101],pp93[101],pp94[101]};
    assign in3325_2 = {pp92[100],pp93[100],pp94[100],pp95[100]};
    CLA_4 KS_3325(s3325, c3325, in3325_1, in3325_2);
    wire[3:0] s3326, in3326_1, in3326_2;
    wire c3326;
    assign in3326_1 = {pp93[99],pp94[99],pp95[99],pp96[99]};
    assign in3326_2 = {pp94[98],pp95[98],pp96[98],pp97[98]};
    CLA_4 KS_3326(s3326, c3326, in3326_1, in3326_2);
    wire[3:0] s3327, in3327_1, in3327_2;
    wire c3327;
    assign in3327_1 = {pp95[97],pp96[97],pp97[97],pp98[97]};
    assign in3327_2 = {pp96[96],pp97[96],pp98[96],pp99[96]};
    CLA_4 KS_3327(s3327, c3327, in3327_1, in3327_2);
    wire[2:0] s3328, in3328_1, in3328_2;
    wire c3328;
    assign in3328_1 = {pp97[95],pp98[95],pp99[95]};
    assign in3328_2 = {pp98[94],pp99[94],pp100[94]};
    CLA_3 KS_3328(s3328, c3328, in3328_1, in3328_2);
    wire[1:0] s3329, in3329_1, in3329_2;
    wire c3329;
    assign in3329_1 = {pp99[93],pp100[93]};
    assign in3329_2 = {pp100[92],pp101[92]};
    CLA_2 KS_3329(s3329, c3329, in3329_1, in3329_2);
    wire[0:0] s3330, in3330_1, in3330_2;
    wire c3330;
    assign in3330_1 = {pp101[91]};
    assign in3330_2 = {pp102[90]};
    Half_Adder KS_3330(s3330, c3330, in3330_1, in3330_2);
    wire[3:0] s3331, in3331_1, in3331_2;
    wire c3331;
    assign in3331_1 = {pp103[89],pp102[91],pp101[93],pp100[95]};
    assign in3331_2 = {pp104[88],pp103[90],pp102[92],pp101[94]};
    CLA_4 KS_3331(s3331, c3331, in3331_1, in3331_2);
    wire[0:0] s3332, in3332_1, in3332_2;
    wire c3332;
    assign in3332_1 = {pp105[87]};
    assign in3332_2 = {pp106[86]};
    Half_Adder KS_3332(s3332, c3332, in3332_1, in3332_2);
    wire[1:0] s3333, in3333_1, in3333_2;
    wire c3333;
    assign in3333_1 = {pp107[85],pp104[89]};
    assign in3333_2 = {pp108[84],pp105[88]};
    CLA_2 KS_3333(s3333, c3333, in3333_1, in3333_2);
    wire[0:0] s3334, in3334_1, in3334_2;
    wire c3334;
    assign in3334_1 = {pp109[83]};
    assign in3334_2 = {pp110[82]};
    Half_Adder KS_3334(s3334, c3334, in3334_1, in3334_2);
    wire[2:0] s3335, in3335_1, in3335_2;
    wire c3335;
    assign in3335_1 = {pp111[81],pp106[87],pp103[91]};
    assign in3335_2 = {pp112[80],pp107[86],pp104[90]};
    CLA_3 KS_3335(s3335, c3335, in3335_1, in3335_2);
    wire[0:0] s3336, in3336_1, in3336_2;
    wire c3336;
    assign in3336_1 = {pp113[79]};
    assign in3336_2 = {pp114[78]};
    Half_Adder KS_3336(s3336, c3336, in3336_1, in3336_2);
    wire[1:0] s3337, in3337_1, in3337_2;
    wire c3337;
    assign in3337_1 = {pp115[77],pp108[85]};
    assign in3337_2 = {pp116[76],pp109[84]};
    CLA_2 KS_3337(s3337, c3337, in3337_1, in3337_2);
    wire[0:0] s3338, in3338_1, in3338_2;
    wire c3338;
    assign in3338_1 = {pp117[75]};
    assign in3338_2 = {pp118[74]};
    Half_Adder KS_3338(s3338, c3338, in3338_1, in3338_2);
    wire[3:0] s3339, in3339_1, in3339_2;
    wire c3339;
    assign in3339_1 = {pp119[73],pp110[83],pp105[89],pp102[93]};
    assign in3339_2 = {pp120[72],pp111[82],pp106[88],pp103[92]};
    CLA_4 KS_3339(s3339, c3339, in3339_1, in3339_2);
    wire[0:0] s3340, in3340_1, in3340_2;
    wire c3340;
    assign in3340_1 = {pp121[71]};
    assign in3340_2 = {pp122[70]};
    Half_Adder KS_3340(s3340, c3340, in3340_1, in3340_2);
    wire[1:0] s3341, in3341_1, in3341_2;
    wire c3341;
    assign in3341_1 = {pp123[69],pp112[81]};
    assign in3341_2 = {pp124[68],pp113[80]};
    CLA_2 KS_3341(s3341, c3341, in3341_1, in3341_2);
    wire[0:0] s3342, in3342_1, in3342_2;
    wire c3342;
    assign in3342_1 = {pp125[67]};
    assign in3342_2 = {pp126[66]};
    Half_Adder KS_3342(s3342, c3342, in3342_1, in3342_2);
    wire[2:0] s3343, in3343_1, in3343_2;
    wire c3343;
    assign in3343_1 = {pp127[65],pp114[79],pp107[87]};
    assign in3343_2 = {c3263,pp115[78],pp108[86]};
    CLA_3 KS_3343(s3343, c3343, in3343_1, in3343_2);
    wire[0:0] s3344, in3344_1, in3344_2;
    wire c3344;
    assign in3344_1 = {c3264};
    assign in3344_2 = {c3265};
    Half_Adder KS_3344(s3344, c3344, in3344_1, in3344_2);
    wire[1:0] s3345, in3345_1, in3345_2;
    wire c3345;
    assign in3345_1 = {c3266,pp116[77]};
    assign in3345_2 = {c3267,pp117[76]};
    CLA_2 KS_3345(s3345, c3345, in3345_1, in3345_2);
    wire[0:0] s3346, in3346_1, in3346_2;
    wire c3346;
    assign in3346_1 = {c3268};
    assign in3346_2 = {c3269};
    Half_Adder KS_3346(s3346, c3346, in3346_1, in3346_2);
    wire[3:0] s3347, in3347_1, in3347_2;
    wire c3347;
    assign in3347_1 = {c3270,pp118[75],pp109[85],pp104[91]};
    assign in3347_2 = {c3271,pp119[74],pp110[84],pp105[90]};
    CLA_4 KS_3347(s3347, c3347, in3347_1, in3347_2);
    wire[0:0] s3348, in3348_1, in3348_2;
    wire c3348;
    assign in3348_1 = {c3272};
    assign in3348_2 = {c3273};
    Half_Adder KS_3348(s3348, c3348, in3348_1, in3348_2);
    wire[1:0] s3349, in3349_1, in3349_2;
    wire c3349;
    assign in3349_1 = {c3274,pp120[73]};
    assign in3349_2 = {c3275,pp121[72]};
    CLA_2 KS_3349(s3349, c3349, in3349_1, in3349_2);
    wire[0:0] s3350, in3350_1, in3350_2;
    wire c3350;
    assign in3350_1 = {c3276};
    assign in3350_2 = {c3277};
    Half_Adder KS_3350(s3350, c3350, in3350_1, in3350_2);
    wire[2:0] s3351, in3351_1, in3351_2;
    wire c3351;
    assign in3351_1 = {c3278,pp122[71],pp111[83]};
    assign in3351_2 = {c3279,pp123[70],pp112[82]};
    CLA_3 KS_3351(s3351, c3351, in3351_1, in3351_2);
    wire[0:0] s3352, in3352_1, in3352_2;
    wire c3352;
    assign in3352_1 = {c3281};
    assign in3352_2 = {c3282};
    Full_Adder KS_3352(s3352, c3352, in3352_1, in3352_2, c3280);
    wire[3:0] s3353, in3353_1, in3353_2;
    wire c3353;
    assign in3353_1 = {pp69[127],pp70[127],pp71[127],pp72[127]};
    assign in3353_2 = {pp70[126],pp71[126],pp72[126],pp73[126]};
    CLA_4 KS_3353(s3353, c3353, in3353_1, in3353_2);
    wire[3:0] s3354, in3354_1, in3354_2;
    wire c3354;
    assign in3354_1 = {pp71[125],pp72[125],pp73[125],pp74[125]};
    assign in3354_2 = {pp72[124],pp73[124],pp74[124],pp75[124]};
    CLA_4 KS_3354(s3354, c3354, in3354_1, in3354_2);
    wire[3:0] s3355, in3355_1, in3355_2;
    wire c3355;
    assign in3355_1 = {pp73[123],pp74[123],pp75[123],pp76[123]};
    assign in3355_2 = {pp74[122],pp75[122],pp76[122],pp77[122]};
    CLA_4 KS_3355(s3355, c3355, in3355_1, in3355_2);
    wire[3:0] s3356, in3356_1, in3356_2;
    wire c3356;
    assign in3356_1 = {pp75[121],pp76[121],pp77[121],pp78[121]};
    assign in3356_2 = {pp76[120],pp77[120],pp78[120],pp79[120]};
    CLA_4 KS_3356(s3356, c3356, in3356_1, in3356_2);
    wire[3:0] s3357, in3357_1, in3357_2;
    wire c3357;
    assign in3357_1 = {pp77[119],pp78[119],pp79[119],pp80[119]};
    assign in3357_2 = {pp78[118],pp79[118],pp80[118],pp81[118]};
    CLA_4 KS_3357(s3357, c3357, in3357_1, in3357_2);
    wire[3:0] s3358, in3358_1, in3358_2;
    wire c3358;
    assign in3358_1 = {pp79[117],pp80[117],pp81[117],pp82[117]};
    assign in3358_2 = {pp80[116],pp81[116],pp82[116],pp83[116]};
    CLA_4 KS_3358(s3358, c3358, in3358_1, in3358_2);
    wire[3:0] s3359, in3359_1, in3359_2;
    wire c3359;
    assign in3359_1 = {pp81[115],pp82[115],pp83[115],pp84[115]};
    assign in3359_2 = {pp82[114],pp83[114],pp84[114],pp85[114]};
    CLA_4 KS_3359(s3359, c3359, in3359_1, in3359_2);
    wire[3:0] s3360, in3360_1, in3360_2;
    wire c3360;
    assign in3360_1 = {pp83[113],pp84[113],pp85[113],pp86[113]};
    assign in3360_2 = {pp84[112],pp85[112],pp86[112],pp87[112]};
    CLA_4 KS_3360(s3360, c3360, in3360_1, in3360_2);
    wire[3:0] s3361, in3361_1, in3361_2;
    wire c3361;
    assign in3361_1 = {pp85[111],pp86[111],pp87[111],pp88[111]};
    assign in3361_2 = {pp86[110],pp87[110],pp88[110],pp89[110]};
    CLA_4 KS_3361(s3361, c3361, in3361_1, in3361_2);
    wire[3:0] s3362, in3362_1, in3362_2;
    wire c3362;
    assign in3362_1 = {pp87[109],pp88[109],pp89[109],pp90[109]};
    assign in3362_2 = {pp88[108],pp89[108],pp90[108],pp91[108]};
    CLA_4 KS_3362(s3362, c3362, in3362_1, in3362_2);
    wire[3:0] s3363, in3363_1, in3363_2;
    wire c3363;
    assign in3363_1 = {pp89[107],pp90[107],pp91[107],pp92[107]};
    assign in3363_2 = {pp90[106],pp91[106],pp92[106],pp93[106]};
    CLA_4 KS_3363(s3363, c3363, in3363_1, in3363_2);
    wire[3:0] s3364, in3364_1, in3364_2;
    wire c3364;
    assign in3364_1 = {pp91[105],pp92[105],pp93[105],pp94[105]};
    assign in3364_2 = {pp92[104],pp93[104],pp94[104],pp95[104]};
    CLA_4 KS_3364(s3364, c3364, in3364_1, in3364_2);
    wire[2:0] s3365, in3365_1, in3365_2;
    wire c3365;
    assign in3365_1 = {pp93[103],pp94[103],pp95[103]};
    assign in3365_2 = {pp94[102],pp95[102],pp96[102]};
    CLA_3 KS_3365(s3365, c3365, in3365_1, in3365_2);
    wire[1:0] s3366, in3366_1, in3366_2;
    wire c3366;
    assign in3366_1 = {pp95[101],pp96[101]};
    assign in3366_2 = {pp96[100],pp97[100]};
    CLA_2 KS_3366(s3366, c3366, in3366_1, in3366_2);
    wire[0:0] s3367, in3367_1, in3367_2;
    wire c3367;
    assign in3367_1 = {pp97[99]};
    assign in3367_2 = {pp98[98]};
    Half_Adder KS_3367(s3367, c3367, in3367_1, in3367_2);
    wire[3:0] s3368, in3368_1, in3368_2;
    wire c3368;
    assign in3368_1 = {pp99[97],pp98[99],pp97[101],pp96[103]};
    assign in3368_2 = {pp100[96],pp99[98],pp98[100],pp97[102]};
    CLA_4 KS_3368(s3368, c3368, in3368_1, in3368_2);
    wire[0:0] s3369, in3369_1, in3369_2;
    wire c3369;
    assign in3369_1 = {pp101[95]};
    assign in3369_2 = {pp102[94]};
    Half_Adder KS_3369(s3369, c3369, in3369_1, in3369_2);
    wire[1:0] s3370, in3370_1, in3370_2;
    wire c3370;
    assign in3370_1 = {pp103[93],pp100[97]};
    assign in3370_2 = {pp104[92],pp101[96]};
    CLA_2 KS_3370(s3370, c3370, in3370_1, in3370_2);
    wire[0:0] s3371, in3371_1, in3371_2;
    wire c3371;
    assign in3371_1 = {pp105[91]};
    assign in3371_2 = {pp106[90]};
    Half_Adder KS_3371(s3371, c3371, in3371_1, in3371_2);
    wire[2:0] s3372, in3372_1, in3372_2;
    wire c3372;
    assign in3372_1 = {pp107[89],pp102[95],pp99[99]};
    assign in3372_2 = {pp108[88],pp103[94],pp100[98]};
    CLA_3 KS_3372(s3372, c3372, in3372_1, in3372_2);
    wire[0:0] s3373, in3373_1, in3373_2;
    wire c3373;
    assign in3373_1 = {pp109[87]};
    assign in3373_2 = {pp110[86]};
    Half_Adder KS_3373(s3373, c3373, in3373_1, in3373_2);
    wire[1:0] s3374, in3374_1, in3374_2;
    wire c3374;
    assign in3374_1 = {pp111[85],pp104[93]};
    assign in3374_2 = {pp112[84],pp105[92]};
    CLA_2 KS_3374(s3374, c3374, in3374_1, in3374_2);
    wire[0:0] s3375, in3375_1, in3375_2;
    wire c3375;
    assign in3375_1 = {pp113[83]};
    assign in3375_2 = {pp114[82]};
    Half_Adder KS_3375(s3375, c3375, in3375_1, in3375_2);
    wire[3:0] s3376, in3376_1, in3376_2;
    wire c3376;
    assign in3376_1 = {pp115[81],pp106[91],pp101[97],pp98[101]};
    assign in3376_2 = {pp116[80],pp107[90],pp102[96],pp99[100]};
    CLA_4 KS_3376(s3376, c3376, in3376_1, in3376_2);
    wire[0:0] s3377, in3377_1, in3377_2;
    wire c3377;
    assign in3377_1 = {pp117[79]};
    assign in3377_2 = {pp118[78]};
    Half_Adder KS_3377(s3377, c3377, in3377_1, in3377_2);
    wire[1:0] s3378, in3378_1, in3378_2;
    wire c3378;
    assign in3378_1 = {pp119[77],pp108[89]};
    assign in3378_2 = {pp120[76],pp109[88]};
    CLA_2 KS_3378(s3378, c3378, in3378_1, in3378_2);
    wire[0:0] s3379, in3379_1, in3379_2;
    wire c3379;
    assign in3379_1 = {pp121[75]};
    assign in3379_2 = {pp122[74]};
    Half_Adder KS_3379(s3379, c3379, in3379_1, in3379_2);
    wire[2:0] s3380, in3380_1, in3380_2;
    wire c3380;
    assign in3380_1 = {pp123[73],pp110[87],pp103[95]};
    assign in3380_2 = {pp124[72],pp111[86],pp104[94]};
    CLA_3 KS_3380(s3380, c3380, in3380_1, in3380_2);
    wire[0:0] s3381, in3381_1, in3381_2;
    wire c3381;
    assign in3381_1 = {pp125[71]};
    assign in3381_2 = {pp126[70]};
    Half_Adder KS_3381(s3381, c3381, in3381_1, in3381_2);
    wire[1:0] s3382, in3382_1, in3382_2;
    wire c3382;
    assign in3382_1 = {pp127[69],pp112[85]};
    assign in3382_2 = {c3312,pp113[84]};
    CLA_2 KS_3382(s3382, c3382, in3382_1, in3382_2);
    wire[0:0] s3383, in3383_1, in3383_2;
    wire c3383;
    assign in3383_1 = {c3313};
    assign in3383_2 = {c3314};
    Half_Adder KS_3383(s3383, c3383, in3383_1, in3383_2);
    wire[3:0] s3384, in3384_1, in3384_2;
    wire c3384;
    assign in3384_1 = {c3316,pp114[83],pp105[93],pp100[99]};
    assign in3384_2 = {c3317,pp115[82],pp106[92],pp101[98]};
    CLA_4_c KS_3384(s3384, c3384, in3384_1, in3384_2, c3315);
    wire[3:0] s3385, in3385_1, in3385_2;
    wire c3385;
    assign in3385_1 = {pp73[127],pp74[127],pp75[127],pp76[127]};
    assign in3385_2 = {pp74[126],pp75[126],pp76[126],pp77[126]};
    CLA_4 KS_3385(s3385, c3385, in3385_1, in3385_2);
    wire[3:0] s3386, in3386_1, in3386_2;
    wire c3386;
    assign in3386_1 = {pp75[125],pp76[125],pp77[125],pp78[125]};
    assign in3386_2 = {pp76[124],pp77[124],pp78[124],pp79[124]};
    CLA_4 KS_3386(s3386, c3386, in3386_1, in3386_2);
    wire[3:0] s3387, in3387_1, in3387_2;
    wire c3387;
    assign in3387_1 = {pp77[123],pp78[123],pp79[123],pp80[123]};
    assign in3387_2 = {pp78[122],pp79[122],pp80[122],pp81[122]};
    CLA_4 KS_3387(s3387, c3387, in3387_1, in3387_2);
    wire[3:0] s3388, in3388_1, in3388_2;
    wire c3388;
    assign in3388_1 = {pp79[121],pp80[121],pp81[121],pp82[121]};
    assign in3388_2 = {pp80[120],pp81[120],pp82[120],pp83[120]};
    CLA_4 KS_3388(s3388, c3388, in3388_1, in3388_2);
    wire[3:0] s3389, in3389_1, in3389_2;
    wire c3389;
    assign in3389_1 = {pp81[119],pp82[119],pp83[119],pp84[119]};
    assign in3389_2 = {pp82[118],pp83[118],pp84[118],pp85[118]};
    CLA_4 KS_3389(s3389, c3389, in3389_1, in3389_2);
    wire[3:0] s3390, in3390_1, in3390_2;
    wire c3390;
    assign in3390_1 = {pp83[117],pp84[117],pp85[117],pp86[117]};
    assign in3390_2 = {pp84[116],pp85[116],pp86[116],pp87[116]};
    CLA_4 KS_3390(s3390, c3390, in3390_1, in3390_2);
    wire[3:0] s3391, in3391_1, in3391_2;
    wire c3391;
    assign in3391_1 = {pp85[115],pp86[115],pp87[115],pp88[115]};
    assign in3391_2 = {pp86[114],pp87[114],pp88[114],pp89[114]};
    CLA_4 KS_3391(s3391, c3391, in3391_1, in3391_2);
    wire[3:0] s3392, in3392_1, in3392_2;
    wire c3392;
    assign in3392_1 = {pp87[113],pp88[113],pp89[113],pp90[113]};
    assign in3392_2 = {pp88[112],pp89[112],pp90[112],pp91[112]};
    CLA_4 KS_3392(s3392, c3392, in3392_1, in3392_2);
    wire[2:0] s3393, in3393_1, in3393_2;
    wire c3393;
    assign in3393_1 = {pp89[111],pp90[111],pp91[111]};
    assign in3393_2 = {pp90[110],pp91[110],pp92[110]};
    CLA_3 KS_3393(s3393, c3393, in3393_1, in3393_2);
    wire[1:0] s3394, in3394_1, in3394_2;
    wire c3394;
    assign in3394_1 = {pp91[109],pp92[109]};
    assign in3394_2 = {pp92[108],pp93[108]};
    CLA_2 KS_3394(s3394, c3394, in3394_1, in3394_2);
    wire[0:0] s3395, in3395_1, in3395_2;
    wire c3395;
    assign in3395_1 = {pp93[107]};
    assign in3395_2 = {pp94[106]};
    Half_Adder KS_3395(s3395, c3395, in3395_1, in3395_2);
    wire[3:0] s3396, in3396_1, in3396_2;
    wire c3396;
    assign in3396_1 = {pp95[105],pp94[107],pp93[109],pp92[111]};
    assign in3396_2 = {pp96[104],pp95[106],pp94[108],pp93[110]};
    CLA_4 KS_3396(s3396, c3396, in3396_1, in3396_2);
    wire[0:0] s3397, in3397_1, in3397_2;
    wire c3397;
    assign in3397_1 = {pp97[103]};
    assign in3397_2 = {pp98[102]};
    Half_Adder KS_3397(s3397, c3397, in3397_1, in3397_2);
    wire[1:0] s3398, in3398_1, in3398_2;
    wire c3398;
    assign in3398_1 = {pp99[101],pp96[105]};
    assign in3398_2 = {pp100[100],pp97[104]};
    CLA_2 KS_3398(s3398, c3398, in3398_1, in3398_2);
    wire[0:0] s3399, in3399_1, in3399_2;
    wire c3399;
    assign in3399_1 = {pp101[99]};
    assign in3399_2 = {pp102[98]};
    Half_Adder KS_3399(s3399, c3399, in3399_1, in3399_2);
    wire[2:0] s3400, in3400_1, in3400_2;
    wire c3400;
    assign in3400_1 = {pp103[97],pp98[103],pp95[107]};
    assign in3400_2 = {pp104[96],pp99[102],pp96[106]};
    CLA_3 KS_3400(s3400, c3400, in3400_1, in3400_2);
    wire[0:0] s3401, in3401_1, in3401_2;
    wire c3401;
    assign in3401_1 = {pp105[95]};
    assign in3401_2 = {pp106[94]};
    Half_Adder KS_3401(s3401, c3401, in3401_1, in3401_2);
    wire[1:0] s3402, in3402_1, in3402_2;
    wire c3402;
    assign in3402_1 = {pp107[93],pp100[101]};
    assign in3402_2 = {pp108[92],pp101[100]};
    CLA_2 KS_3402(s3402, c3402, in3402_1, in3402_2);
    wire[0:0] s3403, in3403_1, in3403_2;
    wire c3403;
    assign in3403_1 = {pp109[91]};
    assign in3403_2 = {pp110[90]};
    Half_Adder KS_3403(s3403, c3403, in3403_1, in3403_2);
    wire[3:0] s3404, in3404_1, in3404_2;
    wire c3404;
    assign in3404_1 = {pp111[89],pp102[99],pp97[105],pp94[109]};
    assign in3404_2 = {pp112[88],pp103[98],pp98[104],pp95[108]};
    CLA_4 KS_3404(s3404, c3404, in3404_1, in3404_2);
    wire[0:0] s3405, in3405_1, in3405_2;
    wire c3405;
    assign in3405_1 = {pp113[87]};
    assign in3405_2 = {pp114[86]};
    Half_Adder KS_3405(s3405, c3405, in3405_1, in3405_2);
    wire[1:0] s3406, in3406_1, in3406_2;
    wire c3406;
    assign in3406_1 = {pp115[85],pp104[97]};
    assign in3406_2 = {pp116[84],pp105[96]};
    CLA_2 KS_3406(s3406, c3406, in3406_1, in3406_2);
    wire[0:0] s3407, in3407_1, in3407_2;
    wire c3407;
    assign in3407_1 = {pp117[83]};
    assign in3407_2 = {pp118[82]};
    Half_Adder KS_3407(s3407, c3407, in3407_1, in3407_2);
    wire[2:0] s3408, in3408_1, in3408_2;
    wire c3408;
    assign in3408_1 = {pp120[80],pp106[95],pp99[103]};
    assign in3408_2 = {pp121[79],pp107[94],pp100[102]};
    CLA_3_c KS_3408(s3408, c3408, in3408_1, in3408_2, pp119[81]);
    wire[3:0] s3409, in3409_1, in3409_2;
    wire c3409;
    assign in3409_1 = {pp77[127],pp78[127],pp79[127],pp80[127]};
    assign in3409_2 = {pp78[126],pp79[126],pp80[126],pp81[126]};
    CLA_4 KS_3409(s3409, c3409, in3409_1, in3409_2);
    wire[3:0] s3410, in3410_1, in3410_2;
    wire c3410;
    assign in3410_1 = {pp79[125],pp80[125],pp81[125],pp82[125]};
    assign in3410_2 = {pp80[124],pp81[124],pp82[124],pp83[124]};
    CLA_4 KS_3410(s3410, c3410, in3410_1, in3410_2);
    wire[3:0] s3411, in3411_1, in3411_2;
    wire c3411;
    assign in3411_1 = {pp81[123],pp82[123],pp83[123],pp84[123]};
    assign in3411_2 = {pp82[122],pp83[122],pp84[122],pp85[122]};
    CLA_4 KS_3411(s3411, c3411, in3411_1, in3411_2);
    wire[3:0] s3412, in3412_1, in3412_2;
    wire c3412;
    assign in3412_1 = {pp83[121],pp84[121],pp85[121],pp86[121]};
    assign in3412_2 = {pp84[120],pp85[120],pp86[120],pp87[120]};
    CLA_4 KS_3412(s3412, c3412, in3412_1, in3412_2);
    wire[2:0] s3413, in3413_1, in3413_2;
    wire c3413;
    assign in3413_1 = {pp85[119],pp86[119],pp87[119]};
    assign in3413_2 = {pp86[118],pp87[118],pp88[118]};
    CLA_3 KS_3413(s3413, c3413, in3413_1, in3413_2);
    wire[1:0] s3414, in3414_1, in3414_2;
    wire c3414;
    assign in3414_1 = {pp87[117],pp88[117]};
    assign in3414_2 = {pp88[116],pp89[116]};
    CLA_2 KS_3414(s3414, c3414, in3414_1, in3414_2);
    wire[0:0] s3415, in3415_1, in3415_2;
    wire c3415;
    assign in3415_1 = {pp89[115]};
    assign in3415_2 = {pp90[114]};
    Half_Adder KS_3415(s3415, c3415, in3415_1, in3415_2);
    wire[3:0] s3416, in3416_1, in3416_2;
    wire c3416;
    assign in3416_1 = {pp91[113],pp90[115],pp89[117],pp88[119]};
    assign in3416_2 = {pp92[112],pp91[114],pp90[116],pp89[118]};
    CLA_4 KS_3416(s3416, c3416, in3416_1, in3416_2);
    wire[0:0] s3417, in3417_1, in3417_2;
    wire c3417;
    assign in3417_1 = {pp93[111]};
    assign in3417_2 = {pp94[110]};
    Half_Adder KS_3417(s3417, c3417, in3417_1, in3417_2);
    wire[1:0] s3418, in3418_1, in3418_2;
    wire c3418;
    assign in3418_1 = {pp95[109],pp92[113]};
    assign in3418_2 = {pp96[108],pp93[112]};
    CLA_2 KS_3418(s3418, c3418, in3418_1, in3418_2);
    wire[0:0] s3419, in3419_1, in3419_2;
    wire c3419;
    assign in3419_1 = {pp97[107]};
    assign in3419_2 = {pp98[106]};
    Half_Adder KS_3419(s3419, c3419, in3419_1, in3419_2);
    wire[2:0] s3420, in3420_1, in3420_2;
    wire c3420;
    assign in3420_1 = {pp99[105],pp94[111],pp91[115]};
    assign in3420_2 = {pp100[104],pp95[110],pp92[114]};
    CLA_3 KS_3420(s3420, c3420, in3420_1, in3420_2);
    wire[0:0] s3421, in3421_1, in3421_2;
    wire c3421;
    assign in3421_1 = {pp101[103]};
    assign in3421_2 = {pp102[102]};
    Half_Adder KS_3421(s3421, c3421, in3421_1, in3421_2);
    wire[1:0] s3422, in3422_1, in3422_2;
    wire c3422;
    assign in3422_1 = {pp103[101],pp96[109]};
    assign in3422_2 = {pp104[100],pp97[108]};
    CLA_2 KS_3422(s3422, c3422, in3422_1, in3422_2);
    wire[0:0] s3423, in3423_1, in3423_2;
    wire c3423;
    assign in3423_1 = {pp106[98]};
    assign in3423_2 = {pp107[97]};
    Full_Adder KS_3423(s3423, c3423, in3423_1, in3423_2, pp105[99]);
    wire[2:0] s3424, in3424_1, in3424_2;
    wire c3424;
    assign in3424_1 = {pp81[127],pp82[127],pp83[127]};
    assign in3424_2 = {pp82[126],pp83[126],pp84[126]};
    CLA_3 KS_3424(s3424, c3424, in3424_1, in3424_2);
    wire[1:0] s3425, in3425_1, in3425_2;
    wire c3425;
    assign in3425_1 = {pp83[125],pp84[125]};
    assign in3425_2 = {pp84[124],pp85[124]};
    CLA_2 KS_3425(s3425, c3425, in3425_1, in3425_2);
    wire[0:0] s3426, in3426_1, in3426_2;
    wire c3426;
    assign in3426_1 = {pp85[123]};
    assign in3426_2 = {pp86[122]};
    Half_Adder KS_3426(s3426, c3426, in3426_1, in3426_2);
    wire[3:0] s3427, in3427_1, in3427_2;
    wire c3427;
    assign in3427_1 = {pp87[121],pp86[123],pp85[125],pp84[127]};
    assign in3427_2 = {pp88[120],pp87[122],pp86[124],pp85[126]};
    CLA_4 KS_3427(s3427, c3427, in3427_1, in3427_2);
    wire[0:0] s3428, in3428_1, in3428_2;
    wire c3428;
    assign in3428_1 = {pp89[119]};
    assign in3428_2 = {pp90[118]};
    Half_Adder KS_3428(s3428, c3428, in3428_1, in3428_2);
    wire[1:0] s3429, in3429_1, in3429_2;
    wire c3429;
    assign in3429_1 = {pp92[116],pp88[121]};
    assign in3429_2 = {pp93[115],pp89[120]};
    CLA_2_c KS_3429(s3429, c3429, in3429_1, in3429_2, pp91[117]);

    /*Stage 3*/
    wire[3:0] s3430, in3430_1, in3430_2;
    wire c3430;
    assign in3430_1 = {pp0[27],pp0[28],pp0[29],pp0[30]};
    assign in3430_2 = {pp1[26],pp1[27],pp1[28],pp1[29]};
    CLA_4 KS_3430(s3430, c3430, in3430_1, in3430_2);
    wire[3:0] s3431, in3431_1, in3431_2;
    wire c3431;
    assign in3431_1 = {pp2[26],pp2[27],pp2[28],pp0[31]};
    assign in3431_2 = {pp3[25],pp3[26],pp3[27],pp1[30]};
    CLA_4 KS_3431(s3431, c3431, in3431_1, in3431_2);
    wire[3:0] s3432, in3432_1, in3432_2;
    wire c3432;
    assign in3432_1 = {pp4[25],pp4[26],pp2[29],pp0[32]};
    assign in3432_2 = {pp5[24],pp5[25],pp3[28],pp1[31]};
    CLA_4 KS_3432(s3432, c3432, in3432_1, in3432_2);
    wire[3:0] s3433, in3433_1, in3433_2;
    wire c3433;
    assign in3433_1 = {pp6[24],pp4[27],pp2[30],pp0[33]};
    assign in3433_2 = {pp7[23],pp5[26],pp3[29],pp1[32]};
    CLA_4 KS_3433(s3433, c3433, in3433_1, in3433_2);
    wire[3:0] s3434, in3434_1, in3434_2;
    wire c3434;
    assign in3434_1 = {pp6[25],pp4[28],pp2[31],pp0[34]};
    assign in3434_2 = {pp7[24],pp5[27],pp3[30],pp1[33]};
    CLA_4 KS_3434(s3434, c3434, in3434_1, in3434_2);
    wire[3:0] s3435, in3435_1, in3435_2;
    wire c3435;
    assign in3435_1 = {pp9[22],pp6[26],pp4[29],pp2[32]};
    assign in3435_2 = {pp10[21],pp7[25],pp5[28],pp3[31]};
    CLA_4_c KS_3435(s3435, c3435, in3435_1, in3435_2, pp8[23]);
    wire[3:0] s3436, in3436_1, in3436_2;
    wire c3436;
    assign in3436_1 = {pp8[24],pp6[27],pp4[30],pp0[35]};
    assign in3436_2 = {pp9[23],pp7[26],pp5[29],pp1[34]};
    CLA_4 KS_3436(s3436, c3436, in3436_1, in3436_2);
    wire[3:0] s3437, in3437_1, in3437_2;
    wire c3437;
    assign in3437_1 = {pp11[21],pp8[25],pp6[28],pp2[33]};
    assign in3437_2 = {pp12[20],pp9[24],pp7[27],pp3[32]};
    CLA_4_c KS_3437(s3437, c3437, in3437_1, in3437_2, pp10[22]);
    wire[3:0] s3438, in3438_1, in3438_2;
    wire c3438;
    assign in3438_1 = {pp10[23],pp8[26],pp4[31],pp0[36]};
    assign in3438_2 = {pp11[22],pp9[25],pp5[30],pp1[35]};
    CLA_4 KS_3438(s3438, c3438, in3438_1, in3438_2);
    wire[3:0] s3439, in3439_1, in3439_2;
    wire c3439;
    assign in3439_1 = {pp13[20],pp10[24],pp6[29],pp2[34]};
    assign in3439_2 = {pp14[19],pp11[23],pp7[28],pp3[33]};
    CLA_4_c KS_3439(s3439, c3439, in3439_1, in3439_2, pp12[21]);
    wire[3:0] s3440, in3440_1, in3440_2;
    wire c3440;
    assign in3440_1 = {pp12[22],pp8[27],pp4[32],pp0[37]};
    assign in3440_2 = {pp13[21],pp9[26],pp5[31],pp1[36]};
    CLA_4 KS_3440(s3440, c3440, in3440_1, in3440_2);
    wire[3:0] s3441, in3441_1, in3441_2;
    wire c3441;
    assign in3441_1 = {pp15[19],pp10[25],pp6[30],pp2[35]};
    assign in3441_2 = {pp16[18],pp11[24],pp7[29],pp3[34]};
    CLA_4_c KS_3441(s3441, c3441, in3441_1, in3441_2, pp14[20]);
    wire[3:0] s3442, in3442_1, in3442_2;
    wire c3442;
    assign in3442_1 = {pp12[23],pp8[28],pp4[33],pp0[38]};
    assign in3442_2 = {pp13[22],pp9[27],pp5[32],pp1[37]};
    CLA_4 KS_3442(s3442, c3442, in3442_1, in3442_2);
    wire[3:0] s3443, in3443_1, in3443_2;
    wire c3443;
    assign in3443_1 = {pp14[21],pp10[26],pp6[31],pp2[36]};
    assign in3443_2 = {pp15[20],pp11[25],pp7[30],pp3[35]};
    CLA_4 KS_3443(s3443, c3443, in3443_1, in3443_2);
    wire[3:0] s3444, in3444_1, in3444_2;
    wire c3444;
    assign in3444_1 = {pp16[19],pp12[24],pp8[29],pp4[34]};
    assign in3444_2 = {pp17[18],pp13[23],pp9[28],pp5[33]};
    CLA_4 KS_3444(s3444, c3444, in3444_1, in3444_2);
    wire[3:0] s3445, in3445_1, in3445_2;
    wire c3445;
    assign in3445_1 = {pp19[16],pp14[22],pp10[27],pp6[32]};
    assign in3445_2 = {pp20[15],pp15[21],pp11[26],pp7[31]};
    CLA_4_c KS_3445(s3445, c3445, in3445_1, in3445_2, pp18[17]);
    wire[3:0] s3446, in3446_1, in3446_2;
    wire c3446;
    assign in3446_1 = {pp16[20],pp12[25],pp8[30],pp0[39]};
    assign in3446_2 = {pp17[19],pp13[24],pp9[29],pp1[38]};
    CLA_4 KS_3446(s3446, c3446, in3446_1, in3446_2);
    wire[3:0] s3447, in3447_1, in3447_2;
    wire c3447;
    assign in3447_1 = {pp18[18],pp14[23],pp10[28],pp2[37]};
    assign in3447_2 = {pp19[17],pp15[22],pp11[27],pp3[36]};
    CLA_4 KS_3447(s3447, c3447, in3447_1, in3447_2);
    wire[3:0] s3448, in3448_1, in3448_2;
    wire c3448;
    assign in3448_1 = {pp21[15],pp16[21],pp12[26],pp4[35]};
    assign in3448_2 = {pp22[14],pp17[20],pp13[25],pp5[34]};
    CLA_4_c KS_3448(s3448, c3448, in3448_1, in3448_2, pp20[16]);
    wire[3:0] s3449, in3449_1, in3449_2;
    wire c3449;
    assign in3449_1 = {pp18[19],pp14[24],pp6[33],pp0[40]};
    assign in3449_2 = {pp19[18],pp15[23],pp7[32],pp1[39]};
    CLA_4 KS_3449(s3449, c3449, in3449_1, in3449_2);
    wire[3:0] s3450, in3450_1, in3450_2;
    wire c3450;
    assign in3450_1 = {pp20[17],pp16[22],pp8[31],pp2[38]};
    assign in3450_2 = {pp21[16],pp17[21],pp9[30],pp3[37]};
    CLA_4 KS_3450(s3450, c3450, in3450_1, in3450_2);
    wire[3:0] s3451, in3451_1, in3451_2;
    wire c3451;
    assign in3451_1 = {pp23[14],pp18[20],pp10[29],pp4[36]};
    assign in3451_2 = {pp24[13],pp19[19],pp11[28],pp5[35]};
    CLA_4_c KS_3451(s3451, c3451, in3451_1, in3451_2, pp22[15]);
    wire[3:0] s3452, in3452_1, in3452_2;
    wire c3452;
    assign in3452_1 = {pp20[18],pp12[27],pp6[34],pp0[41]};
    assign in3452_2 = {pp21[17],pp13[26],pp7[33],pp1[40]};
    CLA_4 KS_3452(s3452, c3452, in3452_1, in3452_2);
    wire[3:0] s3453, in3453_1, in3453_2;
    wire c3453;
    assign in3453_1 = {pp22[16],pp14[25],pp8[32],pp2[39]};
    assign in3453_2 = {pp23[15],pp15[24],pp9[31],pp3[38]};
    CLA_4 KS_3453(s3453, c3453, in3453_1, in3453_2);
    wire[3:0] s3454, in3454_1, in3454_2;
    wire c3454;
    assign in3454_1 = {pp25[13],pp16[23],pp10[30],pp4[37]};
    assign in3454_2 = {pp26[12],pp17[22],pp11[29],pp5[36]};
    CLA_4_c KS_3454(s3454, c3454, in3454_1, in3454_2, pp24[14]);
    wire[3:0] s3455, in3455_1, in3455_2;
    wire c3455;
    assign in3455_1 = {pp18[21],pp12[28],pp6[35],pp0[42]};
    assign in3455_2 = {pp19[20],pp13[27],pp7[34],pp1[41]};
    CLA_4 KS_3455(s3455, c3455, in3455_1, in3455_2);
    wire[3:0] s3456, in3456_1, in3456_2;
    wire c3456;
    assign in3456_1 = {pp20[19],pp14[26],pp8[33],pp2[40]};
    assign in3456_2 = {pp21[18],pp15[25],pp9[32],pp3[39]};
    CLA_4 KS_3456(s3456, c3456, in3456_1, in3456_2);
    wire[3:0] s3457, in3457_1, in3457_2;
    wire c3457;
    assign in3457_1 = {pp22[17],pp16[24],pp10[31],pp4[38]};
    assign in3457_2 = {pp23[16],pp17[23],pp11[30],pp5[37]};
    CLA_4 KS_3457(s3457, c3457, in3457_1, in3457_2);
    wire[3:0] s3458, in3458_1, in3458_2;
    wire c3458;
    assign in3458_1 = {pp24[15],pp18[22],pp12[29],pp6[36]};
    assign in3458_2 = {pp25[14],pp19[21],pp13[28],pp7[35]};
    CLA_4 KS_3458(s3458, c3458, in3458_1, in3458_2);
    wire[3:0] s3459, in3459_1, in3459_2;
    wire c3459;
    assign in3459_1 = {pp26[13],pp20[20],pp14[27],pp8[34]};
    assign in3459_2 = {pp27[12],pp21[19],pp15[26],pp9[33]};
    CLA_4 KS_3459(s3459, c3459, in3459_1, in3459_2);
    wire[3:0] s3460, in3460_1, in3460_2;
    wire c3460;
    assign in3460_1 = {pp28[11],pp22[18],pp16[25],pp10[32]};
    assign in3460_2 = {pp29[10],pp23[17],pp17[24],pp11[31]};
    CLA_4 KS_3460(s3460, c3460, in3460_1, in3460_2);
    wire[3:0] s3461, in3461_1, in3461_2;
    wire c3461;
    assign in3461_1 = {pp31[8],pp24[16],pp18[23],pp12[30]};
    assign in3461_2 = {pp32[7],pp25[15],pp19[22],pp13[29]};
    CLA_4_c KS_3461(s3461, c3461, in3461_1, in3461_2, pp30[9]);
    wire[3:0] s3462, in3462_1, in3462_2;
    wire c3462;
    assign in3462_1 = {pp26[14],pp20[21],pp14[28],pp0[43]};
    assign in3462_2 = {pp27[13],pp21[20],pp15[27],pp1[42]};
    CLA_4 KS_3462(s3462, c3462, in3462_1, in3462_2);
    wire[3:0] s3463, in3463_1, in3463_2;
    wire c3463;
    assign in3463_1 = {pp28[12],pp22[19],pp16[26],pp2[41]};
    assign in3463_2 = {pp29[11],pp23[18],pp17[25],pp3[40]};
    CLA_4 KS_3463(s3463, c3463, in3463_1, in3463_2);
    wire[3:0] s3464, in3464_1, in3464_2;
    wire c3464;
    assign in3464_1 = {pp31[9],pp24[17],pp18[24],pp4[39]};
    assign in3464_2 = {pp32[8],pp25[16],pp19[23],pp5[38]};
    CLA_4_c KS_3464(s3464, c3464, in3464_1, in3464_2, pp30[10]);
    wire[3:0] s3465, in3465_1, in3465_2;
    wire c3465;
    assign in3465_1 = {pp26[15],pp20[22],pp6[37],pp0[44]};
    assign in3465_2 = {pp27[14],pp21[21],pp7[36],pp1[43]};
    CLA_4 KS_3465(s3465, c3465, in3465_1, in3465_2);
    wire[3:0] s3466, in3466_1, in3466_2;
    wire c3466;
    assign in3466_1 = {pp28[13],pp22[20],pp8[35],pp2[42]};
    assign in3466_2 = {pp29[12],pp23[19],pp9[34],pp3[41]};
    CLA_4 KS_3466(s3466, c3466, in3466_1, in3466_2);
    wire[3:0] s3467, in3467_1, in3467_2;
    wire c3467;
    assign in3467_1 = {pp30[11],pp24[18],pp10[33],pp4[40]};
    assign in3467_2 = {pp31[10],pp25[17],pp11[32],pp5[39]};
    CLA_4 KS_3467(s3467, c3467, in3467_1, in3467_2);
    wire[3:0] s3468, in3468_1, in3468_2;
    wire c3468;
    assign in3468_1 = {pp33[8],pp26[16],pp12[31],pp6[38]};
    assign in3468_2 = {pp34[7],pp27[15],pp13[30],pp7[37]};
    CLA_4_c KS_3468(s3468, c3468, in3468_1, in3468_2, pp32[9]);
    wire[3:0] s3469, in3469_1, in3469_2;
    wire c3469;
    assign in3469_1 = {pp28[14],pp14[29],pp8[36],pp2[43]};
    assign in3469_2 = {pp29[13],pp15[28],pp9[35],pp3[42]};
    CLA_4 KS_3469(s3469, c3469, in3469_1, in3469_2);
    wire[3:0] s3470, in3470_1, in3470_2;
    wire c3470;
    assign in3470_1 = {pp30[12],pp16[27],pp10[34],pp4[41]};
    assign in3470_2 = {pp31[11],pp17[26],pp11[33],pp5[40]};
    CLA_4 KS_3470(s3470, c3470, in3470_1, in3470_2);
    wire[3:0] s3471, in3471_1, in3471_2;
    wire c3471;
    assign in3471_1 = {pp32[10],pp18[25],pp12[32],pp6[39]};
    assign in3471_2 = {pp33[9],pp19[24],pp13[31],pp7[38]};
    CLA_4 KS_3471(s3471, c3471, in3471_1, in3471_2);
    wire[3:0] s3472, in3472_1, in3472_2;
    wire c3472;
    assign in3472_1 = {pp35[7],pp20[23],pp14[30],pp8[37]};
    assign in3472_2 = {pp36[6],pp21[22],pp15[29],pp9[36]};
    CLA_4_c KS_3472(s3472, c3472, in3472_1, in3472_2, pp34[8]);
    wire[3:0] s3473, in3473_1, in3473_2;
    wire c3473;
    assign in3473_1 = {pp22[21],pp16[28],pp10[35],pp4[42]};
    assign in3473_2 = {pp23[20],pp17[27],pp11[34],pp5[41]};
    CLA_4 KS_3473(s3473, c3473, in3473_1, in3473_2);
    wire[3:0] s3474, in3474_1, in3474_2;
    wire c3474;
    assign in3474_1 = {pp24[19],pp18[26],pp12[33],pp6[40]};
    assign in3474_2 = {pp25[18],pp19[25],pp13[32],pp7[39]};
    CLA_4 KS_3474(s3474, c3474, in3474_1, in3474_2);
    wire[3:0] s3475, in3475_1, in3475_2;
    wire c3475;
    assign in3475_1 = {pp26[17],pp20[24],pp14[31],pp8[38]};
    assign in3475_2 = {pp27[16],pp21[23],pp15[30],pp9[37]};
    CLA_4 KS_3475(s3475, c3475, in3475_1, in3475_2);
    wire[3:0] s3476, in3476_1, in3476_2;
    wire c3476;
    assign in3476_1 = {pp28[15],pp22[22],pp16[29],pp10[36]};
    assign in3476_2 = {pp29[14],pp23[21],pp17[28],pp11[35]};
    CLA_4 KS_3476(s3476, c3476, in3476_1, in3476_2);
    wire[3:0] s3477, in3477_1, in3477_2;
    wire c3477;
    assign in3477_1 = {pp30[13],pp24[20],pp18[27],pp12[34]};
    assign in3477_2 = {pp31[12],pp25[19],pp19[26],pp13[33]};
    CLA_4 KS_3477(s3477, c3477, in3477_1, in3477_2);
    wire[3:0] s3478, in3478_1, in3478_2;
    wire c3478;
    assign in3478_1 = {pp32[11],pp26[18],pp20[25],pp14[32]};
    assign in3478_2 = {pp33[10],pp27[17],pp21[24],pp15[31]};
    CLA_4 KS_3478(s3478, c3478, in3478_1, in3478_2);
    wire[3:0] s3479, in3479_1, in3479_2;
    wire c3479;
    assign in3479_1 = {pp34[9],pp28[16],pp22[23],pp16[30]};
    assign in3479_2 = {pp35[8],pp29[15],pp23[22],pp17[29]};
    CLA_4 KS_3479(s3479, c3479, in3479_1, in3479_2);
    wire[3:0] s3480, in3480_1, in3480_2;
    wire c3480;
    assign in3480_1 = {pp36[7],pp30[14],pp24[21],pp18[28]};
    assign in3480_2 = {pp37[6],pp31[13],pp25[20],pp19[27]};
    CLA_4 KS_3480(s3480, c3480, in3480_1, in3480_2);
    wire[3:0] s3481, in3481_1, in3481_2;
    wire c3481;
    assign in3481_1 = {pp38[5],pp32[12],pp26[19],pp20[26]};
    assign in3481_2 = {pp39[4],pp33[11],pp27[18],pp21[25]};
    CLA_4 KS_3481(s3481, c3481, in3481_1, in3481_2);
    wire[3:0] s3482, in3482_1, in3482_2;
    wire c3482;
    assign in3482_1 = {pp40[3],pp34[10],pp28[17],pp22[24]};
    assign in3482_2 = {pp41[2],pp35[9],pp29[16],pp23[23]};
    CLA_4 KS_3482(s3482, c3482, in3482_1, in3482_2);
    wire[3:0] s3483, in3483_1, in3483_2;
    wire c3483;
    assign in3483_1 = {pp42[1],pp36[8],pp30[15],pp24[22]};
    assign in3483_2 = {pp43[0],pp37[7],pp31[14],pp25[21]};
    CLA_4 KS_3483(s3483, c3483, in3483_1, in3483_2);
    wire[3:0] s3484, in3484_1, in3484_2;
    wire c3484;
    assign in3484_1 = {c3456,pp38[6],pp32[13],pp26[20]};
    assign in3484_2 = {c3457,pp39[5],pp33[12],pp27[19]};
    CLA_4_c KS_3484(s3484, c3484, in3484_1, in3484_2, c3455);
    wire[3:0] s3485, in3485_1, in3485_2;
    wire c3485;
    assign in3485_1 = {pp40[4],pp34[11],pp28[18],pp6[41]};
    assign in3485_2 = {pp41[3],pp35[10],pp29[17],pp7[40]};
    CLA_4 KS_3485(s3485, c3485, in3485_1, in3485_2);
    wire[3:0] s3486, in3486_1, in3486_2;
    wire c3486;
    assign in3486_1 = {pp36[9],pp30[16],pp8[39],pp8[40]};
    assign in3486_2 = {pp37[8],pp31[15],pp9[38],pp9[39]};
    CLA_4 KS_3486(s3486, c3486, in3486_1, in3486_2);
    wire[3:0] s3487, in3487_1, in3487_2;
    wire c3487;
    assign in3487_1 = {pp38[7],pp32[14],pp10[37],pp10[38]};
    assign in3487_2 = {pp39[6],pp33[13],pp11[36],pp11[37]};
    CLA_4 KS_3487(s3487, c3487, in3487_1, in3487_2);
    wire[3:0] s3488, in3488_1, in3488_2;
    wire c3488;
    assign in3488_1 = {pp40[5],pp34[12],pp12[35],pp12[36]};
    assign in3488_2 = {pp41[4],pp35[11],pp13[34],pp13[35]};
    CLA_4 KS_3488(s3488, c3488, in3488_1, in3488_2);
    wire[3:0] s3489, in3489_1, in3489_2;
    wire c3489;
    assign in3489_1 = {pp43[2],pp36[10],pp14[33],pp14[34]};
    assign in3489_2 = {pp44[1],pp37[9],pp15[32],pp15[33]};
    CLA_4_c KS_3489(s3489, c3489, in3489_1, in3489_2, pp42[3]);
    wire[3:0] s3490, in3490_1, in3490_2;
    wire c3490;
    assign in3490_1 = {pp38[8],pp16[31],pp16[32],pp11[38]};
    assign in3490_2 = {pp39[7],pp17[30],pp17[31],pp12[37]};
    CLA_4 KS_3490(s3490, c3490, in3490_1, in3490_2);
    wire[3:0] s3491, in3491_1, in3491_2;
    wire c3491;
    assign in3491_1 = {pp40[6],pp18[29],pp18[30],pp13[36]};
    assign in3491_2 = {pp41[5],pp19[28],pp19[29],pp14[35]};
    CLA_4 KS_3491(s3491, c3491, in3491_1, in3491_2);
    wire[3:0] s3492, in3492_1, in3492_2;
    wire c3492;
    assign in3492_1 = {pp42[4],pp20[27],pp20[28],pp15[34]};
    assign in3492_2 = {pp43[3],pp21[26],pp21[27],pp16[33]};
    CLA_4 KS_3492(s3492, c3492, in3492_1, in3492_2);
    wire[3:0] s3493, in3493_1, in3493_2;
    wire c3493;
    assign in3493_1 = {pp45[1],pp22[25],pp22[26],pp17[32]};
    assign in3493_2 = {pp46[0],pp23[24],pp23[25],pp18[31]};
    CLA_4_c KS_3493(s3493, c3493, in3493_1, in3493_2, pp44[2]);
    wire[3:0] s3494, in3494_1, in3494_2;
    wire c3494;
    assign in3494_1 = {pp24[23],pp24[24],pp19[30],pp13[37]};
    assign in3494_2 = {pp25[22],pp25[23],pp20[29],pp14[36]};
    CLA_4 KS_3494(s3494, c3494, in3494_1, in3494_2);
    wire[3:0] s3495, in3495_1, in3495_2;
    wire c3495;
    assign in3495_1 = {pp26[21],pp26[22],pp21[28],pp15[35]};
    assign in3495_2 = {pp27[20],pp27[21],pp22[27],pp16[34]};
    CLA_4 KS_3495(s3495, c3495, in3495_1, in3495_2);
    wire[3:0] s3496, in3496_1, in3496_2;
    wire c3496;
    assign in3496_1 = {pp28[19],pp28[20],pp23[26],pp17[33]};
    assign in3496_2 = {pp29[18],pp29[19],pp24[25],pp18[32]};
    CLA_4 KS_3496(s3496, c3496, in3496_1, in3496_2);
    wire[3:0] s3497, in3497_1, in3497_2;
    wire c3497;
    assign in3497_1 = {pp30[17],pp30[18],pp25[24],pp19[31]};
    assign in3497_2 = {pp31[16],pp31[17],pp26[23],pp20[30]};
    CLA_4 KS_3497(s3497, c3497, in3497_1, in3497_2);
    wire[3:0] s3498, in3498_1, in3498_2;
    wire c3498;
    assign in3498_1 = {pp32[15],pp32[16],pp27[22],pp21[29]};
    assign in3498_2 = {pp33[14],pp33[15],pp28[21],pp22[28]};
    CLA_4 KS_3498(s3498, c3498, in3498_1, in3498_2);
    wire[3:0] s3499, in3499_1, in3499_2;
    wire c3499;
    assign in3499_1 = {pp34[13],pp34[14],pp29[20],pp23[27]};
    assign in3499_2 = {pp35[12],pp35[13],pp30[19],pp24[26]};
    CLA_4 KS_3499(s3499, c3499, in3499_1, in3499_2);
    wire[3:0] s3500, in3500_1, in3500_2;
    wire c3500;
    assign in3500_1 = {pp36[11],pp36[12],pp31[18],pp25[25]};
    assign in3500_2 = {pp37[10],pp37[11],pp32[17],pp26[24]};
    CLA_4 KS_3500(s3500, c3500, in3500_1, in3500_2);
    wire[3:0] s3501, in3501_1, in3501_2;
    wire c3501;
    assign in3501_1 = {pp38[9],pp38[10],pp33[16],pp27[23]};
    assign in3501_2 = {pp39[8],pp39[9],pp34[15],pp28[22]};
    CLA_4 KS_3501(s3501, c3501, in3501_1, in3501_2);
    wire[3:0] s3502, in3502_1, in3502_2;
    wire c3502;
    assign in3502_1 = {pp40[7],pp40[8],pp35[14],pp29[21]};
    assign in3502_2 = {pp41[6],pp41[7],pp36[13],pp30[20]};
    CLA_4 KS_3502(s3502, c3502, in3502_1, in3502_2);
    wire[3:0] s3503, in3503_1, in3503_2;
    wire c3503;
    assign in3503_1 = {pp42[5],pp42[6],pp37[12],pp31[19]};
    assign in3503_2 = {pp43[4],pp43[5],pp38[11],pp32[18]};
    CLA_4 KS_3503(s3503, c3503, in3503_1, in3503_2);
    wire[3:0] s3504, in3504_1, in3504_2;
    wire c3504;
    assign in3504_1 = {pp44[3],pp44[4],pp39[10],pp33[17]};
    assign in3504_2 = {pp45[2],pp45[3],pp40[9],pp34[16]};
    CLA_4 KS_3504(s3504, c3504, in3504_1, in3504_2);
    wire[3:0] s3505, in3505_1, in3505_2;
    wire c3505;
    assign in3505_1 = {pp46[1],pp46[2],pp41[8],pp35[15]};
    assign in3505_2 = {pp47[0],pp47[1],pp42[7],pp36[14]};
    CLA_4 KS_3505(s3505, c3505, in3505_1, in3505_2);
    wire[0:0] s3506, in3506_1, in3506_2;
    wire c3506;
    assign in3506_1 = {s1327[2]};
    assign in3506_2 = {s1328[1]};
    Half_Adder KS_3506(s3506, c3506, in3506_1, in3506_2);
    wire[3:0] s3507, in3507_1, in3507_2;
    wire c3507;
    assign in3507_1 = {s1329[0],pp48[0],pp43[6],pp37[13]};
    assign in3507_2 = {c3473,s1327[3],pp44[5],pp38[12]};
    CLA_4 KS_3507(s3507, c3507, in3507_1, in3507_2);
    wire[0:0] s3508, in3508_1, in3508_2;
    wire c3508;
    assign in3508_1 = {c3474};
    assign in3508_2 = {c3475};
    Half_Adder KS_3508(s3508, c3508, in3508_1, in3508_2);
    wire[3:0] s3509, in3509_1, in3509_2;
    wire c3509;
    assign in3509_1 = {c3476,s1328[2],pp45[4],pp39[11]};
    assign in3509_2 = {c3477,s1329[1],pp46[3],pp40[10]};
    CLA_4 KS_3509(s3509, c3509, in3509_1, in3509_2);
    wire[0:0] s3510, in3510_1, in3510_2;
    wire c3510;
    assign in3510_1 = {c3478};
    assign in3510_2 = {c3479};
    Half_Adder KS_3510(s3510, c3510, in3510_1, in3510_2);
    wire[3:0] s3511, in3511_1, in3511_2;
    wire c3511;
    assign in3511_1 = {c3480,s1330[0],pp47[2],pp41[9]};
    assign in3511_2 = {c3481,c3485,pp48[1],pp42[8]};
    CLA_4 KS_3511(s3511, c3511, in3511_1, in3511_2);
    wire[0:0] s3512, in3512_1, in3512_2;
    wire c3512;
    assign in3512_1 = {c3482};
    assign in3512_2 = {c3483};
    Half_Adder KS_3512(s3512, c3512, in3512_1, in3512_2);
    wire[3:0] s3513, in3513_1, in3513_2;
    wire c3513;
    assign in3513_1 = {s3485[3],s3486[3],pp49[0],pp43[7]};
    assign in3513_2 = {s3486[2],s3487[3],c1327,pp44[6]};
    CLA_4_c KS_3513(s3513, c3513, in3513_1, in3513_2, c3484);
    wire[3:0] s3514, in3514_1, in3514_2;
    wire c3514;
    assign in3514_1 = {s1329[2],pp45[5],pp15[36],pp17[35]};
    assign in3514_2 = {s1330[1],pp46[4],pp16[35],pp18[34]};
    CLA_4_c KS_3514(s3514, c3514, in3514_1, in3514_2, s1328[3]);
    wire[3:0] s3515, in3515_1, in3515_2;
    wire c3515;
    assign in3515_1 = {pp47[3],pp17[34],pp19[33],pp21[32]};
    assign in3515_2 = {pp48[2],pp18[33],pp20[32],pp22[31]};
    CLA_4 KS_3515(s3515, c3515, in3515_1, in3515_2);
    wire[3:0] s3516, in3516_1, in3516_2;
    wire c3516;
    assign in3516_1 = {pp49[1],pp19[32],pp21[31],pp23[30]};
    assign in3516_2 = {pp50[0],pp20[31],pp22[30],pp24[29]};
    CLA_4 KS_3516(s3516, c3516, in3516_1, in3516_2);
    wire[3:0] s3517, in3517_1, in3517_2;
    wire c3517;
    assign in3517_1 = {c1328,pp21[30],pp23[29],pp25[28]};
    assign in3517_2 = {s1329[3],pp22[29],pp24[28],pp26[27]};
    CLA_4 KS_3517(s3517, c3517, in3517_1, in3517_2);
    wire[3:0] s3518, in3518_1, in3518_2;
    wire c3518;
    assign in3518_1 = {s1331[1],pp23[28],pp25[27],pp27[26]};
    assign in3518_2 = {s1332[1],pp24[27],pp26[26],pp28[25]};
    CLA_4_c KS_3518(s3518, c3518, in3518_1, in3518_2, s1330[2]);
    wire[3:0] s3519, in3519_1, in3519_2;
    wire c3519;
    assign in3519_1 = {pp25[26],pp27[25],pp29[24],pp23[31]};
    assign in3519_2 = {pp26[25],pp28[24],pp30[23],pp24[30]};
    CLA_4 KS_3519(s3519, c3519, in3519_1, in3519_2);
    wire[3:0] s3520, in3520_1, in3520_2;
    wire c3520;
    assign in3520_1 = {pp27[24],pp29[23],pp31[22],pp25[29]};
    assign in3520_2 = {pp28[23],pp30[22],pp32[21],pp26[28]};
    CLA_4 KS_3520(s3520, c3520, in3520_1, in3520_2);
    wire[3:0] s3521, in3521_1, in3521_2;
    wire c3521;
    assign in3521_1 = {pp29[22],pp31[21],pp33[20],pp27[27]};
    assign in3521_2 = {pp30[21],pp32[20],pp34[19],pp28[26]};
    CLA_4 KS_3521(s3521, c3521, in3521_1, in3521_2);
    wire[3:0] s3522, in3522_1, in3522_2;
    wire c3522;
    assign in3522_1 = {pp31[20],pp33[19],pp35[18],pp29[25]};
    assign in3522_2 = {pp32[19],pp34[18],pp36[17],pp30[24]};
    CLA_4 KS_3522(s3522, c3522, in3522_1, in3522_2);
    wire[3:0] s3523, in3523_1, in3523_2;
    wire c3523;
    assign in3523_1 = {pp33[18],pp35[17],pp37[16],pp31[23]};
    assign in3523_2 = {pp34[17],pp36[16],pp38[15],pp32[22]};
    CLA_4 KS_3523(s3523, c3523, in3523_1, in3523_2);
    wire[3:0] s3524, in3524_1, in3524_2;
    wire c3524;
    assign in3524_1 = {pp35[16],pp37[15],pp39[14],pp33[21]};
    assign in3524_2 = {pp36[15],pp38[14],pp40[13],pp34[20]};
    CLA_4 KS_3524(s3524, c3524, in3524_1, in3524_2);
    wire[3:0] s3525, in3525_1, in3525_2;
    wire c3525;
    assign in3525_1 = {pp37[14],pp39[13],pp41[12],pp35[19]};
    assign in3525_2 = {pp38[13],pp40[12],pp42[11],pp36[18]};
    CLA_4 KS_3525(s3525, c3525, in3525_1, in3525_2);
    wire[3:0] s3526, in3526_1, in3526_2;
    wire c3526;
    assign in3526_1 = {pp39[12],pp41[11],pp43[10],pp37[17]};
    assign in3526_2 = {pp40[11],pp42[10],pp44[9],pp38[16]};
    CLA_4 KS_3526(s3526, c3526, in3526_1, in3526_2);
    wire[3:0] s3527, in3527_1, in3527_2;
    wire c3527;
    assign in3527_1 = {pp41[10],pp43[9],pp45[8],pp39[15]};
    assign in3527_2 = {pp42[9],pp44[8],pp46[7],pp40[14]};
    CLA_4 KS_3527(s3527, c3527, in3527_1, in3527_2);
    wire[3:0] s3528, in3528_1, in3528_2;
    wire c3528;
    assign in3528_1 = {pp43[8],pp45[7],pp47[6],pp41[13]};
    assign in3528_2 = {pp44[7],pp46[6],pp48[5],pp42[12]};
    CLA_4 KS_3528(s3528, c3528, in3528_1, in3528_2);
    wire[3:0] s3529, in3529_1, in3529_2;
    wire c3529;
    assign in3529_1 = {pp45[6],pp47[5],pp49[4],pp43[11]};
    assign in3529_2 = {pp46[5],pp48[4],pp50[3],pp44[10]};
    CLA_4 KS_3529(s3529, c3529, in3529_1, in3529_2);
    wire[3:0] s3530, in3530_1, in3530_2;
    wire c3530;
    assign in3530_1 = {pp47[4],pp49[3],pp51[2],pp45[9]};
    assign in3530_2 = {pp48[3],pp50[2],pp52[1],pp46[8]};
    CLA_4 KS_3530(s3530, c3530, in3530_1, in3530_2);
    wire[3:0] s3531, in3531_1, in3531_2;
    wire c3531;
    assign in3531_1 = {pp49[2],pp51[1],pp53[0],pp47[7]};
    assign in3531_2 = {pp50[1],pp52[0],c1331,pp48[6]};
    CLA_4 KS_3531(s3531, c3531, in3531_1, in3531_2);
    wire[3:0] s3532, in3532_1, in3532_2;
    wire c3532;
    assign in3532_1 = {pp51[0],c1330,c1332,pp49[5]};
    assign in3532_2 = {c1329,s1331[3],s1333[3],pp50[4]};
    CLA_4 KS_3532(s3532, c3532, in3532_1, in3532_2);
    wire[0:0] s3533, in3533_1, in3533_2;
    wire c3533;
    assign in3533_1 = {s1330[3]};
    assign in3533_2 = {s1331[2]};
    Half_Adder KS_3533(s3533, c3533, in3533_1, in3533_2);
    wire[3:0] s3534, in3534_1, in3534_2;
    wire c3534;
    assign in3534_1 = {s1332[2],s1332[3],s1334[3],pp51[3]};
    assign in3534_2 = {s1333[1],s1333[2],s1335[2],pp52[2]};
    CLA_4 KS_3534(s3534, c3534, in3534_1, in3534_2);
    wire[0:0] s3535, in3535_1, in3535_2;
    wire c3535;
    assign in3535_1 = {s1334[1]};
    assign in3535_2 = {s1335[0]};
    Half_Adder KS_3535(s3535, c3535, in3535_1, in3535_2);
    wire[3:0] s3536, in3536_1, in3536_2;
    wire c3536;
    assign in3536_1 = {s1336[0],s1334[2],s1336[2],pp53[1]};
    assign in3536_2 = {c3494,s1335[1],s1337[1],pp54[0]};
    CLA_4 KS_3536(s3536, c3536, in3536_1, in3536_2);
    wire[0:0] s3537, in3537_1, in3537_2;
    wire c3537;
    assign in3537_1 = {c3495};
    assign in3537_2 = {c3496};
    Half_Adder KS_3537(s3537, c3537, in3537_1, in3537_2);
    wire[1:0] s3538, in3538_1, in3538_2;
    wire c3538;
    assign in3538_1 = {c3497,s1336[1]};
    assign in3538_2 = {c3498,s1337[0]};
    CLA_2 KS_3538(s3538, c3538, in3538_1, in3538_2);
    wire[0:0] s3539, in3539_1, in3539_2;
    wire c3539;
    assign in3539_1 = {c3499};
    assign in3539_2 = {c3500};
    Half_Adder KS_3539(s3539, c3539, in3539_1, in3539_2);
    wire[3:0] s3540, in3540_1, in3540_2;
    wire c3540;
    assign in3540_1 = {c3501,s1338[0],s1338[1],c1333};
    assign in3540_2 = {c3502,s3514[3],s1339[0],c1334};
    CLA_4 KS_3540(s3540, c3540, in3540_1, in3540_2);
    wire[0:0] s3541, in3541_1, in3541_2;
    wire c3541;
    assign in3541_1 = {c3503};
    assign in3541_2 = {c3504};
    Half_Adder KS_3541(s3541, c3541, in3541_1, in3541_2);
    wire[1:0] s3542, in3542_1, in3542_2;
    wire c3542;
    assign in3542_1 = {c3505,s3515[2]};
    assign in3542_2 = {c3507,s3516[2]};
    CLA_2 KS_3542(s3542, c3542, in3542_1, in3542_2);
    wire[0:0] s3543, in3543_1, in3543_2;
    wire c3543;
    assign in3543_1 = {c3509};
    assign in3543_2 = {c3511};
    Half_Adder KS_3543(s3543, c3543, in3543_1, in3543_2);
    wire[3:0] s3544, in3544_1, in3544_2;
    wire c3544;
    assign in3544_1 = {c3513,s3517[2],s1340[0],s1335[3]};
    assign in3544_2 = {s3514[2],s3518[2],s1341[0],s1336[3]};
    CLA_4 KS_3544(s3544, c3544, in3544_1, in3544_2);
    wire[0:0] s3545, in3545_1, in3545_2;
    wire c3545;
    assign in3545_1 = {s3515[1]};
    assign in3545_2 = {s3516[1]};
    Half_Adder KS_3545(s3545, c3545, in3545_1, in3545_2);
    wire[1:0] s3546, in3546_1, in3546_2;
    wire c3546;
    assign in3546_1 = {s3518[1],s3519[1]};
    assign in3546_2 = {s3519[0],s3520[1]};
    CLA_2_c KS_3546(s3546, c3546, in3546_1, in3546_2, s3517[1]);
    wire[3:0] s3547, in3547_1, in3547_2;
    wire c3547;
    assign in3547_1 = {s1337[2],pp25[30],pp27[29],pp33[24]};
    assign in3547_2 = {s1338[2],pp26[29],pp28[28],pp34[23]};
    CLA_4 KS_3547(s3547, c3547, in3547_1, in3547_2);
    wire[3:0] s3548, in3548_1, in3548_2;
    wire c3548;
    assign in3548_1 = {s1339[1],pp27[28],pp29[27],pp35[22]};
    assign in3548_2 = {s1340[1],pp28[27],pp30[26],pp36[21]};
    CLA_4 KS_3548(s3548, c3548, in3548_1, in3548_2);
    wire[3:0] s3549, in3549_1, in3549_2;
    wire c3549;
    assign in3549_1 = {s1342[1],pp29[26],pp31[25],pp37[20]};
    assign in3549_2 = {s1343[0],pp30[25],pp32[24],pp38[19]};
    CLA_4_c KS_3549(s3549, c3549, in3549_1, in3549_2, s1341[1]);
    wire[3:0] s3550, in3550_1, in3550_2;
    wire c3550;
    assign in3550_1 = {pp31[24],pp33[23],pp39[18],pp33[25]};
    assign in3550_2 = {pp32[23],pp34[22],pp40[17],pp34[24]};
    CLA_4 KS_3550(s3550, c3550, in3550_1, in3550_2);
    wire[3:0] s3551, in3551_1, in3551_2;
    wire c3551;
    assign in3551_1 = {pp33[22],pp35[21],pp41[16],pp35[23]};
    assign in3551_2 = {pp34[21],pp36[20],pp42[15],pp36[22]};
    CLA_4 KS_3551(s3551, c3551, in3551_1, in3551_2);
    wire[3:0] s3552, in3552_1, in3552_2;
    wire c3552;
    assign in3552_1 = {pp35[20],pp37[19],pp43[14],pp37[21]};
    assign in3552_2 = {pp36[19],pp38[18],pp44[13],pp38[20]};
    CLA_4 KS_3552(s3552, c3552, in3552_1, in3552_2);
    wire[3:0] s3553, in3553_1, in3553_2;
    wire c3553;
    assign in3553_1 = {pp37[18],pp39[17],pp45[12],pp39[19]};
    assign in3553_2 = {pp38[17],pp40[16],pp46[11],pp40[18]};
    CLA_4 KS_3553(s3553, c3553, in3553_1, in3553_2);
    wire[3:0] s3554, in3554_1, in3554_2;
    wire c3554;
    assign in3554_1 = {pp39[16],pp41[15],pp47[10],pp41[17]};
    assign in3554_2 = {pp40[15],pp42[14],pp48[9],pp42[16]};
    CLA_4 KS_3554(s3554, c3554, in3554_1, in3554_2);
    wire[3:0] s3555, in3555_1, in3555_2;
    wire c3555;
    assign in3555_1 = {pp41[14],pp43[13],pp49[8],pp43[15]};
    assign in3555_2 = {pp42[13],pp44[12],pp50[7],pp44[14]};
    CLA_4 KS_3555(s3555, c3555, in3555_1, in3555_2);
    wire[3:0] s3556, in3556_1, in3556_2;
    wire c3556;
    assign in3556_1 = {pp43[12],pp45[11],pp51[6],pp45[13]};
    assign in3556_2 = {pp44[11],pp46[10],pp52[5],pp46[12]};
    CLA_4 KS_3556(s3556, c3556, in3556_1, in3556_2);
    wire[3:0] s3557, in3557_1, in3557_2;
    wire c3557;
    assign in3557_1 = {pp45[10],pp47[9],pp53[4],pp47[11]};
    assign in3557_2 = {pp46[9],pp48[8],pp54[3],pp48[10]};
    CLA_4 KS_3557(s3557, c3557, in3557_1, in3557_2);
    wire[3:0] s3558, in3558_1, in3558_2;
    wire c3558;
    assign in3558_1 = {pp47[8],pp49[7],pp55[2],pp49[9]};
    assign in3558_2 = {pp48[7],pp50[6],pp56[1],pp50[8]};
    CLA_4 KS_3558(s3558, c3558, in3558_1, in3558_2);
    wire[3:0] s3559, in3559_1, in3559_2;
    wire c3559;
    assign in3559_1 = {pp49[6],pp51[5],pp57[0],pp51[7]};
    assign in3559_2 = {pp50[5],pp52[4],c1339,pp52[6]};
    CLA_4 KS_3559(s3559, c3559, in3559_1, in3559_2);
    wire[3:0] s3560, in3560_1, in3560_2;
    wire c3560;
    assign in3560_1 = {pp51[4],pp53[3],c1340,pp53[5]};
    assign in3560_2 = {pp52[3],pp54[2],c1341,pp54[4]};
    CLA_4 KS_3560(s3560, c3560, in3560_1, in3560_2);
    wire[3:0] s3561, in3561_1, in3561_2;
    wire c3561;
    assign in3561_1 = {pp53[2],pp55[1],c1342,pp55[3]};
    assign in3561_2 = {pp54[1],pp56[0],s1343[3],pp56[2]};
    CLA_4 KS_3561(s3561, c3561, in3561_1, in3561_2);
    wire[3:0] s3562, in3562_1, in3562_2;
    wire c3562;
    assign in3562_1 = {pp55[0],c1337,s1344[3],pp57[1]};
    assign in3562_2 = {c1335,c1338,s1345[3],pp58[0]};
    CLA_4 KS_3562(s3562, c3562, in3562_1, in3562_2);
    wire[3:0] s3563, in3563_1, in3563_2;
    wire c3563;
    assign in3563_1 = {c1336,s1339[3],s1346[2],c1343};
    assign in3563_2 = {s1337[3],s1340[3],s1347[2],c1344};
    CLA_4 KS_3563(s3563, c3563, in3563_1, in3563_2);
    wire[3:0] s3564, in3564_1, in3564_2;
    wire c3564;
    assign in3564_1 = {s1338[3],s1341[3],s1348[2],c1345};
    assign in3564_2 = {s1339[2],s1342[3],s1349[1],s1346[3]};
    CLA_4 KS_3564(s3564, c3564, in3564_1, in3564_2);
    wire[3:0] s3565, in3565_1, in3565_2;
    wire c3565;
    assign in3565_1 = {s1340[2],s1343[2],s1350[1],s1347[3]};
    assign in3565_2 = {s1341[2],s1344[2],s1351[1],s1348[3]};
    CLA_4 KS_3565(s3565, c3565, in3565_1, in3565_2);
    wire[0:0] s3566, in3566_1, in3566_2;
    wire c3566;
    assign in3566_1 = {s1342[2]};
    assign in3566_2 = {s1343[1]};
    Half_Adder KS_3566(s3566, c3566, in3566_1, in3566_2);
    wire[1:0] s3567, in3567_1, in3567_2;
    wire c3567;
    assign in3567_1 = {s1344[1],s1345[2]};
    assign in3567_2 = {s1345[1],s1346[1]};
    CLA_2 KS_3567(s3567, c3567, in3567_1, in3567_2);
    wire[0:0] s3568, in3568_1, in3568_2;
    wire c3568;
    assign in3568_1 = {s1346[0]};
    assign in3568_2 = {s1347[0]};
    Half_Adder KS_3568(s3568, c3568, in3568_1, in3568_2);
    wire[3:0] s3569, in3569_1, in3569_2;
    wire c3569;
    assign in3569_1 = {s1348[0],s1347[1],s1352[0],s1349[2]};
    assign in3569_2 = {c3519,s1348[1],s1353[0],s1350[2]};
    CLA_4 KS_3569(s3569, c3569, in3569_1, in3569_2);
    wire[0:0] s3570, in3570_1, in3570_2;
    wire c3570;
    assign in3570_1 = {c3520};
    assign in3570_2 = {c3521};
    Half_Adder KS_3570(s3570, c3570, in3570_1, in3570_2);
    wire[1:0] s3571, in3571_1, in3571_2;
    wire c3571;
    assign in3571_1 = {c3522,s1349[0]};
    assign in3571_2 = {c3523,s1350[0]};
    CLA_2 KS_3571(s3571, c3571, in3571_1, in3571_2);
    wire[0:0] s3572, in3572_1, in3572_2;
    wire c3572;
    assign in3572_1 = {c3524};
    assign in3572_2 = {c3525};
    Half_Adder KS_3572(s3572, c3572, in3572_1, in3572_2);
    wire[3:0] s3573, in3573_1, in3573_2;
    wire c3573;
    assign in3573_1 = {c3526,s1351[0],s1354[0],s1351[2]};
    assign in3573_2 = {c3527,s3547[2],s1355[0],s1352[1]};
    CLA_4 KS_3573(s3573, c3573, in3573_1, in3573_2);
    wire[0:0] s3574, in3574_1, in3574_2;
    wire c3574;
    assign in3574_1 = {c3528};
    assign in3574_2 = {c3529};
    Half_Adder KS_3574(s3574, c3574, in3574_1, in3574_2);
    wire[1:0] s3575, in3575_1, in3575_2;
    wire c3575;
    assign in3575_1 = {c3530,s3548[2]};
    assign in3575_2 = {c3531,s3549[2]};
    CLA_2 KS_3575(s3575, c3575, in3575_1, in3575_2);
    wire[0:0] s3576, in3576_1, in3576_2;
    wire c3576;
    assign in3576_1 = {c3532};
    assign in3576_2 = {c3534};
    Half_Adder KS_3576(s3576, c3576, in3576_1, in3576_2);
    wire[3:0] s3577, in3577_1, in3577_2;
    wire c3577;
    assign in3577_1 = {c3536,s3550[1],s1356[0],s1353[1]};
    assign in3577_2 = {c3540,s3551[1],s1357[0],s1354[1]};
    CLA_4 KS_3577(s3577, c3577, in3577_1, in3577_2);
    wire[0:0] s3578, in3578_1, in3578_2;
    wire c3578;
    assign in3578_1 = {c3544};
    assign in3578_2 = {s3547[1]};
    Half_Adder KS_3578(s3578, c3578, in3578_1, in3578_2);
    wire[1:0] s3579, in3579_1, in3579_2;
    wire c3579;
    assign in3579_1 = {s3548[1],s3552[1]};
    assign in3579_2 = {s3549[1],s3553[1]};
    CLA_2 KS_3579(s3579, c3579, in3579_1, in3579_2);
    wire[0:0] s3580, in3580_1, in3580_2;
    wire c3580;
    assign in3580_1 = {s3550[0]};
    assign in3580_2 = {s3551[0]};
    Half_Adder KS_3580(s3580, c3580, in3580_1, in3580_2);
    wire[3:0] s3581, in3581_1, in3581_2;
    wire c3581;
    assign in3581_1 = {s3553[0],s3554[1],s1358[0],s1355[1]};
    assign in3581_2 = {s3554[0],s3555[1],s3547[3],s1356[1]};
    CLA_4_c KS_3581(s3581, c3581, in3581_1, in3581_2, s3552[0]);
    wire[3:0] s3582, in3582_1, in3582_2;
    wire c3582;
    assign in3582_1 = {s1357[1],pp35[24],pp37[23],pp47[14]};
    assign in3582_2 = {s1358[1],pp36[23],pp38[22],pp48[13]};
    CLA_4 KS_3582(s3582, c3582, in3582_1, in3582_2);
    wire[3:0] s3583, in3583_1, in3583_2;
    wire c3583;
    assign in3583_1 = {pp37[22],pp39[21],pp49[12],pp42[20]};
    assign in3583_2 = {pp38[21],pp40[20],pp50[11],pp43[19]};
    CLA_4 KS_3583(s3583, c3583, in3583_1, in3583_2);
    wire[3:0] s3584, in3584_1, in3584_2;
    wire c3584;
    assign in3584_1 = {pp39[20],pp41[19],pp51[10],pp44[18]};
    assign in3584_2 = {pp40[19],pp42[18],pp52[9],pp45[17]};
    CLA_4 KS_3584(s3584, c3584, in3584_1, in3584_2);
    wire[3:0] s3585, in3585_1, in3585_2;
    wire c3585;
    assign in3585_1 = {pp41[18],pp43[17],pp53[8],pp46[16]};
    assign in3585_2 = {pp42[17],pp44[16],pp54[7],pp47[15]};
    CLA_4 KS_3585(s3585, c3585, in3585_1, in3585_2);
    wire[3:0] s3586, in3586_1, in3586_2;
    wire c3586;
    assign in3586_1 = {pp43[16],pp45[15],pp55[6],pp48[14]};
    assign in3586_2 = {pp44[15],pp46[14],pp56[5],pp49[13]};
    CLA_4 KS_3586(s3586, c3586, in3586_1, in3586_2);
    wire[3:0] s3587, in3587_1, in3587_2;
    wire c3587;
    assign in3587_1 = {pp45[14],pp47[13],pp57[4],pp50[12]};
    assign in3587_2 = {pp46[13],pp48[12],pp58[3],pp51[11]};
    CLA_4 KS_3587(s3587, c3587, in3587_1, in3587_2);
    wire[3:0] s3588, in3588_1, in3588_2;
    wire c3588;
    assign in3588_1 = {pp47[12],pp49[11],pp59[2],pp52[10]};
    assign in3588_2 = {pp48[11],pp50[10],pp60[1],pp53[9]};
    CLA_4 KS_3588(s3588, c3588, in3588_1, in3588_2);
    wire[3:0] s3589, in3589_1, in3589_2;
    wire c3589;
    assign in3589_1 = {pp49[10],pp51[9],pp61[0],pp54[8]};
    assign in3589_2 = {pp50[9],pp52[8],c1352,pp55[7]};
    CLA_4 KS_3589(s3589, c3589, in3589_1, in3589_2);
    wire[3:0] s3590, in3590_1, in3590_2;
    wire c3590;
    assign in3590_1 = {pp51[8],pp53[7],c1353,pp56[6]};
    assign in3590_2 = {pp52[7],pp54[6],c1354,pp57[5]};
    CLA_4 KS_3590(s3590, c3590, in3590_1, in3590_2);
    wire[3:0] s3591, in3591_1, in3591_2;
    wire c3591;
    assign in3591_1 = {pp53[6],pp55[5],c1355,pp58[4]};
    assign in3591_2 = {pp54[5],pp56[4],c1356,pp59[3]};
    CLA_4 KS_3591(s3591, c3591, in3591_1, in3591_2);
    wire[3:0] s3592, in3592_1, in3592_2;
    wire c3592;
    assign in3592_1 = {pp55[4],pp57[3],c1357,pp60[2]};
    assign in3592_2 = {pp56[3],pp58[2],c1358,pp61[1]};
    CLA_4 KS_3592(s3592, c3592, in3592_1, in3592_2);
    wire[3:0] s3593, in3593_1, in3593_2;
    wire c3593;
    assign in3593_1 = {pp57[2],pp59[1],s1359[3],pp62[0]};
    assign in3593_2 = {pp58[1],pp60[0],s1360[3],c1359};
    CLA_4 KS_3593(s3593, c3593, in3593_1, in3593_2);
    wire[3:0] s3594, in3594_1, in3594_2;
    wire c3594;
    assign in3594_1 = {pp59[0],c1349,s1361[3],c1360};
    assign in3594_2 = {c1346,c1350,s1362[2],c1361};
    CLA_4 KS_3594(s3594, c3594, in3594_1, in3594_2);
    wire[3:0] s3595, in3595_1, in3595_2;
    wire c3595;
    assign in3595_1 = {c1347,c1351,s1363[2],s1362[3]};
    assign in3595_2 = {c1348,s1352[3],s1364[2],s1363[3]};
    CLA_4 KS_3595(s3595, c3595, in3595_1, in3595_2);
    wire[3:0] s3596, in3596_1, in3596_2;
    wire c3596;
    assign in3596_1 = {s1349[3],s1353[3],s1365[2],s1364[3]};
    assign in3596_2 = {s1350[3],s1354[3],s1366[1],s1365[3]};
    CLA_4 KS_3596(s3596, c3596, in3596_1, in3596_2);
    wire[3:0] s3597, in3597_1, in3597_2;
    wire c3597;
    assign in3597_1 = {s1351[3],s1355[3],s1367[1],s1366[2]};
    assign in3597_2 = {s1352[2],s1356[3],s1368[1],s1367[2]};
    CLA_4 KS_3597(s3597, c3597, in3597_1, in3597_2);
    wire[3:0] s3598, in3598_1, in3598_2;
    wire c3598;
    assign in3598_1 = {s1353[2],s1357[3],s1369[1],s1368[2]};
    assign in3598_2 = {s1354[2],s1358[3],s1370[0],s1369[2]};
    CLA_4 KS_3598(s3598, c3598, in3598_1, in3598_2);
    wire[3:0] s3599, in3599_1, in3599_2;
    wire c3599;
    assign in3599_1 = {s1355[2],s1359[2],s1371[0],s1370[1]};
    assign in3599_2 = {s1356[2],s1360[2],s1372[0],s1371[1]};
    CLA_4 KS_3599(s3599, c3599, in3599_1, in3599_2);
    wire[3:0] s3600, in3600_1, in3600_2;
    wire c3600;
    assign in3600_1 = {s1357[2],s1361[2],s1373[0],s1372[1]};
    assign in3600_2 = {s1358[2],s1362[1],s1374[0],s1373[1]};
    CLA_4 KS_3600(s3600, c3600, in3600_1, in3600_2);
    wire[0:0] s3601, in3601_1, in3601_2;
    wire c3601;
    assign in3601_1 = {s1359[1]};
    assign in3601_2 = {s1360[1]};
    Half_Adder KS_3601(s3601, c3601, in3601_1, in3601_2);
    wire[1:0] s3602, in3602_1, in3602_2;
    wire c3602;
    assign in3602_1 = {s1361[1],s1363[1]};
    assign in3602_2 = {s1362[0],s1364[1]};
    CLA_2 KS_3602(s3602, c3602, in3602_1, in3602_2);
    wire[0:0] s3603, in3603_1, in3603_2;
    wire c3603;
    assign in3603_1 = {s1363[0]};
    assign in3603_2 = {s1364[0]};
    Half_Adder KS_3603(s3603, c3603, in3603_1, in3603_2);
    wire[3:0] s3604, in3604_1, in3604_2;
    wire c3604;
    assign in3604_1 = {s1365[0],s1365[1],s1375[0],s1374[1]};
    assign in3604_2 = {c3550,s1366[0],s1376[0],s1375[1]};
    CLA_4 KS_3604(s3604, c3604, in3604_1, in3604_2);
    wire[0:0] s3605, in3605_1, in3605_2;
    wire c3605;
    assign in3605_1 = {c3551};
    assign in3605_2 = {c3552};
    Half_Adder KS_3605(s3605, c3605, in3605_1, in3605_2);
    wire[1:0] s3606, in3606_1, in3606_2;
    wire c3606;
    assign in3606_1 = {c3553,s1367[0]};
    assign in3606_2 = {c3554,s1368[0]};
    CLA_2 KS_3606(s3606, c3606, in3606_1, in3606_2);
    wire[0:0] s3607, in3607_1, in3607_2;
    wire c3607;
    assign in3607_1 = {c3555};
    assign in3607_2 = {c3556};
    Half_Adder KS_3607(s3607, c3607, in3607_1, in3607_2);
    wire[3:0] s3608, in3608_1, in3608_2;
    wire c3608;
    assign in3608_1 = {c3557,s1369[0],s1377[0],s1376[1]};
    assign in3608_2 = {c3558,s3582[2],s1378[0],s1377[1]};
    CLA_4 KS_3608(s3608, c3608, in3608_1, in3608_2);
    wire[0:0] s3609, in3609_1, in3609_2;
    wire c3609;
    assign in3609_1 = {c3559};
    assign in3609_2 = {c3560};
    Half_Adder KS_3609(s3609, c3609, in3609_1, in3609_2);
    wire[1:0] s3610, in3610_1, in3610_2;
    wire c3610;
    assign in3610_1 = {c3561,s3583[1]};
    assign in3610_2 = {c3562,s3584[1]};
    CLA_2 KS_3610(s3610, c3610, in3610_1, in3610_2);
    wire[0:0] s3611, in3611_1, in3611_2;
    wire c3611;
    assign in3611_1 = {c3563};
    assign in3611_2 = {c3564};
    Half_Adder KS_3611(s3611, c3611, in3611_1, in3611_2);
    wire[2:0] s3612, in3612_1, in3612_2;
    wire c3612;
    assign in3612_1 = {c3565,s3585[1],s1379[0]};
    assign in3612_2 = {c3569,s3586[1],s1380[0]};
    CLA_3 KS_3612(s3612, c3612, in3612_1, in3612_2);
    wire[0:0] s3613, in3613_1, in3613_2;
    wire c3613;
    assign in3613_1 = {c3573};
    assign in3613_2 = {c3577};
    Half_Adder KS_3613(s3613, c3613, in3613_1, in3613_2);
    wire[1:0] s3614, in3614_1, in3614_2;
    wire c3614;
    assign in3614_1 = {c3581,s3587[1]};
    assign in3614_2 = {s3582[1],s3588[1]};
    CLA_2 KS_3614(s3614, c3614, in3614_1, in3614_2);
    wire[0:0] s3615, in3615_1, in3615_2;
    wire c3615;
    assign in3615_1 = {s3583[0]};
    assign in3615_2 = {s3584[0]};
    Half_Adder KS_3615(s3615, c3615, in3615_1, in3615_2);
    wire[3:0] s3616, in3616_1, in3616_2;
    wire c3616;
    assign in3616_1 = {s3585[0],s3589[1],s1381[0],s1378[1]};
    assign in3616_2 = {s3586[0],s3590[1],s3582[3],s1379[1]};
    CLA_4 KS_3616(s3616, c3616, in3616_1, in3616_2);
    wire[0:0] s3617, in3617_1, in3617_2;
    wire c3617;
    assign in3617_1 = {s3587[0]};
    assign in3617_2 = {s3588[0]};
    Half_Adder KS_3617(s3617, c3617, in3617_1, in3617_2);
    wire[1:0] s3618, in3618_1, in3618_2;
    wire c3618;
    assign in3618_1 = {s3590[0],s3591[1]};
    assign in3618_2 = {s3591[0],s3592[1]};
    CLA_2_c KS_3618(s3618, c3618, in3618_1, in3618_2, s3589[0]);
    wire[3:0] s3619, in3619_1, in3619_2;
    wire c3619;
    assign in3619_1 = {pp45[18],pp47[17],pp65[0],pp54[12]};
    assign in3619_2 = {pp46[17],pp48[16],c1370,pp55[11]};
    CLA_4 KS_3619(s3619, c3619, in3619_1, in3619_2);
    wire[3:0] s3620, in3620_1, in3620_2;
    wire c3620;
    assign in3620_1 = {pp47[16],pp49[15],c1371,pp56[10]};
    assign in3620_2 = {pp48[15],pp50[14],c1372,pp57[9]};
    CLA_4 KS_3620(s3620, c3620, in3620_1, in3620_2);
    wire[3:0] s3621, in3621_1, in3621_2;
    wire c3621;
    assign in3621_1 = {pp49[14],pp51[13],c1373,pp58[8]};
    assign in3621_2 = {pp50[13],pp52[12],c1374,pp59[7]};
    CLA_4 KS_3621(s3621, c3621, in3621_1, in3621_2);
    wire[3:0] s3622, in3622_1, in3622_2;
    wire c3622;
    assign in3622_1 = {pp51[12],pp53[11],c1375,pp60[6]};
    assign in3622_2 = {pp52[11],pp54[10],c1376,pp61[5]};
    CLA_4 KS_3622(s3622, c3622, in3622_1, in3622_2);
    wire[3:0] s3623, in3623_1, in3623_2;
    wire c3623;
    assign in3623_1 = {pp53[10],pp55[9],c1377,pp62[4]};
    assign in3623_2 = {pp54[9],pp56[8],c1378,pp63[3]};
    CLA_4 KS_3623(s3623, c3623, in3623_1, in3623_2);
    wire[3:0] s3624, in3624_1, in3624_2;
    wire c3624;
    assign in3624_1 = {pp55[8],pp57[7],c1379,pp64[2]};
    assign in3624_2 = {pp56[7],pp58[6],c1380,pp65[1]};
    CLA_4 KS_3624(s3624, c3624, in3624_1, in3624_2);
    wire[3:0] s3625, in3625_1, in3625_2;
    wire c3625;
    assign in3625_1 = {pp57[6],pp59[5],c1381,pp66[0]};
    assign in3625_2 = {pp58[5],pp60[4],s1382[3],c1382};
    CLA_4 KS_3625(s3625, c3625, in3625_1, in3625_2);
    wire[3:0] s3626, in3626_1, in3626_2;
    wire c3626;
    assign in3626_1 = {pp59[4],pp61[3],s1383[2],s1383[3]};
    assign in3626_2 = {pp60[3],pp62[2],s1384[2],s1384[3]};
    CLA_4 KS_3626(s3626, c3626, in3626_1, in3626_2);
    wire[3:0] s3627, in3627_1, in3627_2;
    wire c3627;
    assign in3627_1 = {pp61[2],pp63[1],s1385[2],s1385[3]};
    assign in3627_2 = {pp62[1],pp64[0],s1386[2],s1386[3]};
    CLA_4 KS_3627(s3627, c3627, in3627_1, in3627_2);
    wire[3:0] s3628, in3628_1, in3628_2;
    wire c3628;
    assign in3628_1 = {pp63[0],c1366,s1387[2],s1387[3]};
    assign in3628_2 = {c1362,c1367,s1388[1],s1388[2]};
    CLA_4 KS_3628(s3628, c3628, in3628_1, in3628_2);
    wire[3:0] s3629, in3629_1, in3629_2;
    wire c3629;
    assign in3629_1 = {c1363,c1368,s1389[1],s1389[2]};
    assign in3629_2 = {c1364,c1369,s1390[1],s1390[2]};
    CLA_4 KS_3629(s3629, c3629, in3629_1, in3629_2);
    wire[3:0] s3630, in3630_1, in3630_2;
    wire c3630;
    assign in3630_1 = {c1365,s1370[3],s1391[1],s1391[2]};
    assign in3630_2 = {s1366[3],s1371[3],s1392[1],s1392[2]};
    CLA_4 KS_3630(s3630, c3630, in3630_1, in3630_2);
    wire[3:0] s3631, in3631_1, in3631_2;
    wire c3631;
    assign in3631_1 = {s1367[3],s1372[3],s1393[0],s1393[1]};
    assign in3631_2 = {s1368[3],s1373[3],s1394[0],s1394[1]};
    CLA_4 KS_3631(s3631, c3631, in3631_1, in3631_2);
    wire[3:0] s3632, in3632_1, in3632_2;
    wire c3632;
    assign in3632_1 = {s1369[3],s1374[3],s1395[0],s1395[1]};
    assign in3632_2 = {s1370[2],s1375[3],s1396[0],s1396[1]};
    CLA_4 KS_3632(s3632, c3632, in3632_1, in3632_2);
    wire[3:0] s3633, in3633_1, in3633_2;
    wire c3633;
    assign in3633_1 = {s1371[2],s1376[3],s1397[0],s1397[1]};
    assign in3633_2 = {s1372[2],s1377[3],s1398[0],s1398[1]};
    CLA_4 KS_3633(s3633, c3633, in3633_1, in3633_2);
    wire[3:0] s3634, in3634_1, in3634_2;
    wire c3634;
    assign in3634_1 = {s1373[2],s1378[3],s1399[0],s1399[1]};
    assign in3634_2 = {s1374[2],s1379[3],s1400[0],s1400[1]};
    CLA_4 KS_3634(s3634, c3634, in3634_1, in3634_2);
    wire[3:0] s3635, in3635_1, in3635_2;
    wire c3635;
    assign in3635_1 = {s1375[2],s1380[3],s1401[0],s1401[1]};
    assign in3635_2 = {s1376[2],s1381[3],s1402[0],s1402[1]};
    CLA_4 KS_3635(s3635, c3635, in3635_1, in3635_2);
    wire[3:0] s3636, in3636_1, in3636_2;
    wire c3636;
    assign in3636_1 = {s1377[2],s1382[2],s1403[0],s1403[1]};
    assign in3636_2 = {s1378[2],s1383[1],s1404[0],s1404[1]};
    CLA_4 KS_3636(s3636, c3636, in3636_1, in3636_2);
    wire[3:0] s3637, in3637_1, in3637_2;
    wire c3637;
    assign in3637_1 = {s1379[2],s1384[1],s1405[0],s1405[1]};
    assign in3637_2 = {s1380[2],s1385[1],s1406[0],s1406[1]};
    CLA_4 KS_3637(s3637, c3637, in3637_1, in3637_2);
    wire[0:0] s3638, in3638_1, in3638_2;
    wire c3638;
    assign in3638_1 = {s1381[2]};
    assign in3638_2 = {s1382[1]};
    Half_Adder KS_3638(s3638, c3638, in3638_1, in3638_2);
    wire[1:0] s3639, in3639_1, in3639_2;
    wire c3639;
    assign in3639_1 = {s1383[0],s1386[1]};
    assign in3639_2 = {s1384[0],s1387[1]};
    CLA_2 KS_3639(s3639, c3639, in3639_1, in3639_2);
    wire[0:0] s3640, in3640_1, in3640_2;
    wire c3640;
    assign in3640_1 = {s1385[0]};
    assign in3640_2 = {s1386[0]};
    Half_Adder KS_3640(s3640, c3640, in3640_1, in3640_2);
    wire[2:0] s3641, in3641_1, in3641_2;
    wire c3641;
    assign in3641_1 = {s1387[0],s1388[0],s1407[0]};
    assign in3641_2 = {c3583,s1389[0],s1408[0]};
    CLA_3 KS_3641(s3641, c3641, in3641_1, in3641_2);
    wire[0:0] s3642, in3642_1, in3642_2;
    wire c3642;
    assign in3642_1 = {c3584};
    assign in3642_2 = {c3585};
    Half_Adder KS_3642(s3642, c3642, in3642_1, in3642_2);
    wire[1:0] s3643, in3643_1, in3643_2;
    wire c3643;
    assign in3643_1 = {c3586,s1390[0]};
    assign in3643_2 = {c3587,s1391[0]};
    CLA_2 KS_3643(s3643, c3643, in3643_1, in3643_2);
    wire[0:0] s3644, in3644_1, in3644_2;
    wire c3644;
    assign in3644_1 = {c3588};
    assign in3644_2 = {c3589};
    Half_Adder KS_3644(s3644, c3644, in3644_1, in3644_2);
    wire[3:0] s3645, in3645_1, in3645_2;
    wire c3645;
    assign in3645_1 = {c3590,s1392[0],s1409[0],c1407};
    assign in3645_2 = {c3591,s3619[1],s1410[0],s1408[1]};
    CLA_4 KS_3645(s3645, c3645, in3645_1, in3645_2);
    wire[0:0] s3646, in3646_1, in3646_2;
    wire c3646;
    assign in3646_1 = {c3592};
    assign in3646_2 = {c3593};
    Half_Adder KS_3646(s3646, c3646, in3646_1, in3646_2);
    wire[1:0] s3647, in3647_1, in3647_2;
    wire c3647;
    assign in3647_1 = {c3594,s3620[1]};
    assign in3647_2 = {c3595,s3621[1]};
    CLA_2 KS_3647(s3647, c3647, in3647_1, in3647_2);
    wire[0:0] s3648, in3648_1, in3648_2;
    wire c3648;
    assign in3648_1 = {c3596};
    assign in3648_2 = {c3597};
    Half_Adder KS_3648(s3648, c3648, in3648_1, in3648_2);
    wire[2:0] s3649, in3649_1, in3649_2;
    wire c3649;
    assign in3649_1 = {c3598,s3622[1],s1411[0]};
    assign in3649_2 = {c3599,s3623[1],s1412[0]};
    CLA_3 KS_3649(s3649, c3649, in3649_1, in3649_2);
    wire[0:0] s3650, in3650_1, in3650_2;
    wire c3650;
    assign in3650_1 = {c3600};
    assign in3650_2 = {c3604};
    Half_Adder KS_3650(s3650, c3650, in3650_1, in3650_2);
    wire[1:0] s3651, in3651_1, in3651_2;
    wire c3651;
    assign in3651_1 = {c3608,s3624[1]};
    assign in3651_2 = {c3616,s3625[1]};
    CLA_2 KS_3651(s3651, c3651, in3651_1, in3651_2);
    wire[0:0] s3652, in3652_1, in3652_2;
    wire c3652;
    assign in3652_1 = {s3619[0]};
    assign in3652_2 = {s3620[0]};
    Half_Adder KS_3652(s3652, c3652, in3652_1, in3652_2);
    wire[3:0] s3653, in3653_1, in3653_2;
    wire c3653;
    assign in3653_1 = {s3621[0],s3626[1],s1413[0],c1409};
    assign in3653_2 = {s3622[0],s3627[1],s3619[2],s1410[1]};
    CLA_4 KS_3653(s3653, c3653, in3653_1, in3653_2);
    wire[0:0] s3654, in3654_1, in3654_2;
    wire c3654;
    assign in3654_1 = {s3623[0]};
    assign in3654_2 = {s3624[0]};
    Half_Adder KS_3654(s3654, c3654, in3654_1, in3654_2);
    wire[1:0] s3655, in3655_1, in3655_2;
    wire c3655;
    assign in3655_1 = {s3625[0],s3628[1]};
    assign in3655_2 = {s3626[0],s3629[1]};
    CLA_2 KS_3655(s3655, c3655, in3655_1, in3655_2);
    wire[0:0] s3656, in3656_1, in3656_2;
    wire c3656;
    assign in3656_1 = {s3628[0]};
    assign in3656_2 = {s3629[0]};
    Full_Adder KS_3656(s3656, c3656, in3656_1, in3656_2, s3627[0]);
    wire[3:0] s3657, in3657_1, in3657_2;
    wire c3657;
    assign in3657_1 = {pp55[12],pp57[11],c1406,pp68[2]};
    assign in3657_2 = {pp56[11],pp58[10],c1408,pp69[1]};
    CLA_4 KS_3657(s3657, c3657, in3657_1, in3657_2);
    wire[3:0] s3658, in3658_1, in3658_2;
    wire c3658;
    assign in3658_1 = {pp57[10],pp59[9],c1410,pp70[0]};
    assign in3658_2 = {pp58[9],pp60[8],c1412,s1414[3]};
    CLA_4 KS_3658(s3658, c3658, in3658_1, in3658_2);
    wire[3:0] s3659, in3659_1, in3659_2;
    wire c3659;
    assign in3659_1 = {pp59[8],pp61[7],s1414[2],s1415[3]};
    assign in3659_2 = {pp60[7],pp62[6],s1415[2],s1416[3]};
    CLA_4 KS_3659(s3659, c3659, in3659_1, in3659_2);
    wire[3:0] s3660, in3660_1, in3660_2;
    wire c3660;
    assign in3660_1 = {pp61[6],pp63[5],s1416[2],s1417[3]};
    assign in3660_2 = {pp62[5],pp64[4],s1417[2],s1418[3]};
    CLA_4 KS_3660(s3660, c3660, in3660_1, in3660_2);
    wire[3:0] s3661, in3661_1, in3661_2;
    wire c3661;
    assign in3661_1 = {pp63[4],pp65[3],s1418[2],s1419[2]};
    assign in3661_2 = {pp64[3],pp66[2],s1419[1],s1420[2]};
    CLA_4 KS_3661(s3661, c3661, in3661_1, in3661_2);
    wire[3:0] s3662, in3662_1, in3662_2;
    wire c3662;
    assign in3662_1 = {pp65[2],pp67[1],s1420[1],s1421[2]};
    assign in3662_2 = {pp66[1],pp68[0],s1421[1],s1422[2]};
    CLA_4 KS_3662(s3662, c3662, in3662_1, in3662_2);
    wire[3:0] s3663, in3663_1, in3663_2;
    wire c3663;
    assign in3663_1 = {pp67[0],c1388,s1422[1],s1423[2]};
    assign in3663_2 = {c1383,c1389,s1423[1],s1424[2]};
    CLA_4 KS_3663(s3663, c3663, in3663_1, in3663_2);
    wire[3:0] s3664, in3664_1, in3664_2;
    wire c3664;
    assign in3664_1 = {c1384,c1390,s1424[1],s1425[1]};
    assign in3664_2 = {c1385,c1391,s1425[0],s1426[1]};
    CLA_4 KS_3664(s3664, c3664, in3664_1, in3664_2);
    wire[3:0] s3665, in3665_1, in3665_2;
    wire c3665;
    assign in3665_1 = {c1386,c1392,s1426[0],s1427[1]};
    assign in3665_2 = {c1387,s1393[3],s1427[0],s1428[1]};
    CLA_4 KS_3665(s3665, c3665, in3665_1, in3665_2);
    wire[3:0] s3666, in3666_1, in3666_2;
    wire c3666;
    assign in3666_1 = {s1388[3],s1394[3],s1428[0],s1429[1]};
    assign in3666_2 = {s1389[3],s1395[3],s1429[0],s1430[1]};
    CLA_4 KS_3666(s3666, c3666, in3666_1, in3666_2);
    wire[3:0] s3667, in3667_1, in3667_2;
    wire c3667;
    assign in3667_1 = {s1390[3],s1396[3],s1430[0],s1431[1]};
    assign in3667_2 = {s1391[3],s1397[3],s1431[0],s1432[1]};
    CLA_4 KS_3667(s3667, c3667, in3667_1, in3667_2);
    wire[3:0] s3668, in3668_1, in3668_2;
    wire c3668;
    assign in3668_1 = {s1392[3],s1398[3],s1432[0],s1433[1]};
    assign in3668_2 = {s1393[2],s1399[3],s1433[0],s1434[1]};
    CLA_4 KS_3668(s3668, c3668, in3668_1, in3668_2);
    wire[3:0] s3669, in3669_1, in3669_2;
    wire c3669;
    assign in3669_1 = {s1394[2],s1400[3],s1434[0],s1435[1]};
    assign in3669_2 = {s1395[2],s1401[3],s1435[0],s1436[1]};
    CLA_4 KS_3669(s3669, c3669, in3669_1, in3669_2);
    wire[3:0] s3670, in3670_1, in3670_2;
    wire c3670;
    assign in3670_1 = {s1396[2],s1402[3],s1436[0],s1437[1]};
    assign in3670_2 = {s1397[2],s1403[3],s1437[0],s1438[1]};
    CLA_4 KS_3670(s3670, c3670, in3670_1, in3670_2);
    wire[3:0] s3671, in3671_1, in3671_2;
    wire c3671;
    assign in3671_1 = {s1398[2],s1404[3],s1438[0],s1439[1]};
    assign in3671_2 = {s1399[2],s1405[3],s1439[0],s1440[1]};
    CLA_4 KS_3671(s3671, c3671, in3671_1, in3671_2);
    wire[3:0] s3672, in3672_1, in3672_2;
    wire c3672;
    assign in3672_1 = {s1400[2],s1406[3],s1440[0],c1441};
    assign in3672_2 = {s1401[2],s1408[3],s1441[0],s1442[1]};
    CLA_4 KS_3672(s3672, c3672, in3672_1, in3672_2);
    wire[3:0] s3673, in3673_1, in3673_2;
    wire c3673;
    assign in3673_1 = {s1402[2],s1410[3],s1442[0],c1443};
    assign in3673_2 = {s1403[2],s1412[3],s1443[0],s1444[1]};
    CLA_4 KS_3673(s3673, c3673, in3673_1, in3673_2);
    wire[3:0] s3674, in3674_1, in3674_2;
    wire c3674;
    assign in3674_1 = {s1404[2],s1414[1],s1444[0],c1445};
    assign in3674_2 = {s1405[2],s1415[1],s1445[0],s1446[1]};
    CLA_4 KS_3674(s3674, c3674, in3674_1, in3674_2);
    wire[2:0] s3675, in3675_1, in3675_2;
    wire c3675;
    assign in3675_1 = {s1406[2],s1416[1],s1446[0]};
    assign in3675_2 = {s1408[2],s1417[1],s1447[0]};
    CLA_3 KS_3675(s3675, c3675, in3675_1, in3675_2);
    wire[0:0] s3676, in3676_1, in3676_2;
    wire c3676;
    assign in3676_1 = {s1410[2]};
    assign in3676_2 = {s1412[2]};
    Half_Adder KS_3676(s3676, c3676, in3676_1, in3676_2);
    wire[1:0] s3677, in3677_1, in3677_2;
    wire c3677;
    assign in3677_1 = {s1414[0],s1418[1]};
    assign in3677_2 = {s1415[0],s1419[0]};
    CLA_2 KS_3677(s3677, c3677, in3677_1, in3677_2);
    wire[0:0] s3678, in3678_1, in3678_2;
    wire c3678;
    assign in3678_1 = {s1416[0]};
    assign in3678_2 = {s1417[0]};
    Half_Adder KS_3678(s3678, c3678, in3678_1, in3678_2);
    wire[3:0] s3679, in3679_1, in3679_2;
    wire c3679;
    assign in3679_1 = {s1418[0],s1420[0],s1448[0],c1447};
    assign in3679_2 = {c3619,s1421[0],s1449[0],s1448[1]};
    CLA_4 KS_3679(s3679, c3679, in3679_1, in3679_2);
    wire[0:0] s3680, in3680_1, in3680_2;
    wire c3680;
    assign in3680_1 = {c3620};
    assign in3680_2 = {c3621};
    Half_Adder KS_3680(s3680, c3680, in3680_1, in3680_2);
    wire[1:0] s3681, in3681_1, in3681_2;
    wire c3681;
    assign in3681_1 = {c3622,s1422[0]};
    assign in3681_2 = {c3623,s1423[0]};
    CLA_2 KS_3681(s3681, c3681, in3681_1, in3681_2);
    wire[0:0] s3682, in3682_1, in3682_2;
    wire c3682;
    assign in3682_1 = {c3624};
    assign in3682_2 = {c3625};
    Half_Adder KS_3682(s3682, c3682, in3682_1, in3682_2);
    wire[2:0] s3683, in3683_1, in3683_2;
    wire c3683;
    assign in3683_1 = {c3626,s1424[0],s1450[0]};
    assign in3683_2 = {c3627,s3657[1],s1451[0]};
    CLA_3 KS_3683(s3683, c3683, in3683_1, in3683_2);
    wire[0:0] s3684, in3684_1, in3684_2;
    wire c3684;
    assign in3684_1 = {c3628};
    assign in3684_2 = {c3629};
    Half_Adder KS_3684(s3684, c3684, in3684_1, in3684_2);
    wire[1:0] s3685, in3685_1, in3685_2;
    wire c3685;
    assign in3685_1 = {c3630,s3658[1]};
    assign in3685_2 = {c3631,s3659[1]};
    CLA_2 KS_3685(s3685, c3685, in3685_1, in3685_2);
    wire[0:0] s3686, in3686_1, in3686_2;
    wire c3686;
    assign in3686_1 = {c3632};
    assign in3686_2 = {c3633};
    Half_Adder KS_3686(s3686, c3686, in3686_1, in3686_2);
    wire[3:0] s3687, in3687_1, in3687_2;
    wire c3687;
    assign in3687_1 = {c3634,s3660[1],s1452[0],c1449};
    assign in3687_2 = {c3635,s3661[1],s1453[0],s1450[1]};
    CLA_4 KS_3687(s3687, c3687, in3687_1, in3687_2);
    wire[0:0] s3688, in3688_1, in3688_2;
    wire c3688;
    assign in3688_1 = {c3636};
    assign in3688_2 = {c3637};
    Half_Adder KS_3688(s3688, c3688, in3688_1, in3688_2);
    wire[1:0] s3689, in3689_1, in3689_2;
    wire c3689;
    assign in3689_1 = {c3645,s3662[1]};
    assign in3689_2 = {c3653,s3663[1]};
    CLA_2 KS_3689(s3689, c3689, in3689_1, in3689_2);
    wire[0:0] s3690, in3690_1, in3690_2;
    wire c3690;
    assign in3690_1 = {s3657[0]};
    assign in3690_2 = {s3658[0]};
    Half_Adder KS_3690(s3690, c3690, in3690_1, in3690_2);
    wire[2:0] s3691, in3691_1, in3691_2;
    wire c3691;
    assign in3691_1 = {s3659[0],s3664[1],s1454[0]};
    assign in3691_2 = {s3660[0],s3665[1],s3657[2]};
    CLA_3 KS_3691(s3691, c3691, in3691_1, in3691_2);
    wire[0:0] s3692, in3692_1, in3692_2;
    wire c3692;
    assign in3692_1 = {s3661[0]};
    assign in3692_2 = {s3662[0]};
    Half_Adder KS_3692(s3692, c3692, in3692_1, in3692_2);
    wire[1:0] s3693, in3693_1, in3693_2;
    wire c3693;
    assign in3693_1 = {s3663[0],s3666[1]};
    assign in3693_2 = {s3664[0],s3667[1]};
    CLA_2 KS_3693(s3693, c3693, in3693_1, in3693_2);
    wire[0:0] s3694, in3694_1, in3694_2;
    wire c3694;
    assign in3694_1 = {s3666[0]};
    assign in3694_2 = {s3667[0]};
    Full_Adder KS_3694(s3694, c3694, in3694_1, in3694_2, s3665[0]);
    wire[3:0] s3695, in3695_1, in3695_2;
    wire c3695;
    assign in3695_1 = {pp63[8],pp67[5],s1461[1],s1462[2]};
    assign in3695_2 = {pp64[7],pp68[4],s1462[1],s1463[2]};
    CLA_4 KS_3695(s3695, c3695, in3695_1, in3695_2);
    wire[3:0] s3696, in3696_1, in3696_2;
    wire c3696;
    assign in3696_1 = {pp65[6],pp69[3],s1463[1],s1464[2]};
    assign in3696_2 = {pp66[5],pp70[2],s1464[1],s1465[1]};
    CLA_4 KS_3696(s3696, c3696, in3696_1, in3696_2);
    wire[3:0] s3697, in3697_1, in3697_2;
    wire c3697;
    assign in3697_1 = {pp67[4],pp71[1],s1465[0],s1466[1]};
    assign in3697_2 = {pp68[3],pp72[0],s1466[0],s1467[1]};
    CLA_4 KS_3697(s3697, c3697, in3697_1, in3697_2);
    wire[3:0] s3698, in3698_1, in3698_2;
    wire c3698;
    assign in3698_1 = {pp69[2],c1419,s1467[0],s1468[1]};
    assign in3698_2 = {pp70[1],c1420,s1468[0],s1469[1]};
    CLA_4 KS_3698(s3698, c3698, in3698_1, in3698_2);
    wire[3:0] s3699, in3699_1, in3699_2;
    wire c3699;
    assign in3699_1 = {pp71[0],c1421,s1469[0],s1470[1]};
    assign in3699_2 = {c1414,c1422,s1470[0],s1471[1]};
    CLA_4 KS_3699(s3699, c3699, in3699_1, in3699_2);
    wire[3:0] s3700, in3700_1, in3700_2;
    wire c3700;
    assign in3700_1 = {c1415,c1423,s1471[0],s1472[1]};
    assign in3700_2 = {c1416,c1424,s1472[0],s1473[1]};
    CLA_4 KS_3700(s3700, c3700, in3700_1, in3700_2);
    wire[3:0] s3701, in3701_1, in3701_2;
    wire c3701;
    assign in3701_1 = {c1417,s1425[3],s1473[0],s1474[1]};
    assign in3701_2 = {c1418,s1426[3],s1474[0],s1475[1]};
    CLA_4 KS_3701(s3701, c3701, in3701_1, in3701_2);
    wire[3:0] s3702, in3702_1, in3702_2;
    wire c3702;
    assign in3702_1 = {s1419[3],s1427[3],s1475[0],s1476[1]};
    assign in3702_2 = {s1420[3],s1428[3],s1476[0],s1477[1]};
    CLA_4 KS_3702(s3702, c3702, in3702_1, in3702_2);
    wire[3:0] s3703, in3703_1, in3703_2;
    wire c3703;
    assign in3703_1 = {s1421[3],s1429[3],s1477[0],s1478[1]};
    assign in3703_2 = {s1422[3],s1430[3],s1478[0],s1479[1]};
    CLA_4 KS_3703(s3703, c3703, in3703_1, in3703_2);
    wire[3:0] s3704, in3704_1, in3704_2;
    wire c3704;
    assign in3704_1 = {s1423[3],s1431[3],s1479[0],s1480[1]};
    assign in3704_2 = {s1424[3],s1432[3],s1480[0],s1481[1]};
    CLA_4 KS_3704(s3704, c3704, in3704_1, in3704_2);
    wire[3:0] s3705, in3705_1, in3705_2;
    wire c3705;
    assign in3705_1 = {s1425[2],s1433[3],s1481[0],s1482[1]};
    assign in3705_2 = {s1426[2],s1434[3],s1482[0],s1483[1]};
    CLA_4 KS_3705(s3705, c3705, in3705_1, in3705_2);
    wire[3:0] s3706, in3706_1, in3706_2;
    wire c3706;
    assign in3706_1 = {s1427[2],s1435[3],s1483[0],s1484[1]};
    assign in3706_2 = {s1428[2],s1436[3],s1484[0],s1485[1]};
    CLA_4 KS_3706(s3706, c3706, in3706_1, in3706_2);
    wire[3:0] s3707, in3707_1, in3707_2;
    wire c3707;
    assign in3707_1 = {s1429[2],s1437[3],s1485[0],c1486};
    assign in3707_2 = {s1430[2],s1438[3],s1486[0],s1487[1]};
    CLA_4 KS_3707(s3707, c3707, in3707_1, in3707_2);
    wire[3:0] s3708, in3708_1, in3708_2;
    wire c3708;
    assign in3708_1 = {s1431[2],s1439[3],s1487[0],c1488};
    assign in3708_2 = {s1432[2],s1440[3],s1488[0],s1489[1]};
    CLA_4 KS_3708(s3708, c3708, in3708_1, in3708_2);
    wire[3:0] s3709, in3709_1, in3709_2;
    wire c3709;
    assign in3709_1 = {s1433[2],s1442[3],s1489[0],c1490};
    assign in3709_2 = {s1434[2],s1444[3],s1490[0],s1491[1]};
    CLA_4 KS_3709(s3709, c3709, in3709_1, in3709_2);
    wire[3:0] s3710, in3710_1, in3710_2;
    wire c3710;
    assign in3710_1 = {s1435[2],s1446[3],s1491[0],c1492};
    assign in3710_2 = {s1436[2],s1448[3],s1492[0],s1493[1]};
    CLA_4 KS_3710(s3710, c3710, in3710_1, in3710_2);
    wire[3:0] s3711, in3711_1, in3711_2;
    wire c3711;
    assign in3711_1 = {s1437[2],s1450[3],s1493[0],c1494};
    assign in3711_2 = {s1438[2],s1452[3],s1494[0],s1495[1]};
    CLA_4 KS_3711(s3711, c3711, in3711_1, in3711_2);
    wire[3:0] s3712, in3712_1, in3712_2;
    wire c3712;
    assign in3712_1 = {s1439[2],s1454[3],s1495[0],c1496};
    assign in3712_2 = {s1440[2],s1455[1],s1496[0],s1497[1]};
    CLA_4 KS_3712(s3712, c3712, in3712_1, in3712_2);
    wire[2:0] s3713, in3713_1, in3713_2;
    wire c3713;
    assign in3713_1 = {s1442[2],s1456[1],s1497[0]};
    assign in3713_2 = {s1444[2],s1457[0],s1498[0]};
    CLA_3 KS_3713(s3713, c3713, in3713_1, in3713_2);
    wire[0:0] s3714, in3714_1, in3714_2;
    wire c3714;
    assign in3714_1 = {s1446[2]};
    assign in3714_2 = {s1448[2]};
    Half_Adder KS_3714(s3714, c3714, in3714_1, in3714_2);
    wire[1:0] s3715, in3715_1, in3715_2;
    wire c3715;
    assign in3715_1 = {s1450[2],s1458[0]};
    assign in3715_2 = {s1452[2],s1459[0]};
    CLA_2 KS_3715(s3715, c3715, in3715_1, in3715_2);
    wire[0:0] s3716, in3716_1, in3716_2;
    wire c3716;
    assign in3716_1 = {s1454[2]};
    assign in3716_2 = {s1455[0]};
    Half_Adder KS_3716(s3716, c3716, in3716_1, in3716_2);
    wire[3:0] s3717, in3717_1, in3717_2;
    wire c3717;
    assign in3717_1 = {s1456[0],s1460[0],s1499[0],c1498};
    assign in3717_2 = {c3657,s1461[0],s1500[0],s1499[1]};
    CLA_4 KS_3717(s3717, c3717, in3717_1, in3717_2);
    wire[0:0] s3718, in3718_1, in3718_2;
    wire c3718;
    assign in3718_1 = {c3658};
    assign in3718_2 = {c3659};
    Half_Adder KS_3718(s3718, c3718, in3718_1, in3718_2);
    wire[1:0] s3719, in3719_1, in3719_2;
    wire c3719;
    assign in3719_1 = {c3660,s1462[0]};
    assign in3719_2 = {c3661,s1463[0]};
    CLA_2 KS_3719(s3719, c3719, in3719_1, in3719_2);
    wire[0:0] s3720, in3720_1, in3720_2;
    wire c3720;
    assign in3720_1 = {c3662};
    assign in3720_2 = {c3663};
    Half_Adder KS_3720(s3720, c3720, in3720_1, in3720_2);
    wire[2:0] s3721, in3721_1, in3721_2;
    wire c3721;
    assign in3721_1 = {c3664,s1464[0],s1501[0]};
    assign in3721_2 = {c3665,s3695[1],s1502[0]};
    CLA_3 KS_3721(s3721, c3721, in3721_1, in3721_2);
    wire[0:0] s3722, in3722_1, in3722_2;
    wire c3722;
    assign in3722_1 = {c3666};
    assign in3722_2 = {c3667};
    Half_Adder KS_3722(s3722, c3722, in3722_1, in3722_2);
    wire[1:0] s3723, in3723_1, in3723_2;
    wire c3723;
    assign in3723_1 = {c3668,s3696[1]};
    assign in3723_2 = {c3669,s3697[1]};
    CLA_2 KS_3723(s3723, c3723, in3723_1, in3723_2);
    wire[0:0] s3724, in3724_1, in3724_2;
    wire c3724;
    assign in3724_1 = {c3670};
    assign in3724_2 = {c3671};
    Half_Adder KS_3724(s3724, c3724, in3724_1, in3724_2);
    wire[3:0] s3725, in3725_1, in3725_2;
    wire c3725;
    assign in3725_1 = {c3672,s3698[1],s1503[0],c1500};
    assign in3725_2 = {c3673,s3699[1],s1504[0],s1501[1]};
    CLA_4 KS_3725(s3725, c3725, in3725_1, in3725_2);
    wire[0:0] s3726, in3726_1, in3726_2;
    wire c3726;
    assign in3726_1 = {c3674};
    assign in3726_2 = {c3679};
    Half_Adder KS_3726(s3726, c3726, in3726_1, in3726_2);
    wire[1:0] s3727, in3727_1, in3727_2;
    wire c3727;
    assign in3727_1 = {c3687,s3700[1]};
    assign in3727_2 = {s3695[0],s3701[1]};
    CLA_2 KS_3727(s3727, c3727, in3727_1, in3727_2);
    wire[0:0] s3728, in3728_1, in3728_2;
    wire c3728;
    assign in3728_1 = {s3696[0]};
    assign in3728_2 = {s3697[0]};
    Half_Adder KS_3728(s3728, c3728, in3728_1, in3728_2);
    wire[2:0] s3729, in3729_1, in3729_2;
    wire c3729;
    assign in3729_1 = {s3698[0],s3702[1],s1505[0]};
    assign in3729_2 = {s3699[0],s3703[1],s3695[2]};
    CLA_3 KS_3729(s3729, c3729, in3729_1, in3729_2);
    wire[0:0] s3730, in3730_1, in3730_2;
    wire c3730;
    assign in3730_1 = {s3700[0]};
    assign in3730_2 = {s3701[0]};
    Half_Adder KS_3730(s3730, c3730, in3730_1, in3730_2);
    wire[1:0] s3731, in3731_1, in3731_2;
    wire c3731;
    assign in3731_1 = {s3703[0],s3704[1]};
    assign in3731_2 = {s3704[0],s3705[1]};
    CLA_2_c KS_3731(s3731, c3731, in3731_1, in3731_2, s3702[0]);
    wire[3:0] s3732, in3732_1, in3732_2;
    wire c3732;
    assign in3732_1 = {pp72[3],c1458,s1519[0],s1520[1]};
    assign in3732_2 = {pp73[2],c1459,s1520[0],s1521[1]};
    CLA_4 KS_3732(s3732, c3732, in3732_1, in3732_2);
    wire[3:0] s3733, in3733_1, in3733_2;
    wire c3733;
    assign in3733_1 = {pp74[1],c1460,s1521[0],s1522[1]};
    assign in3733_2 = {pp75[0],c1461,s1522[0],s1523[1]};
    CLA_4 KS_3733(s3733, c3733, in3733_1, in3733_2);
    wire[3:0] s3734, in3734_1, in3734_2;
    wire c3734;
    assign in3734_1 = {c1455,c1462,s1523[0],s1524[1]};
    assign in3734_2 = {c1456,c1463,s1524[0],s1525[1]};
    CLA_4 KS_3734(s3734, c3734, in3734_1, in3734_2);
    wire[3:0] s3735, in3735_1, in3735_2;
    wire c3735;
    assign in3735_1 = {s1457[3],c1464,s1525[0],s1526[1]};
    assign in3735_2 = {s1458[3],s1465[3],s1526[0],s1527[1]};
    CLA_4 KS_3735(s3735, c3735, in3735_1, in3735_2);
    wire[3:0] s3736, in3736_1, in3736_2;
    wire c3736;
    assign in3736_1 = {s1459[3],s1466[3],s1527[0],s1528[1]};
    assign in3736_2 = {s1460[3],s1467[3],s1528[0],s1529[1]};
    CLA_4 KS_3736(s3736, c3736, in3736_1, in3736_2);
    wire[3:0] s3737, in3737_1, in3737_2;
    wire c3737;
    assign in3737_1 = {s1461[3],s1468[3],s1529[0],s1530[1]};
    assign in3737_2 = {s1462[3],s1469[3],s1530[0],s1531[1]};
    CLA_4 KS_3737(s3737, c3737, in3737_1, in3737_2);
    wire[3:0] s3738, in3738_1, in3738_2;
    wire c3738;
    assign in3738_1 = {s1463[3],s1470[3],s1531[0],s1532[1]};
    assign in3738_2 = {s1464[3],s1471[3],s1532[0],s1533[1]};
    CLA_4 KS_3738(s3738, c3738, in3738_1, in3738_2);
    wire[3:0] s3739, in3739_1, in3739_2;
    wire c3739;
    assign in3739_1 = {s1465[2],s1472[3],s1533[0],s1534[1]};
    assign in3739_2 = {s1466[2],s1473[3],s1534[0],s1535[1]};
    CLA_4 KS_3739(s3739, c3739, in3739_1, in3739_2);
    wire[3:0] s3740, in3740_1, in3740_2;
    wire c3740;
    assign in3740_1 = {s1467[2],s1474[3],s1535[0],s1536[1]};
    assign in3740_2 = {s1468[2],s1475[3],s1536[0],s1537[1]};
    CLA_4 KS_3740(s3740, c3740, in3740_1, in3740_2);
    wire[3:0] s3741, in3741_1, in3741_2;
    wire c3741;
    assign in3741_1 = {s1469[2],s1476[3],s1537[0],c1538};
    assign in3741_2 = {s1470[2],s1477[3],s1538[0],s1539[1]};
    CLA_4 KS_3741(s3741, c3741, in3741_1, in3741_2);
    wire[3:0] s3742, in3742_1, in3742_2;
    wire c3742;
    assign in3742_1 = {s1471[2],s1478[3],s1539[0],c1540};
    assign in3742_2 = {s1472[2],s1479[3],s1540[0],s1541[1]};
    CLA_4 KS_3742(s3742, c3742, in3742_1, in3742_2);
    wire[3:0] s3743, in3743_1, in3743_2;
    wire c3743;
    assign in3743_1 = {s1473[2],s1480[3],s1541[0],c1542};
    assign in3743_2 = {s1474[2],s1481[3],s1542[0],s1543[1]};
    CLA_4 KS_3743(s3743, c3743, in3743_1, in3743_2);
    wire[3:0] s3744, in3744_1, in3744_2;
    wire c3744;
    assign in3744_1 = {s1475[2],s1482[3],s1543[0],c1544};
    assign in3744_2 = {s1476[2],s1483[3],s1544[0],s1545[1]};
    CLA_4 KS_3744(s3744, c3744, in3744_1, in3744_2);
    wire[3:0] s3745, in3745_1, in3745_2;
    wire c3745;
    assign in3745_1 = {s1477[2],s1484[3],s1545[0],c1546};
    assign in3745_2 = {s1478[2],s1485[3],s1546[0],s1547[1]};
    CLA_4 KS_3745(s3745, c3745, in3745_1, in3745_2);
    wire[3:0] s3746, in3746_1, in3746_2;
    wire c3746;
    assign in3746_1 = {s1479[2],s1487[3],s1547[0],c1548};
    assign in3746_2 = {s1480[2],s1489[3],s1548[0],s1549[1]};
    CLA_4 KS_3746(s3746, c3746, in3746_1, in3746_2);
    wire[3:0] s3747, in3747_1, in3747_2;
    wire c3747;
    assign in3747_1 = {s1481[2],s1491[3],s1549[0],c1550};
    assign in3747_2 = {s1482[2],s1493[3],s1550[0],s1551[1]};
    CLA_4 KS_3747(s3747, c3747, in3747_1, in3747_2);
    wire[3:0] s3748, in3748_1, in3748_2;
    wire c3748;
    assign in3748_1 = {s1483[2],s1495[3],s1551[0],c1552};
    assign in3748_2 = {s1484[2],s1499[3],s1552[0],s1553[1]};
    CLA_4 KS_3748(s3748, c3748, in3748_1, in3748_2);
    wire[3:0] s3749, in3749_1, in3749_2;
    wire c3749;
    assign in3749_1 = {s1485[2],s1503[3],s1553[0],c1554};
    assign in3749_2 = {s1487[2],s1506[0],s1554[0],s1555[1]};
    CLA_4 KS_3749(s3749, c3749, in3749_1, in3749_2);
    wire[2:0] s3750, in3750_1, in3750_2;
    wire c3750;
    assign in3750_1 = {s1489[2],s1507[0],s1555[0]};
    assign in3750_2 = {s1491[2],s1508[0],s1556[0]};
    CLA_3 KS_3750(s3750, c3750, in3750_1, in3750_2);
    wire[0:0] s3751, in3751_1, in3751_2;
    wire c3751;
    assign in3751_1 = {s1493[2]};
    assign in3751_2 = {s1495[2]};
    Half_Adder KS_3751(s3751, c3751, in3751_1, in3751_2);
    wire[1:0] s3752, in3752_1, in3752_2;
    wire c3752;
    assign in3752_1 = {c1497,s1509[0]};
    assign in3752_2 = {s1499[2],s1510[0]};
    CLA_2 KS_3752(s3752, c3752, in3752_1, in3752_2);
    wire[0:0] s3753, in3753_1, in3753_2;
    wire c3753;
    assign in3753_1 = {c1501};
    assign in3753_2 = {s1503[2]};
    Half_Adder KS_3753(s3753, c3753, in3753_1, in3753_2);
    wire[3:0] s3754, in3754_1, in3754_2;
    wire c3754;
    assign in3754_1 = {c1505,s1511[0],s1557[0],c1556};
    assign in3754_2 = {c3695,s1512[0],s1558[0],s1557[1]};
    CLA_4 KS_3754(s3754, c3754, in3754_1, in3754_2);
    wire[0:0] s3755, in3755_1, in3755_2;
    wire c3755;
    assign in3755_1 = {c3696};
    assign in3755_2 = {c3697};
    Half_Adder KS_3755(s3755, c3755, in3755_1, in3755_2);
    wire[1:0] s3756, in3756_1, in3756_2;
    wire c3756;
    assign in3756_1 = {c3698,s1513[0]};
    assign in3756_2 = {c3699,s1514[0]};
    CLA_2 KS_3756(s3756, c3756, in3756_1, in3756_2);
    wire[0:0] s3757, in3757_1, in3757_2;
    wire c3757;
    assign in3757_1 = {c3700};
    assign in3757_2 = {c3701};
    Half_Adder KS_3757(s3757, c3757, in3757_1, in3757_2);
    wire[2:0] s3758, in3758_1, in3758_2;
    wire c3758;
    assign in3758_1 = {c3702,s1515[0],s1559[0]};
    assign in3758_2 = {c3703,s3732[1],s1560[0]};
    CLA_3 KS_3758(s3758, c3758, in3758_1, in3758_2);
    wire[0:0] s3759, in3759_1, in3759_2;
    wire c3759;
    assign in3759_1 = {c3704};
    assign in3759_2 = {c3705};
    Half_Adder KS_3759(s3759, c3759, in3759_1, in3759_2);
    wire[1:0] s3760, in3760_1, in3760_2;
    wire c3760;
    assign in3760_1 = {c3706,s3733[1]};
    assign in3760_2 = {c3707,s3734[1]};
    CLA_2 KS_3760(s3760, c3760, in3760_1, in3760_2);
    wire[0:0] s3761, in3761_1, in3761_2;
    wire c3761;
    assign in3761_1 = {c3708};
    assign in3761_2 = {c3709};
    Half_Adder KS_3761(s3761, c3761, in3761_1, in3761_2);
    wire[3:0] s3762, in3762_1, in3762_2;
    wire c3762;
    assign in3762_1 = {c3710,s3735[1],s1561[0],c1558};
    assign in3762_2 = {c3711,s3736[1],s1562[0],s1559[1]};
    CLA_4 KS_3762(s3762, c3762, in3762_1, in3762_2);
    wire[0:0] s3763, in3763_1, in3763_2;
    wire c3763;
    assign in3763_1 = {c3712};
    assign in3763_2 = {c3717};
    Half_Adder KS_3763(s3763, c3763, in3763_1, in3763_2);
    wire[1:0] s3764, in3764_1, in3764_2;
    wire c3764;
    assign in3764_1 = {c3725,s3737[1]};
    assign in3764_2 = {s3732[0],s3738[1]};
    CLA_2 KS_3764(s3764, c3764, in3764_1, in3764_2);
    wire[0:0] s3765, in3765_1, in3765_2;
    wire c3765;
    assign in3765_1 = {s3733[0]};
    assign in3765_2 = {s3734[0]};
    Half_Adder KS_3765(s3765, c3765, in3765_1, in3765_2);
    wire[2:0] s3766, in3766_1, in3766_2;
    wire c3766;
    assign in3766_1 = {s3735[0],s3739[1],s1563[0]};
    assign in3766_2 = {s3736[0],s3740[1],s3732[2]};
    CLA_3 KS_3766(s3766, c3766, in3766_1, in3766_2);
    wire[0:0] s3767, in3767_1, in3767_2;
    wire c3767;
    assign in3767_1 = {s3737[0]};
    assign in3767_2 = {s3738[0]};
    Half_Adder KS_3767(s3767, c3767, in3767_1, in3767_2);
    wire[1:0] s3768, in3768_1, in3768_2;
    wire c3768;
    assign in3768_1 = {s3740[0],s3741[1]};
    assign in3768_2 = {s3741[0],s3742[1]};
    CLA_2_c KS_3768(s3768, c3768, in3768_1, in3768_2, s3739[0]);
    wire[3:0] s3769, in3769_1, in3769_2;
    wire c3769;
    assign in3769_1 = {s1506[3],c1511,s1577[0],s1578[1]};
    assign in3769_2 = {s1507[3],c1512,s1578[0],s1579[1]};
    CLA_4 KS_3769(s3769, c3769, in3769_1, in3769_2);
    wire[3:0] s3770, in3770_1, in3770_2;
    wire c3770;
    assign in3770_1 = {s1508[3],c1513,s1579[0],s1580[1]};
    assign in3770_2 = {s1509[3],c1514,s1580[0],s1581[1]};
    CLA_4 KS_3770(s3770, c3770, in3770_1, in3770_2);
    wire[3:0] s3771, in3771_1, in3771_2;
    wire c3771;
    assign in3771_1 = {s1510[3],c1515,s1581[0],s1582[1]};
    assign in3771_2 = {s1511[3],s1516[3],s1582[0],s1583[1]};
    CLA_4 KS_3771(s3771, c3771, in3771_1, in3771_2);
    wire[3:0] s3772, in3772_1, in3772_2;
    wire c3772;
    assign in3772_1 = {s1512[3],s1517[3],s1583[0],s1584[1]};
    assign in3772_2 = {s1513[3],s1518[3],s1584[0],s1585[1]};
    CLA_4 KS_3772(s3772, c3772, in3772_1, in3772_2);
    wire[3:0] s3773, in3773_1, in3773_2;
    wire c3773;
    assign in3773_1 = {s1514[3],s1519[3],s1585[0],s1586[1]};
    assign in3773_2 = {s1515[3],s1520[3],s1586[0],s1587[1]};
    CLA_4 KS_3773(s3773, c3773, in3773_1, in3773_2);
    wire[3:0] s3774, in3774_1, in3774_2;
    wire c3774;
    assign in3774_1 = {s1516[2],s1521[3],s1587[0],s1588[1]};
    assign in3774_2 = {s1517[2],s1522[3],s1588[0],s1589[1]};
    CLA_4 KS_3774(s3774, c3774, in3774_1, in3774_2);
    wire[3:0] s3775, in3775_1, in3775_2;
    wire c3775;
    assign in3775_1 = {s1518[2],s1523[3],s1589[0],s1590[1]};
    assign in3775_2 = {s1519[2],s1524[3],s1590[0],s1591[1]};
    CLA_4 KS_3775(s3775, c3775, in3775_1, in3775_2);
    wire[3:0] s3776, in3776_1, in3776_2;
    wire c3776;
    assign in3776_1 = {s1520[2],s1525[3],s1591[0],s1592[1]};
    assign in3776_2 = {s1521[2],s1526[3],s1592[0],s1593[1]};
    CLA_4 KS_3776(s3776, c3776, in3776_1, in3776_2);
    wire[3:0] s3777, in3777_1, in3777_2;
    wire c3777;
    assign in3777_1 = {s1522[2],s1527[3],s1593[0],s1594[1]};
    assign in3777_2 = {s1523[2],s1528[3],s1594[0],s1595[1]};
    CLA_4 KS_3777(s3777, c3777, in3777_1, in3777_2);
    wire[3:0] s3778, in3778_1, in3778_2;
    wire c3778;
    assign in3778_1 = {s1524[2],s1529[3],s1595[0],c1596};
    assign in3778_2 = {s1525[2],s1530[3],s1596[0],s1597[1]};
    CLA_4 KS_3778(s3778, c3778, in3778_1, in3778_2);
    wire[3:0] s3779, in3779_1, in3779_2;
    wire c3779;
    assign in3779_1 = {s1526[2],s1531[3],s1597[0],c1598};
    assign in3779_2 = {s1527[2],s1532[3],s1598[0],s1599[1]};
    CLA_4 KS_3779(s3779, c3779, in3779_1, in3779_2);
    wire[3:0] s3780, in3780_1, in3780_2;
    wire c3780;
    assign in3780_1 = {s1528[2],s1533[3],s1599[0],c1600};
    assign in3780_2 = {s1529[2],s1534[3],s1600[0],s1601[1]};
    CLA_4 KS_3780(s3780, c3780, in3780_1, in3780_2);
    wire[3:0] s3781, in3781_1, in3781_2;
    wire c3781;
    assign in3781_1 = {s1530[2],s1535[3],s1601[0],c1602};
    assign in3781_2 = {s1531[2],s1536[3],s1602[0],s1603[1]};
    CLA_4 KS_3781(s3781, c3781, in3781_1, in3781_2);
    wire[3:0] s3782, in3782_1, in3782_2;
    wire c3782;
    assign in3782_1 = {s1532[2],s1537[3],s1603[0],c1604};
    assign in3782_2 = {s1533[2],s1541[3],s1604[0],s1605[1]};
    CLA_4 KS_3782(s3782, c3782, in3782_1, in3782_2);
    wire[3:0] s3783, in3783_1, in3783_2;
    wire c3783;
    assign in3783_1 = {s1534[2],s1545[3],s1605[0],c1606};
    assign in3783_2 = {s1535[2],s1549[3],s1606[0],s1607[1]};
    CLA_4 KS_3783(s3783, c3783, in3783_1, in3783_2);
    wire[3:0] s3784, in3784_1, in3784_2;
    wire c3784;
    assign in3784_1 = {s1536[2],s1553[3],s1607[0],c1608};
    assign in3784_2 = {s1537[2],s1557[3],s1608[0],s1609[1]};
    CLA_4 KS_3784(s3784, c3784, in3784_1, in3784_2);
    wire[3:0] s3785, in3785_1, in3785_2;
    wire c3785;
    assign in3785_1 = {c1539,s1561[3],s1609[0],c1610};
    assign in3785_2 = {s1541[2],s1564[0],s1610[0],s1611[1]};
    CLA_4 KS_3785(s3785, c3785, in3785_1, in3785_2);
    wire[3:0] s3786, in3786_1, in3786_2;
    wire c3786;
    assign in3786_1 = {c1543,s1565[0],s1611[0],c1612};
    assign in3786_2 = {s1545[2],s1566[0],s1612[0],s1613[1]};
    CLA_4 KS_3786(s3786, c3786, in3786_1, in3786_2);
    wire[2:0] s3787, in3787_1, in3787_2;
    wire c3787;
    assign in3787_1 = {c1547,s1567[0],s1613[0]};
    assign in3787_2 = {s1549[2],s1568[0],s1614[0]};
    CLA_3 KS_3787(s3787, c3787, in3787_1, in3787_2);
    wire[0:0] s3788, in3788_1, in3788_2;
    wire c3788;
    assign in3788_1 = {c1551};
    assign in3788_2 = {s1553[2]};
    Half_Adder KS_3788(s3788, c3788, in3788_1, in3788_2);
    wire[1:0] s3789, in3789_1, in3789_2;
    wire c3789;
    assign in3789_1 = {c1555,s1569[0]};
    assign in3789_2 = {s1557[2],s1570[0]};
    CLA_2 KS_3789(s3789, c3789, in3789_1, in3789_2);
    wire[0:0] s3790, in3790_1, in3790_2;
    wire c3790;
    assign in3790_1 = {c1559};
    assign in3790_2 = {s1561[2]};
    Half_Adder KS_3790(s3790, c3790, in3790_1, in3790_2);
    wire[3:0] s3791, in3791_1, in3791_2;
    wire c3791;
    assign in3791_1 = {c1563,s1571[0],s1615[0],c1614};
    assign in3791_2 = {c3732,s1572[0],s1616[0],s1615[1]};
    CLA_4 KS_3791(s3791, c3791, in3791_1, in3791_2);
    wire[0:0] s3792, in3792_1, in3792_2;
    wire c3792;
    assign in3792_1 = {c3733};
    assign in3792_2 = {c3734};
    Half_Adder KS_3792(s3792, c3792, in3792_1, in3792_2);
    wire[1:0] s3793, in3793_1, in3793_2;
    wire c3793;
    assign in3793_1 = {c3735,s1573[0]};
    assign in3793_2 = {c3736,s1574[0]};
    CLA_2 KS_3793(s3793, c3793, in3793_1, in3793_2);
    wire[0:0] s3794, in3794_1, in3794_2;
    wire c3794;
    assign in3794_1 = {c3737};
    assign in3794_2 = {c3738};
    Half_Adder KS_3794(s3794, c3794, in3794_1, in3794_2);
    wire[2:0] s3795, in3795_1, in3795_2;
    wire c3795;
    assign in3795_1 = {c3739,s1575[0],s1617[0]};
    assign in3795_2 = {c3740,s3769[1],s1618[0]};
    CLA_3 KS_3795(s3795, c3795, in3795_1, in3795_2);
    wire[0:0] s3796, in3796_1, in3796_2;
    wire c3796;
    assign in3796_1 = {c3741};
    assign in3796_2 = {c3742};
    Half_Adder KS_3796(s3796, c3796, in3796_1, in3796_2);
    wire[1:0] s3797, in3797_1, in3797_2;
    wire c3797;
    assign in3797_1 = {c3743,s3770[1]};
    assign in3797_2 = {c3744,s3771[1]};
    CLA_2 KS_3797(s3797, c3797, in3797_1, in3797_2);
    wire[0:0] s3798, in3798_1, in3798_2;
    wire c3798;
    assign in3798_1 = {c3745};
    assign in3798_2 = {c3746};
    Half_Adder KS_3798(s3798, c3798, in3798_1, in3798_2);
    wire[3:0] s3799, in3799_1, in3799_2;
    wire c3799;
    assign in3799_1 = {c3747,s3772[1],s1619[0],c1616};
    assign in3799_2 = {c3748,s3773[1],s1620[0],s1617[1]};
    CLA_4 KS_3799(s3799, c3799, in3799_1, in3799_2);
    wire[0:0] s3800, in3800_1, in3800_2;
    wire c3800;
    assign in3800_1 = {c3749};
    assign in3800_2 = {c3754};
    Half_Adder KS_3800(s3800, c3800, in3800_1, in3800_2);
    wire[1:0] s3801, in3801_1, in3801_2;
    wire c3801;
    assign in3801_1 = {c3762,s3774[1]};
    assign in3801_2 = {s3769[0],s3775[1]};
    CLA_2 KS_3801(s3801, c3801, in3801_1, in3801_2);
    wire[0:0] s3802, in3802_1, in3802_2;
    wire c3802;
    assign in3802_1 = {s3770[0]};
    assign in3802_2 = {s3771[0]};
    Half_Adder KS_3802(s3802, c3802, in3802_1, in3802_2);
    wire[2:0] s3803, in3803_1, in3803_2;
    wire c3803;
    assign in3803_1 = {s3772[0],s3776[1],s1621[0]};
    assign in3803_2 = {s3773[0],s3777[1],s3769[2]};
    CLA_3 KS_3803(s3803, c3803, in3803_1, in3803_2);
    wire[0:0] s3804, in3804_1, in3804_2;
    wire c3804;
    assign in3804_1 = {s3774[0]};
    assign in3804_2 = {s3775[0]};
    Half_Adder KS_3804(s3804, c3804, in3804_1, in3804_2);
    wire[1:0] s3805, in3805_1, in3805_2;
    wire c3805;
    assign in3805_1 = {s3777[0],s3778[1]};
    assign in3805_2 = {s3778[0],s3779[1]};
    CLA_2_c KS_3805(s3805, c3805, in3805_1, in3805_2, s3776[0]);
    wire[3:0] s3806, in3806_1, in3806_2;
    wire c3806;
    assign in3806_1 = {s1564[3],c1573,s1633[1],s1634[2]};
    assign in3806_2 = {s1565[3],c1574,s1634[1],s1635[2]};
    CLA_4 KS_3806(s3806, c3806, in3806_1, in3806_2);
    wire[3:0] s3807, in3807_1, in3807_2;
    wire c3807;
    assign in3807_1 = {s1566[3],c1575,s1635[1],s1636[2]};
    assign in3807_2 = {s1567[3],s1576[3],s1636[1],s1637[2]};
    CLA_4 KS_3807(s3807, c3807, in3807_1, in3807_2);
    wire[3:0] s3808, in3808_1, in3808_2;
    wire c3808;
    assign in3808_1 = {s1568[3],s1577[3],s1637[1],s1638[1]};
    assign in3808_2 = {s1569[3],s1578[3],s1638[0],s1639[1]};
    CLA_4 KS_3808(s3808, c3808, in3808_1, in3808_2);
    wire[3:0] s3809, in3809_1, in3809_2;
    wire c3809;
    assign in3809_1 = {s1570[3],s1579[3],s1639[0],s1640[1]};
    assign in3809_2 = {s1571[3],s1580[3],s1640[0],s1641[1]};
    CLA_4 KS_3809(s3809, c3809, in3809_1, in3809_2);
    wire[3:0] s3810, in3810_1, in3810_2;
    wire c3810;
    assign in3810_1 = {s1572[3],s1581[3],s1641[0],s1642[1]};
    assign in3810_2 = {s1573[3],s1582[3],s1642[0],s1643[1]};
    CLA_4 KS_3810(s3810, c3810, in3810_1, in3810_2);
    wire[3:0] s3811, in3811_1, in3811_2;
    wire c3811;
    assign in3811_1 = {s1574[3],s1583[3],s1643[0],s1644[1]};
    assign in3811_2 = {s1575[3],s1584[3],s1644[0],s1645[1]};
    CLA_4 KS_3811(s3811, c3811, in3811_1, in3811_2);
    wire[3:0] s3812, in3812_1, in3812_2;
    wire c3812;
    assign in3812_1 = {s1576[2],s1585[3],s1645[0],s1646[1]};
    assign in3812_2 = {s1577[2],s1586[3],s1646[0],s1647[1]};
    CLA_4 KS_3812(s3812, c3812, in3812_1, in3812_2);
    wire[3:0] s3813, in3813_1, in3813_2;
    wire c3813;
    assign in3813_1 = {s1578[2],s1587[3],s1647[0],s1648[1]};
    assign in3813_2 = {s1579[2],s1588[3],s1648[0],s1649[1]};
    CLA_4 KS_3813(s3813, c3813, in3813_1, in3813_2);
    wire[3:0] s3814, in3814_1, in3814_2;
    wire c3814;
    assign in3814_1 = {s1580[2],s1589[3],s1649[0],s1650[1]};
    assign in3814_2 = {s1581[2],s1590[3],s1650[0],s1651[1]};
    CLA_4 KS_3814(s3814, c3814, in3814_1, in3814_2);
    wire[3:0] s3815, in3815_1, in3815_2;
    wire c3815;
    assign in3815_1 = {s1582[2],s1591[3],s1651[0],s1652[1]};
    assign in3815_2 = {s1583[2],s1592[3],s1652[0],s1653[1]};
    CLA_4 KS_3815(s3815, c3815, in3815_1, in3815_2);
    wire[3:0] s3816, in3816_1, in3816_2;
    wire c3816;
    assign in3816_1 = {s1584[2],s1593[3],s1653[0],c1654};
    assign in3816_2 = {s1585[2],s1594[3],s1654[0],s1655[1]};
    CLA_4 KS_3816(s3816, c3816, in3816_1, in3816_2);
    wire[3:0] s3817, in3817_1, in3817_2;
    wire c3817;
    assign in3817_1 = {s1586[2],s1595[3],s1655[0],c1656};
    assign in3817_2 = {s1587[2],s1599[3],s1656[0],s1657[1]};
    CLA_4 KS_3817(s3817, c3817, in3817_1, in3817_2);
    wire[3:0] s3818, in3818_1, in3818_2;
    wire c3818;
    assign in3818_1 = {s1588[2],s1603[3],s1657[0],c1658};
    assign in3818_2 = {s1589[2],s1607[3],s1658[0],s1659[1]};
    CLA_4 KS_3818(s3818, c3818, in3818_1, in3818_2);
    wire[3:0] s3819, in3819_1, in3819_2;
    wire c3819;
    assign in3819_1 = {s1590[2],s1611[3],s1659[0],c1660};
    assign in3819_2 = {s1591[2],s1615[3],s1660[0],s1661[1]};
    CLA_4 KS_3819(s3819, c3819, in3819_1, in3819_2);
    wire[3:0] s3820, in3820_1, in3820_2;
    wire c3820;
    assign in3820_1 = {s1592[2],s1619[3],s1661[0],c1662};
    assign in3820_2 = {s1593[2],s1622[0],s1662[0],s1663[1]};
    CLA_4 KS_3820(s3820, c3820, in3820_1, in3820_2);
    wire[3:0] s3821, in3821_1, in3821_2;
    wire c3821;
    assign in3821_1 = {s1594[2],s1623[0],s1663[0],c1664};
    assign in3821_2 = {s1595[2],s1624[0],s1664[0],s1665[1]};
    CLA_4 KS_3821(s3821, c3821, in3821_1, in3821_2);
    wire[3:0] s3822, in3822_1, in3822_2;
    wire c3822;
    assign in3822_1 = {c1597,s1625[0],s1665[0],c1666};
    assign in3822_2 = {s1599[2],s1626[0],s1666[0],s1667[1]};
    CLA_4 KS_3822(s3822, c3822, in3822_1, in3822_2);
    wire[3:0] s3823, in3823_1, in3823_2;
    wire c3823;
    assign in3823_1 = {c1601,s1627[0],s1667[0],c1668};
    assign in3823_2 = {s1603[2],s1628[0],s1668[0],s1669[1]};
    CLA_4 KS_3823(s3823, c3823, in3823_1, in3823_2);
    wire[2:0] s3824, in3824_1, in3824_2;
    wire c3824;
    assign in3824_1 = {c1605,s1629[0],s1669[0]};
    assign in3824_2 = {s1607[2],s1630[0],s1670[0]};
    CLA_3 KS_3824(s3824, c3824, in3824_1, in3824_2);
    wire[0:0] s3825, in3825_1, in3825_2;
    wire c3825;
    assign in3825_1 = {c1609};
    assign in3825_2 = {s1611[2]};
    Half_Adder KS_3825(s3825, c3825, in3825_1, in3825_2);
    wire[1:0] s3826, in3826_1, in3826_2;
    wire c3826;
    assign in3826_1 = {c1613,s1631[0]};
    assign in3826_2 = {s1615[2],s1632[0]};
    CLA_2 KS_3826(s3826, c3826, in3826_1, in3826_2);
    wire[0:0] s3827, in3827_1, in3827_2;
    wire c3827;
    assign in3827_1 = {c1617};
    assign in3827_2 = {s1619[2]};
    Half_Adder KS_3827(s3827, c3827, in3827_1, in3827_2);
    wire[3:0] s3828, in3828_1, in3828_2;
    wire c3828;
    assign in3828_1 = {c1621,s1633[0],s1671[0],c1670};
    assign in3828_2 = {c3769,s1634[0],s1672[0],s1671[1]};
    CLA_4 KS_3828(s3828, c3828, in3828_1, in3828_2);
    wire[0:0] s3829, in3829_1, in3829_2;
    wire c3829;
    assign in3829_1 = {c3770};
    assign in3829_2 = {c3771};
    Half_Adder KS_3829(s3829, c3829, in3829_1, in3829_2);
    wire[1:0] s3830, in3830_1, in3830_2;
    wire c3830;
    assign in3830_1 = {c3772,s1635[0]};
    assign in3830_2 = {c3773,s1636[0]};
    CLA_2 KS_3830(s3830, c3830, in3830_1, in3830_2);
    wire[0:0] s3831, in3831_1, in3831_2;
    wire c3831;
    assign in3831_1 = {c3774};
    assign in3831_2 = {c3775};
    Half_Adder KS_3831(s3831, c3831, in3831_1, in3831_2);
    wire[2:0] s3832, in3832_1, in3832_2;
    wire c3832;
    assign in3832_1 = {c3776,s1637[0],s1673[0]};
    assign in3832_2 = {c3777,s3806[1],s1674[0]};
    CLA_3 KS_3832(s3832, c3832, in3832_1, in3832_2);
    wire[0:0] s3833, in3833_1, in3833_2;
    wire c3833;
    assign in3833_1 = {c3778};
    assign in3833_2 = {c3779};
    Half_Adder KS_3833(s3833, c3833, in3833_1, in3833_2);
    wire[1:0] s3834, in3834_1, in3834_2;
    wire c3834;
    assign in3834_1 = {c3780,s3807[1]};
    assign in3834_2 = {c3781,s3808[1]};
    CLA_2 KS_3834(s3834, c3834, in3834_1, in3834_2);
    wire[0:0] s3835, in3835_1, in3835_2;
    wire c3835;
    assign in3835_1 = {c3782};
    assign in3835_2 = {c3783};
    Half_Adder KS_3835(s3835, c3835, in3835_1, in3835_2);
    wire[3:0] s3836, in3836_1, in3836_2;
    wire c3836;
    assign in3836_1 = {c3784,s3809[1],s1675[0],c1672};
    assign in3836_2 = {c3785,s3810[1],s1676[0],s1673[1]};
    CLA_4 KS_3836(s3836, c3836, in3836_1, in3836_2);
    wire[0:0] s3837, in3837_1, in3837_2;
    wire c3837;
    assign in3837_1 = {c3786};
    assign in3837_2 = {c3791};
    Half_Adder KS_3837(s3837, c3837, in3837_1, in3837_2);
    wire[1:0] s3838, in3838_1, in3838_2;
    wire c3838;
    assign in3838_1 = {c3799,s3811[1]};
    assign in3838_2 = {s3806[0],s3812[1]};
    CLA_2 KS_3838(s3838, c3838, in3838_1, in3838_2);
    wire[0:0] s3839, in3839_1, in3839_2;
    wire c3839;
    assign in3839_1 = {s3807[0]};
    assign in3839_2 = {s3808[0]};
    Half_Adder KS_3839(s3839, c3839, in3839_1, in3839_2);
    wire[2:0] s3840, in3840_1, in3840_2;
    wire c3840;
    assign in3840_1 = {s3809[0],s3813[1],s1677[0]};
    assign in3840_2 = {s3810[0],s3814[1],s3806[2]};
    CLA_3 KS_3840(s3840, c3840, in3840_1, in3840_2);
    wire[0:0] s3841, in3841_1, in3841_2;
    wire c3841;
    assign in3841_1 = {s3811[0]};
    assign in3841_2 = {s3812[0]};
    Half_Adder KS_3841(s3841, c3841, in3841_1, in3841_2);
    wire[1:0] s3842, in3842_1, in3842_2;
    wire c3842;
    assign in3842_1 = {s3814[0],s3815[1]};
    assign in3842_2 = {s3815[0],s3816[1]};
    CLA_2_c KS_3842(s3842, c3842, in3842_1, in3842_2, s3813[0]);
    wire[3:0] s3843, in3843_1, in3843_2;
    wire c3843;
    assign in3843_1 = {s1622[3],s1639[3],s1685[1],s1686[2]};
    assign in3843_2 = {s1623[3],s1640[3],s1686[1],s1687[2]};
    CLA_4 KS_3843(s3843, c3843, in3843_1, in3843_2);
    wire[3:0] s3844, in3844_1, in3844_2;
    wire c3844;
    assign in3844_1 = {s1624[3],s1641[3],s1687[1],s1688[2]};
    assign in3844_2 = {s1625[3],s1642[3],s1688[1],s1689[2]};
    CLA_4 KS_3844(s3844, c3844, in3844_1, in3844_2);
    wire[3:0] s3845, in3845_1, in3845_2;
    wire c3845;
    assign in3845_1 = {s1626[3],s1643[3],s1689[1],s1690[2]};
    assign in3845_2 = {s1627[3],s1644[3],s1690[1],s1691[2]};
    CLA_4 KS_3845(s3845, c3845, in3845_1, in3845_2);
    wire[3:0] s3846, in3846_1, in3846_2;
    wire c3846;
    assign in3846_1 = {s1628[3],s1645[3],s1691[1],s1692[2]};
    assign in3846_2 = {s1629[3],s1646[3],s1692[1],s1693[2]};
    CLA_4 KS_3846(s3846, c3846, in3846_1, in3846_2);
    wire[3:0] s3847, in3847_1, in3847_2;
    wire c3847;
    assign in3847_1 = {s1630[3],s1647[3],s1693[1],s1694[2]};
    assign in3847_2 = {s1631[3],s1648[3],s1694[1],s1695[2]};
    CLA_4 KS_3847(s3847, c3847, in3847_1, in3847_2);
    wire[3:0] s3848, in3848_1, in3848_2;
    wire c3848;
    assign in3848_1 = {s1632[3],s1649[3],s1695[1],s1696[2]};
    assign in3848_2 = {s1633[3],s1650[3],s1696[1],s1697[2]};
    CLA_4 KS_3848(s3848, c3848, in3848_1, in3848_2);
    wire[3:0] s3849, in3849_1, in3849_2;
    wire c3849;
    assign in3849_1 = {s1634[3],s1651[3],s1697[1],s1698[2]};
    assign in3849_2 = {s1635[3],s1652[3],s1698[1],s1699[2]};
    CLA_4 KS_3849(s3849, c3849, in3849_1, in3849_2);
    wire[3:0] s3850, in3850_1, in3850_2;
    wire c3850;
    assign in3850_1 = {s1636[3],s1653[3],s1699[1],s1700[2]};
    assign in3850_2 = {s1637[3],s1657[3],s1700[1],s1701[2]};
    CLA_4 KS_3850(s3850, c3850, in3850_1, in3850_2);
    wire[3:0] s3851, in3851_1, in3851_2;
    wire c3851;
    assign in3851_1 = {s1638[2],s1661[3],s1701[1],s1702[1]};
    assign in3851_2 = {s1639[2],s1665[3],s1702[0],s1703[1]};
    CLA_4 KS_3851(s3851, c3851, in3851_1, in3851_2);
    wire[3:0] s3852, in3852_1, in3852_2;
    wire c3852;
    assign in3852_1 = {s1640[2],s1669[3],s1703[0],s1704[1]};
    assign in3852_2 = {s1641[2],s1673[3],s1704[0],s1705[1]};
    CLA_4 KS_3852(s3852, c3852, in3852_1, in3852_2);
    wire[3:0] s3853, in3853_1, in3853_2;
    wire c3853;
    assign in3853_1 = {s1642[2],s1677[3],s1705[0],s1706[1]};
    assign in3853_2 = {s1643[2],s1678[0],s1706[0],s1707[1]};
    CLA_4 KS_3853(s3853, c3853, in3853_1, in3853_2);
    wire[3:0] s3854, in3854_1, in3854_2;
    wire c3854;
    assign in3854_1 = {s1644[2],s1679[0],s1707[0],s1708[1]};
    assign in3854_2 = {s1645[2],s1680[0],s1708[0],s1709[1]};
    CLA_4 KS_3854(s3854, c3854, in3854_1, in3854_2);
    wire[3:0] s3855, in3855_1, in3855_2;
    wire c3855;
    assign in3855_1 = {s1646[2],s1681[0],s1709[0],c1710};
    assign in3855_2 = {s1647[2],s1682[0],s1710[0],s1711[1]};
    CLA_4 KS_3855(s3855, c3855, in3855_1, in3855_2);
    wire[3:0] s3856, in3856_1, in3856_2;
    wire c3856;
    assign in3856_1 = {s1648[2],s1683[0],s1711[0],c1712};
    assign in3856_2 = {s1649[2],s1684[0],s1712[0],s1713[1]};
    CLA_4 KS_3856(s3856, c3856, in3856_1, in3856_2);
    wire[3:0] s3857, in3857_1, in3857_2;
    wire c3857;
    assign in3857_1 = {s1650[2],s1685[0],s1713[0],c1714};
    assign in3857_2 = {s1651[2],s1686[0],s1714[0],s1715[1]};
    CLA_4 KS_3857(s3857, c3857, in3857_1, in3857_2);
    wire[3:0] s3858, in3858_1, in3858_2;
    wire c3858;
    assign in3858_1 = {s1652[2],s1687[0],s1715[0],c1716};
    assign in3858_2 = {s1653[2],s1688[0],s1716[0],s1717[1]};
    CLA_4 KS_3858(s3858, c3858, in3858_1, in3858_2);
    wire[3:0] s3859, in3859_1, in3859_2;
    wire c3859;
    assign in3859_1 = {c1655,s1689[0],s1717[0],c1718};
    assign in3859_2 = {s1657[2],s1690[0],s1718[0],s1719[1]};
    CLA_4 KS_3859(s3859, c3859, in3859_1, in3859_2);
    wire[3:0] s3860, in3860_1, in3860_2;
    wire c3860;
    assign in3860_1 = {c1659,s1691[0],s1719[0],c1720};
    assign in3860_2 = {s1661[2],s1692[0],s1720[0],s1721[1]};
    CLA_4 KS_3860(s3860, c3860, in3860_1, in3860_2);
    wire[2:0] s3861, in3861_1, in3861_2;
    wire c3861;
    assign in3861_1 = {c1663,s1693[0],s1721[0]};
    assign in3861_2 = {s1665[2],s1694[0],s1722[0]};
    CLA_3 KS_3861(s3861, c3861, in3861_1, in3861_2);
    wire[0:0] s3862, in3862_1, in3862_2;
    wire c3862;
    assign in3862_1 = {c1667};
    assign in3862_2 = {s1669[2]};
    Half_Adder KS_3862(s3862, c3862, in3862_1, in3862_2);
    wire[1:0] s3863, in3863_1, in3863_2;
    wire c3863;
    assign in3863_1 = {c1671,s1695[0]};
    assign in3863_2 = {s1673[2],s1696[0]};
    CLA_2 KS_3863(s3863, c3863, in3863_1, in3863_2);
    wire[0:0] s3864, in3864_1, in3864_2;
    wire c3864;
    assign in3864_1 = {c1675};
    assign in3864_2 = {s1677[2]};
    Half_Adder KS_3864(s3864, c3864, in3864_1, in3864_2);
    wire[3:0] s3865, in3865_1, in3865_2;
    wire c3865;
    assign in3865_1 = {c3806,s1697[0],s1723[0],c1722};
    assign in3865_2 = {c3807,s1698[0],s1724[0],s1723[1]};
    CLA_4 KS_3865(s3865, c3865, in3865_1, in3865_2);
    wire[0:0] s3866, in3866_1, in3866_2;
    wire c3866;
    assign in3866_1 = {c3808};
    assign in3866_2 = {c3809};
    Half_Adder KS_3866(s3866, c3866, in3866_1, in3866_2);
    wire[1:0] s3867, in3867_1, in3867_2;
    wire c3867;
    assign in3867_1 = {c3810,s1699[0]};
    assign in3867_2 = {c3811,s1700[0]};
    CLA_2 KS_3867(s3867, c3867, in3867_1, in3867_2);
    wire[0:0] s3868, in3868_1, in3868_2;
    wire c3868;
    assign in3868_1 = {c3812};
    assign in3868_2 = {c3813};
    Half_Adder KS_3868(s3868, c3868, in3868_1, in3868_2);
    wire[2:0] s3869, in3869_1, in3869_2;
    wire c3869;
    assign in3869_1 = {c3814,s1701[0],s1725[0]};
    assign in3869_2 = {c3815,s3843[1],s1726[0]};
    CLA_3 KS_3869(s3869, c3869, in3869_1, in3869_2);
    wire[0:0] s3870, in3870_1, in3870_2;
    wire c3870;
    assign in3870_1 = {c3816};
    assign in3870_2 = {c3817};
    Half_Adder KS_3870(s3870, c3870, in3870_1, in3870_2);
    wire[1:0] s3871, in3871_1, in3871_2;
    wire c3871;
    assign in3871_1 = {c3818,s3844[1]};
    assign in3871_2 = {c3819,s3845[1]};
    CLA_2 KS_3871(s3871, c3871, in3871_1, in3871_2);
    wire[0:0] s3872, in3872_1, in3872_2;
    wire c3872;
    assign in3872_1 = {c3820};
    assign in3872_2 = {c3821};
    Half_Adder KS_3872(s3872, c3872, in3872_1, in3872_2);
    wire[3:0] s3873, in3873_1, in3873_2;
    wire c3873;
    assign in3873_1 = {c3822,s3846[1],s1727[0],c1724};
    assign in3873_2 = {c3823,s3847[1],s1728[0],s1725[1]};
    CLA_4 KS_3873(s3873, c3873, in3873_1, in3873_2);
    wire[0:0] s3874, in3874_1, in3874_2;
    wire c3874;
    assign in3874_1 = {c3828};
    assign in3874_2 = {c3836};
    Half_Adder KS_3874(s3874, c3874, in3874_1, in3874_2);
    wire[1:0] s3875, in3875_1, in3875_2;
    wire c3875;
    assign in3875_1 = {s3843[0],s3848[1]};
    assign in3875_2 = {s3844[0],s3849[1]};
    CLA_2 KS_3875(s3875, c3875, in3875_1, in3875_2);
    wire[0:0] s3876, in3876_1, in3876_2;
    wire c3876;
    assign in3876_1 = {s3845[0]};
    assign in3876_2 = {s3846[0]};
    Half_Adder KS_3876(s3876, c3876, in3876_1, in3876_2);
    wire[2:0] s3877, in3877_1, in3877_2;
    wire c3877;
    assign in3877_1 = {s3847[0],s3850[1],s1729[0]};
    assign in3877_2 = {s3848[0],s3851[1],s3843[2]};
    CLA_3 KS_3877(s3877, c3877, in3877_1, in3877_2);
    wire[0:0] s3878, in3878_1, in3878_2;
    wire c3878;
    assign in3878_1 = {s3850[0]};
    assign in3878_2 = {s3851[0]};
    Full_Adder KS_3878(s3878, c3878, in3878_1, in3878_2, s3849[0]);
    wire[3:0] s3879, in3879_1, in3879_2;
    wire c3879;
    assign in3879_1 = {s42[0],s1717[3],c1725,s60[0]};
    assign in3879_2 = {s43[0],s1721[3],c1729,s61[0]};
    CLA_4 KS_3879(s3879, c3879, in3879_1, in3879_2);
    wire[3:0] s3880, in3880_1, in3880_2;
    wire c3880;
    assign in3880_1 = {s1678[3],s1725[3],s1730[1],s1730[2]};
    assign in3880_2 = {s1679[3],s1729[3],s1731[1],s1731[2]};
    CLA_4 KS_3880(s3880, c3880, in3880_1, in3880_2);
    wire[3:0] s3881, in3881_1, in3881_2;
    wire c3881;
    assign in3881_1 = {s1680[3],s1730[0],s1732[1],s1732[2]};
    assign in3881_2 = {s1681[3],s1731[0],s1733[1],s1733[2]};
    CLA_4 KS_3881(s3881, c3881, in3881_1, in3881_2);
    wire[3:0] s3882, in3882_1, in3882_2;
    wire c3882;
    assign in3882_1 = {s1682[3],s1732[0],s1734[1],s1734[2]};
    assign in3882_2 = {s1683[3],s1733[0],s1735[1],s1735[2]};
    CLA_4 KS_3882(s3882, c3882, in3882_1, in3882_2);
    wire[3:0] s3883, in3883_1, in3883_2;
    wire c3883;
    assign in3883_1 = {s1684[3],s1734[0],s1736[1],s1736[2]};
    assign in3883_2 = {s1685[3],s1735[0],s1737[1],s1737[2]};
    CLA_4 KS_3883(s3883, c3883, in3883_1, in3883_2);
    wire[3:0] s3884, in3884_1, in3884_2;
    wire c3884;
    assign in3884_1 = {s1686[3],s1736[0],s1738[1],s1738[2]};
    assign in3884_2 = {s1687[3],s1737[0],s1739[1],s1739[2]};
    CLA_4 KS_3884(s3884, c3884, in3884_1, in3884_2);
    wire[3:0] s3885, in3885_1, in3885_2;
    wire c3885;
    assign in3885_1 = {s1688[3],s1738[0],s1740[1],s1740[2]};
    assign in3885_2 = {s1689[3],s1739[0],s1741[1],s1741[2]};
    CLA_4 KS_3885(s3885, c3885, in3885_1, in3885_2);
    wire[3:0] s3886, in3886_1, in3886_2;
    wire c3886;
    assign in3886_1 = {s1690[3],s1740[0],s1742[1],s1742[2]};
    assign in3886_2 = {s1691[3],s1741[0],s1743[1],s1743[2]};
    CLA_4 KS_3886(s3886, c3886, in3886_1, in3886_2);
    wire[3:0] s3887, in3887_1, in3887_2;
    wire c3887;
    assign in3887_1 = {s1692[3],s1742[0],s1744[1],s1744[2]};
    assign in3887_2 = {s1693[3],s1743[0],s1745[1],s1745[2]};
    CLA_4 KS_3887(s3887, c3887, in3887_1, in3887_2);
    wire[3:0] s3888, in3888_1, in3888_2;
    wire c3888;
    assign in3888_1 = {s1694[3],s1744[0],s1746[1],s1746[2]};
    assign in3888_2 = {s1695[3],s1745[0],s1747[1],s1747[2]};
    CLA_4 KS_3888(s3888, c3888, in3888_1, in3888_2);
    wire[3:0] s3889, in3889_1, in3889_2;
    wire c3889;
    assign in3889_1 = {s1696[3],s1746[0],s1748[1],s1748[2]};
    assign in3889_2 = {s1697[3],s1747[0],s1749[1],s1749[2]};
    CLA_4 KS_3889(s3889, c3889, in3889_1, in3889_2);
    wire[3:0] s3890, in3890_1, in3890_2;
    wire c3890;
    assign in3890_1 = {s1698[3],s1748[0],s1750[1],s1750[2]};
    assign in3890_2 = {s1699[3],s1749[0],s1751[1],s1751[2]};
    CLA_4 KS_3890(s3890, c3890, in3890_1, in3890_2);
    wire[3:0] s3891, in3891_1, in3891_2;
    wire c3891;
    assign in3891_1 = {s1700[3],s1750[0],s1752[1],s1752[2]};
    assign in3891_2 = {s1701[3],s1751[0],s1753[1],s1753[2]};
    CLA_4 KS_3891(s3891, c3891, in3891_1, in3891_2);
    wire[3:0] s3892, in3892_1, in3892_2;
    wire c3892;
    assign in3892_1 = {s1702[2],s1752[0],s1754[1],s1754[2]};
    assign in3892_2 = {s1703[2],s1753[0],s1755[1],s1755[2]};
    CLA_4 KS_3892(s3892, c3892, in3892_1, in3892_2);
    wire[3:0] s3893, in3893_1, in3893_2;
    wire c3893;
    assign in3893_1 = {s1704[2],s1754[0],s1756[1],s1756[2]};
    assign in3893_2 = {s1705[2],s1755[0],s1757[1],s1757[2]};
    CLA_4 KS_3893(s3893, c3893, in3893_1, in3893_2);
    wire[3:0] s3894, in3894_1, in3894_2;
    wire c3894;
    assign in3894_1 = {s1706[2],s1756[0],s1758[1],s1758[2]};
    assign in3894_2 = {s1707[2],s1757[0],s1759[1],s1759[2]};
    CLA_4 KS_3894(s3894, c3894, in3894_1, in3894_2);
    wire[3:0] s3895, in3895_1, in3895_2;
    wire c3895;
    assign in3895_1 = {s1708[2],s1758[0],s1760[1],s1760[2]};
    assign in3895_2 = {s1709[2],s1759[0],s1761[1],s1761[2]};
    CLA_4 KS_3895(s3895, c3895, in3895_1, in3895_2);
    wire[3:0] s3896, in3896_1, in3896_2;
    wire c3896;
    assign in3896_1 = {c1711,s1760[0],s1762[1],c1762};
    assign in3896_2 = {s1713[2],s1761[0],s1763[1],s1763[2]};
    CLA_4 KS_3896(s3896, c3896, in3896_1, in3896_2);
    wire[3:0] s3897, in3897_1, in3897_2;
    wire c3897;
    assign in3897_1 = {c1715,s1762[0],s1764[1],c1764};
    assign in3897_2 = {s1717[2],s1763[0],s1765[1],s1765[2]};
    CLA_4 KS_3897(s3897, c3897, in3897_1, in3897_2);
    wire[0:0] s3898, in3898_1, in3898_2;
    wire c3898;
    assign in3898_1 = {c1719};
    assign in3898_2 = {s1721[2]};
    Half_Adder KS_3898(s3898, c3898, in3898_1, in3898_2);
    wire[1:0] s3899, in3899_1, in3899_2;
    wire c3899;
    assign in3899_1 = {c1723,s1764[0]};
    assign in3899_2 = {s1725[2],s1765[0]};
    CLA_2 KS_3899(s3899, c3899, in3899_1, in3899_2);
    wire[0:0] s3900, in3900_1, in3900_2;
    wire c3900;
    assign in3900_1 = {c1727};
    assign in3900_2 = {s1729[2]};
    Half_Adder KS_3900(s3900, c3900, in3900_1, in3900_2);
    wire[2:0] s3901, in3901_1, in3901_2;
    wire c3901;
    assign in3901_1 = {c3843,s1766[0],s1766[1]};
    assign in3901_2 = {c3844,s1767[0],s1767[1]};
    CLA_3 KS_3901(s3901, c3901, in3901_1, in3901_2);
    wire[0:0] s3902, in3902_1, in3902_2;
    wire c3902;
    assign in3902_1 = {c3845};
    assign in3902_2 = {c3846};
    Half_Adder KS_3902(s3902, c3902, in3902_1, in3902_2);
    wire[1:0] s3903, in3903_1, in3903_2;
    wire c3903;
    assign in3903_1 = {c3847,s1768[0]};
    assign in3903_2 = {c3848,s1769[0]};
    CLA_2 KS_3903(s3903, c3903, in3903_1, in3903_2);
    wire[0:0] s3904, in3904_1, in3904_2;
    wire c3904;
    assign in3904_1 = {c3849};
    assign in3904_2 = {c3850};
    Half_Adder KS_3904(s3904, c3904, in3904_1, in3904_2);
    wire[3:0] s3905, in3905_1, in3905_2;
    wire c3905;
    assign in3905_1 = {c3851,s1770[0],s1768[1],c1766};
    assign in3905_2 = {c3852,s3879[1],s1769[1],s1767[2]};
    CLA_4 KS_3905(s3905, c3905, in3905_1, in3905_2);
    wire[0:0] s3906, in3906_1, in3906_2;
    wire c3906;
    assign in3906_1 = {c3853};
    assign in3906_2 = {c3854};
    Half_Adder KS_3906(s3906, c3906, in3906_1, in3906_2);
    wire[1:0] s3907, in3907_1, in3907_2;
    wire c3907;
    assign in3907_1 = {c3855,s3880[1]};
    assign in3907_2 = {c3856,s3881[1]};
    CLA_2 KS_3907(s3907, c3907, in3907_1, in3907_2);
    wire[0:0] s3908, in3908_1, in3908_2;
    wire c3908;
    assign in3908_1 = {c3857};
    assign in3908_2 = {c3858};
    Half_Adder KS_3908(s3908, c3908, in3908_1, in3908_2);
    wire[2:0] s3909, in3909_1, in3909_2;
    wire c3909;
    assign in3909_1 = {c3859,s3882[1],s1770[1]};
    assign in3909_2 = {c3860,s3883[1],s1771[0]};
    CLA_3 KS_3909(s3909, c3909, in3909_1, in3909_2);
    wire[0:0] s3910, in3910_1, in3910_2;
    wire c3910;
    assign in3910_1 = {c3865};
    assign in3910_2 = {c3873};
    Half_Adder KS_3910(s3910, c3910, in3910_1, in3910_2);
    wire[1:0] s3911, in3911_1, in3911_2;
    wire c3911;
    assign in3911_1 = {s3879[0],s3884[1]};
    assign in3911_2 = {s3880[0],s3885[1]};
    CLA_2 KS_3911(s3911, c3911, in3911_1, in3911_2);
    wire[0:0] s3912, in3912_1, in3912_2;
    wire c3912;
    assign in3912_1 = {s3881[0]};
    assign in3912_2 = {s3882[0]};
    Half_Adder KS_3912(s3912, c3912, in3912_1, in3912_2);
    wire[3:0] s3913, in3913_1, in3913_2;
    wire c3913;
    assign in3913_1 = {s3883[0],s3886[1],s1772[0],c1768};
    assign in3913_2 = {s3884[0],s3887[1],s3879[2],s1769[2]};
    CLA_4 KS_3913(s3913, c3913, in3913_1, in3913_2);
    wire[0:0] s3914, in3914_1, in3914_2;
    wire c3914;
    assign in3914_1 = {s3886[0]};
    assign in3914_2 = {s3887[0]};
    Full_Adder KS_3914(s3914, c3914, in3914_1, in3914_2, s3885[0]);
    wire[3:0] s3915, in3915_1, in3915_2;
    wire c3915;
    assign in3915_1 = {s59[1],s1792[0],s1793[1],s1777[2]};
    assign in3915_2 = {s60[1],s1793[0],s1794[1],s1778[2]};
    CLA_4 KS_3915(s3915, c3915, in3915_1, in3915_2);
    wire[3:0] s3916, in3916_1, in3916_2;
    wire c3916;
    assign in3916_1 = {s61[1],s1794[0],s1795[1],s1779[2]};
    assign in3916_2 = {s62[0],s1795[0],s1796[1],s1780[2]};
    CLA_4 KS_3916(s3916, c3916, in3916_1, in3916_2);
    wire[3:0] s3917, in3917_1, in3917_2;
    wire c3917;
    assign in3917_1 = {s63[0],s1796[0],s1797[1],s1781[2]};
    assign in3917_2 = {s64[0],s1797[0],s1798[1],s1782[2]};
    CLA_4 KS_3917(s3917, c3917, in3917_1, in3917_2);
    wire[3:0] s3918, in3918_1, in3918_2;
    wire c3918;
    assign in3918_1 = {s65[0],s1798[0],s1799[1],s1783[2]};
    assign in3918_2 = {s66[0],s1799[0],s1800[1],s1784[2]};
    CLA_4 KS_3918(s3918, c3918, in3918_1, in3918_2);
    wire[3:0] s3919, in3919_1, in3919_2;
    wire c3919;
    assign in3919_1 = {s1730[3],s1800[0],s1801[1],s1785[2]};
    assign in3919_2 = {s1731[3],s1801[0],s1802[1],s1786[2]};
    CLA_4 KS_3919(s3919, c3919, in3919_1, in3919_2);
    wire[3:0] s3920, in3920_1, in3920_2;
    wire c3920;
    assign in3920_1 = {s1732[3],s1802[0],s1803[1],s1787[2]};
    assign in3920_2 = {s1733[3],s1803[0],s1804[1],s1788[2]};
    CLA_4 KS_3920(s3920, c3920, in3920_1, in3920_2);
    wire[3:0] s3921, in3921_1, in3921_2;
    wire c3921;
    assign in3921_1 = {s1734[3],s1804[0],c1805,s1789[2]};
    assign in3921_2 = {s1735[3],s1805[0],s1806[1],s1790[2]};
    CLA_4 KS_3921(s3921, c3921, in3921_1, in3921_2);
    wire[3:0] s3922, in3922_1, in3922_2;
    wire c3922;
    assign in3922_1 = {s1736[3],s1806[0],c1807,s1791[2]};
    assign in3922_2 = {s1737[3],s1807[0],s1808[1],s1792[2]};
    CLA_4 KS_3922(s3922, c3922, in3922_1, in3922_2);
    wire[3:0] s3923, in3923_1, in3923_2;
    wire c3923;
    assign in3923_1 = {s1738[3],s1808[0],c1809,s1793[2]};
    assign in3923_2 = {s1739[3],s1809[0],s1810[1],s1794[2]};
    CLA_4 KS_3923(s3923, c3923, in3923_1, in3923_2);
    wire[3:0] s3924, in3924_1, in3924_2;
    wire c3924;
    assign in3924_1 = {s1740[3],s1810[0],c1811,s1795[2]};
    assign in3924_2 = {s1741[3],s1811[0],s1812[1],s1796[2]};
    CLA_4 KS_3924(s3924, c3924, in3924_1, in3924_2);
    wire[3:0] s3925, in3925_1, in3925_2;
    wire c3925;
    assign in3925_1 = {s1742[3],s1812[0],c1813,s1797[2]};
    assign in3925_2 = {s1743[3],s1813[0],s1814[1],s1798[2]};
    CLA_4 KS_3925(s3925, c3925, in3925_1, in3925_2);
    wire[3:0] s3926, in3926_1, in3926_2;
    wire c3926;
    assign in3926_1 = {s1744[3],s1814[0],c1815,s1799[2]};
    assign in3926_2 = {s1745[3],s1815[0],s1816[1],s1800[2]};
    CLA_4 KS_3926(s3926, c3926, in3926_1, in3926_2);
    wire[3:0] s3927, in3927_1, in3927_2;
    wire c3927;
    assign in3927_1 = {s1746[3],s1816[0],c1817,s1801[2]};
    assign in3927_2 = {s1747[3],s1817[0],s1818[1],s1802[2]};
    CLA_4 KS_3927(s3927, c3927, in3927_1, in3927_2);
    wire[3:0] s3928, in3928_1, in3928_2;
    wire c3928;
    assign in3928_1 = {s1748[3],s1818[0],c1819,s1803[2]};
    assign in3928_2 = {s1749[3],s1819[0],s1820[1],s1804[2]};
    CLA_4 KS_3928(s3928, c3928, in3928_1, in3928_2);
    wire[3:0] s3929, in3929_1, in3929_2;
    wire c3929;
    assign in3929_1 = {s1750[3],s1820[0],c1821,c1806};
    assign in3929_2 = {s1751[3],s1821[0],s1822[1],s1808[2]};
    CLA_4 KS_3929(s3929, c3929, in3929_1, in3929_2);
    wire[3:0] s3930, in3930_1, in3930_2;
    wire c3930;
    assign in3930_1 = {s1752[3],s1822[0],c1823,c1810};
    assign in3930_2 = {s1753[3],s1823[0],s1824[1],s1812[2]};
    CLA_4 KS_3930(s3930, c3930, in3930_1, in3930_2);
    wire[3:0] s3931, in3931_1, in3931_2;
    wire c3931;
    assign in3931_1 = {s1754[3],s1824[0],c1825,c1814};
    assign in3931_2 = {s1755[3],s1825[0],s1826[1],s1816[2]};
    CLA_4 KS_3931(s3931, c3931, in3931_1, in3931_2);
    wire[3:0] s3932, in3932_1, in3932_2;
    wire c3932;
    assign in3932_1 = {s1756[3],s1826[0],c1827,c1818};
    assign in3932_2 = {s1757[3],s1827[0],s1828[1],s1820[2]};
    CLA_4 KS_3932(s3932, c3932, in3932_1, in3932_2);
    wire[1:0] s3933, in3933_1, in3933_2;
    wire c3933;
    assign in3933_1 = {s1758[3],s1828[0]};
    assign in3933_2 = {s1759[3],s1829[0]};
    CLA_2 KS_3933(s3933, c3933, in3933_1, in3933_2);
    wire[0:0] s3934, in3934_1, in3934_2;
    wire c3934;
    assign in3934_1 = {s1760[3]};
    assign in3934_2 = {s1761[3]};
    Half_Adder KS_3934(s3934, c3934, in3934_1, in3934_2);
    wire[2:0] s3935, in3935_1, in3935_2;
    wire c3935;
    assign in3935_1 = {c1763,s1830[0],c1829};
    assign in3935_2 = {s1765[3],s1831[0],s1830[1]};
    CLA_3 KS_3935(s3935, c3935, in3935_1, in3935_2);
    wire[0:0] s3936, in3936_1, in3936_2;
    wire c3936;
    assign in3936_1 = {c1767};
    assign in3936_2 = {s1769[3]};
    Half_Adder KS_3936(s3936, c3936, in3936_1, in3936_2);
    wire[1:0] s3937, in3937_1, in3937_2;
    wire c3937;
    assign in3937_1 = {c1771,s1832[0]};
    assign in3937_2 = {c3879,s1833[0]};
    CLA_2 KS_3937(s3937, c3937, in3937_1, in3937_2);
    wire[0:0] s3938, in3938_1, in3938_2;
    wire c3938;
    assign in3938_1 = {c3880};
    assign in3938_2 = {c3881};
    Half_Adder KS_3938(s3938, c3938, in3938_1, in3938_2);
    wire[3:0] s3939, in3939_1, in3939_2;
    wire c3939;
    assign in3939_1 = {c3882,s1834[0],c1831,c1822};
    assign in3939_2 = {c3883,s1835[0],s1832[1],s1824[2]};
    CLA_4 KS_3939(s3939, c3939, in3939_1, in3939_2);
    wire[0:0] s3940, in3940_1, in3940_2;
    wire c3940;
    assign in3940_1 = {c3884};
    assign in3940_2 = {c3885};
    Half_Adder KS_3940(s3940, c3940, in3940_1, in3940_2);
    wire[1:0] s3941, in3941_1, in3941_2;
    wire c3941;
    assign in3941_1 = {c3886,s1836[0]};
    assign in3941_2 = {c3887,s3915[1]};
    CLA_2 KS_3941(s3941, c3941, in3941_1, in3941_2);
    wire[0:0] s3942, in3942_1, in3942_2;
    wire c3942;
    assign in3942_1 = {c3888};
    assign in3942_2 = {c3889};
    Half_Adder KS_3942(s3942, c3942, in3942_1, in3942_2);
    wire[2:0] s3943, in3943_1, in3943_2;
    wire c3943;
    assign in3943_1 = {c3890,s3916[1],c1833};
    assign in3943_2 = {c3891,s3917[1],s1834[1]};
    CLA_3 KS_3943(s3943, c3943, in3943_1, in3943_2);
    wire[0:0] s3944, in3944_1, in3944_2;
    wire c3944;
    assign in3944_1 = {c3892};
    assign in3944_2 = {c3893};
    Half_Adder KS_3944(s3944, c3944, in3944_1, in3944_2);
    wire[1:0] s3945, in3945_1, in3945_2;
    wire c3945;
    assign in3945_1 = {c3894,s3918[1]};
    assign in3945_2 = {c3895,s3919[1]};
    CLA_2 KS_3945(s3945, c3945, in3945_1, in3945_2);
    wire[0:0] s3946, in3946_1, in3946_2;
    wire c3946;
    assign in3946_1 = {c3896};
    assign in3946_2 = {c3897};
    Half_Adder KS_3946(s3946, c3946, in3946_1, in3946_2);
    wire[3:0] s3947, in3947_1, in3947_2;
    wire c3947;
    assign in3947_1 = {c3905,s3920[1],c1835,c1826};
    assign in3947_2 = {c3913,s3921[1],s1836[1],s1828[2]};
    CLA_4 KS_3947(s3947, c3947, in3947_1, in3947_2);
    wire[0:0] s3948, in3948_1, in3948_2;
    wire c3948;
    assign in3948_1 = {s3915[0]};
    assign in3948_2 = {s3916[0]};
    Half_Adder KS_3948(s3948, c3948, in3948_1, in3948_2);
    wire[1:0] s3949, in3949_1, in3949_2;
    wire c3949;
    assign in3949_1 = {s3917[0],s3922[1]};
    assign in3949_2 = {s3918[0],s3923[1]};
    CLA_2 KS_3949(s3949, c3949, in3949_1, in3949_2);
    wire[0:0] s3950, in3950_1, in3950_2;
    wire c3950;
    assign in3950_1 = {s3919[0]};
    assign in3950_2 = {s3920[0]};
    Half_Adder KS_3950(s3950, c3950, in3950_1, in3950_2);
    wire[2:0] s3951, in3951_1, in3951_2;
    wire c3951;
    assign in3951_1 = {s3921[0],s3924[1],s3915[2]};
    assign in3951_2 = {s3922[0],s3925[1],s3916[2]};
    CLA_3 KS_3951(s3951, c3951, in3951_1, in3951_2);
    wire[0:0] s3952, in3952_1, in3952_2;
    wire c3952;
    assign in3952_1 = {s3924[0]};
    assign in3952_2 = {s3925[0]};
    Full_Adder KS_3952(s3952, c3952, in3952_1, in3952_2, s3923[0]);
    wire[3:0] s3953, in3953_1, in3953_2;
    wire c3953;
    assign in3953_1 = {s95[0],s1858[0],s1858[1],s1841[2]};
    assign in3953_2 = {s96[0],s1859[0],s1859[1],s1842[2]};
    CLA_4 KS_3953(s3953, c3953, in3953_1, in3953_2);
    wire[3:0] s3954, in3954_1, in3954_2;
    wire c3954;
    assign in3954_1 = {s97[0],s1860[0],s1860[1],s1843[2]};
    assign in3954_2 = {s98[0],s1861[0],s1861[1],s1844[2]};
    CLA_4 KS_3954(s3954, c3954, in3954_1, in3954_2);
    wire[3:0] s3955, in3955_1, in3955_2;
    wire c3955;
    assign in3955_1 = {s1773[3],s1862[0],s1862[1],s1845[2]};
    assign in3955_2 = {s1774[3],s1863[0],s1863[1],s1846[2]};
    CLA_4 KS_3955(s3955, c3955, in3955_1, in3955_2);
    wire[3:0] s3956, in3956_1, in3956_2;
    wire c3956;
    assign in3956_1 = {s1775[3],s1864[0],s1864[1],s1847[2]};
    assign in3956_2 = {s1776[3],s1865[0],s1865[1],s1848[2]};
    CLA_4 KS_3956(s3956, c3956, in3956_1, in3956_2);
    wire[3:0] s3957, in3957_1, in3957_2;
    wire c3957;
    assign in3957_1 = {s1777[3],s1866[0],s1866[1],s1849[2]};
    assign in3957_2 = {s1778[3],s1867[0],s1867[1],s1850[2]};
    CLA_4 KS_3957(s3957, c3957, in3957_1, in3957_2);
    wire[3:0] s3958, in3958_1, in3958_2;
    wire c3958;
    assign in3958_1 = {s1779[3],s1868[0],c1868,s1851[2]};
    assign in3958_2 = {s1780[3],s1869[0],s1869[1],s1852[2]};
    CLA_4 KS_3958(s3958, c3958, in3958_1, in3958_2);
    wire[3:0] s3959, in3959_1, in3959_2;
    wire c3959;
    assign in3959_1 = {s1781[3],s1870[0],c1870,s1853[2]};
    assign in3959_2 = {s1782[3],s1871[0],s1871[1],s1854[2]};
    CLA_4 KS_3959(s3959, c3959, in3959_1, in3959_2);
    wire[3:0] s3960, in3960_1, in3960_2;
    wire c3960;
    assign in3960_1 = {s1783[3],s1872[0],c1872,s1855[2]};
    assign in3960_2 = {s1784[3],s1873[0],s1873[1],s1856[2]};
    CLA_4 KS_3960(s3960, c3960, in3960_1, in3960_2);
    wire[3:0] s3961, in3961_1, in3961_2;
    wire c3961;
    assign in3961_1 = {s1785[3],s1874[0],c1874,s1857[2]};
    assign in3961_2 = {s1786[3],s1875[0],s1875[1],s1858[2]};
    CLA_4 KS_3961(s3961, c3961, in3961_1, in3961_2);
    wire[3:0] s3962, in3962_1, in3962_2;
    wire c3962;
    assign in3962_1 = {s1787[3],s1876[0],c1876,s1859[2]};
    assign in3962_2 = {s1788[3],s1877[0],s1877[1],s1860[2]};
    CLA_4 KS_3962(s3962, c3962, in3962_1, in3962_2);
    wire[3:0] s3963, in3963_1, in3963_2;
    wire c3963;
    assign in3963_1 = {s1789[3],s1878[0],c1878,s1861[2]};
    assign in3963_2 = {s1790[3],s1879[0],s1879[1],s1862[2]};
    CLA_4 KS_3963(s3963, c3963, in3963_1, in3963_2);
    wire[3:0] s3964, in3964_1, in3964_2;
    wire c3964;
    assign in3964_1 = {s1791[3],s1880[0],c1880,s1863[2]};
    assign in3964_2 = {s1792[3],s1881[0],s1881[1],s1864[2]};
    CLA_4 KS_3964(s3964, c3964, in3964_1, in3964_2);
    wire[3:0] s3965, in3965_1, in3965_2;
    wire c3965;
    assign in3965_1 = {s1793[3],s1882[0],c1882,s1865[2]};
    assign in3965_2 = {s1794[3],s1883[0],s1883[1],s1866[2]};
    CLA_4 KS_3965(s3965, c3965, in3965_1, in3965_2);
    wire[3:0] s3966, in3966_1, in3966_2;
    wire c3966;
    assign in3966_1 = {s1795[3],s1884[0],c1884,s1867[2]};
    assign in3966_2 = {s1796[3],s1885[0],s1885[1],s1869[2]};
    CLA_4 KS_3966(s3966, c3966, in3966_1, in3966_2);
    wire[3:0] s3967, in3967_1, in3967_2;
    wire c3967;
    assign in3967_1 = {s1797[3],s1886[0],c1886,c1871};
    assign in3967_2 = {s1798[3],s1887[0],s1887[1],s1873[2]};
    CLA_4 KS_3967(s3967, c3967, in3967_1, in3967_2);
    wire[3:0] s3968, in3968_1, in3968_2;
    wire c3968;
    assign in3968_1 = {s1799[3],s1888[0],c1888,c1875};
    assign in3968_2 = {s1800[3],s1889[0],s1889[1],s1877[2]};
    CLA_4 KS_3968(s3968, c3968, in3968_1, in3968_2);
    wire[3:0] s3969, in3969_1, in3969_2;
    wire c3969;
    assign in3969_1 = {s1801[3],s1890[0],c1890,c1879};
    assign in3969_2 = {s1802[3],s1891[0],s1891[1],s1881[2]};
    CLA_4 KS_3969(s3969, c3969, in3969_1, in3969_2);
    wire[3:0] s3970, in3970_1, in3970_2;
    wire c3970;
    assign in3970_1 = {s1803[3],s1892[0],c1892,c1883};
    assign in3970_2 = {s1804[3],s1893[0],s1893[1],s1885[2]};
    CLA_4 KS_3970(s3970, c3970, in3970_1, in3970_2);
    wire[2:0] s3971, in3971_1, in3971_2;
    wire c3971;
    assign in3971_1 = {c1808,s1894[0],c1894};
    assign in3971_2 = {s1812[3],s1895[0],s1895[1]};
    CLA_3 KS_3971(s3971, c3971, in3971_1, in3971_2);
    wire[0:0] s3972, in3972_1, in3972_2;
    wire c3972;
    assign in3972_1 = {c1816};
    assign in3972_2 = {s1820[3]};
    Half_Adder KS_3972(s3972, c3972, in3972_1, in3972_2);
    wire[1:0] s3973, in3973_1, in3973_2;
    wire c3973;
    assign in3973_1 = {c1824,s1896[0]};
    assign in3973_2 = {s1828[3],s1897[0]};
    CLA_2 KS_3973(s3973, c3973, in3973_1, in3973_2);
    wire[0:0] s3974, in3974_1, in3974_2;
    wire c3974;
    assign in3974_1 = {c1832};
    assign in3974_2 = {s1836[3]};
    Half_Adder KS_3974(s3974, c3974, in3974_1, in3974_2);
    wire[3:0] s3975, in3975_1, in3975_2;
    wire c3975;
    assign in3975_1 = {c3915,s1898[0],c1896,c1887};
    assign in3975_2 = {c3916,s1899[0],s1897[1],s1889[2]};
    CLA_4 KS_3975(s3975, c3975, in3975_1, in3975_2);
    wire[0:0] s3976, in3976_1, in3976_2;
    wire c3976;
    assign in3976_1 = {c3917};
    assign in3976_2 = {c3918};
    Half_Adder KS_3976(s3976, c3976, in3976_1, in3976_2);
    wire[1:0] s3977, in3977_1, in3977_2;
    wire c3977;
    assign in3977_1 = {c3919,s1900[0]};
    assign in3977_2 = {c3920,s1901[0]};
    CLA_2 KS_3977(s3977, c3977, in3977_1, in3977_2);
    wire[0:0] s3978, in3978_1, in3978_2;
    wire c3978;
    assign in3978_1 = {c3921};
    assign in3978_2 = {c3922};
    Half_Adder KS_3978(s3978, c3978, in3978_1, in3978_2);
    wire[2:0] s3979, in3979_1, in3979_2;
    wire c3979;
    assign in3979_1 = {c3923,s1902[0],c1898};
    assign in3979_2 = {c3924,s3953[1],s1899[1]};
    CLA_3 KS_3979(s3979, c3979, in3979_1, in3979_2);
    wire[0:0] s3980, in3980_1, in3980_2;
    wire c3980;
    assign in3980_1 = {c3925};
    assign in3980_2 = {c3926};
    Half_Adder KS_3980(s3980, c3980, in3980_1, in3980_2);
    wire[1:0] s3981, in3981_1, in3981_2;
    wire c3981;
    assign in3981_1 = {c3927,s3954[1]};
    assign in3981_2 = {c3928,s3955[1]};
    CLA_2 KS_3981(s3981, c3981, in3981_1, in3981_2);
    wire[0:0] s3982, in3982_1, in3982_2;
    wire c3982;
    assign in3982_1 = {c3929};
    assign in3982_2 = {c3930};
    Half_Adder KS_3982(s3982, c3982, in3982_1, in3982_2);
    wire[3:0] s3983, in3983_1, in3983_2;
    wire c3983;
    assign in3983_1 = {c3931,s3956[1],c1900,c1891};
    assign in3983_2 = {c3932,s3957[1],s1901[1],s1893[2]};
    CLA_4 KS_3983(s3983, c3983, in3983_1, in3983_2);
    wire[0:0] s3984, in3984_1, in3984_2;
    wire c3984;
    assign in3984_1 = {c3939};
    assign in3984_2 = {c3947};
    Half_Adder KS_3984(s3984, c3984, in3984_1, in3984_2);
    wire[1:0] s3985, in3985_1, in3985_2;
    wire c3985;
    assign in3985_1 = {s3953[0],s3958[1]};
    assign in3985_2 = {s3954[0],s3959[1]};
    CLA_2 KS_3985(s3985, c3985, in3985_1, in3985_2);
    wire[0:0] s3986, in3986_1, in3986_2;
    wire c3986;
    assign in3986_1 = {s3955[0]};
    assign in3986_2 = {s3956[0]};
    Half_Adder KS_3986(s3986, c3986, in3986_1, in3986_2);
    wire[2:0] s3987, in3987_1, in3987_2;
    wire c3987;
    assign in3987_1 = {s3957[0],s3960[1],c1902};
    assign in3987_2 = {s3958[0],s3961[1],s3953[2]};
    CLA_3 KS_3987(s3987, c3987, in3987_1, in3987_2);
    wire[0:0] s3988, in3988_1, in3988_2;
    wire c3988;
    assign in3988_1 = {s3960[0]};
    assign in3988_2 = {s3961[0]};
    Full_Adder KS_3988(s3988, c3988, in3988_1, in3988_2, s3959[0]);
    wire[3:0] s3989, in3989_1, in3989_2;
    wire c3989;
    assign in3989_1 = {s135[0],s1924[0],s1924[1],s1907[2]};
    assign in3989_2 = {s136[0],s1925[0],s1925[1],s1908[2]};
    CLA_4 KS_3989(s3989, c3989, in3989_1, in3989_2);
    wire[3:0] s3990, in3990_1, in3990_2;
    wire c3990;
    assign in3990_1 = {s137[0],s1926[0],s1926[1],s1909[2]};
    assign in3990_2 = {s138[0],s1927[0],s1927[1],s1910[2]};
    CLA_4 KS_3990(s3990, c3990, in3990_1, in3990_2);
    wire[3:0] s3991, in3991_1, in3991_2;
    wire c3991;
    assign in3991_1 = {s1837[3],s1928[0],s1928[1],s1911[2]};
    assign in3991_2 = {s1838[3],s1929[0],s1929[1],s1912[2]};
    CLA_4 KS_3991(s3991, c3991, in3991_1, in3991_2);
    wire[3:0] s3992, in3992_1, in3992_2;
    wire c3992;
    assign in3992_1 = {s1839[3],s1930[0],s1930[1],s1913[2]};
    assign in3992_2 = {s1840[3],s1931[0],s1931[1],s1914[2]};
    CLA_4 KS_3992(s3992, c3992, in3992_1, in3992_2);
    wire[3:0] s3993, in3993_1, in3993_2;
    wire c3993;
    assign in3993_1 = {s1841[3],s1932[0],s1932[1],s1915[2]};
    assign in3993_2 = {s1842[3],s1933[0],s1933[1],s1916[2]};
    CLA_4 KS_3993(s3993, c3993, in3993_1, in3993_2);
    wire[3:0] s3994, in3994_1, in3994_2;
    wire c3994;
    assign in3994_1 = {s1843[3],s1934[0],c1934,s1917[2]};
    assign in3994_2 = {s1844[3],s1935[0],s1935[1],s1918[2]};
    CLA_4 KS_3994(s3994, c3994, in3994_1, in3994_2);
    wire[3:0] s3995, in3995_1, in3995_2;
    wire c3995;
    assign in3995_1 = {s1845[3],s1936[0],c1936,s1919[2]};
    assign in3995_2 = {s1846[3],s1937[0],s1937[1],s1920[2]};
    CLA_4 KS_3995(s3995, c3995, in3995_1, in3995_2);
    wire[3:0] s3996, in3996_1, in3996_2;
    wire c3996;
    assign in3996_1 = {s1847[3],s1938[0],c1938,s1921[2]};
    assign in3996_2 = {s1848[3],s1939[0],s1939[1],s1922[2]};
    CLA_4 KS_3996(s3996, c3996, in3996_1, in3996_2);
    wire[3:0] s3997, in3997_1, in3997_2;
    wire c3997;
    assign in3997_1 = {s1849[3],s1940[0],c1940,s1923[2]};
    assign in3997_2 = {s1850[3],s1941[0],s1941[1],s1924[2]};
    CLA_4 KS_3997(s3997, c3997, in3997_1, in3997_2);
    wire[3:0] s3998, in3998_1, in3998_2;
    wire c3998;
    assign in3998_1 = {s1851[3],s1942[0],c1942,s1925[2]};
    assign in3998_2 = {s1852[3],s1943[0],s1943[1],s1926[2]};
    CLA_4 KS_3998(s3998, c3998, in3998_1, in3998_2);
    wire[3:0] s3999, in3999_1, in3999_2;
    wire c3999;
    assign in3999_1 = {s1853[3],s1944[0],c1944,s1927[2]};
    assign in3999_2 = {s1854[3],s1945[0],s1945[1],s1928[2]};
    CLA_4 KS_3999(s3999, c3999, in3999_1, in3999_2);
    wire[3:0] s4000, in4000_1, in4000_2;
    wire c4000;
    assign in4000_1 = {s1855[3],s1946[0],c1946,s1929[2]};
    assign in4000_2 = {s1856[3],s1947[0],s1947[1],s1930[2]};
    CLA_4 KS_4000(s4000, c4000, in4000_1, in4000_2);
    wire[3:0] s4001, in4001_1, in4001_2;
    wire c4001;
    assign in4001_1 = {s1857[3],s1948[0],c1948,s1931[2]};
    assign in4001_2 = {s1858[3],s1949[0],s1949[1],s1932[2]};
    CLA_4 KS_4001(s4001, c4001, in4001_1, in4001_2);
    wire[3:0] s4002, in4002_1, in4002_2;
    wire c4002;
    assign in4002_1 = {s1859[3],s1950[0],c1950,s1933[2]};
    assign in4002_2 = {s1860[3],s1951[0],s1951[1],s1935[2]};
    CLA_4 KS_4002(s4002, c4002, in4002_1, in4002_2);
    wire[3:0] s4003, in4003_1, in4003_2;
    wire c4003;
    assign in4003_1 = {s1861[3],s1952[0],c1952,c1937};
    assign in4003_2 = {s1862[3],s1953[0],s1953[1],s1939[2]};
    CLA_4 KS_4003(s4003, c4003, in4003_1, in4003_2);
    wire[3:0] s4004, in4004_1, in4004_2;
    wire c4004;
    assign in4004_1 = {s1863[3],s1954[0],c1954,c1941};
    assign in4004_2 = {s1864[3],s1955[0],s1955[1],s1943[2]};
    CLA_4 KS_4004(s4004, c4004, in4004_1, in4004_2);
    wire[3:0] s4005, in4005_1, in4005_2;
    wire c4005;
    assign in4005_1 = {s1865[3],s1956[0],c1956,c1945};
    assign in4005_2 = {s1866[3],s1957[0],s1957[1],s1947[2]};
    CLA_4 KS_4005(s4005, c4005, in4005_1, in4005_2);
    wire[3:0] s4006, in4006_1, in4006_2;
    wire c4006;
    assign in4006_1 = {s1867[3],s1958[0],c1958,c1949};
    assign in4006_2 = {s1869[3],s1959[0],s1959[1],s1951[2]};
    CLA_4 KS_4006(s4006, c4006, in4006_1, in4006_2);
    wire[2:0] s4007, in4007_1, in4007_2;
    wire c4007;
    assign in4007_1 = {c1873,s1960[0],c1960};
    assign in4007_2 = {s1877[3],s1961[0],s1961[1]};
    CLA_3 KS_4007(s4007, c4007, in4007_1, in4007_2);
    wire[0:0] s4008, in4008_1, in4008_2;
    wire c4008;
    assign in4008_1 = {c1881};
    assign in4008_2 = {s1885[3]};
    Half_Adder KS_4008(s4008, c4008, in4008_1, in4008_2);
    wire[1:0] s4009, in4009_1, in4009_2;
    wire c4009;
    assign in4009_1 = {c1889,s1962[0]};
    assign in4009_2 = {s1893[3],s1963[0]};
    CLA_2 KS_4009(s4009, c4009, in4009_1, in4009_2);
    wire[0:0] s4010, in4010_1, in4010_2;
    wire c4010;
    assign in4010_1 = {c1897};
    assign in4010_2 = {s1901[3]};
    Half_Adder KS_4010(s4010, c4010, in4010_1, in4010_2);
    wire[3:0] s4011, in4011_1, in4011_2;
    wire c4011;
    assign in4011_1 = {c3953,s1964[0],c1962,c1953};
    assign in4011_2 = {c3954,s1965[0],s1963[1],s1955[2]};
    CLA_4 KS_4011(s4011, c4011, in4011_1, in4011_2);
    wire[0:0] s4012, in4012_1, in4012_2;
    wire c4012;
    assign in4012_1 = {c3955};
    assign in4012_2 = {c3956};
    Half_Adder KS_4012(s4012, c4012, in4012_1, in4012_2);
    wire[1:0] s4013, in4013_1, in4013_2;
    wire c4013;
    assign in4013_1 = {c3957,s1966[0]};
    assign in4013_2 = {c3958,s1967[0]};
    CLA_2 KS_4013(s4013, c4013, in4013_1, in4013_2);
    wire[0:0] s4014, in4014_1, in4014_2;
    wire c4014;
    assign in4014_1 = {c3959};
    assign in4014_2 = {c3960};
    Half_Adder KS_4014(s4014, c4014, in4014_1, in4014_2);
    wire[2:0] s4015, in4015_1, in4015_2;
    wire c4015;
    assign in4015_1 = {c3961,s1968[0],c1964};
    assign in4015_2 = {c3962,s3989[1],s1965[1]};
    CLA_3 KS_4015(s4015, c4015, in4015_1, in4015_2);
    wire[0:0] s4016, in4016_1, in4016_2;
    wire c4016;
    assign in4016_1 = {c3963};
    assign in4016_2 = {c3964};
    Half_Adder KS_4016(s4016, c4016, in4016_1, in4016_2);
    wire[1:0] s4017, in4017_1, in4017_2;
    wire c4017;
    assign in4017_1 = {c3965,s3990[1]};
    assign in4017_2 = {c3966,s3991[1]};
    CLA_2 KS_4017(s4017, c4017, in4017_1, in4017_2);
    wire[0:0] s4018, in4018_1, in4018_2;
    wire c4018;
    assign in4018_1 = {c3967};
    assign in4018_2 = {c3968};
    Half_Adder KS_4018(s4018, c4018, in4018_1, in4018_2);
    wire[3:0] s4019, in4019_1, in4019_2;
    wire c4019;
    assign in4019_1 = {c3969,s3992[1],c1966,c1957};
    assign in4019_2 = {c3970,s3993[1],s1967[1],s1959[2]};
    CLA_4 KS_4019(s4019, c4019, in4019_1, in4019_2);
    wire[0:0] s4020, in4020_1, in4020_2;
    wire c4020;
    assign in4020_1 = {c3975};
    assign in4020_2 = {c3983};
    Half_Adder KS_4020(s4020, c4020, in4020_1, in4020_2);
    wire[1:0] s4021, in4021_1, in4021_2;
    wire c4021;
    assign in4021_1 = {s3989[0],s3994[1]};
    assign in4021_2 = {s3990[0],s3995[1]};
    CLA_2 KS_4021(s4021, c4021, in4021_1, in4021_2);
    wire[0:0] s4022, in4022_1, in4022_2;
    wire c4022;
    assign in4022_1 = {s3991[0]};
    assign in4022_2 = {s3992[0]};
    Half_Adder KS_4022(s4022, c4022, in4022_1, in4022_2);
    wire[2:0] s4023, in4023_1, in4023_2;
    wire c4023;
    assign in4023_1 = {s3993[0],s3996[1],c1968};
    assign in4023_2 = {s3994[0],s3997[1],s3989[2]};
    CLA_3 KS_4023(s4023, c4023, in4023_1, in4023_2);
    wire[0:0] s4024, in4024_1, in4024_2;
    wire c4024;
    assign in4024_1 = {s3996[0]};
    assign in4024_2 = {s3997[0]};
    Full_Adder KS_4024(s4024, c4024, in4024_1, in4024_2, s3995[0]);
    wire[3:0] s4025, in4025_1, in4025_2;
    wire c4025;
    assign in4025_1 = {s187[0],s1990[0],s1991[1],s1973[2]};
    assign in4025_2 = {s188[0],s1991[0],s1992[1],s1974[2]};
    CLA_4 KS_4025(s4025, c4025, in4025_1, in4025_2);
    wire[3:0] s4026, in4026_1, in4026_2;
    wire c4026;
    assign in4026_1 = {s189[0],s1992[0],s1993[1],s1975[2]};
    assign in4026_2 = {s190[0],s1993[0],s1994[1],s1976[2]};
    CLA_4 KS_4026(s4026, c4026, in4026_1, in4026_2);
    wire[3:0] s4027, in4027_1, in4027_2;
    wire c4027;
    assign in4027_1 = {s1903[3],s1994[0],s1995[1],s1977[2]};
    assign in4027_2 = {s1904[3],s1995[0],s1996[1],s1978[2]};
    CLA_4 KS_4027(s4027, c4027, in4027_1, in4027_2);
    wire[3:0] s4028, in4028_1, in4028_2;
    wire c4028;
    assign in4028_1 = {s1905[3],s1996[0],s1997[1],s1979[2]};
    assign in4028_2 = {s1906[3],s1997[0],s1998[1],s1980[2]};
    CLA_4 KS_4028(s4028, c4028, in4028_1, in4028_2);
    wire[3:0] s4029, in4029_1, in4029_2;
    wire c4029;
    assign in4029_1 = {s1907[3],s1998[0],s1999[1],s1981[2]};
    assign in4029_2 = {s1908[3],s1999[0],s2000[1],s1982[2]};
    CLA_4 KS_4029(s4029, c4029, in4029_1, in4029_2);
    wire[3:0] s4030, in4030_1, in4030_2;
    wire c4030;
    assign in4030_1 = {s1909[3],s2000[0],c2001,s1983[2]};
    assign in4030_2 = {s1910[3],s2001[0],s2002[1],s1984[2]};
    CLA_4 KS_4030(s4030, c4030, in4030_1, in4030_2);
    wire[3:0] s4031, in4031_1, in4031_2;
    wire c4031;
    assign in4031_1 = {s1911[3],s2002[0],c2003,s1985[2]};
    assign in4031_2 = {s1912[3],s2003[0],s2004[1],s1986[2]};
    CLA_4 KS_4031(s4031, c4031, in4031_1, in4031_2);
    wire[3:0] s4032, in4032_1, in4032_2;
    wire c4032;
    assign in4032_1 = {s1913[3],s2004[0],c2005,s1987[2]};
    assign in4032_2 = {s1914[3],s2005[0],s2006[1],s1988[2]};
    CLA_4 KS_4032(s4032, c4032, in4032_1, in4032_2);
    wire[3:0] s4033, in4033_1, in4033_2;
    wire c4033;
    assign in4033_1 = {s1915[3],s2006[0],c2007,s1989[2]};
    assign in4033_2 = {s1916[3],s2007[0],s2008[1],s1990[2]};
    CLA_4 KS_4033(s4033, c4033, in4033_1, in4033_2);
    wire[3:0] s4034, in4034_1, in4034_2;
    wire c4034;
    assign in4034_1 = {s1917[3],s2008[0],c2009,s1991[2]};
    assign in4034_2 = {s1918[3],s2009[0],s2010[1],s1992[2]};
    CLA_4 KS_4034(s4034, c4034, in4034_1, in4034_2);
    wire[3:0] s4035, in4035_1, in4035_2;
    wire c4035;
    assign in4035_1 = {s1919[3],s2010[0],c2011,s1993[2]};
    assign in4035_2 = {s1920[3],s2011[0],s2012[1],s1994[2]};
    CLA_4 KS_4035(s4035, c4035, in4035_1, in4035_2);
    wire[3:0] s4036, in4036_1, in4036_2;
    wire c4036;
    assign in4036_1 = {s1921[3],s2012[0],c2013,s1995[2]};
    assign in4036_2 = {s1922[3],s2013[0],s2014[1],s1996[2]};
    CLA_4 KS_4036(s4036, c4036, in4036_1, in4036_2);
    wire[3:0] s4037, in4037_1, in4037_2;
    wire c4037;
    assign in4037_1 = {s1923[3],s2014[0],c2015,s1997[2]};
    assign in4037_2 = {s1924[3],s2015[0],s2016[1],s1998[2]};
    CLA_4 KS_4037(s4037, c4037, in4037_1, in4037_2);
    wire[3:0] s4038, in4038_1, in4038_2;
    wire c4038;
    assign in4038_1 = {s1925[3],s2016[0],c2017,s1999[2]};
    assign in4038_2 = {s1926[3],s2017[0],s2018[1],s2000[2]};
    CLA_4 KS_4038(s4038, c4038, in4038_1, in4038_2);
    wire[3:0] s4039, in4039_1, in4039_2;
    wire c4039;
    assign in4039_1 = {s1927[3],s2018[0],c2019,c2002};
    assign in4039_2 = {s1928[3],s2019[0],s2020[1],s2004[2]};
    CLA_4 KS_4039(s4039, c4039, in4039_1, in4039_2);
    wire[3:0] s4040, in4040_1, in4040_2;
    wire c4040;
    assign in4040_1 = {s1929[3],s2020[0],c2021,c2006};
    assign in4040_2 = {s1930[3],s2021[0],s2022[1],s2008[2]};
    CLA_4 KS_4040(s4040, c4040, in4040_1, in4040_2);
    wire[3:0] s4041, in4041_1, in4041_2;
    wire c4041;
    assign in4041_1 = {s1931[3],s2022[0],c2023,c2010};
    assign in4041_2 = {s1932[3],s2023[0],s2024[1],s2012[2]};
    CLA_4 KS_4041(s4041, c4041, in4041_1, in4041_2);
    wire[3:0] s4042, in4042_1, in4042_2;
    wire c4042;
    assign in4042_1 = {s1933[3],s2024[0],c2025,c2014};
    assign in4042_2 = {s1935[3],s2025[0],s2026[1],s2016[2]};
    CLA_4 KS_4042(s4042, c4042, in4042_1, in4042_2);
    wire[1:0] s4043, in4043_1, in4043_2;
    wire c4043;
    assign in4043_1 = {c1939,s2026[0]};
    assign in4043_2 = {s1943[3],s2027[0]};
    CLA_2 KS_4043(s4043, c4043, in4043_1, in4043_2);
    wire[0:0] s4044, in4044_1, in4044_2;
    wire c4044;
    assign in4044_1 = {c1947};
    assign in4044_2 = {s1951[3]};
    Half_Adder KS_4044(s4044, c4044, in4044_1, in4044_2);
    wire[3:0] s4045, in4045_1, in4045_2;
    wire c4045;
    assign in4045_1 = {c1955,s2028[0],c2027,c2018};
    assign in4045_2 = {s1959[3],s2029[0],s2028[1],s2020[2]};
    CLA_4 KS_4045(s4045, c4045, in4045_1, in4045_2);
    wire[0:0] s4046, in4046_1, in4046_2;
    wire c4046;
    assign in4046_1 = {c1963};
    assign in4046_2 = {s1967[3]};
    Half_Adder KS_4046(s4046, c4046, in4046_1, in4046_2);
    wire[1:0] s4047, in4047_1, in4047_2;
    wire c4047;
    assign in4047_1 = {c3989,s2030[0]};
    assign in4047_2 = {c3990,s2031[0]};
    CLA_2 KS_4047(s4047, c4047, in4047_1, in4047_2);
    wire[0:0] s4048, in4048_1, in4048_2;
    wire c4048;
    assign in4048_1 = {c3991};
    assign in4048_2 = {c3992};
    Half_Adder KS_4048(s4048, c4048, in4048_1, in4048_2);
    wire[2:0] s4049, in4049_1, in4049_2;
    wire c4049;
    assign in4049_1 = {c3993,s2032[0],c2029};
    assign in4049_2 = {c3994,s2033[0],s2030[1]};
    CLA_3 KS_4049(s4049, c4049, in4049_1, in4049_2);
    wire[0:0] s4050, in4050_1, in4050_2;
    wire c4050;
    assign in4050_1 = {c3995};
    assign in4050_2 = {c3996};
    Half_Adder KS_4050(s4050, c4050, in4050_1, in4050_2);
    wire[1:0] s4051, in4051_1, in4051_2;
    wire c4051;
    assign in4051_1 = {c3997,s2034[0]};
    assign in4051_2 = {c3998,s4025[1]};
    CLA_2 KS_4051(s4051, c4051, in4051_1, in4051_2);
    wire[0:0] s4052, in4052_1, in4052_2;
    wire c4052;
    assign in4052_1 = {c3999};
    assign in4052_2 = {c4000};
    Half_Adder KS_4052(s4052, c4052, in4052_1, in4052_2);
    wire[3:0] s4053, in4053_1, in4053_2;
    wire c4053;
    assign in4053_1 = {c4001,s4026[1],c2031,c2022};
    assign in4053_2 = {c4002,s4027[1],s2032[1],s2024[2]};
    CLA_4 KS_4053(s4053, c4053, in4053_1, in4053_2);
    wire[0:0] s4054, in4054_1, in4054_2;
    wire c4054;
    assign in4054_1 = {c4003};
    assign in4054_2 = {c4004};
    Half_Adder KS_4054(s4054, c4054, in4054_1, in4054_2);
    wire[1:0] s4055, in4055_1, in4055_2;
    wire c4055;
    assign in4055_1 = {c4005,s4028[1]};
    assign in4055_2 = {c4006,s4029[1]};
    CLA_2 KS_4055(s4055, c4055, in4055_1, in4055_2);
    wire[0:0] s4056, in4056_1, in4056_2;
    wire c4056;
    assign in4056_1 = {c4011};
    assign in4056_2 = {c4019};
    Half_Adder KS_4056(s4056, c4056, in4056_1, in4056_2);
    wire[2:0] s4057, in4057_1, in4057_2;
    wire c4057;
    assign in4057_1 = {s4025[0],s4030[1],c2033};
    assign in4057_2 = {s4026[0],s4031[1],s2034[1]};
    CLA_3 KS_4057(s4057, c4057, in4057_1, in4057_2);
    wire[0:0] s4058, in4058_1, in4058_2;
    wire c4058;
    assign in4058_1 = {s4027[0]};
    assign in4058_2 = {s4028[0]};
    Half_Adder KS_4058(s4058, c4058, in4058_1, in4058_2);
    wire[1:0] s4059, in4059_1, in4059_2;
    wire c4059;
    assign in4059_1 = {s4029[0],s4032[1]};
    assign in4059_2 = {s4030[0],s4033[1]};
    CLA_2 KS_4059(s4059, c4059, in4059_1, in4059_2);
    wire[0:0] s4060, in4060_1, in4060_2;
    wire c4060;
    assign in4060_1 = {s4032[0]};
    assign in4060_2 = {s4033[0]};
    Full_Adder KS_4060(s4060, c4060, in4060_1, in4060_2, s4031[0]);
    wire[3:0] s4061, in4061_1, in4061_2;
    wire c4061;
    assign in4061_1 = {s252[0],s2056[0],s2057[1],s2040[2]};
    assign in4061_2 = {s253[0],s2057[0],s2058[1],s2041[2]};
    CLA_4 KS_4061(s4061, c4061, in4061_1, in4061_2);
    wire[3:0] s4062, in4062_1, in4062_2;
    wire c4062;
    assign in4062_1 = {s254[0],s2058[0],s2059[1],s2042[2]};
    assign in4062_2 = {s255[0],s2059[0],s2060[1],s2043[2]};
    CLA_4 KS_4062(s4062, c4062, in4062_1, in4062_2);
    wire[3:0] s4063, in4063_1, in4063_2;
    wire c4063;
    assign in4063_1 = {s1969[3],s2060[0],s2061[1],s2044[2]};
    assign in4063_2 = {s1970[3],s2061[0],s2062[1],s2045[2]};
    CLA_4 KS_4063(s4063, c4063, in4063_1, in4063_2);
    wire[3:0] s4064, in4064_1, in4064_2;
    wire c4064;
    assign in4064_1 = {s1971[3],s2062[0],s2063[1],s2046[2]};
    assign in4064_2 = {s1972[3],s2063[0],s2064[1],s2047[2]};
    CLA_4 KS_4064(s4064, c4064, in4064_1, in4064_2);
    wire[3:0] s4065, in4065_1, in4065_2;
    wire c4065;
    assign in4065_1 = {s1973[3],s2064[0],s2065[1],s2048[2]};
    assign in4065_2 = {s1974[3],s2065[0],s2066[1],s2049[2]};
    CLA_4 KS_4065(s4065, c4065, in4065_1, in4065_2);
    wire[3:0] s4066, in4066_1, in4066_2;
    wire c4066;
    assign in4066_1 = {s1975[3],s2066[0],c2067,s2050[2]};
    assign in4066_2 = {s1976[3],s2067[0],s2068[1],s2051[2]};
    CLA_4 KS_4066(s4066, c4066, in4066_1, in4066_2);
    wire[3:0] s4067, in4067_1, in4067_2;
    wire c4067;
    assign in4067_1 = {s1977[3],s2068[0],c2069,s2052[2]};
    assign in4067_2 = {s1978[3],s2069[0],s2070[1],s2053[2]};
    CLA_4 KS_4067(s4067, c4067, in4067_1, in4067_2);
    wire[3:0] s4068, in4068_1, in4068_2;
    wire c4068;
    assign in4068_1 = {s1979[3],s2070[0],c2071,s2054[2]};
    assign in4068_2 = {s1980[3],s2071[0],s2072[1],s2055[2]};
    CLA_4 KS_4068(s4068, c4068, in4068_1, in4068_2);
    wire[3:0] s4069, in4069_1, in4069_2;
    wire c4069;
    assign in4069_1 = {s1981[3],s2072[0],c2073,s2056[2]};
    assign in4069_2 = {s1982[3],s2073[0],s2074[1],s2057[2]};
    CLA_4 KS_4069(s4069, c4069, in4069_1, in4069_2);
    wire[3:0] s4070, in4070_1, in4070_2;
    wire c4070;
    assign in4070_1 = {s1983[3],s2074[0],c2075,s2058[2]};
    assign in4070_2 = {s1984[3],s2075[0],s2076[1],s2059[2]};
    CLA_4 KS_4070(s4070, c4070, in4070_1, in4070_2);
    wire[3:0] s4071, in4071_1, in4071_2;
    wire c4071;
    assign in4071_1 = {s1985[3],s2076[0],c2077,s2060[2]};
    assign in4071_2 = {s1986[3],s2077[0],s2078[1],s2061[2]};
    CLA_4 KS_4071(s4071, c4071, in4071_1, in4071_2);
    wire[3:0] s4072, in4072_1, in4072_2;
    wire c4072;
    assign in4072_1 = {s1987[3],s2078[0],c2079,s2062[2]};
    assign in4072_2 = {s1988[3],s2079[0],s2080[1],s2063[2]};
    CLA_4 KS_4072(s4072, c4072, in4072_1, in4072_2);
    wire[3:0] s4073, in4073_1, in4073_2;
    wire c4073;
    assign in4073_1 = {s1989[3],s2080[0],c2081,s2064[2]};
    assign in4073_2 = {s1990[3],s2081[0],s2082[1],s2065[2]};
    CLA_4 KS_4073(s4073, c4073, in4073_1, in4073_2);
    wire[3:0] s4074, in4074_1, in4074_2;
    wire c4074;
    assign in4074_1 = {s1991[3],s2082[0],c2083,c2066};
    assign in4074_2 = {s1992[3],s2083[0],s2084[1],s2068[2]};
    CLA_4 KS_4074(s4074, c4074, in4074_1, in4074_2);
    wire[3:0] s4075, in4075_1, in4075_2;
    wire c4075;
    assign in4075_1 = {s1993[3],s2084[0],c2085,c2070};
    assign in4075_2 = {s1994[3],s2085[0],s2086[1],s2072[2]};
    CLA_4 KS_4075(s4075, c4075, in4075_1, in4075_2);
    wire[3:0] s4076, in4076_1, in4076_2;
    wire c4076;
    assign in4076_1 = {s1995[3],s2086[0],c2087,c2074};
    assign in4076_2 = {s1996[3],s2087[0],s2088[1],s2076[2]};
    CLA_4 KS_4076(s4076, c4076, in4076_1, in4076_2);
    wire[3:0] s4077, in4077_1, in4077_2;
    wire c4077;
    assign in4077_1 = {s1997[3],s2088[0],c2089,c2078};
    assign in4077_2 = {s1998[3],s2089[0],s2090[1],s2080[2]};
    CLA_4 KS_4077(s4077, c4077, in4077_1, in4077_2);
    wire[3:0] s4078, in4078_1, in4078_2;
    wire c4078;
    assign in4078_1 = {s1999[3],s2090[0],c2091,c2082};
    assign in4078_2 = {s2000[3],s2091[0],s2092[1],s2084[2]};
    CLA_4 KS_4078(s4078, c4078, in4078_1, in4078_2);
    wire[1:0] s4079, in4079_1, in4079_2;
    wire c4079;
    assign in4079_1 = {c2004,s2092[0]};
    assign in4079_2 = {s2008[3],s2093[0]};
    CLA_2 KS_4079(s4079, c4079, in4079_1, in4079_2);
    wire[0:0] s4080, in4080_1, in4080_2;
    wire c4080;
    assign in4080_1 = {c2012};
    assign in4080_2 = {s2016[3]};
    Half_Adder KS_4080(s4080, c4080, in4080_1, in4080_2);
    wire[2:0] s4081, in4081_1, in4081_2;
    wire c4081;
    assign in4081_1 = {c2020,s2094[0],c2093};
    assign in4081_2 = {s2024[3],s2095[0],s2094[1]};
    CLA_3 KS_4081(s4081, c4081, in4081_1, in4081_2);
    wire[0:0] s4082, in4082_1, in4082_2;
    wire c4082;
    assign in4082_1 = {c2028};
    assign in4082_2 = {s2032[3]};
    Half_Adder KS_4082(s4082, c4082, in4082_1, in4082_2);
    wire[1:0] s4083, in4083_1, in4083_2;
    wire c4083;
    assign in4083_1 = {c4025,s2096[0]};
    assign in4083_2 = {c4026,s2097[0]};
    CLA_2 KS_4083(s4083, c4083, in4083_1, in4083_2);
    wire[0:0] s4084, in4084_1, in4084_2;
    wire c4084;
    assign in4084_1 = {c4027};
    assign in4084_2 = {c4028};
    Half_Adder KS_4084(s4084, c4084, in4084_1, in4084_2);
    wire[3:0] s4085, in4085_1, in4085_2;
    wire c4085;
    assign in4085_1 = {c4029,s2098[0],c2095,c2086};
    assign in4085_2 = {c4030,s2099[0],s2096[1],s2088[2]};
    CLA_4 KS_4085(s4085, c4085, in4085_1, in4085_2);
    wire[0:0] s4086, in4086_1, in4086_2;
    wire c4086;
    assign in4086_1 = {c4031};
    assign in4086_2 = {c4032};
    Half_Adder KS_4086(s4086, c4086, in4086_1, in4086_2);
    wire[1:0] s4087, in4087_1, in4087_2;
    wire c4087;
    assign in4087_1 = {c4033,s2100[0]};
    assign in4087_2 = {c4034,s4061[1]};
    CLA_2 KS_4087(s4087, c4087, in4087_1, in4087_2);
    wire[0:0] s4088, in4088_1, in4088_2;
    wire c4088;
    assign in4088_1 = {c4035};
    assign in4088_2 = {c4036};
    Half_Adder KS_4088(s4088, c4088, in4088_1, in4088_2);
    wire[2:0] s4089, in4089_1, in4089_2;
    wire c4089;
    assign in4089_1 = {c4037,s4062[1],c2097};
    assign in4089_2 = {c4038,s4063[1],s2098[1]};
    CLA_3 KS_4089(s4089, c4089, in4089_1, in4089_2);
    wire[0:0] s4090, in4090_1, in4090_2;
    wire c4090;
    assign in4090_1 = {c4039};
    assign in4090_2 = {c4040};
    Half_Adder KS_4090(s4090, c4090, in4090_1, in4090_2);
    wire[1:0] s4091, in4091_1, in4091_2;
    wire c4091;
    assign in4091_1 = {c4041,s4064[1]};
    assign in4091_2 = {c4042,s4065[1]};
    CLA_2 KS_4091(s4091, c4091, in4091_1, in4091_2);
    wire[0:0] s4092, in4092_1, in4092_2;
    wire c4092;
    assign in4092_1 = {c4045};
    assign in4092_2 = {c4053};
    Half_Adder KS_4092(s4092, c4092, in4092_1, in4092_2);
    wire[3:0] s4093, in4093_1, in4093_2;
    wire c4093;
    assign in4093_1 = {s4061[0],s4066[1],c2099,c2090};
    assign in4093_2 = {s4062[0],s4067[1],s2100[1],s2092[2]};
    CLA_4 KS_4093(s4093, c4093, in4093_1, in4093_2);
    wire[0:0] s4094, in4094_1, in4094_2;
    wire c4094;
    assign in4094_1 = {s4063[0]};
    assign in4094_2 = {s4064[0]};
    Half_Adder KS_4094(s4094, c4094, in4094_1, in4094_2);
    wire[1:0] s4095, in4095_1, in4095_2;
    wire c4095;
    assign in4095_1 = {s4065[0],s4068[1]};
    assign in4095_2 = {s4066[0],s4069[1]};
    CLA_2 KS_4095(s4095, c4095, in4095_1, in4095_2);
    wire[0:0] s4096, in4096_1, in4096_2;
    wire c4096;
    assign in4096_1 = {s4068[0]};
    assign in4096_2 = {s4069[0]};
    Full_Adder KS_4096(s4096, c4096, in4096_1, in4096_2, s4067[0]);
    wire[3:0] s4097, in4097_1, in4097_2;
    wire c4097;
    assign in4097_1 = {s327[0],s2122[0],s2123[1],s2106[2]};
    assign in4097_2 = {s328[0],s2123[0],s2124[1],s2107[2]};
    CLA_4 KS_4097(s4097, c4097, in4097_1, in4097_2);
    wire[3:0] s4098, in4098_1, in4098_2;
    wire c4098;
    assign in4098_1 = {s329[0],s2124[0],s2125[1],s2108[2]};
    assign in4098_2 = {s330[0],s2125[0],s2126[1],s2109[2]};
    CLA_4 KS_4098(s4098, c4098, in4098_1, in4098_2);
    wire[3:0] s4099, in4099_1, in4099_2;
    wire c4099;
    assign in4099_1 = {s2035[3],s2126[0],s2127[1],s2110[2]};
    assign in4099_2 = {s2036[3],s2127[0],s2128[1],s2111[2]};
    CLA_4 KS_4099(s4099, c4099, in4099_1, in4099_2);
    wire[3:0] s4100, in4100_1, in4100_2;
    wire c4100;
    assign in4100_1 = {s2037[3],s2128[0],s2129[1],s2112[2]};
    assign in4100_2 = {s2038[3],s2129[0],s2130[1],s2113[2]};
    CLA_4 KS_4100(s4100, c4100, in4100_1, in4100_2);
    wire[3:0] s4101, in4101_1, in4101_2;
    wire c4101;
    assign in4101_1 = {s2039[3],s2130[0],s2131[1],s2114[2]};
    assign in4101_2 = {s2040[3],s2131[0],s2132[1],s2115[2]};
    CLA_4 KS_4101(s4101, c4101, in4101_1, in4101_2);
    wire[3:0] s4102, in4102_1, in4102_2;
    wire c4102;
    assign in4102_1 = {s2041[3],s2132[0],c2133,s2116[2]};
    assign in4102_2 = {s2042[3],s2133[0],s2134[1],s2117[2]};
    CLA_4 KS_4102(s4102, c4102, in4102_1, in4102_2);
    wire[3:0] s4103, in4103_1, in4103_2;
    wire c4103;
    assign in4103_1 = {s2043[3],s2134[0],c2135,s2118[2]};
    assign in4103_2 = {s2044[3],s2135[0],s2136[1],s2119[2]};
    CLA_4 KS_4103(s4103, c4103, in4103_1, in4103_2);
    wire[3:0] s4104, in4104_1, in4104_2;
    wire c4104;
    assign in4104_1 = {s2045[3],s2136[0],c2137,s2120[2]};
    assign in4104_2 = {s2046[3],s2137[0],s2138[1],s2121[2]};
    CLA_4 KS_4104(s4104, c4104, in4104_1, in4104_2);
    wire[3:0] s4105, in4105_1, in4105_2;
    wire c4105;
    assign in4105_1 = {s2047[3],s2138[0],c2139,s2122[2]};
    assign in4105_2 = {s2048[3],s2139[0],s2140[1],s2123[2]};
    CLA_4 KS_4105(s4105, c4105, in4105_1, in4105_2);
    wire[3:0] s4106, in4106_1, in4106_2;
    wire c4106;
    assign in4106_1 = {s2049[3],s2140[0],c2141,s2124[2]};
    assign in4106_2 = {s2050[3],s2141[0],s2142[1],s2125[2]};
    CLA_4 KS_4106(s4106, c4106, in4106_1, in4106_2);
    wire[3:0] s4107, in4107_1, in4107_2;
    wire c4107;
    assign in4107_1 = {s2051[3],s2142[0],c2143,s2126[2]};
    assign in4107_2 = {s2052[3],s2143[0],s2144[1],s2127[2]};
    CLA_4 KS_4107(s4107, c4107, in4107_1, in4107_2);
    wire[3:0] s4108, in4108_1, in4108_2;
    wire c4108;
    assign in4108_1 = {s2053[3],s2144[0],c2145,s2128[2]};
    assign in4108_2 = {s2054[3],s2145[0],s2146[1],s2129[2]};
    CLA_4 KS_4108(s4108, c4108, in4108_1, in4108_2);
    wire[3:0] s4109, in4109_1, in4109_2;
    wire c4109;
    assign in4109_1 = {s2055[3],s2146[0],c2147,s2130[2]};
    assign in4109_2 = {s2056[3],s2147[0],s2148[1],s2131[2]};
    CLA_4 KS_4109(s4109, c4109, in4109_1, in4109_2);
    wire[3:0] s4110, in4110_1, in4110_2;
    wire c4110;
    assign in4110_1 = {s2057[3],s2148[0],c2149,c2132};
    assign in4110_2 = {s2058[3],s2149[0],s2150[1],s2134[2]};
    CLA_4 KS_4110(s4110, c4110, in4110_1, in4110_2);
    wire[3:0] s4111, in4111_1, in4111_2;
    wire c4111;
    assign in4111_1 = {s2059[3],s2150[0],c2151,c2136};
    assign in4111_2 = {s2060[3],s2151[0],s2152[1],s2138[2]};
    CLA_4 KS_4111(s4111, c4111, in4111_1, in4111_2);
    wire[3:0] s4112, in4112_1, in4112_2;
    wire c4112;
    assign in4112_1 = {s2061[3],s2152[0],c2153,c2140};
    assign in4112_2 = {s2062[3],s2153[0],s2154[1],s2142[2]};
    CLA_4 KS_4112(s4112, c4112, in4112_1, in4112_2);
    wire[3:0] s4113, in4113_1, in4113_2;
    wire c4113;
    assign in4113_1 = {s2063[3],s2154[0],c2155,c2144};
    assign in4113_2 = {s2064[3],s2155[0],s2156[1],s2146[2]};
    CLA_4 KS_4113(s4113, c4113, in4113_1, in4113_2);
    wire[3:0] s4114, in4114_1, in4114_2;
    wire c4114;
    assign in4114_1 = {s2065[3],s2156[0],c2157,c2148};
    assign in4114_2 = {s2068[3],s2157[0],s2158[1],s2150[2]};
    CLA_4 KS_4114(s4114, c4114, in4114_1, in4114_2);
    wire[1:0] s4115, in4115_1, in4115_2;
    wire c4115;
    assign in4115_1 = {c2072,s2158[0]};
    assign in4115_2 = {s2076[3],s2159[0]};
    CLA_2 KS_4115(s4115, c4115, in4115_1, in4115_2);
    wire[0:0] s4116, in4116_1, in4116_2;
    wire c4116;
    assign in4116_1 = {c2080};
    assign in4116_2 = {s2084[3]};
    Half_Adder KS_4116(s4116, c4116, in4116_1, in4116_2);
    wire[2:0] s4117, in4117_1, in4117_2;
    wire c4117;
    assign in4117_1 = {c2088,s2160[0],c2159};
    assign in4117_2 = {s2092[3],s2161[0],s2160[1]};
    CLA_3 KS_4117(s4117, c4117, in4117_1, in4117_2);
    wire[0:0] s4118, in4118_1, in4118_2;
    wire c4118;
    assign in4118_1 = {c2096};
    assign in4118_2 = {s2100[3]};
    Half_Adder KS_4118(s4118, c4118, in4118_1, in4118_2);
    wire[1:0] s4119, in4119_1, in4119_2;
    wire c4119;
    assign in4119_1 = {c4061,s2162[0]};
    assign in4119_2 = {c4062,s2163[0]};
    CLA_2 KS_4119(s4119, c4119, in4119_1, in4119_2);
    wire[0:0] s4120, in4120_1, in4120_2;
    wire c4120;
    assign in4120_1 = {c4063};
    assign in4120_2 = {c4064};
    Half_Adder KS_4120(s4120, c4120, in4120_1, in4120_2);
    wire[3:0] s4121, in4121_1, in4121_2;
    wire c4121;
    assign in4121_1 = {c4065,s2164[0],c2161,c2152};
    assign in4121_2 = {c4066,s2165[0],s2162[1],s2154[2]};
    CLA_4 KS_4121(s4121, c4121, in4121_1, in4121_2);
    wire[0:0] s4122, in4122_1, in4122_2;
    wire c4122;
    assign in4122_1 = {c4067};
    assign in4122_2 = {c4068};
    Half_Adder KS_4122(s4122, c4122, in4122_1, in4122_2);
    wire[1:0] s4123, in4123_1, in4123_2;
    wire c4123;
    assign in4123_1 = {c4069,s2166[0]};
    assign in4123_2 = {c4070,s4097[1]};
    CLA_2 KS_4123(s4123, c4123, in4123_1, in4123_2);
    wire[0:0] s4124, in4124_1, in4124_2;
    wire c4124;
    assign in4124_1 = {c4071};
    assign in4124_2 = {c4072};
    Half_Adder KS_4124(s4124, c4124, in4124_1, in4124_2);
    wire[2:0] s4125, in4125_1, in4125_2;
    wire c4125;
    assign in4125_1 = {c4073,s4098[1],c2163};
    assign in4125_2 = {c4074,s4099[1],s2164[1]};
    CLA_3 KS_4125(s4125, c4125, in4125_1, in4125_2);
    wire[0:0] s4126, in4126_1, in4126_2;
    wire c4126;
    assign in4126_1 = {c4075};
    assign in4126_2 = {c4076};
    Half_Adder KS_4126(s4126, c4126, in4126_1, in4126_2);
    wire[1:0] s4127, in4127_1, in4127_2;
    wire c4127;
    assign in4127_1 = {c4077,s4100[1]};
    assign in4127_2 = {c4078,s4101[1]};
    CLA_2 KS_4127(s4127, c4127, in4127_1, in4127_2);
    wire[0:0] s4128, in4128_1, in4128_2;
    wire c4128;
    assign in4128_1 = {c4085};
    assign in4128_2 = {c4093};
    Half_Adder KS_4128(s4128, c4128, in4128_1, in4128_2);
    wire[3:0] s4129, in4129_1, in4129_2;
    wire c4129;
    assign in4129_1 = {s4097[0],s4102[1],c2165,c2156};
    assign in4129_2 = {s4098[0],s4103[1],s2166[1],s2158[2]};
    CLA_4 KS_4129(s4129, c4129, in4129_1, in4129_2);
    wire[0:0] s4130, in4130_1, in4130_2;
    wire c4130;
    assign in4130_1 = {s4099[0]};
    assign in4130_2 = {s4100[0]};
    Half_Adder KS_4130(s4130, c4130, in4130_1, in4130_2);
    wire[1:0] s4131, in4131_1, in4131_2;
    wire c4131;
    assign in4131_1 = {s4101[0],s4104[1]};
    assign in4131_2 = {s4102[0],s4105[1]};
    CLA_2 KS_4131(s4131, c4131, in4131_1, in4131_2);
    wire[0:0] s4132, in4132_1, in4132_2;
    wire c4132;
    assign in4132_1 = {s4104[0]};
    assign in4132_2 = {s4105[0]};
    Full_Adder KS_4132(s4132, c4132, in4132_1, in4132_2, s4103[0]);
    wire[3:0] s4133, in4133_1, in4133_2;
    wire c4133;
    assign in4133_1 = {s415[0],s2188[0],s2188[1],s2170[2]};
    assign in4133_2 = {s416[0],s2189[0],s2189[1],s2171[2]};
    CLA_4 KS_4133(s4133, c4133, in4133_1, in4133_2);
    wire[3:0] s4134, in4134_1, in4134_2;
    wire c4134;
    assign in4134_1 = {s417[0],s2190[0],s2190[1],s2172[2]};
    assign in4134_2 = {s418[0],s2191[0],s2191[1],s2173[2]};
    CLA_4 KS_4134(s4134, c4134, in4134_1, in4134_2);
    wire[3:0] s4135, in4135_1, in4135_2;
    wire c4135;
    assign in4135_1 = {s2101[3],s2192[0],s2192[1],s2174[2]};
    assign in4135_2 = {s2102[3],s2193[0],s2193[1],s2175[2]};
    CLA_4 KS_4135(s4135, c4135, in4135_1, in4135_2);
    wire[3:0] s4136, in4136_1, in4136_2;
    wire c4136;
    assign in4136_1 = {s2103[3],s2194[0],s2194[1],s2176[2]};
    assign in4136_2 = {s2104[3],s2195[0],s2195[1],s2177[2]};
    CLA_4 KS_4136(s4136, c4136, in4136_1, in4136_2);
    wire[3:0] s4137, in4137_1, in4137_2;
    wire c4137;
    assign in4137_1 = {s2105[3],s2196[0],s2196[1],s2178[2]};
    assign in4137_2 = {s2106[3],s2197[0],s2197[1],s2179[2]};
    CLA_4 KS_4137(s4137, c4137, in4137_1, in4137_2);
    wire[3:0] s4138, in4138_1, in4138_2;
    wire c4138;
    assign in4138_1 = {s2107[3],s2198[0],c2198,s2180[2]};
    assign in4138_2 = {s2108[3],s2199[0],s2199[1],s2181[2]};
    CLA_4 KS_4138(s4138, c4138, in4138_1, in4138_2);
    wire[3:0] s4139, in4139_1, in4139_2;
    wire c4139;
    assign in4139_1 = {s2109[3],s2200[0],c2200,s2182[2]};
    assign in4139_2 = {s2110[3],s2201[0],s2201[1],s2183[2]};
    CLA_4 KS_4139(s4139, c4139, in4139_1, in4139_2);
    wire[3:0] s4140, in4140_1, in4140_2;
    wire c4140;
    assign in4140_1 = {s2111[3],s2202[0],c2202,s2184[2]};
    assign in4140_2 = {s2112[3],s2203[0],s2203[1],s2185[2]};
    CLA_4 KS_4140(s4140, c4140, in4140_1, in4140_2);
    wire[3:0] s4141, in4141_1, in4141_2;
    wire c4141;
    assign in4141_1 = {s2113[3],s2204[0],c2204,s2186[2]};
    assign in4141_2 = {s2114[3],s2205[0],s2205[1],s2187[2]};
    CLA_4 KS_4141(s4141, c4141, in4141_1, in4141_2);
    wire[3:0] s4142, in4142_1, in4142_2;
    wire c4142;
    assign in4142_1 = {s2115[3],s2206[0],c2206,s2188[2]};
    assign in4142_2 = {s2116[3],s2207[0],s2207[1],s2189[2]};
    CLA_4 KS_4142(s4142, c4142, in4142_1, in4142_2);
    wire[3:0] s4143, in4143_1, in4143_2;
    wire c4143;
    assign in4143_1 = {s2117[3],s2208[0],c2208,s2190[2]};
    assign in4143_2 = {s2118[3],s2209[0],s2209[1],s2191[2]};
    CLA_4 KS_4143(s4143, c4143, in4143_1, in4143_2);
    wire[3:0] s4144, in4144_1, in4144_2;
    wire c4144;
    assign in4144_1 = {s2119[3],s2210[0],c2210,s2192[2]};
    assign in4144_2 = {s2120[3],s2211[0],s2211[1],s2193[2]};
    CLA_4 KS_4144(s4144, c4144, in4144_1, in4144_2);
    wire[3:0] s4145, in4145_1, in4145_2;
    wire c4145;
    assign in4145_1 = {s2121[3],s2212[0],c2212,s2194[2]};
    assign in4145_2 = {s2122[3],s2213[0],s2213[1],s2195[2]};
    CLA_4 KS_4145(s4145, c4145, in4145_1, in4145_2);
    wire[3:0] s4146, in4146_1, in4146_2;
    wire c4146;
    assign in4146_1 = {s2123[3],s2214[0],c2214,s2196[2]};
    assign in4146_2 = {s2124[3],s2215[0],s2215[1],s2197[2]};
    CLA_4 KS_4146(s4146, c4146, in4146_1, in4146_2);
    wire[3:0] s4147, in4147_1, in4147_2;
    wire c4147;
    assign in4147_1 = {s2125[3],s2216[0],c2216,c2199};
    assign in4147_2 = {s2126[3],s2217[0],s2217[1],s2201[2]};
    CLA_4 KS_4147(s4147, c4147, in4147_1, in4147_2);
    wire[3:0] s4148, in4148_1, in4148_2;
    wire c4148;
    assign in4148_1 = {s2127[3],s2218[0],c2218,c2203};
    assign in4148_2 = {s2128[3],s2219[0],s2219[1],s2205[2]};
    CLA_4 KS_4148(s4148, c4148, in4148_1, in4148_2);
    wire[3:0] s4149, in4149_1, in4149_2;
    wire c4149;
    assign in4149_1 = {s2129[3],s2220[0],c2220,c2207};
    assign in4149_2 = {s2130[3],s2221[0],s2221[1],s2209[2]};
    CLA_4 KS_4149(s4149, c4149, in4149_1, in4149_2);
    wire[3:0] s4150, in4150_1, in4150_2;
    wire c4150;
    assign in4150_1 = {s2131[3],s2222[0],c2222,c2211};
    assign in4150_2 = {s2134[3],s2223[0],s2223[1],s2213[2]};
    CLA_4 KS_4150(s4150, c4150, in4150_1, in4150_2);
    wire[3:0] s4151, in4151_1, in4151_2;
    wire c4151;
    assign in4151_1 = {c2138,s2224[0],c2224,c2215};
    assign in4151_2 = {s2142[3],s2225[0],s2225[1],s2217[2]};
    CLA_4 KS_4151(s4151, c4151, in4151_1, in4151_2);
    wire[0:0] s4152, in4152_1, in4152_2;
    wire c4152;
    assign in4152_1 = {c2146};
    assign in4152_2 = {s2150[3]};
    Half_Adder KS_4152(s4152, c4152, in4152_1, in4152_2);
    wire[1:0] s4153, in4153_1, in4153_2;
    wire c4153;
    assign in4153_1 = {c2154,s2226[0]};
    assign in4153_2 = {s2158[3],s2227[0]};
    CLA_2 KS_4153(s4153, c4153, in4153_1, in4153_2);
    wire[0:0] s4154, in4154_1, in4154_2;
    wire c4154;
    assign in4154_1 = {c2162};
    assign in4154_2 = {s2166[3]};
    Half_Adder KS_4154(s4154, c4154, in4154_1, in4154_2);
    wire[2:0] s4155, in4155_1, in4155_2;
    wire c4155;
    assign in4155_1 = {c4097,s2228[0],c2226};
    assign in4155_2 = {c4098,s2229[0],s2227[1]};
    CLA_3 KS_4155(s4155, c4155, in4155_1, in4155_2);
    wire[0:0] s4156, in4156_1, in4156_2;
    wire c4156;
    assign in4156_1 = {c4099};
    assign in4156_2 = {c4100};
    Half_Adder KS_4156(s4156, c4156, in4156_1, in4156_2);
    wire[1:0] s4157, in4157_1, in4157_2;
    wire c4157;
    assign in4157_1 = {c4101,s2230[0]};
    assign in4157_2 = {c4102,s2231[0]};
    CLA_2 KS_4157(s4157, c4157, in4157_1, in4157_2);
    wire[0:0] s4158, in4158_1, in4158_2;
    wire c4158;
    assign in4158_1 = {c4103};
    assign in4158_2 = {c4104};
    Half_Adder KS_4158(s4158, c4158, in4158_1, in4158_2);
    wire[3:0] s4159, in4159_1, in4159_2;
    wire c4159;
    assign in4159_1 = {c4105,s2232[0],c2228,c2219};
    assign in4159_2 = {c4106,s4133[1],s2229[1],s2221[2]};
    CLA_4 KS_4159(s4159, c4159, in4159_1, in4159_2);
    wire[0:0] s4160, in4160_1, in4160_2;
    wire c4160;
    assign in4160_1 = {c4107};
    assign in4160_2 = {c4108};
    Half_Adder KS_4160(s4160, c4160, in4160_1, in4160_2);
    wire[1:0] s4161, in4161_1, in4161_2;
    wire c4161;
    assign in4161_1 = {c4109,s4134[1]};
    assign in4161_2 = {c4110,s4135[1]};
    CLA_2 KS_4161(s4161, c4161, in4161_1, in4161_2);
    wire[0:0] s4162, in4162_1, in4162_2;
    wire c4162;
    assign in4162_1 = {c4111};
    assign in4162_2 = {c4112};
    Half_Adder KS_4162(s4162, c4162, in4162_1, in4162_2);
    wire[2:0] s4163, in4163_1, in4163_2;
    wire c4163;
    assign in4163_1 = {c4113,s4136[1],c2230};
    assign in4163_2 = {c4114,s4137[1],s2231[1]};
    CLA_3 KS_4163(s4163, c4163, in4163_1, in4163_2);
    wire[0:0] s4164, in4164_1, in4164_2;
    wire c4164;
    assign in4164_1 = {c4121};
    assign in4164_2 = {c4129};
    Half_Adder KS_4164(s4164, c4164, in4164_1, in4164_2);
    wire[1:0] s4165, in4165_1, in4165_2;
    wire c4165;
    assign in4165_1 = {s4133[0],s4138[1]};
    assign in4165_2 = {s4134[0],s4139[1]};
    CLA_2 KS_4165(s4165, c4165, in4165_1, in4165_2);
    wire[0:0] s4166, in4166_1, in4166_2;
    wire c4166;
    assign in4166_1 = {s4135[0]};
    assign in4166_2 = {s4136[0]};
    Half_Adder KS_4166(s4166, c4166, in4166_1, in4166_2);
    wire[3:0] s4167, in4167_1, in4167_2;
    wire c4167;
    assign in4167_1 = {s4137[0],s4140[1],c2232,c2223};
    assign in4167_2 = {s4138[0],s4141[1],s4133[2],s2225[2]};
    CLA_4 KS_4167(s4167, c4167, in4167_1, in4167_2);
    wire[0:0] s4168, in4168_1, in4168_2;
    wire c4168;
    assign in4168_1 = {s4140[0]};
    assign in4168_2 = {s4141[0]};
    Full_Adder KS_4168(s4168, c4168, in4168_1, in4168_2, s4139[0]);
    wire[3:0] s4169, in4169_1, in4169_2;
    wire c4169;
    assign in4169_1 = {s519[0],s2252[0],s2253[1],s2236[2]};
    assign in4169_2 = {s520[0],s2253[0],s2254[1],s2237[2]};
    CLA_4 KS_4169(s4169, c4169, in4169_1, in4169_2);
    wire[3:0] s4170, in4170_1, in4170_2;
    wire c4170;
    assign in4170_1 = {s521[0],s2254[0],s2255[1],s2238[2]};
    assign in4170_2 = {s522[0],s2255[0],s2256[1],s2239[2]};
    CLA_4 KS_4170(s4170, c4170, in4170_1, in4170_2);
    wire[3:0] s4171, in4171_1, in4171_2;
    wire c4171;
    assign in4171_1 = {s523[0],s2256[0],s2257[1],s2240[2]};
    assign in4171_2 = {s524[0],s2257[0],s2258[1],s2241[2]};
    CLA_4 KS_4171(s4171, c4171, in4171_1, in4171_2);
    wire[3:0] s4172, in4172_1, in4172_2;
    wire c4172;
    assign in4172_1 = {s2167[3],s2258[0],s2259[1],s2242[2]};
    assign in4172_2 = {s2168[3],s2259[0],s2260[1],s2243[2]};
    CLA_4 KS_4172(s4172, c4172, in4172_1, in4172_2);
    wire[3:0] s4173, in4173_1, in4173_2;
    wire c4173;
    assign in4173_1 = {s2169[3],s2260[0],s2261[1],s2244[2]};
    assign in4173_2 = {s2170[3],s2261[0],s2262[1],s2245[2]};
    CLA_4 KS_4173(s4173, c4173, in4173_1, in4173_2);
    wire[3:0] s4174, in4174_1, in4174_2;
    wire c4174;
    assign in4174_1 = {s2171[3],s2262[0],s2263[1],s2246[2]};
    assign in4174_2 = {s2172[3],s2263[0],s2264[1],s2247[2]};
    CLA_4 KS_4174(s4174, c4174, in4174_1, in4174_2);
    wire[3:0] s4175, in4175_1, in4175_2;
    wire c4175;
    assign in4175_1 = {s2173[3],s2264[0],c2265,s2248[2]};
    assign in4175_2 = {s2174[3],s2265[0],s2266[1],s2249[2]};
    CLA_4 KS_4175(s4175, c4175, in4175_1, in4175_2);
    wire[3:0] s4176, in4176_1, in4176_2;
    wire c4176;
    assign in4176_1 = {s2175[3],s2266[0],c2267,s2250[2]};
    assign in4176_2 = {s2176[3],s2267[0],s2268[1],s2251[2]};
    CLA_4 KS_4176(s4176, c4176, in4176_1, in4176_2);
    wire[3:0] s4177, in4177_1, in4177_2;
    wire c4177;
    assign in4177_1 = {s2177[3],s2268[0],c2269,s2252[2]};
    assign in4177_2 = {s2178[3],s2269[0],s2270[1],s2253[2]};
    CLA_4 KS_4177(s4177, c4177, in4177_1, in4177_2);
    wire[3:0] s4178, in4178_1, in4178_2;
    wire c4178;
    assign in4178_1 = {s2179[3],s2270[0],c2271,s2254[2]};
    assign in4178_2 = {s2180[3],s2271[0],s2272[1],s2255[2]};
    CLA_4 KS_4178(s4178, c4178, in4178_1, in4178_2);
    wire[3:0] s4179, in4179_1, in4179_2;
    wire c4179;
    assign in4179_1 = {s2181[3],s2272[0],c2273,s2256[2]};
    assign in4179_2 = {s2182[3],s2273[0],s2274[1],s2257[2]};
    CLA_4 KS_4179(s4179, c4179, in4179_1, in4179_2);
    wire[3:0] s4180, in4180_1, in4180_2;
    wire c4180;
    assign in4180_1 = {s2183[3],s2274[0],c2275,s2258[2]};
    assign in4180_2 = {s2184[3],s2275[0],s2276[1],s2259[2]};
    CLA_4 KS_4180(s4180, c4180, in4180_1, in4180_2);
    wire[3:0] s4181, in4181_1, in4181_2;
    wire c4181;
    assign in4181_1 = {s2185[3],s2276[0],c2277,s2260[2]};
    assign in4181_2 = {s2186[3],s2277[0],s2278[1],s2261[2]};
    CLA_4 KS_4181(s4181, c4181, in4181_1, in4181_2);
    wire[3:0] s4182, in4182_1, in4182_2;
    wire c4182;
    assign in4182_1 = {s2187[3],s2278[0],c2279,s2262[2]};
    assign in4182_2 = {s2188[3],s2279[0],s2280[1],s2263[2]};
    CLA_4 KS_4182(s4182, c4182, in4182_1, in4182_2);
    wire[3:0] s4183, in4183_1, in4183_2;
    wire c4183;
    assign in4183_1 = {s2189[3],s2280[0],c2281,c2264};
    assign in4183_2 = {s2190[3],s2281[0],s2282[1],s2266[2]};
    CLA_4 KS_4183(s4183, c4183, in4183_1, in4183_2);
    wire[3:0] s4184, in4184_1, in4184_2;
    wire c4184;
    assign in4184_1 = {s2191[3],s2282[0],c2283,c2268};
    assign in4184_2 = {s2192[3],s2283[0],s2284[1],s2270[2]};
    CLA_4 KS_4184(s4184, c4184, in4184_1, in4184_2);
    wire[3:0] s4185, in4185_1, in4185_2;
    wire c4185;
    assign in4185_1 = {s2193[3],s2284[0],c2285,c2272};
    assign in4185_2 = {s2194[3],s2285[0],s2286[1],s2274[2]};
    CLA_4 KS_4185(s4185, c4185, in4185_1, in4185_2);
    wire[3:0] s4186, in4186_1, in4186_2;
    wire c4186;
    assign in4186_1 = {s2195[3],s2286[0],c2287,c2276};
    assign in4186_2 = {s2196[3],s2287[0],s2288[1],s2278[2]};
    CLA_4 KS_4186(s4186, c4186, in4186_1, in4186_2);
    wire[1:0] s4187, in4187_1, in4187_2;
    wire c4187;
    assign in4187_1 = {s2197[3],s2288[0]};
    assign in4187_2 = {s2201[3],s2289[0]};
    CLA_2 KS_4187(s4187, c4187, in4187_1, in4187_2);
    wire[0:0] s4188, in4188_1, in4188_2;
    wire c4188;
    assign in4188_1 = {c2205};
    assign in4188_2 = {s2209[3]};
    Half_Adder KS_4188(s4188, c4188, in4188_1, in4188_2);
    wire[3:0] s4189, in4189_1, in4189_2;
    wire c4189;
    assign in4189_1 = {c2213,s2290[0],c2289,c2280};
    assign in4189_2 = {s2217[3],s2291[0],s2290[1],s2282[2]};
    CLA_4 KS_4189(s4189, c4189, in4189_1, in4189_2);
    wire[0:0] s4190, in4190_1, in4190_2;
    wire c4190;
    assign in4190_1 = {c2221};
    assign in4190_2 = {s2225[3]};
    Half_Adder KS_4190(s4190, c4190, in4190_1, in4190_2);
    wire[1:0] s4191, in4191_1, in4191_2;
    wire c4191;
    assign in4191_1 = {c2229,s2292[0]};
    assign in4191_2 = {c4133,s2293[0]};
    CLA_2 KS_4191(s4191, c4191, in4191_1, in4191_2);
    wire[0:0] s4192, in4192_1, in4192_2;
    wire c4192;
    assign in4192_1 = {c4134};
    assign in4192_2 = {c4135};
    Half_Adder KS_4192(s4192, c4192, in4192_1, in4192_2);
    wire[2:0] s4193, in4193_1, in4193_2;
    wire c4193;
    assign in4193_1 = {c4136,s2294[0],c2291};
    assign in4193_2 = {c4137,s2295[0],s2292[1]};
    CLA_3 KS_4193(s4193, c4193, in4193_1, in4193_2);
    wire[0:0] s4194, in4194_1, in4194_2;
    wire c4194;
    assign in4194_1 = {c4138};
    assign in4194_2 = {c4139};
    Half_Adder KS_4194(s4194, c4194, in4194_1, in4194_2);
    wire[1:0] s4195, in4195_1, in4195_2;
    wire c4195;
    assign in4195_1 = {c4140,s2296[0]};
    assign in4195_2 = {c4141,s4169[1]};
    CLA_2 KS_4195(s4195, c4195, in4195_1, in4195_2);
    wire[0:0] s4196, in4196_1, in4196_2;
    wire c4196;
    assign in4196_1 = {c4142};
    assign in4196_2 = {c4143};
    Half_Adder KS_4196(s4196, c4196, in4196_1, in4196_2);
    wire[3:0] s4197, in4197_1, in4197_2;
    wire c4197;
    assign in4197_1 = {c4144,s4170[1],c2293,c2284};
    assign in4197_2 = {c4145,s4171[1],s2294[1],s2286[2]};
    CLA_4 KS_4197(s4197, c4197, in4197_1, in4197_2);
    wire[0:0] s4198, in4198_1, in4198_2;
    wire c4198;
    assign in4198_1 = {c4146};
    assign in4198_2 = {c4147};
    Half_Adder KS_4198(s4198, c4198, in4198_1, in4198_2);
    wire[1:0] s4199, in4199_1, in4199_2;
    wire c4199;
    assign in4199_1 = {c4148,s4172[1]};
    assign in4199_2 = {c4149,s4173[1]};
    CLA_2 KS_4199(s4199, c4199, in4199_1, in4199_2);
    wire[0:0] s4200, in4200_1, in4200_2;
    wire c4200;
    assign in4200_1 = {c4150};
    assign in4200_2 = {c4151};
    Half_Adder KS_4200(s4200, c4200, in4200_1, in4200_2);
    wire[2:0] s4201, in4201_1, in4201_2;
    wire c4201;
    assign in4201_1 = {c4159,s4174[1],c2295};
    assign in4201_2 = {c4167,s4175[1],s2296[1]};
    CLA_3 KS_4201(s4201, c4201, in4201_1, in4201_2);
    wire[0:0] s4202, in4202_1, in4202_2;
    wire c4202;
    assign in4202_1 = {s4169[0]};
    assign in4202_2 = {s4170[0]};
    Half_Adder KS_4202(s4202, c4202, in4202_1, in4202_2);
    wire[1:0] s4203, in4203_1, in4203_2;
    wire c4203;
    assign in4203_1 = {s4171[0],s4176[1]};
    assign in4203_2 = {s4172[0],s4177[1]};
    CLA_2 KS_4203(s4203, c4203, in4203_1, in4203_2);
    wire[0:0] s4204, in4204_1, in4204_2;
    wire c4204;
    assign in4204_1 = {s4173[0]};
    assign in4204_2 = {s4174[0]};
    Half_Adder KS_4204(s4204, c4204, in4204_1, in4204_2);
    wire[3:0] s4205, in4205_1, in4205_2;
    wire c4205;
    assign in4205_1 = {s4175[0],s4178[1],s4169[2],c2288};
    assign in4205_2 = {s4176[0],s4179[1],s4170[2],s2290[2]};
    CLA_4 KS_4205(s4205, c4205, in4205_1, in4205_2);
    wire[0:0] s4206, in4206_1, in4206_2;
    wire c4206;
    assign in4206_1 = {s4178[0]};
    assign in4206_2 = {s4179[0]};
    Full_Adder KS_4206(s4206, c4206, in4206_1, in4206_2, s4177[0]);
    wire[3:0] s4207, in4207_1, in4207_2;
    wire c4207;
    assign in4207_1 = {s626[0],s2316[0],s2317[1],s2301[2]};
    assign in4207_2 = {s627[0],s2317[0],s2318[1],s2302[2]};
    CLA_4 KS_4207(s4207, c4207, in4207_1, in4207_2);
    wire[3:0] s4208, in4208_1, in4208_2;
    wire c4208;
    assign in4208_1 = {s628[0],s2318[0],s2319[1],s2303[2]};
    assign in4208_2 = {s629[0],s2319[0],s2320[1],s2304[2]};
    CLA_4 KS_4208(s4208, c4208, in4208_1, in4208_2);
    wire[3:0] s4209, in4209_1, in4209_2;
    wire c4209;
    assign in4209_1 = {s630[0],s2320[0],s2321[1],s2305[2]};
    assign in4209_2 = {s631[0],s2321[0],s2322[1],s2306[2]};
    CLA_4 KS_4209(s4209, c4209, in4209_1, in4209_2);
    wire[3:0] s4210, in4210_1, in4210_2;
    wire c4210;
    assign in4210_1 = {s2233[3],s2322[0],s2323[1],s2307[2]};
    assign in4210_2 = {s2234[3],s2323[0],s2324[1],s2308[2]};
    CLA_4 KS_4210(s4210, c4210, in4210_1, in4210_2);
    wire[3:0] s4211, in4211_1, in4211_2;
    wire c4211;
    assign in4211_1 = {s2235[3],s2324[0],s2325[1],s2309[2]};
    assign in4211_2 = {s2236[3],s2325[0],s2326[1],s2310[2]};
    CLA_4 KS_4211(s4211, c4211, in4211_1, in4211_2);
    wire[3:0] s4212, in4212_1, in4212_2;
    wire c4212;
    assign in4212_1 = {s2237[3],s2326[0],s2327[1],s2311[2]};
    assign in4212_2 = {s2238[3],s2327[0],s2328[1],s2312[2]};
    CLA_4 KS_4212(s4212, c4212, in4212_1, in4212_2);
    wire[3:0] s4213, in4213_1, in4213_2;
    wire c4213;
    assign in4213_1 = {s2239[3],s2328[0],c2329,s2313[2]};
    assign in4213_2 = {s2240[3],s2329[0],s2330[1],s2314[2]};
    CLA_4 KS_4213(s4213, c4213, in4213_1, in4213_2);
    wire[3:0] s4214, in4214_1, in4214_2;
    wire c4214;
    assign in4214_1 = {s2241[3],s2330[0],c2331,s2315[2]};
    assign in4214_2 = {s2242[3],s2331[0],s2332[1],s2316[2]};
    CLA_4 KS_4214(s4214, c4214, in4214_1, in4214_2);
    wire[3:0] s4215, in4215_1, in4215_2;
    wire c4215;
    assign in4215_1 = {s2243[3],s2332[0],c2333,s2317[2]};
    assign in4215_2 = {s2244[3],s2333[0],s2334[1],s2318[2]};
    CLA_4 KS_4215(s4215, c4215, in4215_1, in4215_2);
    wire[3:0] s4216, in4216_1, in4216_2;
    wire c4216;
    assign in4216_1 = {s2245[3],s2334[0],c2335,s2319[2]};
    assign in4216_2 = {s2246[3],s2335[0],s2336[1],s2320[2]};
    CLA_4 KS_4216(s4216, c4216, in4216_1, in4216_2);
    wire[3:0] s4217, in4217_1, in4217_2;
    wire c4217;
    assign in4217_1 = {s2247[3],s2336[0],c2337,s2321[2]};
    assign in4217_2 = {s2248[3],s2337[0],s2338[1],s2322[2]};
    CLA_4 KS_4217(s4217, c4217, in4217_1, in4217_2);
    wire[3:0] s4218, in4218_1, in4218_2;
    wire c4218;
    assign in4218_1 = {s2249[3],s2338[0],c2339,s2323[2]};
    assign in4218_2 = {s2250[3],s2339[0],s2340[1],s2324[2]};
    CLA_4 KS_4218(s4218, c4218, in4218_1, in4218_2);
    wire[3:0] s4219, in4219_1, in4219_2;
    wire c4219;
    assign in4219_1 = {s2251[3],s2340[0],c2341,s2325[2]};
    assign in4219_2 = {s2252[3],s2341[0],s2342[1],s2326[2]};
    CLA_4 KS_4219(s4219, c4219, in4219_1, in4219_2);
    wire[3:0] s4220, in4220_1, in4220_2;
    wire c4220;
    assign in4220_1 = {s2253[3],s2342[0],c2343,s2327[2]};
    assign in4220_2 = {s2254[3],s2343[0],s2344[1],s2328[2]};
    CLA_4 KS_4220(s4220, c4220, in4220_1, in4220_2);
    wire[3:0] s4221, in4221_1, in4221_2;
    wire c4221;
    assign in4221_1 = {s2255[3],s2344[0],c2345,c2330};
    assign in4221_2 = {s2256[3],s2345[0],s2346[1],s2332[2]};
    CLA_4 KS_4221(s4221, c4221, in4221_1, in4221_2);
    wire[3:0] s4222, in4222_1, in4222_2;
    wire c4222;
    assign in4222_1 = {s2257[3],s2346[0],c2347,c2334};
    assign in4222_2 = {s2258[3],s2347[0],s2348[1],s2336[2]};
    CLA_4 KS_4222(s4222, c4222, in4222_1, in4222_2);
    wire[3:0] s4223, in4223_1, in4223_2;
    wire c4223;
    assign in4223_1 = {s2259[3],s2348[0],c2349,c2338};
    assign in4223_2 = {s2260[3],s2349[0],s2350[1],s2340[2]};
    CLA_4 KS_4223(s4223, c4223, in4223_1, in4223_2);
    wire[3:0] s4224, in4224_1, in4224_2;
    wire c4224;
    assign in4224_1 = {s2261[3],s2350[0],c2351,c2342};
    assign in4224_2 = {s2262[3],s2351[0],s2352[1],s2344[2]};
    CLA_4 KS_4224(s4224, c4224, in4224_1, in4224_2);
    wire[1:0] s4225, in4225_1, in4225_2;
    wire c4225;
    assign in4225_1 = {s2263[3],s2352[0]};
    assign in4225_2 = {s2266[3],s2353[0]};
    CLA_2 KS_4225(s4225, c4225, in4225_1, in4225_2);
    wire[0:0] s4226, in4226_1, in4226_2;
    wire c4226;
    assign in4226_1 = {c2270};
    assign in4226_2 = {s2274[3]};
    Half_Adder KS_4226(s4226, c4226, in4226_1, in4226_2);
    wire[2:0] s4227, in4227_1, in4227_2;
    wire c4227;
    assign in4227_1 = {c2278,s2354[0],c2353};
    assign in4227_2 = {s2282[3],s2355[0],s2354[1]};
    CLA_3 KS_4227(s4227, c4227, in4227_1, in4227_2);
    wire[0:0] s4228, in4228_1, in4228_2;
    wire c4228;
    assign in4228_1 = {c2286};
    assign in4228_2 = {s2290[3]};
    Half_Adder KS_4228(s4228, c4228, in4228_1, in4228_2);
    wire[1:0] s4229, in4229_1, in4229_2;
    wire c4229;
    assign in4229_1 = {c2294,s2356[0]};
    assign in4229_2 = {c4169,s2357[0]};
    CLA_2 KS_4229(s4229, c4229, in4229_1, in4229_2);
    wire[0:0] s4230, in4230_1, in4230_2;
    wire c4230;
    assign in4230_1 = {c4170};
    assign in4230_2 = {c4171};
    Half_Adder KS_4230(s4230, c4230, in4230_1, in4230_2);
    wire[3:0] s4231, in4231_1, in4231_2;
    wire c4231;
    assign in4231_1 = {c4172,s2358[0],c2355,c2346};
    assign in4231_2 = {c4173,s2359[0],s2356[1],s2348[2]};
    CLA_4 KS_4231(s4231, c4231, in4231_1, in4231_2);
    wire[0:0] s4232, in4232_1, in4232_2;
    wire c4232;
    assign in4232_1 = {c4174};
    assign in4232_2 = {c4175};
    Half_Adder KS_4232(s4232, c4232, in4232_1, in4232_2);
    wire[1:0] s4233, in4233_1, in4233_2;
    wire c4233;
    assign in4233_1 = {c4176,s2360[0]};
    assign in4233_2 = {c4177,s4207[1]};
    CLA_2 KS_4233(s4233, c4233, in4233_1, in4233_2);
    wire[0:0] s4234, in4234_1, in4234_2;
    wire c4234;
    assign in4234_1 = {c4178};
    assign in4234_2 = {c4179};
    Half_Adder KS_4234(s4234, c4234, in4234_1, in4234_2);
    wire[2:0] s4235, in4235_1, in4235_2;
    wire c4235;
    assign in4235_1 = {c4180,s4208[1],c2357};
    assign in4235_2 = {c4181,s4209[1],s2358[1]};
    CLA_3 KS_4235(s4235, c4235, in4235_1, in4235_2);
    wire[0:0] s4236, in4236_1, in4236_2;
    wire c4236;
    assign in4236_1 = {c4182};
    assign in4236_2 = {c4183};
    Half_Adder KS_4236(s4236, c4236, in4236_1, in4236_2);
    wire[1:0] s4237, in4237_1, in4237_2;
    wire c4237;
    assign in4237_1 = {c4184,s4210[1]};
    assign in4237_2 = {c4185,s4211[1]};
    CLA_2 KS_4237(s4237, c4237, in4237_1, in4237_2);
    wire[0:0] s4238, in4238_1, in4238_2;
    wire c4238;
    assign in4238_1 = {c4186};
    assign in4238_2 = {c4189};
    Half_Adder KS_4238(s4238, c4238, in4238_1, in4238_2);
    wire[3:0] s4239, in4239_1, in4239_2;
    wire c4239;
    assign in4239_1 = {c4197,s4212[1],c2359,c2350};
    assign in4239_2 = {c4205,s4213[1],s2360[1],s2352[2]};
    CLA_4 KS_4239(s4239, c4239, in4239_1, in4239_2);
    wire[0:0] s4240, in4240_1, in4240_2;
    wire c4240;
    assign in4240_1 = {s4207[0]};
    assign in4240_2 = {s4208[0]};
    Half_Adder KS_4240(s4240, c4240, in4240_1, in4240_2);
    wire[1:0] s4241, in4241_1, in4241_2;
    wire c4241;
    assign in4241_1 = {s4209[0],s4214[1]};
    assign in4241_2 = {s4210[0],s4215[1]};
    CLA_2 KS_4241(s4241, c4241, in4241_1, in4241_2);
    wire[0:0] s4242, in4242_1, in4242_2;
    wire c4242;
    assign in4242_1 = {s4211[0]};
    assign in4242_2 = {s4212[0]};
    Half_Adder KS_4242(s4242, c4242, in4242_1, in4242_2);
    wire[2:0] s4243, in4243_1, in4243_2;
    wire c4243;
    assign in4243_1 = {s4213[0],s4216[1],s4207[2]};
    assign in4243_2 = {s4214[0],s4217[1],s4208[2]};
    CLA_3 KS_4243(s4243, c4243, in4243_1, in4243_2);
    wire[0:0] s4244, in4244_1, in4244_2;
    wire c4244;
    assign in4244_1 = {s4216[0]};
    assign in4244_2 = {s4217[0]};
    Full_Adder KS_4244(s4244, c4244, in4244_1, in4244_2, s4215[0]);
    wire[3:0] s4245, in4245_1, in4245_2;
    wire c4245;
    assign in4245_1 = {s732[0],s2381[0],s2381[1],s2365[2]};
    assign in4245_2 = {s733[0],s2382[0],s2382[1],s2366[2]};
    CLA_4 KS_4245(s4245, c4245, in4245_1, in4245_2);
    wire[3:0] s4246, in4246_1, in4246_2;
    wire c4246;
    assign in4246_1 = {s734[0],s2383[0],s2383[1],s2367[2]};
    assign in4246_2 = {s735[0],s2384[0],s2384[1],s2368[2]};
    CLA_4 KS_4246(s4246, c4246, in4246_1, in4246_2);
    wire[3:0] s4247, in4247_1, in4247_2;
    wire c4247;
    assign in4247_1 = {s2297[3],s2385[0],s2385[1],s2369[2]};
    assign in4247_2 = {s2298[3],s2386[0],s2386[1],s2370[2]};
    CLA_4 KS_4247(s4247, c4247, in4247_1, in4247_2);
    wire[3:0] s4248, in4248_1, in4248_2;
    wire c4248;
    assign in4248_1 = {s2299[3],s2387[0],s2387[1],s2371[2]};
    assign in4248_2 = {s2300[3],s2388[0],s2388[1],s2372[2]};
    CLA_4 KS_4248(s4248, c4248, in4248_1, in4248_2);
    wire[3:0] s4249, in4249_1, in4249_2;
    wire c4249;
    assign in4249_1 = {s2301[3],s2389[0],s2389[1],s2373[2]};
    assign in4249_2 = {s2302[3],s2390[0],s2390[1],s2374[2]};
    CLA_4 KS_4249(s4249, c4249, in4249_1, in4249_2);
    wire[3:0] s4250, in4250_1, in4250_2;
    wire c4250;
    assign in4250_1 = {s2303[3],s2391[0],s2391[1],s2375[2]};
    assign in4250_2 = {s2304[3],s2392[0],s2392[1],s2376[2]};
    CLA_4 KS_4250(s4250, c4250, in4250_1, in4250_2);
    wire[3:0] s4251, in4251_1, in4251_2;
    wire c4251;
    assign in4251_1 = {s2305[3],s2393[0],c2393,s2377[2]};
    assign in4251_2 = {s2306[3],s2394[0],s2394[1],s2378[2]};
    CLA_4 KS_4251(s4251, c4251, in4251_1, in4251_2);
    wire[3:0] s4252, in4252_1, in4252_2;
    wire c4252;
    assign in4252_1 = {s2307[3],s2395[0],c2395,s2379[2]};
    assign in4252_2 = {s2308[3],s2396[0],s2396[1],s2380[2]};
    CLA_4 KS_4252(s4252, c4252, in4252_1, in4252_2);
    wire[3:0] s4253, in4253_1, in4253_2;
    wire c4253;
    assign in4253_1 = {s2309[3],s2397[0],c2397,s2381[2]};
    assign in4253_2 = {s2310[3],s2398[0],s2398[1],s2382[2]};
    CLA_4 KS_4253(s4253, c4253, in4253_1, in4253_2);
    wire[3:0] s4254, in4254_1, in4254_2;
    wire c4254;
    assign in4254_1 = {s2311[3],s2399[0],c2399,s2383[2]};
    assign in4254_2 = {s2312[3],s2400[0],s2400[1],s2384[2]};
    CLA_4 KS_4254(s4254, c4254, in4254_1, in4254_2);
    wire[3:0] s4255, in4255_1, in4255_2;
    wire c4255;
    assign in4255_1 = {s2313[3],s2401[0],c2401,s2385[2]};
    assign in4255_2 = {s2314[3],s2402[0],s2402[1],s2386[2]};
    CLA_4 KS_4255(s4255, c4255, in4255_1, in4255_2);
    wire[3:0] s4256, in4256_1, in4256_2;
    wire c4256;
    assign in4256_1 = {s2315[3],s2403[0],c2403,s2387[2]};
    assign in4256_2 = {s2316[3],s2404[0],s2404[1],s2388[2]};
    CLA_4 KS_4256(s4256, c4256, in4256_1, in4256_2);
    wire[3:0] s4257, in4257_1, in4257_2;
    wire c4257;
    assign in4257_1 = {s2317[3],s2405[0],c2405,s2389[2]};
    assign in4257_2 = {s2318[3],s2406[0],s2406[1],s2390[2]};
    CLA_4 KS_4257(s4257, c4257, in4257_1, in4257_2);
    wire[3:0] s4258, in4258_1, in4258_2;
    wire c4258;
    assign in4258_1 = {s2319[3],s2407[0],c2407,s2391[2]};
    assign in4258_2 = {s2320[3],s2408[0],s2408[1],s2392[2]};
    CLA_4 KS_4258(s4258, c4258, in4258_1, in4258_2);
    wire[3:0] s4259, in4259_1, in4259_2;
    wire c4259;
    assign in4259_1 = {s2321[3],s2409[0],c2409,c2394};
    assign in4259_2 = {s2322[3],s2410[0],s2410[1],s2396[2]};
    CLA_4 KS_4259(s4259, c4259, in4259_1, in4259_2);
    wire[3:0] s4260, in4260_1, in4260_2;
    wire c4260;
    assign in4260_1 = {s2323[3],s2411[0],c2411,c2398};
    assign in4260_2 = {s2324[3],s2412[0],s2412[1],s2400[2]};
    CLA_4 KS_4260(s4260, c4260, in4260_1, in4260_2);
    wire[3:0] s4261, in4261_1, in4261_2;
    wire c4261;
    assign in4261_1 = {s2325[3],s2413[0],c2413,c2402};
    assign in4261_2 = {s2326[3],s2414[0],s2414[1],s2404[2]};
    CLA_4 KS_4261(s4261, c4261, in4261_1, in4261_2);
    wire[3:0] s4262, in4262_1, in4262_2;
    wire c4262;
    assign in4262_1 = {s2327[3],s2415[0],c2415,c2406};
    assign in4262_2 = {s2328[3],s2416[0],s2416[1],s2408[2]};
    CLA_4 KS_4262(s4262, c4262, in4262_1, in4262_2);
    wire[2:0] s4263, in4263_1, in4263_2;
    wire c4263;
    assign in4263_1 = {c2332,s2417[0],c2417};
    assign in4263_2 = {s2336[3],s2418[0],s2418[1]};
    CLA_3 KS_4263(s4263, c4263, in4263_1, in4263_2);
    wire[0:0] s4264, in4264_1, in4264_2;
    wire c4264;
    assign in4264_1 = {c2340};
    assign in4264_2 = {s2344[3]};
    Half_Adder KS_4264(s4264, c4264, in4264_1, in4264_2);
    wire[1:0] s4265, in4265_1, in4265_2;
    wire c4265;
    assign in4265_1 = {c2348,s2419[0]};
    assign in4265_2 = {s2352[3],s2420[0]};
    CLA_2 KS_4265(s4265, c4265, in4265_1, in4265_2);
    wire[0:0] s4266, in4266_1, in4266_2;
    wire c4266;
    assign in4266_1 = {c2356};
    assign in4266_2 = {s2360[3]};
    Half_Adder KS_4266(s4266, c4266, in4266_1, in4266_2);
    wire[3:0] s4267, in4267_1, in4267_2;
    wire c4267;
    assign in4267_1 = {c4207,s2421[0],c2419,c2410};
    assign in4267_2 = {c4208,s2422[0],s2420[1],s2412[2]};
    CLA_4 KS_4267(s4267, c4267, in4267_1, in4267_2);
    wire[0:0] s4268, in4268_1, in4268_2;
    wire c4268;
    assign in4268_1 = {c4209};
    assign in4268_2 = {c4210};
    Half_Adder KS_4268(s4268, c4268, in4268_1, in4268_2);
    wire[1:0] s4269, in4269_1, in4269_2;
    wire c4269;
    assign in4269_1 = {c4211,s2423[0]};
    assign in4269_2 = {c4212,s2424[0]};
    CLA_2 KS_4269(s4269, c4269, in4269_1, in4269_2);
    wire[0:0] s4270, in4270_1, in4270_2;
    wire c4270;
    assign in4270_1 = {c4213};
    assign in4270_2 = {c4214};
    Half_Adder KS_4270(s4270, c4270, in4270_1, in4270_2);
    wire[2:0] s4271, in4271_1, in4271_2;
    wire c4271;
    assign in4271_1 = {c4215,s2425[0],c2421};
    assign in4271_2 = {c4216,s4245[1],s2422[1]};
    CLA_3 KS_4271(s4271, c4271, in4271_1, in4271_2);
    wire[0:0] s4272, in4272_1, in4272_2;
    wire c4272;
    assign in4272_1 = {c4217};
    assign in4272_2 = {c4218};
    Half_Adder KS_4272(s4272, c4272, in4272_1, in4272_2);
    wire[1:0] s4273, in4273_1, in4273_2;
    wire c4273;
    assign in4273_1 = {c4219,s4246[1]};
    assign in4273_2 = {c4220,s4247[1]};
    CLA_2 KS_4273(s4273, c4273, in4273_1, in4273_2);
    wire[0:0] s4274, in4274_1, in4274_2;
    wire c4274;
    assign in4274_1 = {c4221};
    assign in4274_2 = {c4222};
    Half_Adder KS_4274(s4274, c4274, in4274_1, in4274_2);
    wire[3:0] s4275, in4275_1, in4275_2;
    wire c4275;
    assign in4275_1 = {c4223,s4248[1],c2423,c2414};
    assign in4275_2 = {c4224,s4249[1],s2424[1],s2416[2]};
    CLA_4 KS_4275(s4275, c4275, in4275_1, in4275_2);
    wire[0:0] s4276, in4276_1, in4276_2;
    wire c4276;
    assign in4276_1 = {c4231};
    assign in4276_2 = {c4239};
    Half_Adder KS_4276(s4276, c4276, in4276_1, in4276_2);
    wire[1:0] s4277, in4277_1, in4277_2;
    wire c4277;
    assign in4277_1 = {s4245[0],s4250[1]};
    assign in4277_2 = {s4246[0],s4251[1]};
    CLA_2 KS_4277(s4277, c4277, in4277_1, in4277_2);
    wire[0:0] s4278, in4278_1, in4278_2;
    wire c4278;
    assign in4278_1 = {s4247[0]};
    assign in4278_2 = {s4248[0]};
    Half_Adder KS_4278(s4278, c4278, in4278_1, in4278_2);
    wire[2:0] s4279, in4279_1, in4279_2;
    wire c4279;
    assign in4279_1 = {s4249[0],s4252[1],c2425};
    assign in4279_2 = {s4250[0],s4253[1],s4245[2]};
    CLA_3 KS_4279(s4279, c4279, in4279_1, in4279_2);
    wire[0:0] s4280, in4280_1, in4280_2;
    wire c4280;
    assign in4280_1 = {s4252[0]};
    assign in4280_2 = {s4253[0]};
    Full_Adder KS_4280(s4280, c4280, in4280_1, in4280_2, s4251[0]);
    wire[3:0] s4281, in4281_1, in4281_2;
    wire c4281;
    assign in4281_1 = {s828[0],s2446[0],s2446[1],s2429[2]};
    assign in4281_2 = {s829[0],s2447[0],s2447[1],s2430[2]};
    CLA_4 KS_4281(s4281, c4281, in4281_1, in4281_2);
    wire[3:0] s4282, in4282_1, in4282_2;
    wire c4282;
    assign in4282_1 = {s830[0],s2448[0],s2448[1],s2431[2]};
    assign in4282_2 = {s831[0],s2449[0],s2449[1],s2432[2]};
    CLA_4 KS_4282(s4282, c4282, in4282_1, in4282_2);
    wire[3:0] s4283, in4283_1, in4283_2;
    wire c4283;
    assign in4283_1 = {s2361[3],s2450[0],s2450[1],s2433[2]};
    assign in4283_2 = {s2362[3],s2451[0],s2451[1],s2434[2]};
    CLA_4 KS_4283(s4283, c4283, in4283_1, in4283_2);
    wire[3:0] s4284, in4284_1, in4284_2;
    wire c4284;
    assign in4284_1 = {s2363[3],s2452[0],s2452[1],s2435[2]};
    assign in4284_2 = {s2364[3],s2453[0],s2453[1],s2436[2]};
    CLA_4 KS_4284(s4284, c4284, in4284_1, in4284_2);
    wire[3:0] s4285, in4285_1, in4285_2;
    wire c4285;
    assign in4285_1 = {s2365[3],s2454[0],s2454[1],s2437[2]};
    assign in4285_2 = {s2366[3],s2455[0],s2455[1],s2438[2]};
    CLA_4 KS_4285(s4285, c4285, in4285_1, in4285_2);
    wire[3:0] s4286, in4286_1, in4286_2;
    wire c4286;
    assign in4286_1 = {s2367[3],s2456[0],s2456[1],s2439[2]};
    assign in4286_2 = {s2368[3],s2457[0],s2457[1],s2440[2]};
    CLA_4 KS_4286(s4286, c4286, in4286_1, in4286_2);
    wire[3:0] s4287, in4287_1, in4287_2;
    wire c4287;
    assign in4287_1 = {s2369[3],s2458[0],c2458,s2441[2]};
    assign in4287_2 = {s2370[3],s2459[0],s2459[1],s2442[2]};
    CLA_4 KS_4287(s4287, c4287, in4287_1, in4287_2);
    wire[3:0] s4288, in4288_1, in4288_2;
    wire c4288;
    assign in4288_1 = {s2371[3],s2460[0],c2460,s2443[2]};
    assign in4288_2 = {s2372[3],s2461[0],s2461[1],s2444[2]};
    CLA_4 KS_4288(s4288, c4288, in4288_1, in4288_2);
    wire[3:0] s4289, in4289_1, in4289_2;
    wire c4289;
    assign in4289_1 = {s2373[3],s2462[0],c2462,s2445[2]};
    assign in4289_2 = {s2374[3],s2463[0],s2463[1],s2446[2]};
    CLA_4 KS_4289(s4289, c4289, in4289_1, in4289_2);
    wire[3:0] s4290, in4290_1, in4290_2;
    wire c4290;
    assign in4290_1 = {s2375[3],s2464[0],c2464,s2447[2]};
    assign in4290_2 = {s2376[3],s2465[0],s2465[1],s2448[2]};
    CLA_4 KS_4290(s4290, c4290, in4290_1, in4290_2);
    wire[3:0] s4291, in4291_1, in4291_2;
    wire c4291;
    assign in4291_1 = {s2377[3],s2466[0],c2466,s2449[2]};
    assign in4291_2 = {s2378[3],s2467[0],s2467[1],s2450[2]};
    CLA_4 KS_4291(s4291, c4291, in4291_1, in4291_2);
    wire[3:0] s4292, in4292_1, in4292_2;
    wire c4292;
    assign in4292_1 = {s2379[3],s2468[0],c2468,s2451[2]};
    assign in4292_2 = {s2380[3],s2469[0],s2469[1],s2452[2]};
    CLA_4 KS_4292(s4292, c4292, in4292_1, in4292_2);
    wire[3:0] s4293, in4293_1, in4293_2;
    wire c4293;
    assign in4293_1 = {s2381[3],s2470[0],c2470,s2453[2]};
    assign in4293_2 = {s2382[3],s2471[0],s2471[1],s2454[2]};
    CLA_4 KS_4293(s4293, c4293, in4293_1, in4293_2);
    wire[3:0] s4294, in4294_1, in4294_2;
    wire c4294;
    assign in4294_1 = {s2383[3],s2472[0],c2472,s2455[2]};
    assign in4294_2 = {s2384[3],s2473[0],s2473[1],s2456[2]};
    CLA_4 KS_4294(s4294, c4294, in4294_1, in4294_2);
    wire[3:0] s4295, in4295_1, in4295_2;
    wire c4295;
    assign in4295_1 = {s2385[3],s2474[0],c2474,c2457};
    assign in4295_2 = {s2386[3],s2475[0],s2475[1],s2459[2]};
    CLA_4 KS_4295(s4295, c4295, in4295_1, in4295_2);
    wire[3:0] s4296, in4296_1, in4296_2;
    wire c4296;
    assign in4296_1 = {s2387[3],s2476[0],c2476,c2461};
    assign in4296_2 = {s2388[3],s2477[0],s2477[1],s2463[2]};
    CLA_4 KS_4296(s4296, c4296, in4296_1, in4296_2);
    wire[3:0] s4297, in4297_1, in4297_2;
    wire c4297;
    assign in4297_1 = {s2389[3],s2478[0],c2478,c2465};
    assign in4297_2 = {s2390[3],s2479[0],s2479[1],s2467[2]};
    CLA_4 KS_4297(s4297, c4297, in4297_1, in4297_2);
    wire[3:0] s4298, in4298_1, in4298_2;
    wire c4298;
    assign in4298_1 = {s2391[3],s2480[0],c2480,c2469};
    assign in4298_2 = {s2392[3],s2481[0],s2481[1],s2471[2]};
    CLA_4 KS_4298(s4298, c4298, in4298_1, in4298_2);
    wire[3:0] s4299, in4299_1, in4299_2;
    wire c4299;
    assign in4299_1 = {c2396,s2482[0],c2482,c2473};
    assign in4299_2 = {s2400[3],s2483[0],s2483[1],s2475[2]};
    CLA_4 KS_4299(s4299, c4299, in4299_1, in4299_2);
    wire[0:0] s4300, in4300_1, in4300_2;
    wire c4300;
    assign in4300_1 = {c2404};
    assign in4300_2 = {s2408[3]};
    Half_Adder KS_4300(s4300, c4300, in4300_1, in4300_2);
    wire[1:0] s4301, in4301_1, in4301_2;
    wire c4301;
    assign in4301_1 = {c2412,s2484[0]};
    assign in4301_2 = {s2416[3],s2485[0]};
    CLA_2 KS_4301(s4301, c4301, in4301_1, in4301_2);
    wire[0:0] s4302, in4302_1, in4302_2;
    wire c4302;
    assign in4302_1 = {c2420};
    assign in4302_2 = {s2424[3]};
    Half_Adder KS_4302(s4302, c4302, in4302_1, in4302_2);
    wire[2:0] s4303, in4303_1, in4303_2;
    wire c4303;
    assign in4303_1 = {c4245,s2486[0],c2484};
    assign in4303_2 = {c4246,s2487[0],s2485[1]};
    CLA_3 KS_4303(s4303, c4303, in4303_1, in4303_2);
    wire[0:0] s4304, in4304_1, in4304_2;
    wire c4304;
    assign in4304_1 = {c4247};
    assign in4304_2 = {c4248};
    Half_Adder KS_4304(s4304, c4304, in4304_1, in4304_2);
    wire[1:0] s4305, in4305_1, in4305_2;
    wire c4305;
    assign in4305_1 = {c4249,s2488[0]};
    assign in4305_2 = {c4250,s2489[0]};
    CLA_2 KS_4305(s4305, c4305, in4305_1, in4305_2);
    wire[0:0] s4306, in4306_1, in4306_2;
    wire c4306;
    assign in4306_1 = {c4251};
    assign in4306_2 = {c4252};
    Half_Adder KS_4306(s4306, c4306, in4306_1, in4306_2);
    wire[3:0] s4307, in4307_1, in4307_2;
    wire c4307;
    assign in4307_1 = {c4253,s2490[0],c2486,c2477};
    assign in4307_2 = {c4254,s4281[1],s2487[1],s2479[2]};
    CLA_4 KS_4307(s4307, c4307, in4307_1, in4307_2);
    wire[0:0] s4308, in4308_1, in4308_2;
    wire c4308;
    assign in4308_1 = {c4255};
    assign in4308_2 = {c4256};
    Half_Adder KS_4308(s4308, c4308, in4308_1, in4308_2);
    wire[1:0] s4309, in4309_1, in4309_2;
    wire c4309;
    assign in4309_1 = {c4257,s4282[1]};
    assign in4309_2 = {c4258,s4283[1]};
    CLA_2 KS_4309(s4309, c4309, in4309_1, in4309_2);
    wire[0:0] s4310, in4310_1, in4310_2;
    wire c4310;
    assign in4310_1 = {c4259};
    assign in4310_2 = {c4260};
    Half_Adder KS_4310(s4310, c4310, in4310_1, in4310_2);
    wire[2:0] s4311, in4311_1, in4311_2;
    wire c4311;
    assign in4311_1 = {c4261,s4284[1],c2488};
    assign in4311_2 = {c4262,s4285[1],s2489[1]};
    CLA_3 KS_4311(s4311, c4311, in4311_1, in4311_2);
    wire[0:0] s4312, in4312_1, in4312_2;
    wire c4312;
    assign in4312_1 = {c4267};
    assign in4312_2 = {c4275};
    Half_Adder KS_4312(s4312, c4312, in4312_1, in4312_2);
    wire[1:0] s4313, in4313_1, in4313_2;
    wire c4313;
    assign in4313_1 = {s4281[0],s4286[1]};
    assign in4313_2 = {s4282[0],s4287[1]};
    CLA_2 KS_4313(s4313, c4313, in4313_1, in4313_2);
    wire[0:0] s4314, in4314_1, in4314_2;
    wire c4314;
    assign in4314_1 = {s4283[0]};
    assign in4314_2 = {s4284[0]};
    Half_Adder KS_4314(s4314, c4314, in4314_1, in4314_2);
    wire[3:0] s4315, in4315_1, in4315_2;
    wire c4315;
    assign in4315_1 = {s4285[0],s4288[1],c2490,c2481};
    assign in4315_2 = {s4286[0],s4289[1],s4281[2],s2483[2]};
    CLA_4 KS_4315(s4315, c4315, in4315_1, in4315_2);
    wire[0:0] s4316, in4316_1, in4316_2;
    wire c4316;
    assign in4316_1 = {s4288[0]};
    assign in4316_2 = {s4289[0]};
    Full_Adder KS_4316(s4316, c4316, in4316_1, in4316_2, s4287[0]);
    wire[3:0] s4317, in4317_1, in4317_2;
    wire c4317;
    assign in4317_1 = {s914[0],s2510[0],s2511[1],s2495[2]};
    assign in4317_2 = {s915[0],s2511[0],s2512[1],s2496[2]};
    CLA_4 KS_4317(s4317, c4317, in4317_1, in4317_2);
    wire[3:0] s4318, in4318_1, in4318_2;
    wire c4318;
    assign in4318_1 = {s916[0],s2512[0],s2513[1],s2497[2]};
    assign in4318_2 = {s917[0],s2513[0],s2514[1],s2498[2]};
    CLA_4 KS_4318(s4318, c4318, in4318_1, in4318_2);
    wire[3:0] s4319, in4319_1, in4319_2;
    wire c4319;
    assign in4319_1 = {s918[0],s2514[0],s2515[1],s2499[2]};
    assign in4319_2 = {s919[0],s2515[0],s2516[1],s2500[2]};
    CLA_4 KS_4319(s4319, c4319, in4319_1, in4319_2);
    wire[3:0] s4320, in4320_1, in4320_2;
    wire c4320;
    assign in4320_1 = {s2426[3],s2516[0],s2517[1],s2501[2]};
    assign in4320_2 = {s2427[3],s2517[0],s2518[1],s2502[2]};
    CLA_4 KS_4320(s4320, c4320, in4320_1, in4320_2);
    wire[3:0] s4321, in4321_1, in4321_2;
    wire c4321;
    assign in4321_1 = {s2428[3],s2518[0],s2519[1],s2503[2]};
    assign in4321_2 = {s2429[3],s2519[0],s2520[1],s2504[2]};
    CLA_4 KS_4321(s4321, c4321, in4321_1, in4321_2);
    wire[3:0] s4322, in4322_1, in4322_2;
    wire c4322;
    assign in4322_1 = {s2430[3],s2520[0],s2521[1],s2505[2]};
    assign in4322_2 = {s2431[3],s2521[0],s2522[1],s2506[2]};
    CLA_4 KS_4322(s4322, c4322, in4322_1, in4322_2);
    wire[3:0] s4323, in4323_1, in4323_2;
    wire c4323;
    assign in4323_1 = {s2432[3],s2522[0],c2523,s2507[2]};
    assign in4323_2 = {s2433[3],s2523[0],s2524[1],s2508[2]};
    CLA_4 KS_4323(s4323, c4323, in4323_1, in4323_2);
    wire[3:0] s4324, in4324_1, in4324_2;
    wire c4324;
    assign in4324_1 = {s2434[3],s2524[0],c2525,s2509[2]};
    assign in4324_2 = {s2435[3],s2525[0],s2526[1],s2510[2]};
    CLA_4 KS_4324(s4324, c4324, in4324_1, in4324_2);
    wire[3:0] s4325, in4325_1, in4325_2;
    wire c4325;
    assign in4325_1 = {s2436[3],s2526[0],c2527,s2511[2]};
    assign in4325_2 = {s2437[3],s2527[0],s2528[1],s2512[2]};
    CLA_4 KS_4325(s4325, c4325, in4325_1, in4325_2);
    wire[3:0] s4326, in4326_1, in4326_2;
    wire c4326;
    assign in4326_1 = {s2438[3],s2528[0],c2529,s2513[2]};
    assign in4326_2 = {s2439[3],s2529[0],s2530[1],s2514[2]};
    CLA_4 KS_4326(s4326, c4326, in4326_1, in4326_2);
    wire[3:0] s4327, in4327_1, in4327_2;
    wire c4327;
    assign in4327_1 = {s2440[3],s2530[0],c2531,s2515[2]};
    assign in4327_2 = {s2441[3],s2531[0],s2532[1],s2516[2]};
    CLA_4 KS_4327(s4327, c4327, in4327_1, in4327_2);
    wire[3:0] s4328, in4328_1, in4328_2;
    wire c4328;
    assign in4328_1 = {s2442[3],s2532[0],c2533,s2517[2]};
    assign in4328_2 = {s2443[3],s2533[0],s2534[1],s2518[2]};
    CLA_4 KS_4328(s4328, c4328, in4328_1, in4328_2);
    wire[3:0] s4329, in4329_1, in4329_2;
    wire c4329;
    assign in4329_1 = {s2444[3],s2534[0],c2535,s2519[2]};
    assign in4329_2 = {s2445[3],s2535[0],s2536[1],s2520[2]};
    CLA_4 KS_4329(s4329, c4329, in4329_1, in4329_2);
    wire[3:0] s4330, in4330_1, in4330_2;
    wire c4330;
    assign in4330_1 = {s2446[3],s2536[0],c2537,s2521[2]};
    assign in4330_2 = {s2447[3],s2537[0],s2538[1],s2522[2]};
    CLA_4 KS_4330(s4330, c4330, in4330_1, in4330_2);
    wire[3:0] s4331, in4331_1, in4331_2;
    wire c4331;
    assign in4331_1 = {s2448[3],s2538[0],c2539,c2524};
    assign in4331_2 = {s2449[3],s2539[0],s2540[1],s2526[2]};
    CLA_4 KS_4331(s4331, c4331, in4331_1, in4331_2);
    wire[3:0] s4332, in4332_1, in4332_2;
    wire c4332;
    assign in4332_1 = {s2450[3],s2540[0],c2541,c2528};
    assign in4332_2 = {s2451[3],s2541[0],s2542[1],s2530[2]};
    CLA_4 KS_4332(s4332, c4332, in4332_1, in4332_2);
    wire[3:0] s4333, in4333_1, in4333_2;
    wire c4333;
    assign in4333_1 = {s2452[3],s2542[0],c2543,c2532};
    assign in4333_2 = {s2453[3],s2543[0],s2544[1],s2534[2]};
    CLA_4 KS_4333(s4333, c4333, in4333_1, in4333_2);
    wire[3:0] s4334, in4334_1, in4334_2;
    wire c4334;
    assign in4334_1 = {s2454[3],s2544[0],c2545,c2536};
    assign in4334_2 = {s2455[3],s2545[0],s2546[1],s2538[2]};
    CLA_4 KS_4334(s4334, c4334, in4334_1, in4334_2);
    wire[1:0] s4335, in4335_1, in4335_2;
    wire c4335;
    assign in4335_1 = {s2456[3],s2546[0]};
    assign in4335_2 = {s2459[3],s2547[0]};
    CLA_2 KS_4335(s4335, c4335, in4335_1, in4335_2);
    wire[0:0] s4336, in4336_1, in4336_2;
    wire c4336;
    assign in4336_1 = {c2463};
    assign in4336_2 = {s2467[3]};
    Half_Adder KS_4336(s4336, c4336, in4336_1, in4336_2);
    wire[2:0] s4337, in4337_1, in4337_2;
    wire c4337;
    assign in4337_1 = {c2471,s2548[0],c2547};
    assign in4337_2 = {s2475[3],s2549[0],s2548[1]};
    CLA_3 KS_4337(s4337, c4337, in4337_1, in4337_2);
    wire[0:0] s4338, in4338_1, in4338_2;
    wire c4338;
    assign in4338_1 = {c2479};
    assign in4338_2 = {s2483[3]};
    Half_Adder KS_4338(s4338, c4338, in4338_1, in4338_2);
    wire[1:0] s4339, in4339_1, in4339_2;
    wire c4339;
    assign in4339_1 = {c2487,s2550[0]};
    assign in4339_2 = {c4281,s2551[0]};
    CLA_2 KS_4339(s4339, c4339, in4339_1, in4339_2);
    wire[0:0] s4340, in4340_1, in4340_2;
    wire c4340;
    assign in4340_1 = {c4282};
    assign in4340_2 = {c4283};
    Half_Adder KS_4340(s4340, c4340, in4340_1, in4340_2);
    wire[3:0] s4341, in4341_1, in4341_2;
    wire c4341;
    assign in4341_1 = {c4284,s2552[0],c2549,c2540};
    assign in4341_2 = {c4285,s2553[0],s2550[1],s2542[2]};
    CLA_4 KS_4341(s4341, c4341, in4341_1, in4341_2);
    wire[0:0] s4342, in4342_1, in4342_2;
    wire c4342;
    assign in4342_1 = {c4286};
    assign in4342_2 = {c4287};
    Half_Adder KS_4342(s4342, c4342, in4342_1, in4342_2);
    wire[1:0] s4343, in4343_1, in4343_2;
    wire c4343;
    assign in4343_1 = {c4288,s2554[0]};
    assign in4343_2 = {c4289,s4317[1]};
    CLA_2 KS_4343(s4343, c4343, in4343_1, in4343_2);
    wire[0:0] s4344, in4344_1, in4344_2;
    wire c4344;
    assign in4344_1 = {c4290};
    assign in4344_2 = {c4291};
    Half_Adder KS_4344(s4344, c4344, in4344_1, in4344_2);
    wire[2:0] s4345, in4345_1, in4345_2;
    wire c4345;
    assign in4345_1 = {c4292,s4318[1],c2551};
    assign in4345_2 = {c4293,s4319[1],s2552[1]};
    CLA_3 KS_4345(s4345, c4345, in4345_1, in4345_2);
    wire[0:0] s4346, in4346_1, in4346_2;
    wire c4346;
    assign in4346_1 = {c4294};
    assign in4346_2 = {c4295};
    Half_Adder KS_4346(s4346, c4346, in4346_1, in4346_2);
    wire[1:0] s4347, in4347_1, in4347_2;
    wire c4347;
    assign in4347_1 = {c4296,s4320[1]};
    assign in4347_2 = {c4297,s4321[1]};
    CLA_2 KS_4347(s4347, c4347, in4347_1, in4347_2);
    wire[0:0] s4348, in4348_1, in4348_2;
    wire c4348;
    assign in4348_1 = {c4298};
    assign in4348_2 = {c4299};
    Half_Adder KS_4348(s4348, c4348, in4348_1, in4348_2);
    wire[3:0] s4349, in4349_1, in4349_2;
    wire c4349;
    assign in4349_1 = {c4307,s4322[1],c2553,c2544};
    assign in4349_2 = {c4315,s4323[1],s2554[1],s2546[2]};
    CLA_4 KS_4349(s4349, c4349, in4349_1, in4349_2);
    wire[0:0] s4350, in4350_1, in4350_2;
    wire c4350;
    assign in4350_1 = {s4317[0]};
    assign in4350_2 = {s4318[0]};
    Half_Adder KS_4350(s4350, c4350, in4350_1, in4350_2);
    wire[1:0] s4351, in4351_1, in4351_2;
    wire c4351;
    assign in4351_1 = {s4319[0],s4324[1]};
    assign in4351_2 = {s4320[0],s4325[1]};
    CLA_2 KS_4351(s4351, c4351, in4351_1, in4351_2);
    wire[0:0] s4352, in4352_1, in4352_2;
    wire c4352;
    assign in4352_1 = {s4321[0]};
    assign in4352_2 = {s4322[0]};
    Half_Adder KS_4352(s4352, c4352, in4352_1, in4352_2);
    wire[2:0] s4353, in4353_1, in4353_2;
    wire c4353;
    assign in4353_1 = {s4323[0],s4326[1],s4317[2]};
    assign in4353_2 = {s4324[0],s4327[1],s4318[2]};
    CLA_3 KS_4353(s4353, c4353, in4353_1, in4353_2);
    wire[0:0] s4354, in4354_1, in4354_2;
    wire c4354;
    assign in4354_1 = {s4326[0]};
    assign in4354_2 = {s4327[0]};
    Full_Adder KS_4354(s4354, c4354, in4354_1, in4354_2, s4325[0]);
    wire[3:0] s4355, in4355_1, in4355_2;
    wire c4355;
    assign in4355_1 = {s995[0],s2576[0],s2576[1],s2558[2]};
    assign in4355_2 = {s996[0],s2577[0],s2577[1],s2559[2]};
    CLA_4 KS_4355(s4355, c4355, in4355_1, in4355_2);
    wire[3:0] s4356, in4356_1, in4356_2;
    wire c4356;
    assign in4356_1 = {s997[0],s2578[0],s2578[1],s2560[2]};
    assign in4356_2 = {s998[0],s2579[0],s2579[1],s2561[2]};
    CLA_4 KS_4356(s4356, c4356, in4356_1, in4356_2);
    wire[3:0] s4357, in4357_1, in4357_2;
    wire c4357;
    assign in4357_1 = {s2491[3],s2580[0],s2580[1],s2562[2]};
    assign in4357_2 = {s2492[3],s2581[0],s2581[1],s2563[2]};
    CLA_4 KS_4357(s4357, c4357, in4357_1, in4357_2);
    wire[3:0] s4358, in4358_1, in4358_2;
    wire c4358;
    assign in4358_1 = {s2493[3],s2582[0],s2582[1],s2564[2]};
    assign in4358_2 = {s2494[3],s2583[0],s2583[1],s2565[2]};
    CLA_4 KS_4358(s4358, c4358, in4358_1, in4358_2);
    wire[3:0] s4359, in4359_1, in4359_2;
    wire c4359;
    assign in4359_1 = {s2495[3],s2584[0],s2584[1],s2566[2]};
    assign in4359_2 = {s2496[3],s2585[0],s2585[1],s2567[2]};
    CLA_4 KS_4359(s4359, c4359, in4359_1, in4359_2);
    wire[3:0] s4360, in4360_1, in4360_2;
    wire c4360;
    assign in4360_1 = {s2497[3],s2586[0],c2586,s2568[2]};
    assign in4360_2 = {s2498[3],s2587[0],s2587[1],s2569[2]};
    CLA_4 KS_4360(s4360, c4360, in4360_1, in4360_2);
    wire[3:0] s4361, in4361_1, in4361_2;
    wire c4361;
    assign in4361_1 = {s2499[3],s2588[0],c2588,s2570[2]};
    assign in4361_2 = {s2500[3],s2589[0],s2589[1],s2571[2]};
    CLA_4 KS_4361(s4361, c4361, in4361_1, in4361_2);
    wire[3:0] s4362, in4362_1, in4362_2;
    wire c4362;
    assign in4362_1 = {s2501[3],s2590[0],c2590,s2572[2]};
    assign in4362_2 = {s2502[3],s2591[0],s2591[1],s2573[2]};
    CLA_4 KS_4362(s4362, c4362, in4362_1, in4362_2);
    wire[3:0] s4363, in4363_1, in4363_2;
    wire c4363;
    assign in4363_1 = {s2503[3],s2592[0],c2592,s2574[2]};
    assign in4363_2 = {s2504[3],s2593[0],s2593[1],s2575[2]};
    CLA_4 KS_4363(s4363, c4363, in4363_1, in4363_2);
    wire[3:0] s4364, in4364_1, in4364_2;
    wire c4364;
    assign in4364_1 = {s2505[3],s2594[0],c2594,s2576[2]};
    assign in4364_2 = {s2506[3],s2595[0],s2595[1],s2577[2]};
    CLA_4 KS_4364(s4364, c4364, in4364_1, in4364_2);
    wire[3:0] s4365, in4365_1, in4365_2;
    wire c4365;
    assign in4365_1 = {s2507[3],s2596[0],c2596,s2578[2]};
    assign in4365_2 = {s2508[3],s2597[0],s2597[1],s2579[2]};
    CLA_4 KS_4365(s4365, c4365, in4365_1, in4365_2);
    wire[3:0] s4366, in4366_1, in4366_2;
    wire c4366;
    assign in4366_1 = {s2509[3],s2598[0],c2598,s2580[2]};
    assign in4366_2 = {s2510[3],s2599[0],s2599[1],s2581[2]};
    CLA_4 KS_4366(s4366, c4366, in4366_1, in4366_2);
    wire[3:0] s4367, in4367_1, in4367_2;
    wire c4367;
    assign in4367_1 = {s2511[3],s2600[0],c2600,s2582[2]};
    assign in4367_2 = {s2512[3],s2601[0],s2601[1],s2583[2]};
    CLA_4 KS_4367(s4367, c4367, in4367_1, in4367_2);
    wire[3:0] s4368, in4368_1, in4368_2;
    wire c4368;
    assign in4368_1 = {s2513[3],s2602[0],c2602,s2584[2]};
    assign in4368_2 = {s2514[3],s2603[0],s2603[1],s2585[2]};
    CLA_4 KS_4368(s4368, c4368, in4368_1, in4368_2);
    wire[3:0] s4369, in4369_1, in4369_2;
    wire c4369;
    assign in4369_1 = {s2515[3],s2604[0],c2604,c2587};
    assign in4369_2 = {s2516[3],s2605[0],s2605[1],s2589[2]};
    CLA_4 KS_4369(s4369, c4369, in4369_1, in4369_2);
    wire[3:0] s4370, in4370_1, in4370_2;
    wire c4370;
    assign in4370_1 = {s2517[3],s2606[0],c2606,c2591};
    assign in4370_2 = {s2518[3],s2607[0],s2607[1],s2593[2]};
    CLA_4 KS_4370(s4370, c4370, in4370_1, in4370_2);
    wire[3:0] s4371, in4371_1, in4371_2;
    wire c4371;
    assign in4371_1 = {s2519[3],s2608[0],c2608,c2595};
    assign in4371_2 = {s2520[3],s2609[0],s2609[1],s2597[2]};
    CLA_4 KS_4371(s4371, c4371, in4371_1, in4371_2);
    wire[3:0] s4372, in4372_1, in4372_2;
    wire c4372;
    assign in4372_1 = {s2521[3],s2610[0],c2610,c2599};
    assign in4372_2 = {s2522[3],s2611[0],s2611[1],s2601[2]};
    CLA_4 KS_4372(s4372, c4372, in4372_1, in4372_2);
    wire[3:0] s4373, in4373_1, in4373_2;
    wire c4373;
    assign in4373_1 = {c2526,s2612[0],c2612,c2603};
    assign in4373_2 = {s2530[3],s2613[0],s2613[1],s2605[2]};
    CLA_4 KS_4373(s4373, c4373, in4373_1, in4373_2);
    wire[0:0] s4374, in4374_1, in4374_2;
    wire c4374;
    assign in4374_1 = {c2534};
    assign in4374_2 = {s2538[3]};
    Half_Adder KS_4374(s4374, c4374, in4374_1, in4374_2);
    wire[1:0] s4375, in4375_1, in4375_2;
    wire c4375;
    assign in4375_1 = {c2542,s2614[0]};
    assign in4375_2 = {s2546[3],s2615[0]};
    CLA_2 KS_4375(s4375, c4375, in4375_1, in4375_2);
    wire[0:0] s4376, in4376_1, in4376_2;
    wire c4376;
    assign in4376_1 = {c2550};
    assign in4376_2 = {s2554[3]};
    Half_Adder KS_4376(s4376, c4376, in4376_1, in4376_2);
    wire[2:0] s4377, in4377_1, in4377_2;
    wire c4377;
    assign in4377_1 = {c4317,s2616[0],c2614};
    assign in4377_2 = {c4318,s2617[0],s2615[1]};
    CLA_3 KS_4377(s4377, c4377, in4377_1, in4377_2);
    wire[0:0] s4378, in4378_1, in4378_2;
    wire c4378;
    assign in4378_1 = {c4319};
    assign in4378_2 = {c4320};
    Half_Adder KS_4378(s4378, c4378, in4378_1, in4378_2);
    wire[1:0] s4379, in4379_1, in4379_2;
    wire c4379;
    assign in4379_1 = {c4321,s2618[0]};
    assign in4379_2 = {c4322,s2619[0]};
    CLA_2 KS_4379(s4379, c4379, in4379_1, in4379_2);
    wire[0:0] s4380, in4380_1, in4380_2;
    wire c4380;
    assign in4380_1 = {c4323};
    assign in4380_2 = {c4324};
    Half_Adder KS_4380(s4380, c4380, in4380_1, in4380_2);
    wire[3:0] s4381, in4381_1, in4381_2;
    wire c4381;
    assign in4381_1 = {c4325,s2620[0],c2616,c2607};
    assign in4381_2 = {c4326,s4355[1],s2617[1],s2609[2]};
    CLA_4 KS_4381(s4381, c4381, in4381_1, in4381_2);
    wire[0:0] s4382, in4382_1, in4382_2;
    wire c4382;
    assign in4382_1 = {c4327};
    assign in4382_2 = {c4328};
    Half_Adder KS_4382(s4382, c4382, in4382_1, in4382_2);
    wire[1:0] s4383, in4383_1, in4383_2;
    wire c4383;
    assign in4383_1 = {c4329,s4356[1]};
    assign in4383_2 = {c4330,s4357[1]};
    CLA_2 KS_4383(s4383, c4383, in4383_1, in4383_2);
    wire[0:0] s4384, in4384_1, in4384_2;
    wire c4384;
    assign in4384_1 = {c4331};
    assign in4384_2 = {c4332};
    Half_Adder KS_4384(s4384, c4384, in4384_1, in4384_2);
    wire[2:0] s4385, in4385_1, in4385_2;
    wire c4385;
    assign in4385_1 = {c4333,s4358[1],c2618};
    assign in4385_2 = {c4334,s4359[1],s2619[1]};
    CLA_3 KS_4385(s4385, c4385, in4385_1, in4385_2);
    wire[0:0] s4386, in4386_1, in4386_2;
    wire c4386;
    assign in4386_1 = {c4341};
    assign in4386_2 = {c4349};
    Half_Adder KS_4386(s4386, c4386, in4386_1, in4386_2);
    wire[1:0] s4387, in4387_1, in4387_2;
    wire c4387;
    assign in4387_1 = {s4355[0],s4360[1]};
    assign in4387_2 = {s4356[0],s4361[1]};
    CLA_2 KS_4387(s4387, c4387, in4387_1, in4387_2);
    wire[0:0] s4388, in4388_1, in4388_2;
    wire c4388;
    assign in4388_1 = {s4357[0]};
    assign in4388_2 = {s4358[0]};
    Half_Adder KS_4388(s4388, c4388, in4388_1, in4388_2);
    wire[3:0] s4389, in4389_1, in4389_2;
    wire c4389;
    assign in4389_1 = {s4359[0],s4362[1],c2620,c2611};
    assign in4389_2 = {s4360[0],s4363[1],s4355[2],s2613[2]};
    CLA_4 KS_4389(s4389, c4389, in4389_1, in4389_2);
    wire[0:0] s4390, in4390_1, in4390_2;
    wire c4390;
    assign in4390_1 = {s4362[0]};
    assign in4390_2 = {s4363[0]};
    Full_Adder KS_4390(s4390, c4390, in4390_1, in4390_2, s4361[0]);
    wire[3:0] s4391, in4391_1, in4391_2;
    wire c4391;
    assign in4391_1 = {s1064[0],s2641[0],s2642[1],s2625[2]};
    assign in4391_2 = {s1065[0],s2642[0],s2643[1],s2626[2]};
    CLA_4 KS_4391(s4391, c4391, in4391_1, in4391_2);
    wire[3:0] s4392, in4392_1, in4392_2;
    wire c4392;
    assign in4392_1 = {s1066[0],s2643[0],s2644[1],s2627[2]};
    assign in4392_2 = {s1067[0],s2644[0],s2645[1],s2628[2]};
    CLA_4 KS_4392(s4392, c4392, in4392_1, in4392_2);
    wire[3:0] s4393, in4393_1, in4393_2;
    wire c4393;
    assign in4393_1 = {s1068[0],s2645[0],s2646[1],s2629[2]};
    assign in4393_2 = {s1069[0],s2646[0],s2647[1],s2630[2]};
    CLA_4 KS_4393(s4393, c4393, in4393_1, in4393_2);
    wire[3:0] s4394, in4394_1, in4394_2;
    wire c4394;
    assign in4394_1 = {s2555[3],s2647[0],s2648[1],s2631[2]};
    assign in4394_2 = {s2556[3],s2648[0],s2649[1],s2632[2]};
    CLA_4 KS_4394(s4394, c4394, in4394_1, in4394_2);
    wire[3:0] s4395, in4395_1, in4395_2;
    wire c4395;
    assign in4395_1 = {s2557[3],s2649[0],s2650[1],s2633[2]};
    assign in4395_2 = {s2558[3],s2650[0],s2651[1],s2634[2]};
    CLA_4 KS_4395(s4395, c4395, in4395_1, in4395_2);
    wire[3:0] s4396, in4396_1, in4396_2;
    wire c4396;
    assign in4396_1 = {s2559[3],s2651[0],c2652,s2635[2]};
    assign in4396_2 = {s2560[3],s2652[0],s2653[1],s2636[2]};
    CLA_4 KS_4396(s4396, c4396, in4396_1, in4396_2);
    wire[3:0] s4397, in4397_1, in4397_2;
    wire c4397;
    assign in4397_1 = {s2561[3],s2653[0],c2654,s2637[2]};
    assign in4397_2 = {s2562[3],s2654[0],s2655[1],s2638[2]};
    CLA_4 KS_4397(s4397, c4397, in4397_1, in4397_2);
    wire[3:0] s4398, in4398_1, in4398_2;
    wire c4398;
    assign in4398_1 = {s2563[3],s2655[0],c2656,s2639[2]};
    assign in4398_2 = {s2564[3],s2656[0],s2657[1],s2640[2]};
    CLA_4 KS_4398(s4398, c4398, in4398_1, in4398_2);
    wire[3:0] s4399, in4399_1, in4399_2;
    wire c4399;
    assign in4399_1 = {s2565[3],s2657[0],c2658,s2641[2]};
    assign in4399_2 = {s2566[3],s2658[0],s2659[1],s2642[2]};
    CLA_4 KS_4399(s4399, c4399, in4399_1, in4399_2);
    wire[3:0] s4400, in4400_1, in4400_2;
    wire c4400;
    assign in4400_1 = {s2567[3],s2659[0],c2660,s2643[2]};
    assign in4400_2 = {s2568[3],s2660[0],s2661[1],s2644[2]};
    CLA_4 KS_4400(s4400, c4400, in4400_1, in4400_2);
    wire[3:0] s4401, in4401_1, in4401_2;
    wire c4401;
    assign in4401_1 = {s2569[3],s2661[0],c2662,s2645[2]};
    assign in4401_2 = {s2570[3],s2662[0],s2663[1],s2646[2]};
    CLA_4 KS_4401(s4401, c4401, in4401_1, in4401_2);
    wire[3:0] s4402, in4402_1, in4402_2;
    wire c4402;
    assign in4402_1 = {s2571[3],s2663[0],c2664,s2647[2]};
    assign in4402_2 = {s2572[3],s2664[0],s2665[1],s2648[2]};
    CLA_4 KS_4402(s4402, c4402, in4402_1, in4402_2);
    wire[3:0] s4403, in4403_1, in4403_2;
    wire c4403;
    assign in4403_1 = {s2573[3],s2665[0],c2666,s2649[2]};
    assign in4403_2 = {s2574[3],s2666[0],s2667[1],s2650[2]};
    CLA_4 KS_4403(s4403, c4403, in4403_1, in4403_2);
    wire[3:0] s4404, in4404_1, in4404_2;
    wire c4404;
    assign in4404_1 = {s2575[3],s2667[0],c2668,s2651[2]};
    assign in4404_2 = {s2576[3],s2668[0],s2669[1],s2653[2]};
    CLA_4 KS_4404(s4404, c4404, in4404_1, in4404_2);
    wire[3:0] s4405, in4405_1, in4405_2;
    wire c4405;
    assign in4405_1 = {s2577[3],s2669[0],c2670,c2655};
    assign in4405_2 = {s2578[3],s2670[0],s2671[1],s2657[2]};
    CLA_4 KS_4405(s4405, c4405, in4405_1, in4405_2);
    wire[3:0] s4406, in4406_1, in4406_2;
    wire c4406;
    assign in4406_1 = {s2579[3],s2671[0],c2672,c2659};
    assign in4406_2 = {s2580[3],s2672[0],s2673[1],s2661[2]};
    CLA_4 KS_4406(s4406, c4406, in4406_1, in4406_2);
    wire[3:0] s4407, in4407_1, in4407_2;
    wire c4407;
    assign in4407_1 = {s2581[3],s2673[0],c2674,c2663};
    assign in4407_2 = {s2582[3],s2674[0],s2675[1],s2665[2]};
    CLA_4 KS_4407(s4407, c4407, in4407_1, in4407_2);
    wire[3:0] s4408, in4408_1, in4408_2;
    wire c4408;
    assign in4408_1 = {s2583[3],s2675[0],c2676,c2667};
    assign in4408_2 = {s2584[3],s2676[0],s2677[1],s2669[2]};
    CLA_4 KS_4408(s4408, c4408, in4408_1, in4408_2);
    wire[1:0] s4409, in4409_1, in4409_2;
    wire c4409;
    assign in4409_1 = {s2585[3],s2677[0]};
    assign in4409_2 = {s2589[3],s2678[0]};
    CLA_2 KS_4409(s4409, c4409, in4409_1, in4409_2);
    wire[0:0] s4410, in4410_1, in4410_2;
    wire c4410;
    assign in4410_1 = {c2593};
    assign in4410_2 = {s2597[3]};
    Half_Adder KS_4410(s4410, c4410, in4410_1, in4410_2);
    wire[2:0] s4411, in4411_1, in4411_2;
    wire c4411;
    assign in4411_1 = {c2601,s2679[0],c2678};
    assign in4411_2 = {s2605[3],s2680[0],s2679[1]};
    CLA_3 KS_4411(s4411, c4411, in4411_1, in4411_2);
    wire[0:0] s4412, in4412_1, in4412_2;
    wire c4412;
    assign in4412_1 = {c2609};
    assign in4412_2 = {s2613[3]};
    Half_Adder KS_4412(s4412, c4412, in4412_1, in4412_2);
    wire[1:0] s4413, in4413_1, in4413_2;
    wire c4413;
    assign in4413_1 = {c2617,s2681[0]};
    assign in4413_2 = {c4355,s2682[0]};
    CLA_2 KS_4413(s4413, c4413, in4413_1, in4413_2);
    wire[0:0] s4414, in4414_1, in4414_2;
    wire c4414;
    assign in4414_1 = {c4356};
    assign in4414_2 = {c4357};
    Half_Adder KS_4414(s4414, c4414, in4414_1, in4414_2);
    wire[3:0] s4415, in4415_1, in4415_2;
    wire c4415;
    assign in4415_1 = {c4358,s2683[0],c2680,c2671};
    assign in4415_2 = {c4359,s2684[0],s2681[1],s2673[2]};
    CLA_4 KS_4415(s4415, c4415, in4415_1, in4415_2);
    wire[0:0] s4416, in4416_1, in4416_2;
    wire c4416;
    assign in4416_1 = {c4360};
    assign in4416_2 = {c4361};
    Half_Adder KS_4416(s4416, c4416, in4416_1, in4416_2);
    wire[1:0] s4417, in4417_1, in4417_2;
    wire c4417;
    assign in4417_1 = {c4362,s2685[0]};
    assign in4417_2 = {c4363,s4391[1]};
    CLA_2 KS_4417(s4417, c4417, in4417_1, in4417_2);
    wire[0:0] s4418, in4418_1, in4418_2;
    wire c4418;
    assign in4418_1 = {c4364};
    assign in4418_2 = {c4365};
    Half_Adder KS_4418(s4418, c4418, in4418_1, in4418_2);
    wire[2:0] s4419, in4419_1, in4419_2;
    wire c4419;
    assign in4419_1 = {c4366,s4392[1],c2682};
    assign in4419_2 = {c4367,s4393[1],s2683[1]};
    CLA_3 KS_4419(s4419, c4419, in4419_1, in4419_2);
    wire[0:0] s4420, in4420_1, in4420_2;
    wire c4420;
    assign in4420_1 = {c4368};
    assign in4420_2 = {c4369};
    Half_Adder KS_4420(s4420, c4420, in4420_1, in4420_2);
    wire[1:0] s4421, in4421_1, in4421_2;
    wire c4421;
    assign in4421_1 = {c4370,s4394[1]};
    assign in4421_2 = {c4371,s4395[1]};
    CLA_2 KS_4421(s4421, c4421, in4421_1, in4421_2);
    wire[0:0] s4422, in4422_1, in4422_2;
    wire c4422;
    assign in4422_1 = {c4372};
    assign in4422_2 = {c4373};
    Half_Adder KS_4422(s4422, c4422, in4422_1, in4422_2);
    wire[3:0] s4423, in4423_1, in4423_2;
    wire c4423;
    assign in4423_1 = {c4381,s4396[1],c2684,c2675};
    assign in4423_2 = {c4389,s4397[1],s2685[1],s2677[2]};
    CLA_4 KS_4423(s4423, c4423, in4423_1, in4423_2);
    wire[0:0] s4424, in4424_1, in4424_2;
    wire c4424;
    assign in4424_1 = {s4391[0]};
    assign in4424_2 = {s4392[0]};
    Half_Adder KS_4424(s4424, c4424, in4424_1, in4424_2);
    wire[1:0] s4425, in4425_1, in4425_2;
    wire c4425;
    assign in4425_1 = {s4393[0],s4398[1]};
    assign in4425_2 = {s4394[0],s4399[1]};
    CLA_2 KS_4425(s4425, c4425, in4425_1, in4425_2);
    wire[0:0] s4426, in4426_1, in4426_2;
    wire c4426;
    assign in4426_1 = {s4395[0]};
    assign in4426_2 = {s4396[0]};
    Half_Adder KS_4426(s4426, c4426, in4426_1, in4426_2);
    wire[2:0] s4427, in4427_1, in4427_2;
    wire c4427;
    assign in4427_1 = {s4397[0],s4400[1],s4391[2]};
    assign in4427_2 = {s4398[0],s4401[1],s4392[2]};
    CLA_3 KS_4427(s4427, c4427, in4427_1, in4427_2);
    wire[0:0] s4428, in4428_1, in4428_2;
    wire c4428;
    assign in4428_1 = {s4400[0]};
    assign in4428_2 = {s4401[0]};
    Full_Adder KS_4428(s4428, c4428, in4428_1, in4428_2, s4399[0]);
    wire[3:0] s4429, in4429_1, in4429_2;
    wire c4429;
    assign in4429_1 = {s1128[0],s2706[0],s2707[1],s2689[2]};
    assign in4429_2 = {s1129[0],s2707[0],s2708[1],s2690[2]};
    CLA_4 KS_4429(s4429, c4429, in4429_1, in4429_2);
    wire[3:0] s4430, in4430_1, in4430_2;
    wire c4430;
    assign in4430_1 = {s1130[0],s2708[0],s2709[1],s2691[2]};
    assign in4430_2 = {s1131[0],s2709[0],s2710[1],s2692[2]};
    CLA_4 KS_4430(s4430, c4430, in4430_1, in4430_2);
    wire[3:0] s4431, in4431_1, in4431_2;
    wire c4431;
    assign in4431_1 = {s2621[3],s2710[0],s2711[1],s2693[2]};
    assign in4431_2 = {s2622[3],s2711[0],s2712[1],s2694[2]};
    CLA_4 KS_4431(s4431, c4431, in4431_1, in4431_2);
    wire[3:0] s4432, in4432_1, in4432_2;
    wire c4432;
    assign in4432_1 = {s2623[3],s2712[0],s2713[1],s2695[2]};
    assign in4432_2 = {s2624[3],s2713[0],s2714[1],s2696[2]};
    CLA_4 KS_4432(s4432, c4432, in4432_1, in4432_2);
    wire[3:0] s4433, in4433_1, in4433_2;
    wire c4433;
    assign in4433_1 = {s2625[3],s2714[0],s2715[1],s2697[2]};
    assign in4433_2 = {s2626[3],s2715[0],s2716[1],s2698[2]};
    CLA_4 KS_4433(s4433, c4433, in4433_1, in4433_2);
    wire[3:0] s4434, in4434_1, in4434_2;
    wire c4434;
    assign in4434_1 = {s2627[3],s2716[0],c2717,s2699[2]};
    assign in4434_2 = {s2628[3],s2717[0],s2718[1],s2700[2]};
    CLA_4 KS_4434(s4434, c4434, in4434_1, in4434_2);
    wire[3:0] s4435, in4435_1, in4435_2;
    wire c4435;
    assign in4435_1 = {s2629[3],s2718[0],c2719,s2701[2]};
    assign in4435_2 = {s2630[3],s2719[0],s2720[1],s2702[2]};
    CLA_4 KS_4435(s4435, c4435, in4435_1, in4435_2);
    wire[3:0] s4436, in4436_1, in4436_2;
    wire c4436;
    assign in4436_1 = {s2631[3],s2720[0],c2721,s2703[2]};
    assign in4436_2 = {s2632[3],s2721[0],s2722[1],s2704[2]};
    CLA_4 KS_4436(s4436, c4436, in4436_1, in4436_2);
    wire[3:0] s4437, in4437_1, in4437_2;
    wire c4437;
    assign in4437_1 = {s2633[3],s2722[0],c2723,s2705[2]};
    assign in4437_2 = {s2634[3],s2723[0],s2724[1],s2706[2]};
    CLA_4 KS_4437(s4437, c4437, in4437_1, in4437_2);
    wire[3:0] s4438, in4438_1, in4438_2;
    wire c4438;
    assign in4438_1 = {s2635[3],s2724[0],c2725,s2707[2]};
    assign in4438_2 = {s2636[3],s2725[0],s2726[1],s2708[2]};
    CLA_4 KS_4438(s4438, c4438, in4438_1, in4438_2);
    wire[3:0] s4439, in4439_1, in4439_2;
    wire c4439;
    assign in4439_1 = {s2637[3],s2726[0],c2727,s2709[2]};
    assign in4439_2 = {s2638[3],s2727[0],s2728[1],s2710[2]};
    CLA_4 KS_4439(s4439, c4439, in4439_1, in4439_2);
    wire[3:0] s4440, in4440_1, in4440_2;
    wire c4440;
    assign in4440_1 = {s2639[3],s2728[0],c2729,s2711[2]};
    assign in4440_2 = {s2640[3],s2729[0],s2730[1],s2712[2]};
    CLA_4 KS_4440(s4440, c4440, in4440_1, in4440_2);
    wire[3:0] s4441, in4441_1, in4441_2;
    wire c4441;
    assign in4441_1 = {s2641[3],s2730[0],c2731,s2713[2]};
    assign in4441_2 = {s2642[3],s2731[0],s2732[1],s2714[2]};
    CLA_4 KS_4441(s4441, c4441, in4441_1, in4441_2);
    wire[3:0] s4442, in4442_1, in4442_2;
    wire c4442;
    assign in4442_1 = {s2643[3],s2732[0],c2733,s2715[2]};
    assign in4442_2 = {s2644[3],s2733[0],s2734[1],s2716[2]};
    CLA_4 KS_4442(s4442, c4442, in4442_1, in4442_2);
    wire[3:0] s4443, in4443_1, in4443_2;
    wire c4443;
    assign in4443_1 = {s2645[3],s2734[0],c2735,c2718};
    assign in4443_2 = {s2646[3],s2735[0],s2736[1],s2720[2]};
    CLA_4 KS_4443(s4443, c4443, in4443_1, in4443_2);
    wire[3:0] s4444, in4444_1, in4444_2;
    wire c4444;
    assign in4444_1 = {s2647[3],s2736[0],c2737,c2722};
    assign in4444_2 = {s2648[3],s2737[0],s2738[1],s2724[2]};
    CLA_4 KS_4444(s4444, c4444, in4444_1, in4444_2);
    wire[3:0] s4445, in4445_1, in4445_2;
    wire c4445;
    assign in4445_1 = {s2649[3],s2738[0],c2739,c2726};
    assign in4445_2 = {s2650[3],s2739[0],s2740[1],s2728[2]};
    CLA_4 KS_4445(s4445, c4445, in4445_1, in4445_2);
    wire[3:0] s4446, in4446_1, in4446_2;
    wire c4446;
    assign in4446_1 = {s2651[3],s2740[0],c2741,c2730};
    assign in4446_2 = {s2653[3],s2741[0],s2742[1],s2732[2]};
    CLA_4 KS_4446(s4446, c4446, in4446_1, in4446_2);
    wire[1:0] s4447, in4447_1, in4447_2;
    wire c4447;
    assign in4447_1 = {c2657,s2742[0]};
    assign in4447_2 = {s2661[3],s2743[0]};
    CLA_2 KS_4447(s4447, c4447, in4447_1, in4447_2);
    wire[0:0] s4448, in4448_1, in4448_2;
    wire c4448;
    assign in4448_1 = {c2665};
    assign in4448_2 = {s2669[3]};
    Half_Adder KS_4448(s4448, c4448, in4448_1, in4448_2);
    wire[3:0] s4449, in4449_1, in4449_2;
    wire c4449;
    assign in4449_1 = {c2673,s2744[0],c2743,c2734};
    assign in4449_2 = {s2677[3],s2745[0],s2744[1],s2736[2]};
    CLA_4 KS_4449(s4449, c4449, in4449_1, in4449_2);
    wire[0:0] s4450, in4450_1, in4450_2;
    wire c4450;
    assign in4450_1 = {c2681};
    assign in4450_2 = {s2685[3]};
    Half_Adder KS_4450(s4450, c4450, in4450_1, in4450_2);
    wire[1:0] s4451, in4451_1, in4451_2;
    wire c4451;
    assign in4451_1 = {c4391,s2746[0]};
    assign in4451_2 = {c4392,s2747[0]};
    CLA_2 KS_4451(s4451, c4451, in4451_1, in4451_2);
    wire[0:0] s4452, in4452_1, in4452_2;
    wire c4452;
    assign in4452_1 = {c4393};
    assign in4452_2 = {c4394};
    Half_Adder KS_4452(s4452, c4452, in4452_1, in4452_2);
    wire[2:0] s4453, in4453_1, in4453_2;
    wire c4453;
    assign in4453_1 = {c4395,s2748[0],c2745};
    assign in4453_2 = {c4396,s2749[0],s2746[1]};
    CLA_3 KS_4453(s4453, c4453, in4453_1, in4453_2);
    wire[0:0] s4454, in4454_1, in4454_2;
    wire c4454;
    assign in4454_1 = {c4397};
    assign in4454_2 = {c4398};
    Half_Adder KS_4454(s4454, c4454, in4454_1, in4454_2);
    wire[1:0] s4455, in4455_1, in4455_2;
    wire c4455;
    assign in4455_1 = {c4399,s2750[0]};
    assign in4455_2 = {c4400,s4429[1]};
    CLA_2 KS_4455(s4455, c4455, in4455_1, in4455_2);
    wire[0:0] s4456, in4456_1, in4456_2;
    wire c4456;
    assign in4456_1 = {c4401};
    assign in4456_2 = {c4402};
    Half_Adder KS_4456(s4456, c4456, in4456_1, in4456_2);
    wire[3:0] s4457, in4457_1, in4457_2;
    wire c4457;
    assign in4457_1 = {c4403,s4430[1],c2747,c2738};
    assign in4457_2 = {c4404,s4431[1],s2748[1],s2740[2]};
    CLA_4 KS_4457(s4457, c4457, in4457_1, in4457_2);
    wire[0:0] s4458, in4458_1, in4458_2;
    wire c4458;
    assign in4458_1 = {c4405};
    assign in4458_2 = {c4406};
    Half_Adder KS_4458(s4458, c4458, in4458_1, in4458_2);
    wire[1:0] s4459, in4459_1, in4459_2;
    wire c4459;
    assign in4459_1 = {c4407,s4432[1]};
    assign in4459_2 = {c4408,s4433[1]};
    CLA_2 KS_4459(s4459, c4459, in4459_1, in4459_2);
    wire[0:0] s4460, in4460_1, in4460_2;
    wire c4460;
    assign in4460_1 = {c4415};
    assign in4460_2 = {c4423};
    Half_Adder KS_4460(s4460, c4460, in4460_1, in4460_2);
    wire[2:0] s4461, in4461_1, in4461_2;
    wire c4461;
    assign in4461_1 = {s4429[0],s4434[1],c2749};
    assign in4461_2 = {s4430[0],s4435[1],s2750[1]};
    CLA_3 KS_4461(s4461, c4461, in4461_1, in4461_2);
    wire[0:0] s4462, in4462_1, in4462_2;
    wire c4462;
    assign in4462_1 = {s4431[0]};
    assign in4462_2 = {s4432[0]};
    Half_Adder KS_4462(s4462, c4462, in4462_1, in4462_2);
    wire[1:0] s4463, in4463_1, in4463_2;
    wire c4463;
    assign in4463_1 = {s4433[0],s4436[1]};
    assign in4463_2 = {s4434[0],s4437[1]};
    CLA_2 KS_4463(s4463, c4463, in4463_1, in4463_2);
    wire[0:0] s4464, in4464_1, in4464_2;
    wire c4464;
    assign in4464_1 = {s4436[0]};
    assign in4464_2 = {s4437[0]};
    Full_Adder KS_4464(s4464, c4464, in4464_1, in4464_2, s4435[0]);
    wire[3:0] s4465, in4465_1, in4465_2;
    wire c4465;
    assign in4465_1 = {s1180[0],s2770[0],s2770[1],s2753[2]};
    assign in4465_2 = {s1181[0],s2771[0],s2771[1],s2754[2]};
    CLA_4 KS_4465(s4465, c4465, in4465_1, in4465_2);
    wire[3:0] s4466, in4466_1, in4466_2;
    wire c4466;
    assign in4466_1 = {s1182[0],s2772[0],s2772[1],s2755[2]};
    assign in4466_2 = {s1183[0],s2773[0],s2773[1],s2756[2]};
    CLA_4 KS_4466(s4466, c4466, in4466_1, in4466_2);
    wire[3:0] s4467, in4467_1, in4467_2;
    wire c4467;
    assign in4467_1 = {s1184[0],s2774[0],s2774[1],s2757[2]};
    assign in4467_2 = {s1185[0],s2775[0],s2775[1],s2758[2]};
    CLA_4 KS_4467(s4467, c4467, in4467_1, in4467_2);
    wire[3:0] s4468, in4468_1, in4468_2;
    wire c4468;
    assign in4468_1 = {s2686[3],s2776[0],s2776[1],s2759[2]};
    assign in4468_2 = {s2687[3],s2777[0],s2777[1],s2760[2]};
    CLA_4 KS_4468(s4468, c4468, in4468_1, in4468_2);
    wire[3:0] s4469, in4469_1, in4469_2;
    wire c4469;
    assign in4469_1 = {s2688[3],s2778[0],s2778[1],s2761[2]};
    assign in4469_2 = {s2689[3],s2779[0],s2779[1],s2762[2]};
    CLA_4 KS_4469(s4469, c4469, in4469_1, in4469_2);
    wire[3:0] s4470, in4470_1, in4470_2;
    wire c4470;
    assign in4470_1 = {s2690[3],s2780[0],s2780[1],s2763[2]};
    assign in4470_2 = {s2691[3],s2781[0],s2781[1],s2764[2]};
    CLA_4 KS_4470(s4470, c4470, in4470_1, in4470_2);
    wire[3:0] s4471, in4471_1, in4471_2;
    wire c4471;
    assign in4471_1 = {s2692[3],s2782[0],c2782,s2765[2]};
    assign in4471_2 = {s2693[3],s2783[0],s2783[1],s2766[2]};
    CLA_4 KS_4471(s4471, c4471, in4471_1, in4471_2);
    wire[3:0] s4472, in4472_1, in4472_2;
    wire c4472;
    assign in4472_1 = {s2694[3],s2784[0],c2784,s2767[2]};
    assign in4472_2 = {s2695[3],s2785[0],s2785[1],s2768[2]};
    CLA_4 KS_4472(s4472, c4472, in4472_1, in4472_2);
    wire[3:0] s4473, in4473_1, in4473_2;
    wire c4473;
    assign in4473_1 = {s2696[3],s2786[0],c2786,s2769[2]};
    assign in4473_2 = {s2697[3],s2787[0],s2787[1],s2770[2]};
    CLA_4 KS_4473(s4473, c4473, in4473_1, in4473_2);
    wire[3:0] s4474, in4474_1, in4474_2;
    wire c4474;
    assign in4474_1 = {s2698[3],s2788[0],c2788,s2771[2]};
    assign in4474_2 = {s2699[3],s2789[0],s2789[1],s2772[2]};
    CLA_4 KS_4474(s4474, c4474, in4474_1, in4474_2);
    wire[3:0] s4475, in4475_1, in4475_2;
    wire c4475;
    assign in4475_1 = {s2700[3],s2790[0],c2790,s2773[2]};
    assign in4475_2 = {s2701[3],s2791[0],s2791[1],s2774[2]};
    CLA_4 KS_4475(s4475, c4475, in4475_1, in4475_2);
    wire[3:0] s4476, in4476_1, in4476_2;
    wire c4476;
    assign in4476_1 = {s2702[3],s2792[0],c2792,s2775[2]};
    assign in4476_2 = {s2703[3],s2793[0],s2793[1],s2776[2]};
    CLA_4 KS_4476(s4476, c4476, in4476_1, in4476_2);
    wire[3:0] s4477, in4477_1, in4477_2;
    wire c4477;
    assign in4477_1 = {s2704[3],s2794[0],c2794,s2777[2]};
    assign in4477_2 = {s2705[3],s2795[0],s2795[1],s2778[2]};
    CLA_4 KS_4477(s4477, c4477, in4477_1, in4477_2);
    wire[3:0] s4478, in4478_1, in4478_2;
    wire c4478;
    assign in4478_1 = {s2706[3],s2796[0],c2796,s2779[2]};
    assign in4478_2 = {s2707[3],s2797[0],s2797[1],s2780[2]};
    CLA_4 KS_4478(s4478, c4478, in4478_1, in4478_2);
    wire[3:0] s4479, in4479_1, in4479_2;
    wire c4479;
    assign in4479_1 = {s2708[3],s2798[0],c2798,s2781[2]};
    assign in4479_2 = {s2709[3],s2799[0],s2799[1],s2783[2]};
    CLA_4 KS_4479(s4479, c4479, in4479_1, in4479_2);
    wire[3:0] s4480, in4480_1, in4480_2;
    wire c4480;
    assign in4480_1 = {s2710[3],s2800[0],c2800,c2785};
    assign in4480_2 = {s2711[3],s2801[0],s2801[1],s2787[2]};
    CLA_4 KS_4480(s4480, c4480, in4480_1, in4480_2);
    wire[3:0] s4481, in4481_1, in4481_2;
    wire c4481;
    assign in4481_1 = {s2712[3],s2802[0],c2802,c2789};
    assign in4481_2 = {s2713[3],s2803[0],s2803[1],s2791[2]};
    CLA_4 KS_4481(s4481, c4481, in4481_1, in4481_2);
    wire[3:0] s4482, in4482_1, in4482_2;
    wire c4482;
    assign in4482_1 = {s2714[3],s2804[0],c2804,c2793};
    assign in4482_2 = {s2715[3],s2805[0],s2805[1],s2795[2]};
    CLA_4 KS_4482(s4482, c4482, in4482_1, in4482_2);
    wire[3:0] s4483, in4483_1, in4483_2;
    wire c4483;
    assign in4483_1 = {s2716[3],s2806[0],c2806,c2797};
    assign in4483_2 = {s2720[3],s2807[0],s2807[1],s2799[2]};
    CLA_4 KS_4483(s4483, c4483, in4483_1, in4483_2);
    wire[0:0] s4484, in4484_1, in4484_2;
    wire c4484;
    assign in4484_1 = {c2724};
    assign in4484_2 = {s2728[3]};
    Half_Adder KS_4484(s4484, c4484, in4484_1, in4484_2);
    wire[1:0] s4485, in4485_1, in4485_2;
    wire c4485;
    assign in4485_1 = {c2732,s2808[0]};
    assign in4485_2 = {s2736[3],s2809[0]};
    CLA_2 KS_4485(s4485, c4485, in4485_1, in4485_2);
    wire[0:0] s4486, in4486_1, in4486_2;
    wire c4486;
    assign in4486_1 = {c2740};
    assign in4486_2 = {s2744[3]};
    Half_Adder KS_4486(s4486, c4486, in4486_1, in4486_2);
    wire[2:0] s4487, in4487_1, in4487_2;
    wire c4487;
    assign in4487_1 = {c2748,s2810[0],c2808};
    assign in4487_2 = {c4429,s2811[0],s2809[1]};
    CLA_3 KS_4487(s4487, c4487, in4487_1, in4487_2);
    wire[0:0] s4488, in4488_1, in4488_2;
    wire c4488;
    assign in4488_1 = {c4430};
    assign in4488_2 = {c4431};
    Half_Adder KS_4488(s4488, c4488, in4488_1, in4488_2);
    wire[1:0] s4489, in4489_1, in4489_2;
    wire c4489;
    assign in4489_1 = {c4432,s2812[0]};
    assign in4489_2 = {c4433,s2813[0]};
    CLA_2 KS_4489(s4489, c4489, in4489_1, in4489_2);
    wire[0:0] s4490, in4490_1, in4490_2;
    wire c4490;
    assign in4490_1 = {c4434};
    assign in4490_2 = {c4435};
    Half_Adder KS_4490(s4490, c4490, in4490_1, in4490_2);
    wire[3:0] s4491, in4491_1, in4491_2;
    wire c4491;
    assign in4491_1 = {c4436,s2814[0],c2810,c2801};
    assign in4491_2 = {c4437,s4465[1],s2811[1],s2803[2]};
    CLA_4 KS_4491(s4491, c4491, in4491_1, in4491_2);
    wire[0:0] s4492, in4492_1, in4492_2;
    wire c4492;
    assign in4492_1 = {c4438};
    assign in4492_2 = {c4439};
    Half_Adder KS_4492(s4492, c4492, in4492_1, in4492_2);
    wire[1:0] s4493, in4493_1, in4493_2;
    wire c4493;
    assign in4493_1 = {c4440,s4466[1]};
    assign in4493_2 = {c4441,s4467[1]};
    CLA_2 KS_4493(s4493, c4493, in4493_1, in4493_2);
    wire[0:0] s4494, in4494_1, in4494_2;
    wire c4494;
    assign in4494_1 = {c4442};
    assign in4494_2 = {c4443};
    Half_Adder KS_4494(s4494, c4494, in4494_1, in4494_2);
    wire[2:0] s4495, in4495_1, in4495_2;
    wire c4495;
    assign in4495_1 = {c4444,s4468[1],c2812};
    assign in4495_2 = {c4445,s4469[1],s2813[1]};
    CLA_3 KS_4495(s4495, c4495, in4495_1, in4495_2);
    wire[0:0] s4496, in4496_1, in4496_2;
    wire c4496;
    assign in4496_1 = {c4446};
    assign in4496_2 = {c4449};
    Half_Adder KS_4496(s4496, c4496, in4496_1, in4496_2);
    wire[1:0] s4497, in4497_1, in4497_2;
    wire c4497;
    assign in4497_1 = {c4457,s4470[1]};
    assign in4497_2 = {s4465[0],s4471[1]};
    CLA_2 KS_4497(s4497, c4497, in4497_1, in4497_2);
    wire[0:0] s4498, in4498_1, in4498_2;
    wire c4498;
    assign in4498_1 = {s4466[0]};
    assign in4498_2 = {s4467[0]};
    Half_Adder KS_4498(s4498, c4498, in4498_1, in4498_2);
    wire[3:0] s4499, in4499_1, in4499_2;
    wire c4499;
    assign in4499_1 = {s4468[0],s4472[1],c2814,c2805};
    assign in4499_2 = {s4469[0],s4473[1],s4465[2],s2807[2]};
    CLA_4 KS_4499(s4499, c4499, in4499_1, in4499_2);
    wire[0:0] s4500, in4500_1, in4500_2;
    wire c4500;
    assign in4500_1 = {s4470[0]};
    assign in4500_2 = {s4471[0]};
    Half_Adder KS_4500(s4500, c4500, in4500_1, in4500_2);
    wire[1:0] s4501, in4501_1, in4501_2;
    wire c4501;
    assign in4501_1 = {s4473[0],s4474[1]};
    assign in4501_2 = {s4474[0],s4475[1]};
    CLA_2_c KS_4501(s4501, c4501, in4501_1, in4501_2, s4472[0]);
    wire[3:0] s4502, in4502_1, in4502_2;
    wire c4502;
    assign in4502_1 = {s1225[0],s2835[0],s2835[1],s2819[2]};
    assign in4502_2 = {s1226[0],s2836[0],s2836[1],s2820[2]};
    CLA_4 KS_4502(s4502, c4502, in4502_1, in4502_2);
    wire[3:0] s4503, in4503_1, in4503_2;
    wire c4503;
    assign in4503_1 = {s1227[0],s2837[0],s2837[1],s2821[2]};
    assign in4503_2 = {s1228[0],s2838[0],s2838[1],s2822[2]};
    CLA_4 KS_4503(s4503, c4503, in4503_1, in4503_2);
    wire[3:0] s4504, in4504_1, in4504_2;
    wire c4504;
    assign in4504_1 = {s1229[0],s2839[0],s2839[1],s2823[2]};
    assign in4504_2 = {s1230[0],s2840[0],s2840[1],s2824[2]};
    CLA_4 KS_4504(s4504, c4504, in4504_1, in4504_2);
    wire[3:0] s4505, in4505_1, in4505_2;
    wire c4505;
    assign in4505_1 = {s2751[3],s2841[0],s2841[1],s2825[2]};
    assign in4505_2 = {s2752[3],s2842[0],s2842[1],s2826[2]};
    CLA_4 KS_4505(s4505, c4505, in4505_1, in4505_2);
    wire[3:0] s4506, in4506_1, in4506_2;
    wire c4506;
    assign in4506_1 = {s2753[3],s2843[0],s2843[1],s2827[2]};
    assign in4506_2 = {s2754[3],s2844[0],s2844[1],s2828[2]};
    CLA_4 KS_4506(s4506, c4506, in4506_1, in4506_2);
    wire[3:0] s4507, in4507_1, in4507_2;
    wire c4507;
    assign in4507_1 = {s2755[3],s2845[0],s2845[1],s2829[2]};
    assign in4507_2 = {s2756[3],s2846[0],s2846[1],s2830[2]};
    CLA_4 KS_4507(s4507, c4507, in4507_1, in4507_2);
    wire[3:0] s4508, in4508_1, in4508_2;
    wire c4508;
    assign in4508_1 = {s2757[3],s2847[0],c2847,s2831[2]};
    assign in4508_2 = {s2758[3],s2848[0],s2848[1],s2832[2]};
    CLA_4 KS_4508(s4508, c4508, in4508_1, in4508_2);
    wire[3:0] s4509, in4509_1, in4509_2;
    wire c4509;
    assign in4509_1 = {s2759[3],s2849[0],c2849,s2833[2]};
    assign in4509_2 = {s2760[3],s2850[0],s2850[1],s2834[2]};
    CLA_4 KS_4509(s4509, c4509, in4509_1, in4509_2);
    wire[3:0] s4510, in4510_1, in4510_2;
    wire c4510;
    assign in4510_1 = {s2761[3],s2851[0],c2851,s2835[2]};
    assign in4510_2 = {s2762[3],s2852[0],s2852[1],s2836[2]};
    CLA_4 KS_4510(s4510, c4510, in4510_1, in4510_2);
    wire[3:0] s4511, in4511_1, in4511_2;
    wire c4511;
    assign in4511_1 = {s2763[3],s2853[0],c2853,s2837[2]};
    assign in4511_2 = {s2764[3],s2854[0],s2854[1],s2838[2]};
    CLA_4 KS_4511(s4511, c4511, in4511_1, in4511_2);
    wire[3:0] s4512, in4512_1, in4512_2;
    wire c4512;
    assign in4512_1 = {s2765[3],s2855[0],c2855,s2839[2]};
    assign in4512_2 = {s2766[3],s2856[0],s2856[1],s2840[2]};
    CLA_4 KS_4512(s4512, c4512, in4512_1, in4512_2);
    wire[3:0] s4513, in4513_1, in4513_2;
    wire c4513;
    assign in4513_1 = {s2767[3],s2857[0],c2857,s2841[2]};
    assign in4513_2 = {s2768[3],s2858[0],s2858[1],s2842[2]};
    CLA_4 KS_4513(s4513, c4513, in4513_1, in4513_2);
    wire[3:0] s4514, in4514_1, in4514_2;
    wire c4514;
    assign in4514_1 = {s2769[3],s2859[0],c2859,s2843[2]};
    assign in4514_2 = {s2770[3],s2860[0],s2860[1],s2844[2]};
    CLA_4 KS_4514(s4514, c4514, in4514_1, in4514_2);
    wire[3:0] s4515, in4515_1, in4515_2;
    wire c4515;
    assign in4515_1 = {s2771[3],s2861[0],c2861,s2845[2]};
    assign in4515_2 = {s2772[3],s2862[0],s2862[1],s2846[2]};
    CLA_4 KS_4515(s4515, c4515, in4515_1, in4515_2);
    wire[3:0] s4516, in4516_1, in4516_2;
    wire c4516;
    assign in4516_1 = {s2773[3],s2863[0],c2863,c2848};
    assign in4516_2 = {s2774[3],s2864[0],s2864[1],s2850[2]};
    CLA_4 KS_4516(s4516, c4516, in4516_1, in4516_2);
    wire[3:0] s4517, in4517_1, in4517_2;
    wire c4517;
    assign in4517_1 = {s2775[3],s2865[0],c2865,c2852};
    assign in4517_2 = {s2776[3],s2866[0],s2866[1],s2854[2]};
    CLA_4 KS_4517(s4517, c4517, in4517_1, in4517_2);
    wire[3:0] s4518, in4518_1, in4518_2;
    wire c4518;
    assign in4518_1 = {s2777[3],s2867[0],c2867,c2856};
    assign in4518_2 = {s2778[3],s2868[0],s2868[1],s2858[2]};
    CLA_4 KS_4518(s4518, c4518, in4518_1, in4518_2);
    wire[3:0] s4519, in4519_1, in4519_2;
    wire c4519;
    assign in4519_1 = {s2779[3],s2869[0],c2869,c2860};
    assign in4519_2 = {s2780[3],s2870[0],s2870[1],s2862[2]};
    CLA_4 KS_4519(s4519, c4519, in4519_1, in4519_2);
    wire[2:0] s4520, in4520_1, in4520_2;
    wire c4520;
    assign in4520_1 = {s2781[3],s2871[0],c2871};
    assign in4520_2 = {s2783[3],s2872[0],s2872[1]};
    CLA_3 KS_4520(s4520, c4520, in4520_1, in4520_2);
    wire[0:0] s4521, in4521_1, in4521_2;
    wire c4521;
    assign in4521_1 = {c2787};
    assign in4521_2 = {s2791[3]};
    Half_Adder KS_4521(s4521, c4521, in4521_1, in4521_2);
    wire[1:0] s4522, in4522_1, in4522_2;
    wire c4522;
    assign in4522_1 = {c2795,s2873[0]};
    assign in4522_2 = {s2799[3],s2874[0]};
    CLA_2 KS_4522(s4522, c4522, in4522_1, in4522_2);
    wire[0:0] s4523, in4523_1, in4523_2;
    wire c4523;
    assign in4523_1 = {c2803};
    assign in4523_2 = {s2807[3]};
    Half_Adder KS_4523(s4523, c4523, in4523_1, in4523_2);
    wire[3:0] s4524, in4524_1, in4524_2;
    wire c4524;
    assign in4524_1 = {c2811,s2875[0],c2873,c2864};
    assign in4524_2 = {c4465,s2876[0],s2874[1],s2866[2]};
    CLA_4 KS_4524(s4524, c4524, in4524_1, in4524_2);
    wire[0:0] s4525, in4525_1, in4525_2;
    wire c4525;
    assign in4525_1 = {c4466};
    assign in4525_2 = {c4467};
    Half_Adder KS_4525(s4525, c4525, in4525_1, in4525_2);
    wire[1:0] s4526, in4526_1, in4526_2;
    wire c4526;
    assign in4526_1 = {c4468,s2877[0]};
    assign in4526_2 = {c4469,s2878[0]};
    CLA_2 KS_4526(s4526, c4526, in4526_1, in4526_2);
    wire[0:0] s4527, in4527_1, in4527_2;
    wire c4527;
    assign in4527_1 = {c4470};
    assign in4527_2 = {c4471};
    Half_Adder KS_4527(s4527, c4527, in4527_1, in4527_2);
    wire[2:0] s4528, in4528_1, in4528_2;
    wire c4528;
    assign in4528_1 = {c4472,s2879[0],c2875};
    assign in4528_2 = {c4473,s4502[1],s2876[1]};
    CLA_3 KS_4528(s4528, c4528, in4528_1, in4528_2);
    wire[0:0] s4529, in4529_1, in4529_2;
    wire c4529;
    assign in4529_1 = {c4474};
    assign in4529_2 = {c4475};
    Half_Adder KS_4529(s4529, c4529, in4529_1, in4529_2);
    wire[1:0] s4530, in4530_1, in4530_2;
    wire c4530;
    assign in4530_1 = {c4476,s4503[1]};
    assign in4530_2 = {c4477,s4504[1]};
    CLA_2 KS_4530(s4530, c4530, in4530_1, in4530_2);
    wire[0:0] s4531, in4531_1, in4531_2;
    wire c4531;
    assign in4531_1 = {c4478};
    assign in4531_2 = {c4479};
    Half_Adder KS_4531(s4531, c4531, in4531_1, in4531_2);
    wire[3:0] s4532, in4532_1, in4532_2;
    wire c4532;
    assign in4532_1 = {c4480,s4505[1],c2877,c2868};
    assign in4532_2 = {c4481,s4506[1],s2878[1],s2870[2]};
    CLA_4 KS_4532(s4532, c4532, in4532_1, in4532_2);
    wire[0:0] s4533, in4533_1, in4533_2;
    wire c4533;
    assign in4533_1 = {c4482};
    assign in4533_2 = {c4483};
    Half_Adder KS_4533(s4533, c4533, in4533_1, in4533_2);
    wire[1:0] s4534, in4534_1, in4534_2;
    wire c4534;
    assign in4534_1 = {c4491,s4507[1]};
    assign in4534_2 = {c4499,s4508[1]};
    CLA_2 KS_4534(s4534, c4534, in4534_1, in4534_2);
    wire[0:0] s4535, in4535_1, in4535_2;
    wire c4535;
    assign in4535_1 = {s4502[0]};
    assign in4535_2 = {s4503[0]};
    Half_Adder KS_4535(s4535, c4535, in4535_1, in4535_2);
    wire[2:0] s4536, in4536_1, in4536_2;
    wire c4536;
    assign in4536_1 = {s4504[0],s4509[1],c2879};
    assign in4536_2 = {s4505[0],s4510[1],s4502[2]};
    CLA_3 KS_4536(s4536, c4536, in4536_1, in4536_2);
    wire[0:0] s4537, in4537_1, in4537_2;
    wire c4537;
    assign in4537_1 = {s4506[0]};
    assign in4537_2 = {s4507[0]};
    Half_Adder KS_4537(s4537, c4537, in4537_1, in4537_2);
    wire[1:0] s4538, in4538_1, in4538_2;
    wire c4538;
    assign in4538_1 = {s4508[0],s4511[1]};
    assign in4538_2 = {s4509[0],s4512[1]};
    CLA_2 KS_4538(s4538, c4538, in4538_1, in4538_2);
    wire[0:0] s4539, in4539_1, in4539_2;
    wire c4539;
    assign in4539_1 = {s4511[0]};
    assign in4539_2 = {s4512[0]};
    Full_Adder KS_4539(s4539, c4539, in4539_1, in4539_2, s4510[0]);
    wire[3:0] s4540, in4540_1, in4540_2;
    wire c4540;
    assign in4540_1 = {s1263[0],s2900[0],s2900[1],s2883[2]};
    assign in4540_2 = {s1264[0],s2901[0],s2901[1],s2884[2]};
    CLA_4 KS_4540(s4540, c4540, in4540_1, in4540_2);
    wire[3:0] s4541, in4541_1, in4541_2;
    wire c4541;
    assign in4541_1 = {s1265[0],s2902[0],s2902[1],s2885[2]};
    assign in4541_2 = {s1266[0],s2903[0],s2903[1],s2886[2]};
    CLA_4 KS_4541(s4541, c4541, in4541_1, in4541_2);
    wire[3:0] s4542, in4542_1, in4542_2;
    wire c4542;
    assign in4542_1 = {s2815[3],s2904[0],s2904[1],s2887[2]};
    assign in4542_2 = {s2816[3],s2905[0],s2905[1],s2888[2]};
    CLA_4 KS_4542(s4542, c4542, in4542_1, in4542_2);
    wire[3:0] s4543, in4543_1, in4543_2;
    wire c4543;
    assign in4543_1 = {s2817[3],s2906[0],s2906[1],s2889[2]};
    assign in4543_2 = {s2818[3],s2907[0],s2907[1],s2890[2]};
    CLA_4 KS_4543(s4543, c4543, in4543_1, in4543_2);
    wire[3:0] s4544, in4544_1, in4544_2;
    wire c4544;
    assign in4544_1 = {s2819[3],s2908[0],s2908[1],s2891[2]};
    assign in4544_2 = {s2820[3],s2909[0],s2909[1],s2892[2]};
    CLA_4 KS_4544(s4544, c4544, in4544_1, in4544_2);
    wire[3:0] s4545, in4545_1, in4545_2;
    wire c4545;
    assign in4545_1 = {s2821[3],s2910[0],s2910[1],s2893[2]};
    assign in4545_2 = {s2822[3],s2911[0],s2911[1],s2894[2]};
    CLA_4 KS_4545(s4545, c4545, in4545_1, in4545_2);
    wire[3:0] s4546, in4546_1, in4546_2;
    wire c4546;
    assign in4546_1 = {s2823[3],s2912[0],c2912,s2895[2]};
    assign in4546_2 = {s2824[3],s2913[0],s2913[1],s2896[2]};
    CLA_4 KS_4546(s4546, c4546, in4546_1, in4546_2);
    wire[3:0] s4547, in4547_1, in4547_2;
    wire c4547;
    assign in4547_1 = {s2825[3],s2914[0],c2914,s2897[2]};
    assign in4547_2 = {s2826[3],s2915[0],s2915[1],s2898[2]};
    CLA_4 KS_4547(s4547, c4547, in4547_1, in4547_2);
    wire[3:0] s4548, in4548_1, in4548_2;
    wire c4548;
    assign in4548_1 = {s2827[3],s2916[0],c2916,s2899[2]};
    assign in4548_2 = {s2828[3],s2917[0],s2917[1],s2900[2]};
    CLA_4 KS_4548(s4548, c4548, in4548_1, in4548_2);
    wire[3:0] s4549, in4549_1, in4549_2;
    wire c4549;
    assign in4549_1 = {s2829[3],s2918[0],c2918,s2901[2]};
    assign in4549_2 = {s2830[3],s2919[0],s2919[1],s2902[2]};
    CLA_4 KS_4549(s4549, c4549, in4549_1, in4549_2);
    wire[3:0] s4550, in4550_1, in4550_2;
    wire c4550;
    assign in4550_1 = {s2831[3],s2920[0],c2920,s2903[2]};
    assign in4550_2 = {s2832[3],s2921[0],s2921[1],s2904[2]};
    CLA_4 KS_4550(s4550, c4550, in4550_1, in4550_2);
    wire[3:0] s4551, in4551_1, in4551_2;
    wire c4551;
    assign in4551_1 = {s2833[3],s2922[0],c2922,s2905[2]};
    assign in4551_2 = {s2834[3],s2923[0],s2923[1],s2906[2]};
    CLA_4 KS_4551(s4551, c4551, in4551_1, in4551_2);
    wire[3:0] s4552, in4552_1, in4552_2;
    wire c4552;
    assign in4552_1 = {s2835[3],s2924[0],c2924,s2907[2]};
    assign in4552_2 = {s2836[3],s2925[0],s2925[1],s2908[2]};
    CLA_4 KS_4552(s4552, c4552, in4552_1, in4552_2);
    wire[3:0] s4553, in4553_1, in4553_2;
    wire c4553;
    assign in4553_1 = {s2837[3],s2926[0],c2926,s2909[2]};
    assign in4553_2 = {s2838[3],s2927[0],s2927[1],s2910[2]};
    CLA_4 KS_4553(s4553, c4553, in4553_1, in4553_2);
    wire[3:0] s4554, in4554_1, in4554_2;
    wire c4554;
    assign in4554_1 = {s2839[3],s2928[0],c2928,c2911};
    assign in4554_2 = {s2840[3],s2929[0],s2929[1],s2913[2]};
    CLA_4 KS_4554(s4554, c4554, in4554_1, in4554_2);
    wire[3:0] s4555, in4555_1, in4555_2;
    wire c4555;
    assign in4555_1 = {s2841[3],s2930[0],c2930,c2915};
    assign in4555_2 = {s2842[3],s2931[0],s2931[1],s2917[2]};
    CLA_4 KS_4555(s4555, c4555, in4555_1, in4555_2);
    wire[3:0] s4556, in4556_1, in4556_2;
    wire c4556;
    assign in4556_1 = {s2843[3],s2932[0],c2932,c2919};
    assign in4556_2 = {s2844[3],s2933[0],s2933[1],s2921[2]};
    CLA_4 KS_4556(s4556, c4556, in4556_1, in4556_2);
    wire[3:0] s4557, in4557_1, in4557_2;
    wire c4557;
    assign in4557_1 = {s2845[3],s2934[0],c2934,c2923};
    assign in4557_2 = {s2846[3],s2935[0],s2935[1],s2925[2]};
    CLA_4 KS_4557(s4557, c4557, in4557_1, in4557_2);
    wire[3:0] s4558, in4558_1, in4558_2;
    wire c4558;
    assign in4558_1 = {c2850,s2936[0],c2936,c2927};
    assign in4558_2 = {s2854[3],s2937[0],s2937[1],s2929[2]};
    CLA_4 KS_4558(s4558, c4558, in4558_1, in4558_2);
    wire[0:0] s4559, in4559_1, in4559_2;
    wire c4559;
    assign in4559_1 = {c2858};
    assign in4559_2 = {s2862[3]};
    Half_Adder KS_4559(s4559, c4559, in4559_1, in4559_2);
    wire[1:0] s4560, in4560_1, in4560_2;
    wire c4560;
    assign in4560_1 = {c2866,s2938[0]};
    assign in4560_2 = {s2870[3],s2939[0]};
    CLA_2 KS_4560(s4560, c4560, in4560_1, in4560_2);
    wire[0:0] s4561, in4561_1, in4561_2;
    wire c4561;
    assign in4561_1 = {c2874};
    assign in4561_2 = {s2878[3]};
    Half_Adder KS_4561(s4561, c4561, in4561_1, in4561_2);
    wire[2:0] s4562, in4562_1, in4562_2;
    wire c4562;
    assign in4562_1 = {c4502,s2940[0],c2938};
    assign in4562_2 = {c4503,s2941[0],s2939[1]};
    CLA_3 KS_4562(s4562, c4562, in4562_1, in4562_2);
    wire[0:0] s4563, in4563_1, in4563_2;
    wire c4563;
    assign in4563_1 = {c4504};
    assign in4563_2 = {c4505};
    Half_Adder KS_4563(s4563, c4563, in4563_1, in4563_2);
    wire[1:0] s4564, in4564_1, in4564_2;
    wire c4564;
    assign in4564_1 = {c4506,s2942[0]};
    assign in4564_2 = {c4507,s2943[0]};
    CLA_2 KS_4564(s4564, c4564, in4564_1, in4564_2);
    wire[0:0] s4565, in4565_1, in4565_2;
    wire c4565;
    assign in4565_1 = {c4508};
    assign in4565_2 = {c4509};
    Half_Adder KS_4565(s4565, c4565, in4565_1, in4565_2);
    wire[3:0] s4566, in4566_1, in4566_2;
    wire c4566;
    assign in4566_1 = {c4510,s2944[0],c2940,c2931};
    assign in4566_2 = {c4511,s4540[1],s2941[1],s2933[2]};
    CLA_4 KS_4566(s4566, c4566, in4566_1, in4566_2);
    wire[0:0] s4567, in4567_1, in4567_2;
    wire c4567;
    assign in4567_1 = {c4512};
    assign in4567_2 = {c4513};
    Half_Adder KS_4567(s4567, c4567, in4567_1, in4567_2);
    wire[1:0] s4568, in4568_1, in4568_2;
    wire c4568;
    assign in4568_1 = {c4514,s4541[1]};
    assign in4568_2 = {c4515,s4542[1]};
    CLA_2 KS_4568(s4568, c4568, in4568_1, in4568_2);
    wire[0:0] s4569, in4569_1, in4569_2;
    wire c4569;
    assign in4569_1 = {c4516};
    assign in4569_2 = {c4517};
    Half_Adder KS_4569(s4569, c4569, in4569_1, in4569_2);
    wire[2:0] s4570, in4570_1, in4570_2;
    wire c4570;
    assign in4570_1 = {c4518,s4543[1],c2942};
    assign in4570_2 = {c4519,s4544[1],s2943[1]};
    CLA_3 KS_4570(s4570, c4570, in4570_1, in4570_2);
    wire[0:0] s4571, in4571_1, in4571_2;
    wire c4571;
    assign in4571_1 = {c4524};
    assign in4571_2 = {c4532};
    Half_Adder KS_4571(s4571, c4571, in4571_1, in4571_2);
    wire[1:0] s4572, in4572_1, in4572_2;
    wire c4572;
    assign in4572_1 = {s4540[0],s4545[1]};
    assign in4572_2 = {s4541[0],s4546[1]};
    CLA_2 KS_4572(s4572, c4572, in4572_1, in4572_2);
    wire[0:0] s4573, in4573_1, in4573_2;
    wire c4573;
    assign in4573_1 = {s4542[0]};
    assign in4573_2 = {s4543[0]};
    Half_Adder KS_4573(s4573, c4573, in4573_1, in4573_2);
    wire[3:0] s4574, in4574_1, in4574_2;
    wire c4574;
    assign in4574_1 = {s4544[0],s4547[1],c2944,c2935};
    assign in4574_2 = {s4545[0],s4548[1],s4540[2],s2937[2]};
    CLA_4 KS_4574(s4574, c4574, in4574_1, in4574_2);
    wire[0:0] s4575, in4575_1, in4575_2;
    wire c4575;
    assign in4575_1 = {s4547[0]};
    assign in4575_2 = {s4548[0]};
    Full_Adder KS_4575(s4575, c4575, in4575_1, in4575_2, s4546[0]);
    wire[3:0] s4576, in4576_1, in4576_2;
    wire c4576;
    assign in4576_1 = {s1289[0],s2964[0],s2965[1],s2949[2]};
    assign in4576_2 = {s1290[0],s2965[0],s2966[1],s2950[2]};
    CLA_4 KS_4576(s4576, c4576, in4576_1, in4576_2);
    wire[3:0] s4577, in4577_1, in4577_2;
    wire c4577;
    assign in4577_1 = {s1291[0],s2966[0],s2967[1],s2951[2]};
    assign in4577_2 = {s1292[0],s2967[0],s2968[1],s2952[2]};
    CLA_4 KS_4577(s4577, c4577, in4577_1, in4577_2);
    wire[3:0] s4578, in4578_1, in4578_2;
    wire c4578;
    assign in4578_1 = {s1293[0],s2968[0],s2969[1],s2953[2]};
    assign in4578_2 = {s1294[0],s2969[0],s2970[1],s2954[2]};
    CLA_4 KS_4578(s4578, c4578, in4578_1, in4578_2);
    wire[3:0] s4579, in4579_1, in4579_2;
    wire c4579;
    assign in4579_1 = {s2880[3],s2970[0],s2971[1],s2955[2]};
    assign in4579_2 = {s2881[3],s2971[0],s2972[1],s2956[2]};
    CLA_4 KS_4579(s4579, c4579, in4579_1, in4579_2);
    wire[3:0] s4580, in4580_1, in4580_2;
    wire c4580;
    assign in4580_1 = {s2882[3],s2972[0],s2973[1],s2957[2]};
    assign in4580_2 = {s2883[3],s2973[0],s2974[1],s2958[2]};
    CLA_4 KS_4580(s4580, c4580, in4580_1, in4580_2);
    wire[3:0] s4581, in4581_1, in4581_2;
    wire c4581;
    assign in4581_1 = {s2884[3],s2974[0],s2975[1],s2959[2]};
    assign in4581_2 = {s2885[3],s2975[0],s2976[1],s2960[2]};
    CLA_4 KS_4581(s4581, c4581, in4581_1, in4581_2);
    wire[3:0] s4582, in4582_1, in4582_2;
    wire c4582;
    assign in4582_1 = {s2886[3],s2976[0],c2977,s2961[2]};
    assign in4582_2 = {s2887[3],s2977[0],s2978[1],s2962[2]};
    CLA_4 KS_4582(s4582, c4582, in4582_1, in4582_2);
    wire[3:0] s4583, in4583_1, in4583_2;
    wire c4583;
    assign in4583_1 = {s2888[3],s2978[0],c2979,s2963[2]};
    assign in4583_2 = {s2889[3],s2979[0],s2980[1],s2964[2]};
    CLA_4 KS_4583(s4583, c4583, in4583_1, in4583_2);
    wire[3:0] s4584, in4584_1, in4584_2;
    wire c4584;
    assign in4584_1 = {s2890[3],s2980[0],c2981,s2965[2]};
    assign in4584_2 = {s2891[3],s2981[0],s2982[1],s2966[2]};
    CLA_4 KS_4584(s4584, c4584, in4584_1, in4584_2);
    wire[3:0] s4585, in4585_1, in4585_2;
    wire c4585;
    assign in4585_1 = {s2892[3],s2982[0],c2983,s2967[2]};
    assign in4585_2 = {s2893[3],s2983[0],s2984[1],s2968[2]};
    CLA_4 KS_4585(s4585, c4585, in4585_1, in4585_2);
    wire[3:0] s4586, in4586_1, in4586_2;
    wire c4586;
    assign in4586_1 = {s2894[3],s2984[0],c2985,s2969[2]};
    assign in4586_2 = {s2895[3],s2985[0],s2986[1],s2970[2]};
    CLA_4 KS_4586(s4586, c4586, in4586_1, in4586_2);
    wire[3:0] s4587, in4587_1, in4587_2;
    wire c4587;
    assign in4587_1 = {s2896[3],s2986[0],c2987,s2971[2]};
    assign in4587_2 = {s2897[3],s2987[0],s2988[1],s2972[2]};
    CLA_4 KS_4587(s4587, c4587, in4587_1, in4587_2);
    wire[3:0] s4588, in4588_1, in4588_2;
    wire c4588;
    assign in4588_1 = {s2898[3],s2988[0],c2989,s2973[2]};
    assign in4588_2 = {s2899[3],s2989[0],s2990[1],s2974[2]};
    CLA_4 KS_4588(s4588, c4588, in4588_1, in4588_2);
    wire[3:0] s4589, in4589_1, in4589_2;
    wire c4589;
    assign in4589_1 = {s2900[3],s2990[0],c2991,s2975[2]};
    assign in4589_2 = {s2901[3],s2991[0],s2992[1],s2976[2]};
    CLA_4 KS_4589(s4589, c4589, in4589_1, in4589_2);
    wire[3:0] s4590, in4590_1, in4590_2;
    wire c4590;
    assign in4590_1 = {s2902[3],s2992[0],c2993,c2978};
    assign in4590_2 = {s2903[3],s2993[0],s2994[1],s2980[2]};
    CLA_4 KS_4590(s4590, c4590, in4590_1, in4590_2);
    wire[3:0] s4591, in4591_1, in4591_2;
    wire c4591;
    assign in4591_1 = {s2904[3],s2994[0],c2995,c2982};
    assign in4591_2 = {s2905[3],s2995[0],s2996[1],s2984[2]};
    CLA_4 KS_4591(s4591, c4591, in4591_1, in4591_2);
    wire[3:0] s4592, in4592_1, in4592_2;
    wire c4592;
    assign in4592_1 = {s2906[3],s2996[0],c2997,c2986};
    assign in4592_2 = {s2907[3],s2997[0],s2998[1],s2988[2]};
    CLA_4 KS_4592(s4592, c4592, in4592_1, in4592_2);
    wire[3:0] s4593, in4593_1, in4593_2;
    wire c4593;
    assign in4593_1 = {s2908[3],s2998[0],c2999,c2990};
    assign in4593_2 = {s2909[3],s2999[0],s3000[1],s2992[2]};
    CLA_4 KS_4593(s4593, c4593, in4593_1, in4593_2);
    wire[1:0] s4594, in4594_1, in4594_2;
    wire c4594;
    assign in4594_1 = {s2910[3],s3000[0]};
    assign in4594_2 = {s2913[3],s3001[0]};
    CLA_2 KS_4594(s4594, c4594, in4594_1, in4594_2);
    wire[0:0] s4595, in4595_1, in4595_2;
    wire c4595;
    assign in4595_1 = {c2917};
    assign in4595_2 = {s2921[3]};
    Half_Adder KS_4595(s4595, c4595, in4595_1, in4595_2);
    wire[2:0] s4596, in4596_1, in4596_2;
    wire c4596;
    assign in4596_1 = {c2925,s3002[0],c3001};
    assign in4596_2 = {s2929[3],s3003[0],s3002[1]};
    CLA_3 KS_4596(s4596, c4596, in4596_1, in4596_2);
    wire[0:0] s4597, in4597_1, in4597_2;
    wire c4597;
    assign in4597_1 = {c2933};
    assign in4597_2 = {s2937[3]};
    Half_Adder KS_4597(s4597, c4597, in4597_1, in4597_2);
    wire[1:0] s4598, in4598_1, in4598_2;
    wire c4598;
    assign in4598_1 = {c2941,s3004[0]};
    assign in4598_2 = {c4540,s3005[0]};
    CLA_2 KS_4598(s4598, c4598, in4598_1, in4598_2);
    wire[0:0] s4599, in4599_1, in4599_2;
    wire c4599;
    assign in4599_1 = {c4541};
    assign in4599_2 = {c4542};
    Half_Adder KS_4599(s4599, c4599, in4599_1, in4599_2);
    wire[3:0] s4600, in4600_1, in4600_2;
    wire c4600;
    assign in4600_1 = {c4543,s3006[0],c3003,c2994};
    assign in4600_2 = {c4544,s3007[0],s3004[1],s2996[2]};
    CLA_4 KS_4600(s4600, c4600, in4600_1, in4600_2);
    wire[0:0] s4601, in4601_1, in4601_2;
    wire c4601;
    assign in4601_1 = {c4545};
    assign in4601_2 = {c4546};
    Half_Adder KS_4601(s4601, c4601, in4601_1, in4601_2);
    wire[1:0] s4602, in4602_1, in4602_2;
    wire c4602;
    assign in4602_1 = {c4547,s3008[0]};
    assign in4602_2 = {c4548,s4576[1]};
    CLA_2 KS_4602(s4602, c4602, in4602_1, in4602_2);
    wire[0:0] s4603, in4603_1, in4603_2;
    wire c4603;
    assign in4603_1 = {c4549};
    assign in4603_2 = {c4550};
    Half_Adder KS_4603(s4603, c4603, in4603_1, in4603_2);
    wire[2:0] s4604, in4604_1, in4604_2;
    wire c4604;
    assign in4604_1 = {c4551,s4577[1],c3005};
    assign in4604_2 = {c4552,s4578[1],s3006[1]};
    CLA_3 KS_4604(s4604, c4604, in4604_1, in4604_2);
    wire[0:0] s4605, in4605_1, in4605_2;
    wire c4605;
    assign in4605_1 = {c4553};
    assign in4605_2 = {c4554};
    Half_Adder KS_4605(s4605, c4605, in4605_1, in4605_2);
    wire[1:0] s4606, in4606_1, in4606_2;
    wire c4606;
    assign in4606_1 = {c4555,s4579[1]};
    assign in4606_2 = {c4556,s4580[1]};
    CLA_2 KS_4606(s4606, c4606, in4606_1, in4606_2);
    wire[0:0] s4607, in4607_1, in4607_2;
    wire c4607;
    assign in4607_1 = {c4557};
    assign in4607_2 = {c4558};
    Half_Adder KS_4607(s4607, c4607, in4607_1, in4607_2);
    wire[3:0] s4608, in4608_1, in4608_2;
    wire c4608;
    assign in4608_1 = {c4566,s4581[1],c3007,c2998};
    assign in4608_2 = {c4574,s4582[1],s3008[1],s3000[2]};
    CLA_4 KS_4608(s4608, c4608, in4608_1, in4608_2);
    wire[0:0] s4609, in4609_1, in4609_2;
    wire c4609;
    assign in4609_1 = {s4576[0]};
    assign in4609_2 = {s4577[0]};
    Half_Adder KS_4609(s4609, c4609, in4609_1, in4609_2);
    wire[1:0] s4610, in4610_1, in4610_2;
    wire c4610;
    assign in4610_1 = {s4578[0],s4583[1]};
    assign in4610_2 = {s4579[0],s4584[1]};
    CLA_2 KS_4610(s4610, c4610, in4610_1, in4610_2);
    wire[0:0] s4611, in4611_1, in4611_2;
    wire c4611;
    assign in4611_1 = {s4580[0]};
    assign in4611_2 = {s4581[0]};
    Half_Adder KS_4611(s4611, c4611, in4611_1, in4611_2);
    wire[2:0] s4612, in4612_1, in4612_2;
    wire c4612;
    assign in4612_1 = {s4582[0],s4585[1],s4576[2]};
    assign in4612_2 = {s4583[0],s4586[1],s4577[2]};
    CLA_3 KS_4612(s4612, c4612, in4612_1, in4612_2);
    wire[0:0] s4613, in4613_1, in4613_2;
    wire c4613;
    assign in4613_1 = {s4585[0]};
    assign in4613_2 = {s4586[0]};
    Full_Adder KS_4613(s4613, c4613, in4613_1, in4613_2, s4584[0]);
    wire[3:0] s4614, in4614_1, in4614_2;
    wire c4614;
    assign in4614_1 = {s1310[0],s3030[0],s3030[1],s3012[2]};
    assign in4614_2 = {s1311[0],s3031[0],s3031[1],s3013[2]};
    CLA_4 KS_4614(s4614, c4614, in4614_1, in4614_2);
    wire[3:0] s4615, in4615_1, in4615_2;
    wire c4615;
    assign in4615_1 = {s1312[0],s3032[0],s3032[1],s3014[2]};
    assign in4615_2 = {s1313[0],s3033[0],s3033[1],s3015[2]};
    CLA_4 KS_4615(s4615, c4615, in4615_1, in4615_2);
    wire[3:0] s4616, in4616_1, in4616_2;
    wire c4616;
    assign in4616_1 = {s2945[3],s3034[0],s3034[1],s3016[2]};
    assign in4616_2 = {s2946[3],s3035[0],s3035[1],s3017[2]};
    CLA_4 KS_4616(s4616, c4616, in4616_1, in4616_2);
    wire[3:0] s4617, in4617_1, in4617_2;
    wire c4617;
    assign in4617_1 = {s2947[3],s3036[0],s3036[1],s3018[2]};
    assign in4617_2 = {s2948[3],s3037[0],s3037[1],s3019[2]};
    CLA_4 KS_4617(s4617, c4617, in4617_1, in4617_2);
    wire[3:0] s4618, in4618_1, in4618_2;
    wire c4618;
    assign in4618_1 = {s2949[3],s3038[0],s3038[1],s3020[2]};
    assign in4618_2 = {s2950[3],s3039[0],s3039[1],s3021[2]};
    CLA_4 KS_4618(s4618, c4618, in4618_1, in4618_2);
    wire[3:0] s4619, in4619_1, in4619_2;
    wire c4619;
    assign in4619_1 = {s2951[3],s3040[0],c3040,s3022[2]};
    assign in4619_2 = {s2952[3],s3041[0],s3041[1],s3023[2]};
    CLA_4 KS_4619(s4619, c4619, in4619_1, in4619_2);
    wire[3:0] s4620, in4620_1, in4620_2;
    wire c4620;
    assign in4620_1 = {s2953[3],s3042[0],c3042,s3024[2]};
    assign in4620_2 = {s2954[3],s3043[0],s3043[1],s3025[2]};
    CLA_4 KS_4620(s4620, c4620, in4620_1, in4620_2);
    wire[3:0] s4621, in4621_1, in4621_2;
    wire c4621;
    assign in4621_1 = {s2955[3],s3044[0],c3044,s3026[2]};
    assign in4621_2 = {s2956[3],s3045[0],s3045[1],s3027[2]};
    CLA_4 KS_4621(s4621, c4621, in4621_1, in4621_2);
    wire[3:0] s4622, in4622_1, in4622_2;
    wire c4622;
    assign in4622_1 = {s2957[3],s3046[0],c3046,s3028[2]};
    assign in4622_2 = {s2958[3],s3047[0],s3047[1],s3029[2]};
    CLA_4 KS_4622(s4622, c4622, in4622_1, in4622_2);
    wire[3:0] s4623, in4623_1, in4623_2;
    wire c4623;
    assign in4623_1 = {s2959[3],s3048[0],c3048,s3030[2]};
    assign in4623_2 = {s2960[3],s3049[0],s3049[1],s3031[2]};
    CLA_4 KS_4623(s4623, c4623, in4623_1, in4623_2);
    wire[3:0] s4624, in4624_1, in4624_2;
    wire c4624;
    assign in4624_1 = {s2961[3],s3050[0],c3050,s3032[2]};
    assign in4624_2 = {s2962[3],s3051[0],s3051[1],s3033[2]};
    CLA_4 KS_4624(s4624, c4624, in4624_1, in4624_2);
    wire[3:0] s4625, in4625_1, in4625_2;
    wire c4625;
    assign in4625_1 = {s2963[3],s3052[0],c3052,s3034[2]};
    assign in4625_2 = {s2964[3],s3053[0],s3053[1],s3035[2]};
    CLA_4 KS_4625(s4625, c4625, in4625_1, in4625_2);
    wire[3:0] s4626, in4626_1, in4626_2;
    wire c4626;
    assign in4626_1 = {s2965[3],s3054[0],c3054,s3036[2]};
    assign in4626_2 = {s2966[3],s3055[0],s3055[1],s3037[2]};
    CLA_4 KS_4626(s4626, c4626, in4626_1, in4626_2);
    wire[3:0] s4627, in4627_1, in4627_2;
    wire c4627;
    assign in4627_1 = {s2967[3],s3056[0],c3056,s3038[2]};
    assign in4627_2 = {s2968[3],s3057[0],s3057[1],s3039[2]};
    CLA_4 KS_4627(s4627, c4627, in4627_1, in4627_2);
    wire[3:0] s4628, in4628_1, in4628_2;
    wire c4628;
    assign in4628_1 = {s2969[3],s3058[0],c3058,c3041};
    assign in4628_2 = {s2970[3],s3059[0],s3059[1],s3043[2]};
    CLA_4 KS_4628(s4628, c4628, in4628_1, in4628_2);
    wire[3:0] s4629, in4629_1, in4629_2;
    wire c4629;
    assign in4629_1 = {s2971[3],s3060[0],c3060,c3045};
    assign in4629_2 = {s2972[3],s3061[0],s3061[1],s3047[2]};
    CLA_4 KS_4629(s4629, c4629, in4629_1, in4629_2);
    wire[3:0] s4630, in4630_1, in4630_2;
    wire c4630;
    assign in4630_1 = {s2973[3],s3062[0],c3062,c3049};
    assign in4630_2 = {s2974[3],s3063[0],s3063[1],s3051[2]};
    CLA_4 KS_4630(s4630, c4630, in4630_1, in4630_2);
    wire[3:0] s4631, in4631_1, in4631_2;
    wire c4631;
    assign in4631_1 = {s2975[3],s3064[0],c3064,c3053};
    assign in4631_2 = {s2976[3],s3065[0],s3065[1],s3055[2]};
    CLA_4 KS_4631(s4631, c4631, in4631_1, in4631_2);
    wire[3:0] s4632, in4632_1, in4632_2;
    wire c4632;
    assign in4632_1 = {c2980,s3066[0],c3066,c3057};
    assign in4632_2 = {s2984[3],s3067[0],s3067[1],s3059[2]};
    CLA_4 KS_4632(s4632, c4632, in4632_1, in4632_2);
    wire[0:0] s4633, in4633_1, in4633_2;
    wire c4633;
    assign in4633_1 = {c2988};
    assign in4633_2 = {s2992[3]};
    Half_Adder KS_4633(s4633, c4633, in4633_1, in4633_2);
    wire[1:0] s4634, in4634_1, in4634_2;
    wire c4634;
    assign in4634_1 = {c2996,s3068[0]};
    assign in4634_2 = {s3000[3],s3069[0]};
    CLA_2 KS_4634(s4634, c4634, in4634_1, in4634_2);
    wire[0:0] s4635, in4635_1, in4635_2;
    wire c4635;
    assign in4635_1 = {c3004};
    assign in4635_2 = {s3008[3]};
    Half_Adder KS_4635(s4635, c4635, in4635_1, in4635_2);
    wire[2:0] s4636, in4636_1, in4636_2;
    wire c4636;
    assign in4636_1 = {c4576,s3070[0],c3068};
    assign in4636_2 = {c4577,s3071[0],s3069[1]};
    CLA_3 KS_4636(s4636, c4636, in4636_1, in4636_2);
    wire[0:0] s4637, in4637_1, in4637_2;
    wire c4637;
    assign in4637_1 = {c4578};
    assign in4637_2 = {c4579};
    Half_Adder KS_4637(s4637, c4637, in4637_1, in4637_2);
    wire[1:0] s4638, in4638_1, in4638_2;
    wire c4638;
    assign in4638_1 = {c4580,s3072[0]};
    assign in4638_2 = {c4581,s3073[0]};
    CLA_2 KS_4638(s4638, c4638, in4638_1, in4638_2);
    wire[0:0] s4639, in4639_1, in4639_2;
    wire c4639;
    assign in4639_1 = {c4582};
    assign in4639_2 = {c4583};
    Half_Adder KS_4639(s4639, c4639, in4639_1, in4639_2);
    wire[3:0] s4640, in4640_1, in4640_2;
    wire c4640;
    assign in4640_1 = {c4584,s3074[0],c3070,c3061};
    assign in4640_2 = {c4585,s4614[1],s3071[1],s3063[2]};
    CLA_4 KS_4640(s4640, c4640, in4640_1, in4640_2);
    wire[0:0] s4641, in4641_1, in4641_2;
    wire c4641;
    assign in4641_1 = {c4586};
    assign in4641_2 = {c4587};
    Half_Adder KS_4641(s4641, c4641, in4641_1, in4641_2);
    wire[1:0] s4642, in4642_1, in4642_2;
    wire c4642;
    assign in4642_1 = {c4588,s4615[1]};
    assign in4642_2 = {c4589,s4616[1]};
    CLA_2 KS_4642(s4642, c4642, in4642_1, in4642_2);
    wire[0:0] s4643, in4643_1, in4643_2;
    wire c4643;
    assign in4643_1 = {c4590};
    assign in4643_2 = {c4591};
    Half_Adder KS_4643(s4643, c4643, in4643_1, in4643_2);
    wire[2:0] s4644, in4644_1, in4644_2;
    wire c4644;
    assign in4644_1 = {c4592,s4617[1],c3072};
    assign in4644_2 = {c4593,s4618[1],s3073[1]};
    CLA_3 KS_4644(s4644, c4644, in4644_1, in4644_2);
    wire[0:0] s4645, in4645_1, in4645_2;
    wire c4645;
    assign in4645_1 = {c4600};
    assign in4645_2 = {c4608};
    Half_Adder KS_4645(s4645, c4645, in4645_1, in4645_2);
    wire[1:0] s4646, in4646_1, in4646_2;
    wire c4646;
    assign in4646_1 = {s4614[0],s4619[1]};
    assign in4646_2 = {s4615[0],s4620[1]};
    CLA_2 KS_4646(s4646, c4646, in4646_1, in4646_2);
    wire[0:0] s4647, in4647_1, in4647_2;
    wire c4647;
    assign in4647_1 = {s4616[0]};
    assign in4647_2 = {s4617[0]};
    Half_Adder KS_4647(s4647, c4647, in4647_1, in4647_2);
    wire[3:0] s4648, in4648_1, in4648_2;
    wire c4648;
    assign in4648_1 = {s4618[0],s4621[1],c3074,c3065};
    assign in4648_2 = {s4619[0],s4622[1],s4614[2],s3067[2]};
    CLA_4 KS_4648(s4648, c4648, in4648_1, in4648_2);
    wire[0:0] s4649, in4649_1, in4649_2;
    wire c4649;
    assign in4649_1 = {s4621[0]};
    assign in4649_2 = {s4622[0]};
    Full_Adder KS_4649(s4649, c4649, in4649_1, in4649_2, s4620[0]);
    wire[3:0] s4650, in4650_1, in4650_2;
    wire c4650;
    assign in4650_1 = {s1319[0],s3095[0],s3096[1],s3079[2]};
    assign in4650_2 = {s1320[0],s3096[0],s3097[1],s3080[2]};
    CLA_4 KS_4650(s4650, c4650, in4650_1, in4650_2);
    wire[3:0] s4651, in4651_1, in4651_2;
    wire c4651;
    assign in4651_1 = {s1321[0],s3097[0],s3098[1],s3081[2]};
    assign in4651_2 = {s1322[0],s3098[0],s3099[1],s3082[2]};
    CLA_4 KS_4651(s4651, c4651, in4651_1, in4651_2);
    wire[3:0] s4652, in4652_1, in4652_2;
    wire c4652;
    assign in4652_1 = {s1323[0],s3099[0],s3100[1],s3083[2]};
    assign in4652_2 = {s1324[0],s3100[0],s3101[1],s3084[2]};
    CLA_4 KS_4652(s4652, c4652, in4652_1, in4652_2);
    wire[3:0] s4653, in4653_1, in4653_2;
    wire c4653;
    assign in4653_1 = {s3009[3],s3101[0],s3102[1],s3085[2]};
    assign in4653_2 = {s3010[3],s3102[0],s3103[1],s3086[2]};
    CLA_4 KS_4653(s4653, c4653, in4653_1, in4653_2);
    wire[3:0] s4654, in4654_1, in4654_2;
    wire c4654;
    assign in4654_1 = {s3011[3],s3103[0],s3104[1],s3087[2]};
    assign in4654_2 = {s3012[3],s3104[0],s3105[1],s3088[2]};
    CLA_4 KS_4654(s4654, c4654, in4654_1, in4654_2);
    wire[3:0] s4655, in4655_1, in4655_2;
    wire c4655;
    assign in4655_1 = {s3013[3],s3105[0],c3106,s3089[2]};
    assign in4655_2 = {s3014[3],s3106[0],s3107[1],s3090[2]};
    CLA_4 KS_4655(s4655, c4655, in4655_1, in4655_2);
    wire[3:0] s4656, in4656_1, in4656_2;
    wire c4656;
    assign in4656_1 = {s3015[3],s3107[0],c3108,s3091[2]};
    assign in4656_2 = {s3016[3],s3108[0],s3109[1],s3092[2]};
    CLA_4 KS_4656(s4656, c4656, in4656_1, in4656_2);
    wire[3:0] s4657, in4657_1, in4657_2;
    wire c4657;
    assign in4657_1 = {s3017[3],s3109[0],c3110,s3093[2]};
    assign in4657_2 = {s3018[3],s3110[0],s3111[1],s3094[2]};
    CLA_4 KS_4657(s4657, c4657, in4657_1, in4657_2);
    wire[3:0] s4658, in4658_1, in4658_2;
    wire c4658;
    assign in4658_1 = {s3019[3],s3111[0],c3112,s3095[2]};
    assign in4658_2 = {s3020[3],s3112[0],s3113[1],s3096[2]};
    CLA_4 KS_4658(s4658, c4658, in4658_1, in4658_2);
    wire[3:0] s4659, in4659_1, in4659_2;
    wire c4659;
    assign in4659_1 = {s3021[3],s3113[0],c3114,s3097[2]};
    assign in4659_2 = {s3022[3],s3114[0],s3115[1],s3098[2]};
    CLA_4 KS_4659(s4659, c4659, in4659_1, in4659_2);
    wire[3:0] s4660, in4660_1, in4660_2;
    wire c4660;
    assign in4660_1 = {s3023[3],s3115[0],c3116,s3099[2]};
    assign in4660_2 = {s3024[3],s3116[0],s3117[1],s3100[2]};
    CLA_4 KS_4660(s4660, c4660, in4660_1, in4660_2);
    wire[3:0] s4661, in4661_1, in4661_2;
    wire c4661;
    assign in4661_1 = {s3025[3],s3117[0],c3118,s3101[2]};
    assign in4661_2 = {s3026[3],s3118[0],s3119[1],s3102[2]};
    CLA_4 KS_4661(s4661, c4661, in4661_1, in4661_2);
    wire[3:0] s4662, in4662_1, in4662_2;
    wire c4662;
    assign in4662_1 = {s3027[3],s3119[0],c3120,s3103[2]};
    assign in4662_2 = {s3028[3],s3120[0],s3121[1],s3104[2]};
    CLA_4 KS_4662(s4662, c4662, in4662_1, in4662_2);
    wire[3:0] s4663, in4663_1, in4663_2;
    wire c4663;
    assign in4663_1 = {s3029[3],s3121[0],c3122,s3105[2]};
    assign in4663_2 = {s3030[3],s3122[0],s3123[1],s3107[2]};
    CLA_4 KS_4663(s4663, c4663, in4663_1, in4663_2);
    wire[3:0] s4664, in4664_1, in4664_2;
    wire c4664;
    assign in4664_1 = {s3031[3],s3123[0],c3124,c3109};
    assign in4664_2 = {s3032[3],s3124[0],s3125[1],s3111[2]};
    CLA_4 KS_4664(s4664, c4664, in4664_1, in4664_2);
    wire[3:0] s4665, in4665_1, in4665_2;
    wire c4665;
    assign in4665_1 = {s3033[3],s3125[0],c3126,c3113};
    assign in4665_2 = {s3034[3],s3126[0],s3127[1],s3115[2]};
    CLA_4 KS_4665(s4665, c4665, in4665_1, in4665_2);
    wire[3:0] s4666, in4666_1, in4666_2;
    wire c4666;
    assign in4666_1 = {s3035[3],s3127[0],c3128,c3117};
    assign in4666_2 = {s3036[3],s3128[0],s3129[1],s3119[2]};
    CLA_4 KS_4666(s4666, c4666, in4666_1, in4666_2);
    wire[3:0] s4667, in4667_1, in4667_2;
    wire c4667;
    assign in4667_1 = {s3037[3],s3129[0],c3130,c3121};
    assign in4667_2 = {s3038[3],s3130[0],s3131[1],s3123[2]};
    CLA_4 KS_4667(s4667, c4667, in4667_1, in4667_2);
    wire[1:0] s4668, in4668_1, in4668_2;
    wire c4668;
    assign in4668_1 = {s3039[3],s3131[0]};
    assign in4668_2 = {s3043[3],s3132[0]};
    CLA_2 KS_4668(s4668, c4668, in4668_1, in4668_2);
    wire[0:0] s4669, in4669_1, in4669_2;
    wire c4669;
    assign in4669_1 = {c3047};
    assign in4669_2 = {s3051[3]};
    Half_Adder KS_4669(s4669, c4669, in4669_1, in4669_2);
    wire[2:0] s4670, in4670_1, in4670_2;
    wire c4670;
    assign in4670_1 = {c3055,s3133[0],c3132};
    assign in4670_2 = {s3059[3],s3134[0],s3133[1]};
    CLA_3 KS_4670(s4670, c4670, in4670_1, in4670_2);
    wire[0:0] s4671, in4671_1, in4671_2;
    wire c4671;
    assign in4671_1 = {c3063};
    assign in4671_2 = {s3067[3]};
    Half_Adder KS_4671(s4671, c4671, in4671_1, in4671_2);
    wire[1:0] s4672, in4672_1, in4672_2;
    wire c4672;
    assign in4672_1 = {c3071,s3135[0]};
    assign in4672_2 = {c4614,s3136[0]};
    CLA_2 KS_4672(s4672, c4672, in4672_1, in4672_2);
    wire[0:0] s4673, in4673_1, in4673_2;
    wire c4673;
    assign in4673_1 = {c4615};
    assign in4673_2 = {c4616};
    Half_Adder KS_4673(s4673, c4673, in4673_1, in4673_2);
    wire[3:0] s4674, in4674_1, in4674_2;
    wire c4674;
    assign in4674_1 = {c4617,s3137[0],c3134,c3125};
    assign in4674_2 = {c4618,s3138[0],s3135[1],s3127[2]};
    CLA_4 KS_4674(s4674, c4674, in4674_1, in4674_2);
    wire[0:0] s4675, in4675_1, in4675_2;
    wire c4675;
    assign in4675_1 = {c4619};
    assign in4675_2 = {c4620};
    Half_Adder KS_4675(s4675, c4675, in4675_1, in4675_2);
    wire[1:0] s4676, in4676_1, in4676_2;
    wire c4676;
    assign in4676_1 = {c4621,s3139[0]};
    assign in4676_2 = {c4622,s4650[1]};
    CLA_2 KS_4676(s4676, c4676, in4676_1, in4676_2);
    wire[0:0] s4677, in4677_1, in4677_2;
    wire c4677;
    assign in4677_1 = {c4623};
    assign in4677_2 = {c4624};
    Half_Adder KS_4677(s4677, c4677, in4677_1, in4677_2);
    wire[2:0] s4678, in4678_1, in4678_2;
    wire c4678;
    assign in4678_1 = {c4625,s4651[1],c3136};
    assign in4678_2 = {c4626,s4652[1],s3137[1]};
    CLA_3 KS_4678(s4678, c4678, in4678_1, in4678_2);
    wire[0:0] s4679, in4679_1, in4679_2;
    wire c4679;
    assign in4679_1 = {c4627};
    assign in4679_2 = {c4628};
    Half_Adder KS_4679(s4679, c4679, in4679_1, in4679_2);
    wire[1:0] s4680, in4680_1, in4680_2;
    wire c4680;
    assign in4680_1 = {c4629,s4653[1]};
    assign in4680_2 = {c4630,s4654[1]};
    CLA_2 KS_4680(s4680, c4680, in4680_1, in4680_2);
    wire[0:0] s4681, in4681_1, in4681_2;
    wire c4681;
    assign in4681_1 = {c4631};
    assign in4681_2 = {c4632};
    Half_Adder KS_4681(s4681, c4681, in4681_1, in4681_2);
    wire[3:0] s4682, in4682_1, in4682_2;
    wire c4682;
    assign in4682_1 = {c4640,s4655[1],c3138,c3129};
    assign in4682_2 = {c4648,s4656[1],s3139[1],s3131[2]};
    CLA_4 KS_4682(s4682, c4682, in4682_1, in4682_2);
    wire[0:0] s4683, in4683_1, in4683_2;
    wire c4683;
    assign in4683_1 = {s4650[0]};
    assign in4683_2 = {s4651[0]};
    Half_Adder KS_4683(s4683, c4683, in4683_1, in4683_2);
    wire[1:0] s4684, in4684_1, in4684_2;
    wire c4684;
    assign in4684_1 = {s4652[0],s4657[1]};
    assign in4684_2 = {s4653[0],s4658[1]};
    CLA_2 KS_4684(s4684, c4684, in4684_1, in4684_2);
    wire[0:0] s4685, in4685_1, in4685_2;
    wire c4685;
    assign in4685_1 = {s4654[0]};
    assign in4685_2 = {s4655[0]};
    Half_Adder KS_4685(s4685, c4685, in4685_1, in4685_2);
    wire[2:0] s4686, in4686_1, in4686_2;
    wire c4686;
    assign in4686_1 = {s4656[0],s4659[1],s4650[2]};
    assign in4686_2 = {s4657[0],s4660[1],s4651[2]};
    CLA_3 KS_4686(s4686, c4686, in4686_1, in4686_2);
    wire[0:0] s4687, in4687_1, in4687_2;
    wire c4687;
    assign in4687_1 = {s4659[0]};
    assign in4687_2 = {s4660[0]};
    Full_Adder KS_4687(s4687, c4687, in4687_1, in4687_2, s4658[0]);
    wire[3:0] s4688, in4688_1, in4688_2;
    wire c4688;
    assign in4688_1 = {c1315,s3160[0],s3161[1],s3143[2]};
    assign in4688_2 = {c1319,s3161[0],s3162[1],s3144[2]};
    CLA_4 KS_4688(s4688, c4688, in4688_1, in4688_2);
    wire[3:0] s4689, in4689_1, in4689_2;
    wire c4689;
    assign in4689_1 = {s1325[0],s3162[0],s3163[1],s3145[2]};
    assign in4689_2 = {s1326[0],s3163[0],s3164[1],s3146[2]};
    CLA_4 KS_4689(s4689, c4689, in4689_1, in4689_2);
    wire[3:0] s4690, in4690_1, in4690_2;
    wire c4690;
    assign in4690_1 = {s3075[3],s3164[0],s3165[1],s3147[2]};
    assign in4690_2 = {s3076[3],s3165[0],s3166[1],s3148[2]};
    CLA_4 KS_4690(s4690, c4690, in4690_1, in4690_2);
    wire[3:0] s4691, in4691_1, in4691_2;
    wire c4691;
    assign in4691_1 = {s3077[3],s3166[0],s3167[1],s3149[2]};
    assign in4691_2 = {s3078[3],s3167[0],s3168[1],s3150[2]};
    CLA_4 KS_4691(s4691, c4691, in4691_1, in4691_2);
    wire[3:0] s4692, in4692_1, in4692_2;
    wire c4692;
    assign in4692_1 = {s3079[3],s3168[0],s3169[1],s3151[2]};
    assign in4692_2 = {s3080[3],s3169[0],s3170[1],s3152[2]};
    CLA_4 KS_4692(s4692, c4692, in4692_1, in4692_2);
    wire[3:0] s4693, in4693_1, in4693_2;
    wire c4693;
    assign in4693_1 = {s3081[3],s3170[0],c3171,s3153[2]};
    assign in4693_2 = {s3082[3],s3171[0],s3172[1],s3154[2]};
    CLA_4 KS_4693(s4693, c4693, in4693_1, in4693_2);
    wire[3:0] s4694, in4694_1, in4694_2;
    wire c4694;
    assign in4694_1 = {s3083[3],s3172[0],c3173,s3155[2]};
    assign in4694_2 = {s3084[3],s3173[0],s3174[1],s3156[2]};
    CLA_4 KS_4694(s4694, c4694, in4694_1, in4694_2);
    wire[3:0] s4695, in4695_1, in4695_2;
    wire c4695;
    assign in4695_1 = {s3085[3],s3174[0],c3175,s3157[2]};
    assign in4695_2 = {s3086[3],s3175[0],s3176[1],s3158[2]};
    CLA_4 KS_4695(s4695, c4695, in4695_1, in4695_2);
    wire[3:0] s4696, in4696_1, in4696_2;
    wire c4696;
    assign in4696_1 = {s3087[3],s3176[0],c3177,s3159[2]};
    assign in4696_2 = {s3088[3],s3177[0],s3178[1],s3160[2]};
    CLA_4 KS_4696(s4696, c4696, in4696_1, in4696_2);
    wire[3:0] s4697, in4697_1, in4697_2;
    wire c4697;
    assign in4697_1 = {s3089[3],s3178[0],c3179,s3161[2]};
    assign in4697_2 = {s3090[3],s3179[0],s3180[1],s3162[2]};
    CLA_4 KS_4697(s4697, c4697, in4697_1, in4697_2);
    wire[3:0] s4698, in4698_1, in4698_2;
    wire c4698;
    assign in4698_1 = {s3091[3],s3180[0],c3181,s3163[2]};
    assign in4698_2 = {s3092[3],s3181[0],s3182[1],s3164[2]};
    CLA_4 KS_4698(s4698, c4698, in4698_1, in4698_2);
    wire[3:0] s4699, in4699_1, in4699_2;
    wire c4699;
    assign in4699_1 = {s3093[3],s3182[0],c3183,s3165[2]};
    assign in4699_2 = {s3094[3],s3183[0],s3184[1],s3166[2]};
    CLA_4 KS_4699(s4699, c4699, in4699_1, in4699_2);
    wire[3:0] s4700, in4700_1, in4700_2;
    wire c4700;
    assign in4700_1 = {s3095[3],s3184[0],c3185,s3167[2]};
    assign in4700_2 = {s3096[3],s3185[0],s3186[1],s3168[2]};
    CLA_4 KS_4700(s4700, c4700, in4700_1, in4700_2);
    wire[3:0] s4701, in4701_1, in4701_2;
    wire c4701;
    assign in4701_1 = {s3097[3],s3186[0],c3187,c3169};
    assign in4701_2 = {s3098[3],s3187[0],s3188[1],s3170[2]};
    CLA_4 KS_4701(s4701, c4701, in4701_1, in4701_2);
    wire[3:0] s4702, in4702_1, in4702_2;
    wire c4702;
    assign in4702_1 = {s3099[3],s3188[0],c3189,c3172};
    assign in4702_2 = {s3100[3],s3189[0],s3190[1],s3174[2]};
    CLA_4 KS_4702(s4702, c4702, in4702_1, in4702_2);
    wire[3:0] s4703, in4703_1, in4703_2;
    wire c4703;
    assign in4703_1 = {s3101[3],s3190[0],c3191,c3176};
    assign in4703_2 = {s3102[3],s3191[0],s3192[1],s3178[2]};
    CLA_4 KS_4703(s4703, c4703, in4703_1, in4703_2);
    wire[3:0] s4704, in4704_1, in4704_2;
    wire c4704;
    assign in4704_1 = {s3103[3],s3192[0],c3193,c3180};
    assign in4704_2 = {s3104[3],s3193[0],s3194[1],s3182[2]};
    CLA_4 KS_4704(s4704, c4704, in4704_1, in4704_2);
    wire[3:0] s4705, in4705_1, in4705_2;
    wire c4705;
    assign in4705_1 = {s3105[3],s3194[0],c3195,c3184};
    assign in4705_2 = {s3107[3],s3195[0],s3196[1],s3186[2]};
    CLA_4 KS_4705(s4705, c4705, in4705_1, in4705_2);
    wire[1:0] s4706, in4706_1, in4706_2;
    wire c4706;
    assign in4706_1 = {c3111,s3196[0]};
    assign in4706_2 = {s3115[3],s3197[0]};
    CLA_2 KS_4706(s4706, c4706, in4706_1, in4706_2);
    wire[0:0] s4707, in4707_1, in4707_2;
    wire c4707;
    assign in4707_1 = {c3119};
    assign in4707_2 = {s3123[3]};
    Half_Adder KS_4707(s4707, c4707, in4707_1, in4707_2);
    wire[3:0] s4708, in4708_1, in4708_2;
    wire c4708;
    assign in4708_1 = {c3127,s3198[0],c3197,c3188};
    assign in4708_2 = {s3131[3],s3199[0],s3198[1],s3190[2]};
    CLA_4 KS_4708(s4708, c4708, in4708_1, in4708_2);
    wire[0:0] s4709, in4709_1, in4709_2;
    wire c4709;
    assign in4709_1 = {c3135};
    assign in4709_2 = {s3139[3]};
    Half_Adder KS_4709(s4709, c4709, in4709_1, in4709_2);
    wire[1:0] s4710, in4710_1, in4710_2;
    wire c4710;
    assign in4710_1 = {c4650,s3200[0]};
    assign in4710_2 = {c4651,s3201[0]};
    CLA_2 KS_4710(s4710, c4710, in4710_1, in4710_2);
    wire[0:0] s4711, in4711_1, in4711_2;
    wire c4711;
    assign in4711_1 = {c4652};
    assign in4711_2 = {c4653};
    Half_Adder KS_4711(s4711, c4711, in4711_1, in4711_2);
    wire[2:0] s4712, in4712_1, in4712_2;
    wire c4712;
    assign in4712_1 = {c4654,s3202[0],c3199};
    assign in4712_2 = {c4655,s3203[0],s3200[1]};
    CLA_3 KS_4712(s4712, c4712, in4712_1, in4712_2);
    wire[0:0] s4713, in4713_1, in4713_2;
    wire c4713;
    assign in4713_1 = {c4656};
    assign in4713_2 = {c4657};
    Half_Adder KS_4713(s4713, c4713, in4713_1, in4713_2);
    wire[1:0] s4714, in4714_1, in4714_2;
    wire c4714;
    assign in4714_1 = {c4658,s3204[0]};
    assign in4714_2 = {c4659,s4688[1]};
    CLA_2 KS_4714(s4714, c4714, in4714_1, in4714_2);
    wire[0:0] s4715, in4715_1, in4715_2;
    wire c4715;
    assign in4715_1 = {c4660};
    assign in4715_2 = {c4661};
    Half_Adder KS_4715(s4715, c4715, in4715_1, in4715_2);
    wire[3:0] s4716, in4716_1, in4716_2;
    wire c4716;
    assign in4716_1 = {c4662,s4689[1],c3201,c3192};
    assign in4716_2 = {c4663,s4690[1],s3202[1],s3194[2]};
    CLA_4 KS_4716(s4716, c4716, in4716_1, in4716_2);
    wire[0:0] s4717, in4717_1, in4717_2;
    wire c4717;
    assign in4717_1 = {c4664};
    assign in4717_2 = {c4665};
    Half_Adder KS_4717(s4717, c4717, in4717_1, in4717_2);
    wire[1:0] s4718, in4718_1, in4718_2;
    wire c4718;
    assign in4718_1 = {c4666,s4691[1]};
    assign in4718_2 = {c4667,s4692[1]};
    CLA_2 KS_4718(s4718, c4718, in4718_1, in4718_2);
    wire[0:0] s4719, in4719_1, in4719_2;
    wire c4719;
    assign in4719_1 = {c4674};
    assign in4719_2 = {c4682};
    Half_Adder KS_4719(s4719, c4719, in4719_1, in4719_2);
    wire[2:0] s4720, in4720_1, in4720_2;
    wire c4720;
    assign in4720_1 = {s4688[0],s4693[1],c3203};
    assign in4720_2 = {s4689[0],s4694[1],s3204[1]};
    CLA_3 KS_4720(s4720, c4720, in4720_1, in4720_2);
    wire[0:0] s4721, in4721_1, in4721_2;
    wire c4721;
    assign in4721_1 = {s4690[0]};
    assign in4721_2 = {s4691[0]};
    Half_Adder KS_4721(s4721, c4721, in4721_1, in4721_2);
    wire[1:0] s4722, in4722_1, in4722_2;
    wire c4722;
    assign in4722_1 = {s4692[0],s4695[1]};
    assign in4722_2 = {s4693[0],s4696[1]};
    CLA_2 KS_4722(s4722, c4722, in4722_1, in4722_2);
    wire[0:0] s4723, in4723_1, in4723_2;
    wire c4723;
    assign in4723_1 = {s4695[0]};
    assign in4723_2 = {s4696[0]};
    Full_Adder KS_4723(s4723, c4723, in4723_1, in4723_2, s4694[0]);
    wire[3:0] s4724, in4724_1, in4724_2;
    wire c4724;
    assign in4724_1 = {pp122[61],s3218[0],s3219[1],pp125[61]};
    assign in4724_2 = {pp123[60],s3219[0],s3220[1],pp126[60]};
    CLA_4 KS_4724(s4724, c4724, in4724_1, in4724_2);
    wire[3:0] s4725, in4725_1, in4725_2;
    wire c4725;
    assign in4725_1 = {pp124[59],s3220[0],s3221[1],pp127[59]};
    assign in4725_2 = {pp125[58],s3221[0],s3222[1],s3205[2]};
    CLA_4 KS_4725(s4725, c4725, in4725_1, in4725_2);
    wire[3:0] s4726, in4726_1, in4726_2;
    wire c4726;
    assign in4726_1 = {pp126[57],s3222[0],s3223[1],s3206[2]};
    assign in4726_2 = {pp127[56],s3223[0],s3224[1],s3207[2]};
    CLA_4 KS_4726(s4726, c4726, in4726_1, in4726_2);
    wire[3:0] s4727, in4727_1, in4727_2;
    wire c4727;
    assign in4727_1 = {s3140[3],s3224[0],s3225[1],s3208[2]};
    assign in4727_2 = {s3141[3],s3225[0],s3226[1],s3209[2]};
    CLA_4 KS_4727(s4727, c4727, in4727_1, in4727_2);
    wire[3:0] s4728, in4728_1, in4728_2;
    wire c4728;
    assign in4728_1 = {s3142[3],s3226[0],s3227[1],s3210[2]};
    assign in4728_2 = {s3143[3],s3227[0],s3228[1],s3211[2]};
    CLA_4 KS_4728(s4728, c4728, in4728_1, in4728_2);
    wire[3:0] s4729, in4729_1, in4729_2;
    wire c4729;
    assign in4729_1 = {s3144[3],s3228[0],s3229[1],s3212[2]};
    assign in4729_2 = {s3145[3],s3229[0],s3230[1],s3213[2]};
    CLA_4 KS_4729(s4729, c4729, in4729_1, in4729_2);
    wire[3:0] s4730, in4730_1, in4730_2;
    wire c4730;
    assign in4730_1 = {s3146[3],s3230[0],c3231,s3214[2]};
    assign in4730_2 = {s3147[3],s3231[0],s3232[1],s3215[2]};
    CLA_4 KS_4730(s4730, c4730, in4730_1, in4730_2);
    wire[3:0] s4731, in4731_1, in4731_2;
    wire c4731;
    assign in4731_1 = {s3148[3],s3232[0],c3233,s3216[2]};
    assign in4731_2 = {s3149[3],s3233[0],s3234[1],s3217[2]};
    CLA_4 KS_4731(s4731, c4731, in4731_1, in4731_2);
    wire[3:0] s4732, in4732_1, in4732_2;
    wire c4732;
    assign in4732_1 = {s3150[3],s3234[0],c3235,s3218[2]};
    assign in4732_2 = {s3151[3],s3235[0],s3236[1],s3219[2]};
    CLA_4 KS_4732(s4732, c4732, in4732_1, in4732_2);
    wire[3:0] s4733, in4733_1, in4733_2;
    wire c4733;
    assign in4733_1 = {s3152[3],s3236[0],c3237,s3220[2]};
    assign in4733_2 = {s3153[3],s3237[0],s3238[1],s3221[2]};
    CLA_4 KS_4733(s4733, c4733, in4733_1, in4733_2);
    wire[3:0] s4734, in4734_1, in4734_2;
    wire c4734;
    assign in4734_1 = {s3154[3],s3238[0],c3239,s3222[2]};
    assign in4734_2 = {s3155[3],s3239[0],s3240[1],s3223[2]};
    CLA_4 KS_4734(s4734, c4734, in4734_1, in4734_2);
    wire[3:0] s4735, in4735_1, in4735_2;
    wire c4735;
    assign in4735_1 = {s3156[3],s3240[0],c3241,s3224[2]};
    assign in4735_2 = {s3157[3],s3241[0],s3242[1],s3225[2]};
    CLA_4 KS_4735(s4735, c4735, in4735_1, in4735_2);
    wire[3:0] s4736, in4736_1, in4736_2;
    wire c4736;
    assign in4736_1 = {s3158[3],s3242[0],c3243,s3226[2]};
    assign in4736_2 = {s3159[3],s3243[0],s3244[1],s3227[2]};
    CLA_4 KS_4736(s4736, c4736, in4736_1, in4736_2);
    wire[3:0] s4737, in4737_1, in4737_2;
    wire c4737;
    assign in4737_1 = {s3160[3],s3244[0],c3245,s3228[2]};
    assign in4737_2 = {s3161[3],s3245[0],s3246[1],s3229[2]};
    CLA_4 KS_4737(s4737, c4737, in4737_1, in4737_2);
    wire[3:0] s4738, in4738_1, in4738_2;
    wire c4738;
    assign in4738_1 = {s3162[3],s3246[0],c3247,c3230};
    assign in4738_2 = {s3163[3],s3247[0],s3248[1],s3232[2]};
    CLA_4 KS_4738(s4738, c4738, in4738_1, in4738_2);
    wire[3:0] s4739, in4739_1, in4739_2;
    wire c4739;
    assign in4739_1 = {s3164[3],s3248[0],c3249,c3234};
    assign in4739_2 = {s3165[3],s3249[0],s3250[1],s3236[2]};
    CLA_4 KS_4739(s4739, c4739, in4739_1, in4739_2);
    wire[3:0] s4740, in4740_1, in4740_2;
    wire c4740;
    assign in4740_1 = {s3166[3],s3250[0],c3251,c3238};
    assign in4740_2 = {s3167[3],s3251[0],s3252[1],s3240[2]};
    CLA_4 KS_4740(s4740, c4740, in4740_1, in4740_2);
    wire[3:0] s4741, in4741_1, in4741_2;
    wire c4741;
    assign in4741_1 = {c3168,s3252[0],c3253,c3242};
    assign in4741_2 = {s3170[3],s3253[0],s3254[1],s3244[2]};
    CLA_4 KS_4741(s4741, c4741, in4741_1, in4741_2);
    wire[1:0] s4742, in4742_1, in4742_2;
    wire c4742;
    assign in4742_1 = {c3174,s3254[0]};
    assign in4742_2 = {s3178[3],s3255[0]};
    CLA_2 KS_4742(s4742, c4742, in4742_1, in4742_2);
    wire[0:0] s4743, in4743_1, in4743_2;
    wire c4743;
    assign in4743_1 = {c3182};
    assign in4743_2 = {s3186[3]};
    Half_Adder KS_4743(s4743, c4743, in4743_1, in4743_2);
    wire[3:0] s4744, in4744_1, in4744_2;
    wire c4744;
    assign in4744_1 = {c3190,s3256[0],c3255,c3246};
    assign in4744_2 = {s3194[3],s3257[0],s3256[1],s3248[2]};
    CLA_4 KS_4744(s4744, c4744, in4744_1, in4744_2);
    wire[0:0] s4745, in4745_1, in4745_2;
    wire c4745;
    assign in4745_1 = {c3198};
    assign in4745_2 = {s3202[3]};
    Half_Adder KS_4745(s4745, c4745, in4745_1, in4745_2);
    wire[1:0] s4746, in4746_1, in4746_2;
    wire c4746;
    assign in4746_1 = {c4688,s3258[0]};
    assign in4746_2 = {c4689,s3259[0]};
    CLA_2 KS_4746(s4746, c4746, in4746_1, in4746_2);
    wire[0:0] s4747, in4747_1, in4747_2;
    wire c4747;
    assign in4747_1 = {c4690};
    assign in4747_2 = {c4691};
    Half_Adder KS_4747(s4747, c4747, in4747_1, in4747_2);
    wire[2:0] s4748, in4748_1, in4748_2;
    wire c4748;
    assign in4748_1 = {c4692,s3260[0],c3257};
    assign in4748_2 = {c4693,s3261[0],s3258[1]};
    CLA_3 KS_4748(s4748, c4748, in4748_1, in4748_2);
    wire[0:0] s4749, in4749_1, in4749_2;
    wire c4749;
    assign in4749_1 = {c4694};
    assign in4749_2 = {c4695};
    Half_Adder KS_4749(s4749, c4749, in4749_1, in4749_2);
    wire[1:0] s4750, in4750_1, in4750_2;
    wire c4750;
    assign in4750_1 = {c4696,s3262[0]};
    assign in4750_2 = {c4697,s4724[1]};
    CLA_2 KS_4750(s4750, c4750, in4750_1, in4750_2);
    wire[0:0] s4751, in4751_1, in4751_2;
    wire c4751;
    assign in4751_1 = {c4698};
    assign in4751_2 = {c4699};
    Half_Adder KS_4751(s4751, c4751, in4751_1, in4751_2);
    wire[3:0] s4752, in4752_1, in4752_2;
    wire c4752;
    assign in4752_1 = {c4700,s4725[1],c3259,c3250};
    assign in4752_2 = {c4701,s4726[1],s3260[1],s3252[2]};
    CLA_4 KS_4752(s4752, c4752, in4752_1, in4752_2);
    wire[0:0] s4753, in4753_1, in4753_2;
    wire c4753;
    assign in4753_1 = {c4702};
    assign in4753_2 = {c4703};
    Half_Adder KS_4753(s4753, c4753, in4753_1, in4753_2);
    wire[1:0] s4754, in4754_1, in4754_2;
    wire c4754;
    assign in4754_1 = {c4704,s4727[1]};
    assign in4754_2 = {c4705,s4728[1]};
    CLA_2 KS_4754(s4754, c4754, in4754_1, in4754_2);
    wire[0:0] s4755, in4755_1, in4755_2;
    wire c4755;
    assign in4755_1 = {c4708};
    assign in4755_2 = {c4716};
    Half_Adder KS_4755(s4755, c4755, in4755_1, in4755_2);
    wire[2:0] s4756, in4756_1, in4756_2;
    wire c4756;
    assign in4756_1 = {s4724[0],s4729[1],c3261};
    assign in4756_2 = {s4725[0],s4730[1],s3262[1]};
    CLA_3 KS_4756(s4756, c4756, in4756_1, in4756_2);
    wire[0:0] s4757, in4757_1, in4757_2;
    wire c4757;
    assign in4757_1 = {s4726[0]};
    assign in4757_2 = {s4727[0]};
    Half_Adder KS_4757(s4757, c4757, in4757_1, in4757_2);
    wire[1:0] s4758, in4758_1, in4758_2;
    wire c4758;
    assign in4758_1 = {s4728[0],s4731[1]};
    assign in4758_2 = {s4729[0],s4732[1]};
    CLA_2 KS_4758(s4758, c4758, in4758_1, in4758_2);
    wire[0:0] s4759, in4759_1, in4759_2;
    wire c4759;
    assign in4759_1 = {s4731[0]};
    assign in4759_2 = {s4732[0]};
    Full_Adder KS_4759(s4759, c4759, in4759_1, in4759_2, s4730[0]);
    wire[3:0] s4760, in4760_1, in4760_2;
    wire c4760;
    assign in4760_1 = {pp116[71],s3267[0],s3267[1],pp119[71]};
    assign in4760_2 = {pp117[70],s3268[0],s3268[1],pp120[70]};
    CLA_4 KS_4760(s4760, c4760, in4760_1, in4760_2);
    wire[3:0] s4761, in4761_1, in4761_2;
    wire c4761;
    assign in4761_1 = {pp118[69],s3269[0],s3269[1],pp121[69]};
    assign in4761_2 = {pp119[68],s3270[0],s3270[1],pp122[68]};
    CLA_4 KS_4761(s4761, c4761, in4761_1, in4761_2);
    wire[3:0] s4762, in4762_1, in4762_2;
    wire c4762;
    assign in4762_1 = {pp120[67],s3271[0],s3271[1],pp123[67]};
    assign in4762_2 = {pp121[66],s3272[0],s3272[1],pp124[66]};
    CLA_4 KS_4762(s4762, c4762, in4762_1, in4762_2);
    wire[3:0] s4763, in4763_1, in4763_2;
    wire c4763;
    assign in4763_1 = {pp122[65],s3273[0],s3273[1],pp125[65]};
    assign in4763_2 = {pp123[64],s3274[0],s3274[1],pp126[64]};
    CLA_4 KS_4763(s4763, c4763, in4763_1, in4763_2);
    wire[3:0] s4764, in4764_1, in4764_2;
    wire c4764;
    assign in4764_1 = {pp124[63],s3275[0],s3275[1],pp127[63]};
    assign in4764_2 = {pp125[62],s3276[0],s3276[1],s3263[2]};
    CLA_4 KS_4764(s4764, c4764, in4764_1, in4764_2);
    wire[3:0] s4765, in4765_1, in4765_2;
    wire c4765;
    assign in4765_1 = {pp126[61],s3277[0],s3277[1],s3264[2]};
    assign in4765_2 = {pp127[60],s3278[0],s3278[1],s3265[2]};
    CLA_4 KS_4765(s4765, c4765, in4765_1, in4765_2);
    wire[3:0] s4766, in4766_1, in4766_2;
    wire c4766;
    assign in4766_1 = {s3205[3],s3279[0],s3279[1],s3266[2]};
    assign in4766_2 = {s3206[3],s3280[0],s3280[1],s3267[2]};
    CLA_4 KS_4766(s4766, c4766, in4766_1, in4766_2);
    wire[3:0] s4767, in4767_1, in4767_2;
    wire c4767;
    assign in4767_1 = {s3207[3],s3281[0],s3281[1],s3268[2]};
    assign in4767_2 = {s3208[3],s3282[0],s3282[1],s3269[2]};
    CLA_4 KS_4767(s4767, c4767, in4767_1, in4767_2);
    wire[3:0] s4768, in4768_1, in4768_2;
    wire c4768;
    assign in4768_1 = {s3209[3],s3283[0],s3283[1],s3270[2]};
    assign in4768_2 = {s3210[3],s3284[0],s3284[1],s3271[2]};
    CLA_4 KS_4768(s4768, c4768, in4768_1, in4768_2);
    wire[3:0] s4769, in4769_1, in4769_2;
    wire c4769;
    assign in4769_1 = {s3211[3],s3285[0],c3285,s3272[2]};
    assign in4769_2 = {s3212[3],s3286[0],s3286[1],s3273[2]};
    CLA_4 KS_4769(s4769, c4769, in4769_1, in4769_2);
    wire[3:0] s4770, in4770_1, in4770_2;
    wire c4770;
    assign in4770_1 = {s3213[3],s3287[0],c3287,s3274[2]};
    assign in4770_2 = {s3214[3],s3288[0],s3288[1],s3275[2]};
    CLA_4 KS_4770(s4770, c4770, in4770_1, in4770_2);
    wire[3:0] s4771, in4771_1, in4771_2;
    wire c4771;
    assign in4771_1 = {s3215[3],s3289[0],c3289,s3276[2]};
    assign in4771_2 = {s3216[3],s3290[0],s3290[1],s3277[2]};
    CLA_4 KS_4771(s4771, c4771, in4771_1, in4771_2);
    wire[3:0] s4772, in4772_1, in4772_2;
    wire c4772;
    assign in4772_1 = {s3217[3],s3291[0],c3291,s3278[2]};
    assign in4772_2 = {s3218[3],s3292[0],s3292[1],s3279[2]};
    CLA_4 KS_4772(s4772, c4772, in4772_1, in4772_2);
    wire[3:0] s4773, in4773_1, in4773_2;
    wire c4773;
    assign in4773_1 = {s3219[3],s3293[0],c3293,s3280[2]};
    assign in4773_2 = {s3220[3],s3294[0],s3294[1],s3281[2]};
    CLA_4 KS_4773(s4773, c4773, in4773_1, in4773_2);
    wire[3:0] s4774, in4774_1, in4774_2;
    wire c4774;
    assign in4774_1 = {s3221[3],s3295[0],c3295,s3282[2]};
    assign in4774_2 = {s3222[3],s3296[0],s3296[1],s3283[2]};
    CLA_4 KS_4774(s4774, c4774, in4774_1, in4774_2);
    wire[3:0] s4775, in4775_1, in4775_2;
    wire c4775;
    assign in4775_1 = {s3223[3],s3297[0],c3297,c3284};
    assign in4775_2 = {s3224[3],s3298[0],s3298[1],s3286[2]};
    CLA_4 KS_4775(s4775, c4775, in4775_1, in4775_2);
    wire[3:0] s4776, in4776_1, in4776_2;
    wire c4776;
    assign in4776_1 = {s3225[3],s3299[0],c3299,c3288};
    assign in4776_2 = {s3226[3],s3300[0],s3300[1],s3290[2]};
    CLA_4 KS_4776(s4776, c4776, in4776_1, in4776_2);
    wire[3:0] s4777, in4777_1, in4777_2;
    wire c4777;
    assign in4777_1 = {s3227[3],s3301[0],c3301,c3292};
    assign in4777_2 = {s3228[3],s3302[0],s3302[1],s3294[2]};
    CLA_4 KS_4777(s4777, c4777, in4777_1, in4777_2);
    wire[2:0] s4778, in4778_1, in4778_2;
    wire c4778;
    assign in4778_1 = {c3229,s3303[0],c3303};
    assign in4778_2 = {s3232[3],s3304[0],s3304[1]};
    CLA_3 KS_4778(s4778, c4778, in4778_1, in4778_2);
    wire[0:0] s4779, in4779_1, in4779_2;
    wire c4779;
    assign in4779_1 = {c3236};
    assign in4779_2 = {s3240[3]};
    Half_Adder KS_4779(s4779, c4779, in4779_1, in4779_2);
    wire[1:0] s4780, in4780_1, in4780_2;
    wire c4780;
    assign in4780_1 = {c3244,s3305[0]};
    assign in4780_2 = {s3248[3],s3306[0]};
    CLA_2 KS_4780(s4780, c4780, in4780_1, in4780_2);
    wire[0:0] s4781, in4781_1, in4781_2;
    wire c4781;
    assign in4781_1 = {c3252};
    assign in4781_2 = {s3256[3]};
    Half_Adder KS_4781(s4781, c4781, in4781_1, in4781_2);
    wire[3:0] s4782, in4782_1, in4782_2;
    wire c4782;
    assign in4782_1 = {c3260,s3307[0],c3305,c3296};
    assign in4782_2 = {c4724,s3308[0],s3306[1],s3298[2]};
    CLA_4 KS_4782(s4782, c4782, in4782_1, in4782_2);
    wire[0:0] s4783, in4783_1, in4783_2;
    wire c4783;
    assign in4783_1 = {c4725};
    assign in4783_2 = {c4726};
    Half_Adder KS_4783(s4783, c4783, in4783_1, in4783_2);
    wire[1:0] s4784, in4784_1, in4784_2;
    wire c4784;
    assign in4784_1 = {c4727,s3309[0]};
    assign in4784_2 = {c4728,s3310[0]};
    CLA_2 KS_4784(s4784, c4784, in4784_1, in4784_2);
    wire[0:0] s4785, in4785_1, in4785_2;
    wire c4785;
    assign in4785_1 = {c4729};
    assign in4785_2 = {c4730};
    Half_Adder KS_4785(s4785, c4785, in4785_1, in4785_2);
    wire[2:0] s4786, in4786_1, in4786_2;
    wire c4786;
    assign in4786_1 = {c4731,s3311[0],c3307};
    assign in4786_2 = {c4732,s4760[1],s3308[1]};
    CLA_3 KS_4786(s4786, c4786, in4786_1, in4786_2);
    wire[0:0] s4787, in4787_1, in4787_2;
    wire c4787;
    assign in4787_1 = {c4733};
    assign in4787_2 = {c4734};
    Half_Adder KS_4787(s4787, c4787, in4787_1, in4787_2);
    wire[1:0] s4788, in4788_1, in4788_2;
    wire c4788;
    assign in4788_1 = {c4735,s4761[1]};
    assign in4788_2 = {c4736,s4762[1]};
    CLA_2 KS_4788(s4788, c4788, in4788_1, in4788_2);
    wire[0:0] s4789, in4789_1, in4789_2;
    wire c4789;
    assign in4789_1 = {c4737};
    assign in4789_2 = {c4738};
    Half_Adder KS_4789(s4789, c4789, in4789_1, in4789_2);
    wire[3:0] s4790, in4790_1, in4790_2;
    wire c4790;
    assign in4790_1 = {c4739,s4763[1],c3309,c3300};
    assign in4790_2 = {c4740,s4764[1],s3310[1],s3302[2]};
    CLA_4 KS_4790(s4790, c4790, in4790_1, in4790_2);
    wire[0:0] s4791, in4791_1, in4791_2;
    wire c4791;
    assign in4791_1 = {c4741};
    assign in4791_2 = {c4744};
    Half_Adder KS_4791(s4791, c4791, in4791_1, in4791_2);
    wire[1:0] s4792, in4792_1, in4792_2;
    wire c4792;
    assign in4792_1 = {c4752,s4765[1]};
    assign in4792_2 = {s4760[0],s4766[1]};
    CLA_2 KS_4792(s4792, c4792, in4792_1, in4792_2);
    wire[0:0] s4793, in4793_1, in4793_2;
    wire c4793;
    assign in4793_1 = {s4761[0]};
    assign in4793_2 = {s4762[0]};
    Half_Adder KS_4793(s4793, c4793, in4793_1, in4793_2);
    wire[2:0] s4794, in4794_1, in4794_2;
    wire c4794;
    assign in4794_1 = {s4763[0],s4767[1],c3311};
    assign in4794_2 = {s4764[0],s4768[1],s4760[2]};
    CLA_3 KS_4794(s4794, c4794, in4794_1, in4794_2);
    wire[0:0] s4795, in4795_1, in4795_2;
    wire c4795;
    assign in4795_1 = {s4765[0]};
    assign in4795_2 = {s4766[0]};
    Half_Adder KS_4795(s4795, c4795, in4795_1, in4795_2);
    wire[1:0] s4796, in4796_1, in4796_2;
    wire c4796;
    assign in4796_1 = {s4768[0],s4769[1]};
    assign in4796_2 = {s4769[0],s4770[1]};
    CLA_2_c KS_4796(s4796, c4796, in4796_1, in4796_2, s4767[0]);
    wire[3:0] s4797, in4797_1, in4797_2;
    wire c4797;
    assign in4797_1 = {pp112[79],c3286,pp124[69],pp113[81]};
    assign in4797_2 = {pp113[78],c3294,pp125[68],pp114[80]};
    CLA_4 KS_4797(s4797, c4797, in4797_1, in4797_2);
    wire[3:0] s4798, in4798_1, in4798_2;
    wire c4798;
    assign in4798_1 = {pp114[77],c3302,pp126[67],pp115[79]};
    assign in4798_2 = {pp115[76],c3310,pp127[66],pp116[78]};
    CLA_4 KS_4798(s4798, c4798, in4798_1, in4798_2);
    wire[3:0] s4799, in4799_1, in4799_2;
    wire c4799;
    assign in4799_1 = {pp116[75],s3312[0],s3312[1],pp117[77]};
    assign in4799_2 = {pp117[74],s3313[0],s3313[1],pp118[76]};
    CLA_4 KS_4799(s4799, c4799, in4799_1, in4799_2);
    wire[3:0] s4800, in4800_1, in4800_2;
    wire c4800;
    assign in4800_1 = {pp118[73],s3314[0],s3314[1],pp119[75]};
    assign in4800_2 = {pp119[72],s3315[0],s3315[1],pp120[74]};
    CLA_4 KS_4800(s4800, c4800, in4800_1, in4800_2);
    wire[3:0] s4801, in4801_1, in4801_2;
    wire c4801;
    assign in4801_1 = {pp120[71],s3316[0],s3316[1],pp121[73]};
    assign in4801_2 = {pp121[70],s3317[0],s3317[1],pp122[72]};
    CLA_4 KS_4801(s4801, c4801, in4801_1, in4801_2);
    wire[3:0] s4802, in4802_1, in4802_2;
    wire c4802;
    assign in4802_1 = {pp122[69],s3318[0],s3318[1],pp123[71]};
    assign in4802_2 = {pp123[68],s3319[0],s3319[1],pp124[70]};
    CLA_4 KS_4802(s4802, c4802, in4802_1, in4802_2);
    wire[3:0] s4803, in4803_1, in4803_2;
    wire c4803;
    assign in4803_1 = {pp124[67],s3320[0],s3320[1],pp125[69]};
    assign in4803_2 = {pp125[66],s3321[0],s3321[1],pp126[68]};
    CLA_4 KS_4803(s4803, c4803, in4803_1, in4803_2);
    wire[3:0] s4804, in4804_1, in4804_2;
    wire c4804;
    assign in4804_1 = {pp126[65],s3322[0],s3322[1],pp127[67]};
    assign in4804_2 = {pp127[64],s3323[0],s3323[1],s3312[2]};
    CLA_4 KS_4804(s4804, c4804, in4804_1, in4804_2);
    wire[3:0] s4805, in4805_1, in4805_2;
    wire c4805;
    assign in4805_1 = {s3263[3],s3324[0],s3324[1],s3313[2]};
    assign in4805_2 = {s3264[3],s3325[0],s3325[1],s3314[2]};
    CLA_4 KS_4805(s4805, c4805, in4805_1, in4805_2);
    wire[3:0] s4806, in4806_1, in4806_2;
    wire c4806;
    assign in4806_1 = {s3265[3],s3326[0],s3326[1],s3315[2]};
    assign in4806_2 = {s3266[3],s3327[0],s3327[1],s3316[2]};
    CLA_4 KS_4806(s4806, c4806, in4806_1, in4806_2);
    wire[3:0] s4807, in4807_1, in4807_2;
    wire c4807;
    assign in4807_1 = {s3267[3],s3328[0],s3328[1],s3317[2]};
    assign in4807_2 = {s3268[3],s3329[0],s3329[1],s3318[2]};
    CLA_4 KS_4807(s4807, c4807, in4807_1, in4807_2);
    wire[3:0] s4808, in4808_1, in4808_2;
    wire c4808;
    assign in4808_1 = {s3269[3],s3330[0],c3330,s3319[2]};
    assign in4808_2 = {s3270[3],s3331[0],s3331[1],s3320[2]};
    CLA_4 KS_4808(s4808, c4808, in4808_1, in4808_2);
    wire[3:0] s4809, in4809_1, in4809_2;
    wire c4809;
    assign in4809_1 = {s3271[3],s3332[0],c3332,s3321[2]};
    assign in4809_2 = {s3272[3],s3333[0],s3333[1],s3322[2]};
    CLA_4 KS_4809(s4809, c4809, in4809_1, in4809_2);
    wire[3:0] s4810, in4810_1, in4810_2;
    wire c4810;
    assign in4810_1 = {s3273[3],s3334[0],c3334,s3323[2]};
    assign in4810_2 = {s3274[3],s3335[0],s3335[1],s3324[2]};
    CLA_4 KS_4810(s4810, c4810, in4810_1, in4810_2);
    wire[3:0] s4811, in4811_1, in4811_2;
    wire c4811;
    assign in4811_1 = {s3275[3],s3336[0],c3336,s3325[2]};
    assign in4811_2 = {s3276[3],s3337[0],s3337[1],s3326[2]};
    CLA_4 KS_4811(s4811, c4811, in4811_1, in4811_2);
    wire[3:0] s4812, in4812_1, in4812_2;
    wire c4812;
    assign in4812_1 = {s3277[3],s3338[0],c3338,s3327[2]};
    assign in4812_2 = {s3278[3],s3339[0],s3339[1],s3328[2]};
    CLA_4 KS_4812(s4812, c4812, in4812_1, in4812_2);
    wire[3:0] s4813, in4813_1, in4813_2;
    wire c4813;
    assign in4813_1 = {s3279[3],s3340[0],c3340,c3329};
    assign in4813_2 = {s3280[3],s3341[0],s3341[1],s3331[2]};
    CLA_4 KS_4813(s4813, c4813, in4813_1, in4813_2);
    wire[3:0] s4814, in4814_1, in4814_2;
    wire c4814;
    assign in4814_1 = {s3281[3],s3342[0],c3342,c3333};
    assign in4814_2 = {s3282[3],s3343[0],s3343[1],s3335[2]};
    CLA_4 KS_4814(s4814, c4814, in4814_1, in4814_2);
    wire[2:0] s4815, in4815_1, in4815_2;
    wire c4815;
    assign in4815_1 = {c3283,s3344[0],c3344};
    assign in4815_2 = {s3286[3],s3345[0],s3345[1]};
    CLA_3 KS_4815(s4815, c4815, in4815_1, in4815_2);
    wire[0:0] s4816, in4816_1, in4816_2;
    wire c4816;
    assign in4816_1 = {c3290};
    assign in4816_2 = {s3294[3]};
    Half_Adder KS_4816(s4816, c4816, in4816_1, in4816_2);
    wire[1:0] s4817, in4817_1, in4817_2;
    wire c4817;
    assign in4817_1 = {c3298,s3346[0]};
    assign in4817_2 = {s3302[3],s3347[0]};
    CLA_2 KS_4817(s4817, c4817, in4817_1, in4817_2);
    wire[0:0] s4818, in4818_1, in4818_2;
    wire c4818;
    assign in4818_1 = {c3306};
    assign in4818_2 = {s3310[3]};
    Half_Adder KS_4818(s4818, c4818, in4818_1, in4818_2);
    wire[3:0] s4819, in4819_1, in4819_2;
    wire c4819;
    assign in4819_1 = {c4760,s3348[0],c3346,c3337};
    assign in4819_2 = {c4761,s3349[0],s3347[1],s3339[2]};
    CLA_4 KS_4819(s4819, c4819, in4819_1, in4819_2);
    wire[0:0] s4820, in4820_1, in4820_2;
    wire c4820;
    assign in4820_1 = {c4762};
    assign in4820_2 = {c4763};
    Half_Adder KS_4820(s4820, c4820, in4820_1, in4820_2);
    wire[1:0] s4821, in4821_1, in4821_2;
    wire c4821;
    assign in4821_1 = {c4764,s3350[0]};
    assign in4821_2 = {c4765,s3351[0]};
    CLA_2 KS_4821(s4821, c4821, in4821_1, in4821_2);
    wire[0:0] s4822, in4822_1, in4822_2;
    wire c4822;
    assign in4822_1 = {c4766};
    assign in4822_2 = {c4767};
    Half_Adder KS_4822(s4822, c4822, in4822_1, in4822_2);
    wire[2:0] s4823, in4823_1, in4823_2;
    wire c4823;
    assign in4823_1 = {c4768,s3352[0],c3348};
    assign in4823_2 = {c4769,s4797[1],s3349[1]};
    CLA_3 KS_4823(s4823, c4823, in4823_1, in4823_2);
    wire[0:0] s4824, in4824_1, in4824_2;
    wire c4824;
    assign in4824_1 = {c4770};
    assign in4824_2 = {c4771};
    Half_Adder KS_4824(s4824, c4824, in4824_1, in4824_2);
    wire[1:0] s4825, in4825_1, in4825_2;
    wire c4825;
    assign in4825_1 = {c4772,s4798[1]};
    assign in4825_2 = {c4773,s4799[1]};
    CLA_2 KS_4825(s4825, c4825, in4825_1, in4825_2);
    wire[0:0] s4826, in4826_1, in4826_2;
    wire c4826;
    assign in4826_1 = {c4774};
    assign in4826_2 = {c4775};
    Half_Adder KS_4826(s4826, c4826, in4826_1, in4826_2);
    wire[3:0] s4827, in4827_1, in4827_2;
    wire c4827;
    assign in4827_1 = {c4776,s4800[1],c3350,c3341};
    assign in4827_2 = {c4777,s4801[1],s3351[1],s3343[2]};
    CLA_4 KS_4827(s4827, c4827, in4827_1, in4827_2);
    wire[0:0] s4828, in4828_1, in4828_2;
    wire c4828;
    assign in4828_1 = {c4782};
    assign in4828_2 = {c4790};
    Half_Adder KS_4828(s4828, c4828, in4828_1, in4828_2);
    wire[1:0] s4829, in4829_1, in4829_2;
    wire c4829;
    assign in4829_1 = {s4797[0],s4802[1]};
    assign in4829_2 = {s4798[0],s4803[1]};
    CLA_2 KS_4829(s4829, c4829, in4829_1, in4829_2);
    wire[0:0] s4830, in4830_1, in4830_2;
    wire c4830;
    assign in4830_1 = {s4799[0]};
    assign in4830_2 = {s4800[0]};
    Half_Adder KS_4830(s4830, c4830, in4830_1, in4830_2);
    wire[2:0] s4831, in4831_1, in4831_2;
    wire c4831;
    assign in4831_1 = {s4801[0],s4804[1],c3352};
    assign in4831_2 = {s4802[0],s4805[1],s4797[2]};
    CLA_3 KS_4831(s4831, c4831, in4831_1, in4831_2);
    wire[0:0] s4832, in4832_1, in4832_2;
    wire c4832;
    assign in4832_1 = {s4804[0]};
    assign in4832_2 = {s4805[0]};
    Full_Adder KS_4832(s4832, c4832, in4832_1, in4832_2, s4803[0]);
    wire[3:0] s4833, in4833_1, in4833_2;
    wire c4833;
    assign in4833_1 = {pp106[89],c3318,pp116[81],pp107[91]};
    assign in4833_2 = {pp107[88],c3319,pp117[80],pp108[90]};
    CLA_4 KS_4833(s4833, c4833, in4833_1, in4833_2);
    wire[3:0] s4834, in4834_1, in4834_2;
    wire c4834;
    assign in4834_1 = {pp108[87],c3320,pp118[79],pp109[89]};
    assign in4834_2 = {pp109[86],c3321,pp119[78],pp110[88]};
    CLA_4 KS_4834(s4834, c4834, in4834_1, in4834_2);
    wire[3:0] s4835, in4835_1, in4835_2;
    wire c4835;
    assign in4835_1 = {pp110[85],c3322,pp120[77],pp111[87]};
    assign in4835_2 = {pp111[84],c3323,pp121[76],pp112[86]};
    CLA_4 KS_4835(s4835, c4835, in4835_1, in4835_2);
    wire[3:0] s4836, in4836_1, in4836_2;
    wire c4836;
    assign in4836_1 = {pp112[83],c3324,pp122[75],pp113[85]};
    assign in4836_2 = {pp113[82],c3325,pp123[74],pp114[84]};
    CLA_4 KS_4836(s4836, c4836, in4836_1, in4836_2);
    wire[3:0] s4837, in4837_1, in4837_2;
    wire c4837;
    assign in4837_1 = {pp114[81],c3326,pp124[73],pp115[83]};
    assign in4837_2 = {pp115[80],c3327,pp125[72],pp116[82]};
    CLA_4 KS_4837(s4837, c4837, in4837_1, in4837_2);
    wire[3:0] s4838, in4838_1, in4838_2;
    wire c4838;
    assign in4838_1 = {pp116[79],c3331,pp126[71],pp117[81]};
    assign in4838_2 = {pp117[78],c3339,pp127[70],pp118[80]};
    CLA_4 KS_4838(s4838, c4838, in4838_1, in4838_2);
    wire[3:0] s4839, in4839_1, in4839_2;
    wire c4839;
    assign in4839_1 = {pp118[77],c3347,s3353[1],pp119[79]};
    assign in4839_2 = {pp119[76],s3353[0],s3354[1],pp120[78]};
    CLA_4 KS_4839(s4839, c4839, in4839_1, in4839_2);
    wire[3:0] s4840, in4840_1, in4840_2;
    wire c4840;
    assign in4840_1 = {pp120[75],s3354[0],s3355[1],pp121[77]};
    assign in4840_2 = {pp121[74],s3355[0],s3356[1],pp122[76]};
    CLA_4 KS_4840(s4840, c4840, in4840_1, in4840_2);
    wire[3:0] s4841, in4841_1, in4841_2;
    wire c4841;
    assign in4841_1 = {pp122[73],s3356[0],s3357[1],pp123[75]};
    assign in4841_2 = {pp123[72],s3357[0],s3358[1],pp124[74]};
    CLA_4 KS_4841(s4841, c4841, in4841_1, in4841_2);
    wire[3:0] s4842, in4842_1, in4842_2;
    wire c4842;
    assign in4842_1 = {pp124[71],s3358[0],s3359[1],pp125[73]};
    assign in4842_2 = {pp125[70],s3359[0],s3360[1],pp126[72]};
    CLA_4 KS_4842(s4842, c4842, in4842_1, in4842_2);
    wire[3:0] s4843, in4843_1, in4843_2;
    wire c4843;
    assign in4843_1 = {pp126[69],s3360[0],s3361[1],pp127[71]};
    assign in4843_2 = {pp127[68],s3361[0],s3362[1],s3353[2]};
    CLA_4 KS_4843(s4843, c4843, in4843_1, in4843_2);
    wire[3:0] s4844, in4844_1, in4844_2;
    wire c4844;
    assign in4844_1 = {s3312[3],s3362[0],s3363[1],s3354[2]};
    assign in4844_2 = {s3313[3],s3363[0],s3364[1],s3355[2]};
    CLA_4 KS_4844(s4844, c4844, in4844_1, in4844_2);
    wire[3:0] s4845, in4845_1, in4845_2;
    wire c4845;
    assign in4845_1 = {s3314[3],s3364[0],s3365[1],s3356[2]};
    assign in4845_2 = {s3315[3],s3365[0],s3366[1],s3357[2]};
    CLA_4 KS_4845(s4845, c4845, in4845_1, in4845_2);
    wire[3:0] s4846, in4846_1, in4846_2;
    wire c4846;
    assign in4846_1 = {s3316[3],s3366[0],c3367,s3358[2]};
    assign in4846_2 = {s3317[3],s3367[0],s3368[1],s3359[2]};
    CLA_4 KS_4846(s4846, c4846, in4846_1, in4846_2);
    wire[3:0] s4847, in4847_1, in4847_2;
    wire c4847;
    assign in4847_1 = {s3318[3],s3368[0],c3369,s3360[2]};
    assign in4847_2 = {s3319[3],s3369[0],s3370[1],s3361[2]};
    CLA_4 KS_4847(s4847, c4847, in4847_1, in4847_2);
    wire[3:0] s4848, in4848_1, in4848_2;
    wire c4848;
    assign in4848_1 = {s3320[3],s3370[0],c3371,s3362[2]};
    assign in4848_2 = {s3321[3],s3371[0],s3372[1],s3363[2]};
    CLA_4 KS_4848(s4848, c4848, in4848_1, in4848_2);
    wire[3:0] s4849, in4849_1, in4849_2;
    wire c4849;
    assign in4849_1 = {s3322[3],s3372[0],c3373,s3364[2]};
    assign in4849_2 = {s3323[3],s3373[0],s3374[1],s3365[2]};
    CLA_4 KS_4849(s4849, c4849, in4849_1, in4849_2);
    wire[3:0] s4850, in4850_1, in4850_2;
    wire c4850;
    assign in4850_1 = {s3324[3],s3374[0],c3375,c3366};
    assign in4850_2 = {s3325[3],s3375[0],s3376[1],s3368[2]};
    CLA_4 KS_4850(s4850, c4850, in4850_1, in4850_2);
    wire[1:0] s4851, in4851_1, in4851_2;
    wire c4851;
    assign in4851_1 = {s3326[3],s3376[0]};
    assign in4851_2 = {s3327[3],s3377[0]};
    CLA_2 KS_4851(s4851, c4851, in4851_1, in4851_2);
    wire[0:0] s4852, in4852_1, in4852_2;
    wire c4852;
    assign in4852_1 = {c3328};
    assign in4852_2 = {s3331[3]};
    Half_Adder KS_4852(s4852, c4852, in4852_1, in4852_2);
    wire[2:0] s4853, in4853_1, in4853_2;
    wire c4853;
    assign in4853_1 = {c3335,s3378[0],c3377};
    assign in4853_2 = {s3339[3],s3379[0],s3378[1]};
    CLA_3 KS_4853(s4853, c4853, in4853_1, in4853_2);
    wire[0:0] s4854, in4854_1, in4854_2;
    wire c4854;
    assign in4854_1 = {c3343};
    assign in4854_2 = {s3347[3]};
    Half_Adder KS_4854(s4854, c4854, in4854_1, in4854_2);
    wire[1:0] s4855, in4855_1, in4855_2;
    wire c4855;
    assign in4855_1 = {c3351,s3380[0]};
    assign in4855_2 = {c4797,s3381[0]};
    CLA_2 KS_4855(s4855, c4855, in4855_1, in4855_2);
    wire[0:0] s4856, in4856_1, in4856_2;
    wire c4856;
    assign in4856_1 = {c4798};
    assign in4856_2 = {c4799};
    Half_Adder KS_4856(s4856, c4856, in4856_1, in4856_2);
    wire[3:0] s4857, in4857_1, in4857_2;
    wire c4857;
    assign in4857_1 = {c4800,s3382[0],c3379,c3370};
    assign in4857_2 = {c4801,s3383[0],s3380[1],s3372[2]};
    CLA_4 KS_4857(s4857, c4857, in4857_1, in4857_2);
    wire[0:0] s4858, in4858_1, in4858_2;
    wire c4858;
    assign in4858_1 = {c4802};
    assign in4858_2 = {c4803};
    Half_Adder KS_4858(s4858, c4858, in4858_1, in4858_2);
    wire[1:0] s4859, in4859_1, in4859_2;
    wire c4859;
    assign in4859_1 = {c4804,s3384[0]};
    assign in4859_2 = {c4805,s4833[1]};
    CLA_2 KS_4859(s4859, c4859, in4859_1, in4859_2);
    wire[0:0] s4860, in4860_1, in4860_2;
    wire c4860;
    assign in4860_1 = {c4806};
    assign in4860_2 = {c4807};
    Half_Adder KS_4860(s4860, c4860, in4860_1, in4860_2);
    wire[2:0] s4861, in4861_1, in4861_2;
    wire c4861;
    assign in4861_1 = {c4808,s4834[1],c3381};
    assign in4861_2 = {c4809,s4835[1],s3382[1]};
    CLA_3 KS_4861(s4861, c4861, in4861_1, in4861_2);
    wire[0:0] s4862, in4862_1, in4862_2;
    wire c4862;
    assign in4862_1 = {c4810};
    assign in4862_2 = {c4811};
    Half_Adder KS_4862(s4862, c4862, in4862_1, in4862_2);
    wire[1:0] s4863, in4863_1, in4863_2;
    wire c4863;
    assign in4863_1 = {c4812,s4836[1]};
    assign in4863_2 = {c4813,s4837[1]};
    CLA_2 KS_4863(s4863, c4863, in4863_1, in4863_2);
    wire[0:0] s4864, in4864_1, in4864_2;
    wire c4864;
    assign in4864_1 = {c4814};
    assign in4864_2 = {c4819};
    Half_Adder KS_4864(s4864, c4864, in4864_1, in4864_2);
    wire[3:0] s4865, in4865_1, in4865_2;
    wire c4865;
    assign in4865_1 = {c4827,s4838[1],c3383,c3374};
    assign in4865_2 = {s4833[0],s4839[1],s3384[1],s3376[2]};
    CLA_4 KS_4865(s4865, c4865, in4865_1, in4865_2);
    wire[0:0] s4866, in4866_1, in4866_2;
    wire c4866;
    assign in4866_1 = {s4834[0]};
    assign in4866_2 = {s4835[0]};
    Half_Adder KS_4866(s4866, c4866, in4866_1, in4866_2);
    wire[1:0] s4867, in4867_1, in4867_2;
    wire c4867;
    assign in4867_1 = {s4836[0],s4840[1]};
    assign in4867_2 = {s4837[0],s4841[1]};
    CLA_2 KS_4867(s4867, c4867, in4867_1, in4867_2);
    wire[0:0] s4868, in4868_1, in4868_2;
    wire c4868;
    assign in4868_1 = {s4838[0]};
    assign in4868_2 = {s4839[0]};
    Half_Adder KS_4868(s4868, c4868, in4868_1, in4868_2);
    wire[2:0] s4869, in4869_1, in4869_2;
    wire c4869;
    assign in4869_1 = {s4841[0],s4842[1],s4833[2]};
    assign in4869_2 = {s4842[0],s4843[1],s4834[2]};
    CLA_3_c KS_4869(s4869, c4869, in4869_1, in4869_2, s4840[0]);
    wire[3:0] s4870, in4870_1, in4870_2;
    wire c4870;
    assign in4870_1 = {pp102[97],pp122[78],pp108[93],pp101[101]};
    assign in4870_2 = {pp103[96],pp123[77],pp109[92],pp102[100]};
    CLA_4 KS_4870(s4870, c4870, in4870_1, in4870_2);
    wire[3:0] s4871, in4871_1, in4871_2;
    wire c4871;
    assign in4871_1 = {pp104[95],pp124[76],pp110[91],pp103[99]};
    assign in4871_2 = {pp105[94],pp125[75],pp111[90],pp104[98]};
    CLA_4 KS_4871(s4871, c4871, in4871_1, in4871_2);
    wire[3:0] s4872, in4872_1, in4872_2;
    wire c4872;
    assign in4872_1 = {pp106[93],pp126[74],pp112[89],pp105[97]};
    assign in4872_2 = {pp107[92],pp127[73],pp113[88],pp106[96]};
    CLA_4 KS_4872(s4872, c4872, in4872_1, in4872_2);
    wire[3:0] s4873, in4873_1, in4873_2;
    wire c4873;
    assign in4873_1 = {pp108[91],c3353,pp114[87],pp107[95]};
    assign in4873_2 = {pp109[90],c3354,pp115[86],pp108[94]};
    CLA_4 KS_4873(s4873, c4873, in4873_1, in4873_2);
    wire[3:0] s4874, in4874_1, in4874_2;
    wire c4874;
    assign in4874_1 = {pp110[89],c3355,pp116[85],pp109[93]};
    assign in4874_2 = {pp111[88],c3356,pp117[84],pp110[92]};
    CLA_4 KS_4874(s4874, c4874, in4874_1, in4874_2);
    wire[3:0] s4875, in4875_1, in4875_2;
    wire c4875;
    assign in4875_1 = {pp112[87],c3357,pp118[83],pp111[91]};
    assign in4875_2 = {pp113[86],c3358,pp119[82],pp112[90]};
    CLA_4 KS_4875(s4875, c4875, in4875_1, in4875_2);
    wire[3:0] s4876, in4876_1, in4876_2;
    wire c4876;
    assign in4876_1 = {pp114[85],c3359,pp120[81],pp113[89]};
    assign in4876_2 = {pp115[84],c3360,pp121[80],pp114[88]};
    CLA_4 KS_4876(s4876, c4876, in4876_1, in4876_2);
    wire[3:0] s4877, in4877_1, in4877_2;
    wire c4877;
    assign in4877_1 = {pp116[83],c3361,pp122[79],pp115[87]};
    assign in4877_2 = {pp117[82],c3362,pp123[78],pp116[86]};
    CLA_4 KS_4877(s4877, c4877, in4877_1, in4877_2);
    wire[3:0] s4878, in4878_1, in4878_2;
    wire c4878;
    assign in4878_1 = {pp118[81],c3363,pp124[77],pp117[85]};
    assign in4878_2 = {pp119[80],c3364,pp125[76],pp118[84]};
    CLA_4 KS_4878(s4878, c4878, in4878_1, in4878_2);
    wire[3:0] s4879, in4879_1, in4879_2;
    wire c4879;
    assign in4879_1 = {pp120[79],c3368,pp126[75],pp119[83]};
    assign in4879_2 = {pp121[78],c3376,pp127[74],pp120[82]};
    CLA_4 KS_4879(s4879, c4879, in4879_1, in4879_2);
    wire[3:0] s4880, in4880_1, in4880_2;
    wire c4880;
    assign in4880_1 = {pp122[77],c3384,s3385[1],pp121[81]};
    assign in4880_2 = {pp123[76],s3385[0],s3386[1],pp122[80]};
    CLA_4 KS_4880(s4880, c4880, in4880_1, in4880_2);
    wire[3:0] s4881, in4881_1, in4881_2;
    wire c4881;
    assign in4881_1 = {pp124[75],s3386[0],s3387[1],pp123[79]};
    assign in4881_2 = {pp125[74],s3387[0],s3388[1],pp124[78]};
    CLA_4 KS_4881(s4881, c4881, in4881_1, in4881_2);
    wire[3:0] s4882, in4882_1, in4882_2;
    wire c4882;
    assign in4882_1 = {pp126[73],s3388[0],s3389[1],pp125[77]};
    assign in4882_2 = {pp127[72],s3389[0],s3390[1],pp126[76]};
    CLA_4 KS_4882(s4882, c4882, in4882_1, in4882_2);
    wire[3:0] s4883, in4883_1, in4883_2;
    wire c4883;
    assign in4883_1 = {s3353[3],s3390[0],s3391[1],pp127[75]};
    assign in4883_2 = {s3354[3],s3391[0],s3392[1],s3385[2]};
    CLA_4 KS_4883(s4883, c4883, in4883_1, in4883_2);
    wire[3:0] s4884, in4884_1, in4884_2;
    wire c4884;
    assign in4884_1 = {s3355[3],s3392[0],s3393[1],s3386[2]};
    assign in4884_2 = {s3356[3],s3393[0],s3394[1],s3387[2]};
    CLA_4 KS_4884(s4884, c4884, in4884_1, in4884_2);
    wire[3:0] s4885, in4885_1, in4885_2;
    wire c4885;
    assign in4885_1 = {s3357[3],s3394[0],c3395,s3388[2]};
    assign in4885_2 = {s3358[3],s3395[0],s3396[1],s3389[2]};
    CLA_4 KS_4885(s4885, c4885, in4885_1, in4885_2);
    wire[3:0] s4886, in4886_1, in4886_2;
    wire c4886;
    assign in4886_1 = {s3359[3],s3396[0],c3397,s3390[2]};
    assign in4886_2 = {s3360[3],s3397[0],s3398[1],s3391[2]};
    CLA_4 KS_4886(s4886, c4886, in4886_1, in4886_2);
    wire[3:0] s4887, in4887_1, in4887_2;
    wire c4887;
    assign in4887_1 = {s3361[3],s3398[0],c3399,s3392[2]};
    assign in4887_2 = {s3362[3],s3399[0],s3400[1],s3393[2]};
    CLA_4 KS_4887(s4887, c4887, in4887_1, in4887_2);
    wire[1:0] s4888, in4888_1, in4888_2;
    wire c4888;
    assign in4888_1 = {s3363[3],s3400[0]};
    assign in4888_2 = {s3364[3],s3401[0]};
    CLA_2 KS_4888(s4888, c4888, in4888_1, in4888_2);
    wire[0:0] s4889, in4889_1, in4889_2;
    wire c4889;
    assign in4889_1 = {c3365};
    assign in4889_2 = {s3368[3]};
    Half_Adder KS_4889(s4889, c4889, in4889_1, in4889_2);
    wire[2:0] s4890, in4890_1, in4890_2;
    wire c4890;
    assign in4890_1 = {c3372,s3402[0],c3401};
    assign in4890_2 = {s3376[3],s3403[0],s3402[1]};
    CLA_3 KS_4890(s4890, c4890, in4890_1, in4890_2);
    wire[0:0] s4891, in4891_1, in4891_2;
    wire c4891;
    assign in4891_1 = {c3380};
    assign in4891_2 = {s3384[3]};
    Half_Adder KS_4891(s4891, c4891, in4891_1, in4891_2);
    wire[1:0] s4892, in4892_1, in4892_2;
    wire c4892;
    assign in4892_1 = {c4833,s3404[0]};
    assign in4892_2 = {c4834,s3405[0]};
    CLA_2 KS_4892(s4892, c4892, in4892_1, in4892_2);
    wire[0:0] s4893, in4893_1, in4893_2;
    wire c4893;
    assign in4893_1 = {c4835};
    assign in4893_2 = {c4836};
    Half_Adder KS_4893(s4893, c4893, in4893_1, in4893_2);
    wire[3:0] s4894, in4894_1, in4894_2;
    wire c4894;
    assign in4894_1 = {c4837,s3406[0],c3403,c3394};
    assign in4894_2 = {c4838,s3407[0],s3404[1],s3396[2]};
    CLA_4 KS_4894(s4894, c4894, in4894_1, in4894_2);
    wire[0:0] s4895, in4895_1, in4895_2;
    wire c4895;
    assign in4895_1 = {c4839};
    assign in4895_2 = {c4840};
    Half_Adder KS_4895(s4895, c4895, in4895_1, in4895_2);
    wire[1:0] s4896, in4896_1, in4896_2;
    wire c4896;
    assign in4896_1 = {c4841,s3408[0]};
    assign in4896_2 = {c4842,s4870[1]};
    CLA_2 KS_4896(s4896, c4896, in4896_1, in4896_2);
    wire[0:0] s4897, in4897_1, in4897_2;
    wire c4897;
    assign in4897_1 = {c4843};
    assign in4897_2 = {c4844};
    Half_Adder KS_4897(s4897, c4897, in4897_1, in4897_2);
    wire[2:0] s4898, in4898_1, in4898_2;
    wire c4898;
    assign in4898_1 = {c4845,s4871[1],c3405};
    assign in4898_2 = {c4846,s4872[1],s3406[1]};
    CLA_3 KS_4898(s4898, c4898, in4898_1, in4898_2);
    wire[0:0] s4899, in4899_1, in4899_2;
    wire c4899;
    assign in4899_1 = {c4847};
    assign in4899_2 = {c4848};
    Half_Adder KS_4899(s4899, c4899, in4899_1, in4899_2);
    wire[1:0] s4900, in4900_1, in4900_2;
    wire c4900;
    assign in4900_1 = {c4849,s4873[1]};
    assign in4900_2 = {c4850,s4874[1]};
    CLA_2 KS_4900(s4900, c4900, in4900_1, in4900_2);
    wire[0:0] s4901, in4901_1, in4901_2;
    wire c4901;
    assign in4901_1 = {c4857};
    assign in4901_2 = {c4865};
    Half_Adder KS_4901(s4901, c4901, in4901_1, in4901_2);
    wire[3:0] s4902, in4902_1, in4902_2;
    wire c4902;
    assign in4902_1 = {s4870[0],s4875[1],c3407,c3398};
    assign in4902_2 = {s4871[0],s4876[1],s3408[1],s3400[2]};
    CLA_4 KS_4902(s4902, c4902, in4902_1, in4902_2);
    wire[0:0] s4903, in4903_1, in4903_2;
    wire c4903;
    assign in4903_1 = {s4872[0]};
    assign in4903_2 = {s4873[0]};
    Half_Adder KS_4903(s4903, c4903, in4903_1, in4903_2);
    wire[1:0] s4904, in4904_1, in4904_2;
    wire c4904;
    assign in4904_1 = {s4874[0],s4877[1]};
    assign in4904_2 = {s4875[0],s4878[1]};
    CLA_2 KS_4904(s4904, c4904, in4904_1, in4904_2);
    wire[0:0] s4905, in4905_1, in4905_2;
    wire c4905;
    assign in4905_1 = {s4877[0]};
    assign in4905_2 = {s4878[0]};
    Full_Adder KS_4905(s4905, c4905, in4905_1, in4905_2, s4876[0]);
    wire[3:0] s4906, in4906_1, in4906_2;
    wire c4906;
    assign in4906_1 = {pp96[107],pp108[96],pp98[107],pp93[113]};
    assign in4906_2 = {pp97[106],pp109[95],pp99[106],pp94[112]};
    CLA_4 KS_4906(s4906, c4906, in4906_1, in4906_2);
    wire[3:0] s4907, in4907_1, in4907_2;
    wire c4907;
    assign in4907_1 = {pp98[105],pp110[94],pp100[105],pp95[111]};
    assign in4907_2 = {pp99[104],pp111[93],pp101[104],pp96[110]};
    CLA_4 KS_4907(s4907, c4907, in4907_1, in4907_2);
    wire[3:0] s4908, in4908_1, in4908_2;
    wire c4908;
    assign in4908_1 = {pp100[103],pp112[92],pp102[103],pp97[109]};
    assign in4908_2 = {pp101[102],pp113[91],pp103[102],pp98[108]};
    CLA_4 KS_4908(s4908, c4908, in4908_1, in4908_2);
    wire[3:0] s4909, in4909_1, in4909_2;
    wire c4909;
    assign in4909_1 = {pp102[101],pp114[90],pp104[101],pp99[107]};
    assign in4909_2 = {pp103[100],pp115[89],pp105[100],pp100[106]};
    CLA_4 KS_4909(s4909, c4909, in4909_1, in4909_2);
    wire[3:0] s4910, in4910_1, in4910_2;
    wire c4910;
    assign in4910_1 = {pp104[99],pp116[88],pp106[99],pp101[105]};
    assign in4910_2 = {pp105[98],pp117[87],pp107[98],pp102[104]};
    CLA_4 KS_4910(s4910, c4910, in4910_1, in4910_2);
    wire[3:0] s4911, in4911_1, in4911_2;
    wire c4911;
    assign in4911_1 = {pp106[97],pp118[86],pp108[97],pp103[103]};
    assign in4911_2 = {pp107[96],pp119[85],pp109[96],pp104[102]};
    CLA_4 KS_4911(s4911, c4911, in4911_1, in4911_2);
    wire[3:0] s4912, in4912_1, in4912_2;
    wire c4912;
    assign in4912_1 = {pp108[95],pp120[84],pp110[95],pp105[101]};
    assign in4912_2 = {pp109[94],pp121[83],pp111[94],pp106[100]};
    CLA_4 KS_4912(s4912, c4912, in4912_1, in4912_2);
    wire[3:0] s4913, in4913_1, in4913_2;
    wire c4913;
    assign in4913_1 = {pp110[93],pp122[82],pp112[93],pp107[99]};
    assign in4913_2 = {pp111[92],pp123[81],pp113[92],pp108[98]};
    CLA_4 KS_4913(s4913, c4913, in4913_1, in4913_2);
    wire[3:0] s4914, in4914_1, in4914_2;
    wire c4914;
    assign in4914_1 = {pp112[91],pp124[80],pp114[91],pp109[97]};
    assign in4914_2 = {pp113[90],pp125[79],pp115[90],pp110[96]};
    CLA_4 KS_4914(s4914, c4914, in4914_1, in4914_2);
    wire[3:0] s4915, in4915_1, in4915_2;
    wire c4915;
    assign in4915_1 = {pp114[89],pp126[78],pp116[89],pp111[95]};
    assign in4915_2 = {pp115[88],pp127[77],pp117[88],pp112[94]};
    CLA_4 KS_4915(s4915, c4915, in4915_1, in4915_2);
    wire[3:0] s4916, in4916_1, in4916_2;
    wire c4916;
    assign in4916_1 = {pp116[87],c3385,pp118[87],pp113[93]};
    assign in4916_2 = {pp117[86],c3386,pp119[86],pp114[92]};
    CLA_4 KS_4916(s4916, c4916, in4916_1, in4916_2);
    wire[3:0] s4917, in4917_1, in4917_2;
    wire c4917;
    assign in4917_1 = {pp118[85],c3387,pp120[85],pp115[91]};
    assign in4917_2 = {pp119[84],c3388,pp121[84],pp116[90]};
    CLA_4 KS_4917(s4917, c4917, in4917_1, in4917_2);
    wire[3:0] s4918, in4918_1, in4918_2;
    wire c4918;
    assign in4918_1 = {pp120[83],c3389,pp122[83],pp117[89]};
    assign in4918_2 = {pp121[82],c3390,pp123[82],pp118[88]};
    CLA_4 KS_4918(s4918, c4918, in4918_1, in4918_2);
    wire[3:0] s4919, in4919_1, in4919_2;
    wire c4919;
    assign in4919_1 = {pp122[81],c3391,pp124[81],pp119[87]};
    assign in4919_2 = {pp123[80],c3392,pp125[80],pp120[86]};
    CLA_4 KS_4919(s4919, c4919, in4919_1, in4919_2);
    wire[3:0] s4920, in4920_1, in4920_2;
    wire c4920;
    assign in4920_1 = {pp124[79],c3396,pp126[79],pp121[85]};
    assign in4920_2 = {pp125[78],c3404,pp127[78],pp122[84]};
    CLA_4 KS_4920(s4920, c4920, in4920_1, in4920_2);
    wire[3:0] s4921, in4921_1, in4921_2;
    wire c4921;
    assign in4921_1 = {pp126[77],s3409[0],s3409[1],pp123[83]};
    assign in4921_2 = {pp127[76],s3410[0],s3410[1],pp124[82]};
    CLA_4 KS_4921(s4921, c4921, in4921_1, in4921_2);
    wire[3:0] s4922, in4922_1, in4922_2;
    wire c4922;
    assign in4922_1 = {s3385[3],s3411[0],s3411[1],pp125[81]};
    assign in4922_2 = {s3386[3],s3412[0],s3412[1],pp126[80]};
    CLA_4 KS_4922(s4922, c4922, in4922_1, in4922_2);
    wire[3:0] s4923, in4923_1, in4923_2;
    wire c4923;
    assign in4923_1 = {s3387[3],s3413[0],s3413[1],pp127[79]};
    assign in4923_2 = {s3388[3],s3414[0],s3414[1],s3409[2]};
    CLA_4 KS_4923(s4923, c4923, in4923_1, in4923_2);
    wire[3:0] s4924, in4924_1, in4924_2;
    wire c4924;
    assign in4924_1 = {s3389[3],s3415[0],c3415,s3410[2]};
    assign in4924_2 = {s3390[3],s3416[0],s3416[1],s3411[2]};
    CLA_4 KS_4924(s4924, c4924, in4924_1, in4924_2);
    wire[0:0] s4925, in4925_1, in4925_2;
    wire c4925;
    assign in4925_1 = {s3391[3]};
    assign in4925_2 = {s3392[3]};
    Half_Adder KS_4925(s4925, c4925, in4925_1, in4925_2);
    wire[1:0] s4926, in4926_1, in4926_2;
    wire c4926;
    assign in4926_1 = {c3393,s3417[0]};
    assign in4926_2 = {s3396[3],s3418[0]};
    CLA_2 KS_4926(s4926, c4926, in4926_1, in4926_2);
    wire[0:0] s4927, in4927_1, in4927_2;
    wire c4927;
    assign in4927_1 = {c3400};
    assign in4927_2 = {s3404[3]};
    Half_Adder KS_4927(s4927, c4927, in4927_1, in4927_2);
    wire[2:0] s4928, in4928_1, in4928_2;
    wire c4928;
    assign in4928_1 = {c3408,s3419[0],c3417};
    assign in4928_2 = {c4870,s3420[0],s3418[1]};
    CLA_3 KS_4928(s4928, c4928, in4928_1, in4928_2);
    wire[0:0] s4929, in4929_1, in4929_2;
    wire c4929;
    assign in4929_1 = {c4871};
    assign in4929_2 = {c4872};
    Half_Adder KS_4929(s4929, c4929, in4929_1, in4929_2);
    wire[1:0] s4930, in4930_1, in4930_2;
    wire c4930;
    assign in4930_1 = {c4873,s3421[0]};
    assign in4930_2 = {c4874,s3422[0]};
    CLA_2 KS_4930(s4930, c4930, in4930_1, in4930_2);
    wire[0:0] s4931, in4931_1, in4931_2;
    wire c4931;
    assign in4931_1 = {c4875};
    assign in4931_2 = {c4876};
    Half_Adder KS_4931(s4931, c4931, in4931_1, in4931_2);
    wire[3:0] s4932, in4932_1, in4932_2;
    wire c4932;
    assign in4932_1 = {c4877,s3423[0],c3419,s3412[2]};
    assign in4932_2 = {c4878,s4906[1],s3420[1],s3413[2]};
    CLA_4 KS_4932(s4932, c4932, in4932_1, in4932_2);
    wire[0:0] s4933, in4933_1, in4933_2;
    wire c4933;
    assign in4933_1 = {c4879};
    assign in4933_2 = {c4880};
    Half_Adder KS_4933(s4933, c4933, in4933_1, in4933_2);
    wire[1:0] s4934, in4934_1, in4934_2;
    wire c4934;
    assign in4934_1 = {c4881,s4907[1]};
    assign in4934_2 = {c4882,s4908[1]};
    CLA_2 KS_4934(s4934, c4934, in4934_1, in4934_2);
    wire[0:0] s4935, in4935_1, in4935_2;
    wire c4935;
    assign in4935_1 = {c4883};
    assign in4935_2 = {c4884};
    Half_Adder KS_4935(s4935, c4935, in4935_1, in4935_2);
    wire[2:0] s4936, in4936_1, in4936_2;
    wire c4936;
    assign in4936_1 = {c4885,s4909[1],c3421};
    assign in4936_2 = {c4886,s4910[1],s3422[1]};
    CLA_3 KS_4936(s4936, c4936, in4936_1, in4936_2);
    wire[0:0] s4937, in4937_1, in4937_2;
    wire c4937;
    assign in4937_1 = {c4887};
    assign in4937_2 = {c4894};
    Half_Adder KS_4937(s4937, c4937, in4937_1, in4937_2);
    wire[1:0] s4938, in4938_1, in4938_2;
    wire c4938;
    assign in4938_1 = {c4902,s4911[1]};
    assign in4938_2 = {s4906[0],s4912[1]};
    CLA_2 KS_4938(s4938, c4938, in4938_1, in4938_2);
    wire[0:0] s4939, in4939_1, in4939_2;
    wire c4939;
    assign in4939_1 = {s4907[0]};
    assign in4939_2 = {s4908[0]};
    Half_Adder KS_4939(s4939, c4939, in4939_1, in4939_2);
    wire[3:0] s4940, in4940_1, in4940_2;
    wire c4940;
    assign in4940_1 = {s4909[0],s4913[1],c3423,c3414};
    assign in4940_2 = {s4910[0],s4914[1],s4906[2],s3416[2]};
    CLA_4 KS_4940(s4940, c4940, in4940_1, in4940_2);
    wire[0:0] s4941, in4941_1, in4941_2;
    wire c4941;
    assign in4941_1 = {s4911[0]};
    assign in4941_2 = {s4912[0]};
    Half_Adder KS_4941(s4941, c4941, in4941_1, in4941_2);
    wire[1:0] s4942, in4942_1, in4942_2;
    wire c4942;
    assign in4942_1 = {s4914[0],s4915[1]};
    assign in4942_2 = {s4915[0],s4916[1]};
    CLA_2_c KS_4942(s4942, c4942, in4942_1, in4942_2, s4913[0]);
    wire[3:0] s4943, in4943_1, in4943_2;
    wire c4943;
    assign in4943_1 = {pp90[117],pp94[114],pp90[119],pp87[123]};
    assign in4943_2 = {pp91[116],pp95[113],pp91[118],pp88[122]};
    CLA_4 KS_4943(s4943, c4943, in4943_1, in4943_2);
    wire[3:0] s4944, in4944_1, in4944_2;
    wire c4944;
    assign in4944_1 = {pp92[115],pp96[112],pp92[117],pp89[121]};
    assign in4944_2 = {pp93[114],pp97[111],pp93[116],pp90[120]};
    CLA_4 KS_4944(s4944, c4944, in4944_1, in4944_2);
    wire[3:0] s4945, in4945_1, in4945_2;
    wire c4945;
    assign in4945_1 = {pp94[113],pp98[110],pp94[115],pp91[119]};
    assign in4945_2 = {pp95[112],pp99[109],pp95[114],pp92[118]};
    CLA_4 KS_4945(s4945, c4945, in4945_1, in4945_2);
    wire[3:0] s4946, in4946_1, in4946_2;
    wire c4946;
    assign in4946_1 = {pp96[111],pp100[108],pp96[113],pp93[117]};
    assign in4946_2 = {pp97[110],pp101[107],pp97[112],pp94[116]};
    CLA_4 KS_4946(s4946, c4946, in4946_1, in4946_2);
    wire[3:0] s4947, in4947_1, in4947_2;
    wire c4947;
    assign in4947_1 = {pp98[109],pp102[106],pp98[111],pp95[115]};
    assign in4947_2 = {pp99[108],pp103[105],pp99[110],pp96[114]};
    CLA_4 KS_4947(s4947, c4947, in4947_1, in4947_2);
    wire[3:0] s4948, in4948_1, in4948_2;
    wire c4948;
    assign in4948_1 = {pp100[107],pp104[104],pp100[109],pp97[113]};
    assign in4948_2 = {pp101[106],pp105[103],pp101[108],pp98[112]};
    CLA_4 KS_4948(s4948, c4948, in4948_1, in4948_2);
    wire[3:0] s4949, in4949_1, in4949_2;
    wire c4949;
    assign in4949_1 = {pp102[105],pp106[102],pp102[107],pp99[111]};
    assign in4949_2 = {pp103[104],pp107[101],pp103[106],pp100[110]};
    CLA_4 KS_4949(s4949, c4949, in4949_1, in4949_2);
    wire[3:0] s4950, in4950_1, in4950_2;
    wire c4950;
    assign in4950_1 = {pp104[103],pp108[100],pp104[105],pp101[109]};
    assign in4950_2 = {pp105[102],pp109[99],pp105[104],pp102[108]};
    CLA_4 KS_4950(s4950, c4950, in4950_1, in4950_2);
    wire[3:0] s4951, in4951_1, in4951_2;
    wire c4951;
    assign in4951_1 = {pp106[101],pp110[98],pp106[103],pp103[107]};
    assign in4951_2 = {pp107[100],pp111[97],pp107[102],pp104[106]};
    CLA_4 KS_4951(s4951, c4951, in4951_1, in4951_2);
    wire[3:0] s4952, in4952_1, in4952_2;
    wire c4952;
    assign in4952_1 = {pp108[99],pp112[96],pp108[101],pp105[105]};
    assign in4952_2 = {pp109[98],pp113[95],pp109[100],pp106[104]};
    CLA_4 KS_4952(s4952, c4952, in4952_1, in4952_2);
    wire[3:0] s4953, in4953_1, in4953_2;
    wire c4953;
    assign in4953_1 = {pp110[97],pp114[94],pp110[99],pp107[103]};
    assign in4953_2 = {pp111[96],pp115[93],pp111[98],pp108[102]};
    CLA_4 KS_4953(s4953, c4953, in4953_1, in4953_2);
    wire[3:0] s4954, in4954_1, in4954_2;
    wire c4954;
    assign in4954_1 = {pp112[95],pp116[92],pp112[97],pp109[101]};
    assign in4954_2 = {pp113[94],pp117[91],pp113[96],pp110[100]};
    CLA_4 KS_4954(s4954, c4954, in4954_1, in4954_2);
    wire[3:0] s4955, in4955_1, in4955_2;
    wire c4955;
    assign in4955_1 = {pp114[93],pp118[90],pp114[95],pp111[99]};
    assign in4955_2 = {pp115[92],pp119[89],pp115[94],pp112[98]};
    CLA_4 KS_4955(s4955, c4955, in4955_1, in4955_2);
    wire[3:0] s4956, in4956_1, in4956_2;
    wire c4956;
    assign in4956_1 = {pp116[91],pp120[88],pp116[93],pp113[97]};
    assign in4956_2 = {pp117[90],pp121[87],pp117[92],pp114[96]};
    CLA_4 KS_4956(s4956, c4956, in4956_1, in4956_2);
    wire[3:0] s4957, in4957_1, in4957_2;
    wire c4957;
    assign in4957_1 = {pp118[89],pp122[86],pp118[91],pp115[95]};
    assign in4957_2 = {pp119[88],pp123[85],pp119[90],pp116[94]};
    CLA_4 KS_4957(s4957, c4957, in4957_1, in4957_2);
    wire[3:0] s4958, in4958_1, in4958_2;
    wire c4958;
    assign in4958_1 = {pp120[87],pp124[84],pp120[89],pp117[93]};
    assign in4958_2 = {pp121[86],pp125[83],pp121[88],pp118[92]};
    CLA_4 KS_4958(s4958, c4958, in4958_1, in4958_2);
    wire[3:0] s4959, in4959_1, in4959_2;
    wire c4959;
    assign in4959_1 = {pp122[85],pp126[82],pp122[87],pp119[91]};
    assign in4959_2 = {pp123[84],pp127[81],pp123[86],pp120[90]};
    CLA_4 KS_4959(s4959, c4959, in4959_1, in4959_2);
    wire[3:0] s4960, in4960_1, in4960_2;
    wire c4960;
    assign in4960_1 = {pp124[83],c3409,pp124[85],pp121[89]};
    assign in4960_2 = {pp125[82],c3410,pp125[84],pp122[88]};
    CLA_4 KS_4960(s4960, c4960, in4960_1, in4960_2);
    wire[1:0] s4961, in4961_1, in4961_2;
    wire c4961;
    assign in4961_1 = {pp126[81],c3411};
    assign in4961_2 = {pp127[80],c3412};
    CLA_2 KS_4961(s4961, c4961, in4961_1, in4961_2);
    wire[0:0] s4962, in4962_1, in4962_2;
    wire c4962;
    assign in4962_1 = {s3409[3]};
    assign in4962_2 = {s3410[3]};
    Half_Adder KS_4962(s4962, c4962, in4962_1, in4962_2);
    wire[3:0] s4963, in4963_1, in4963_2;
    wire c4963;
    assign in4963_1 = {s3411[3],c3416,pp126[83],pp123[87]};
    assign in4963_2 = {s3412[3],s3424[0],pp127[82],pp124[86]};
    CLA_4 KS_4963(s4963, c4963, in4963_1, in4963_2);
    wire[0:0] s4964, in4964_1, in4964_2;
    wire c4964;
    assign in4964_1 = {c3413};
    assign in4964_2 = {s3416[3]};
    Half_Adder KS_4964(s4964, c4964, in4964_1, in4964_2);
    wire[1:0] s4965, in4965_1, in4965_2;
    wire c4965;
    assign in4965_1 = {c3420,s3425[0]};
    assign in4965_2 = {c4906,s3426[0]};
    CLA_2 KS_4965(s4965, c4965, in4965_1, in4965_2);
    wire[0:0] s4966, in4966_1, in4966_2;
    wire c4966;
    assign in4966_1 = {c4907};
    assign in4966_2 = {c4908};
    Half_Adder KS_4966(s4966, c4966, in4966_1, in4966_2);
    wire[2:0] s4967, in4967_1, in4967_2;
    wire c4967;
    assign in4967_1 = {c4909,s3427[0],s3424[1]};
    assign in4967_2 = {c4910,s3428[0],s3425[1]};
    CLA_3 KS_4967(s4967, c4967, in4967_1, in4967_2);
    wire[0:0] s4968, in4968_1, in4968_2;
    wire c4968;
    assign in4968_1 = {c4911};
    assign in4968_2 = {c4912};
    Half_Adder KS_4968(s4968, c4968, in4968_1, in4968_2);
    wire[1:0] s4969, in4969_1, in4969_2;
    wire c4969;
    assign in4969_1 = {c4913,s3429[0]};
    assign in4969_2 = {c4914,s4943[1]};
    CLA_2 KS_4969(s4969, c4969, in4969_1, in4969_2);
    wire[0:0] s4970, in4970_1, in4970_2;
    wire c4970;
    assign in4970_1 = {c4915};
    assign in4970_2 = {c4916};
    Half_Adder KS_4970(s4970, c4970, in4970_1, in4970_2);
    wire[3:0] s4971, in4971_1, in4971_2;
    wire c4971;
    assign in4971_1 = {c4917,s4944[1],c3426,pp125[85]};
    assign in4971_2 = {c4918,s4945[1],s3427[1],pp126[84]};
    CLA_4 KS_4971(s4971, c4971, in4971_1, in4971_2);
    wire[0:0] s4972, in4972_1, in4972_2;
    wire c4972;
    assign in4972_1 = {c4919};
    assign in4972_2 = {c4920};
    Half_Adder KS_4972(s4972, c4972, in4972_1, in4972_2);
    wire[1:0] s4973, in4973_1, in4973_2;
    wire c4973;
    assign in4973_1 = {c4921,s4946[1]};
    assign in4973_2 = {c4922,s4947[1]};
    CLA_2 KS_4973(s4973, c4973, in4973_1, in4973_2);
    wire[0:0] s4974, in4974_1, in4974_2;
    wire c4974;
    assign in4974_1 = {c4923};
    assign in4974_2 = {c4924};
    Half_Adder KS_4974(s4974, c4974, in4974_1, in4974_2);
    wire[2:0] s4975, in4975_1, in4975_2;
    wire c4975;
    assign in4975_1 = {c4932,s4948[1],c3428};
    assign in4975_2 = {c4940,s4949[1],s3429[1]};
    CLA_3 KS_4975(s4975, c4975, in4975_1, in4975_2);
    wire[0:0] s4976, in4976_1, in4976_2;
    wire c4976;
    assign in4976_1 = {s4943[0]};
    assign in4976_2 = {s4944[0]};
    Half_Adder KS_4976(s4976, c4976, in4976_1, in4976_2);
    wire[1:0] s4977, in4977_1, in4977_2;
    wire c4977;
    assign in4977_1 = {s4945[0],s4950[1]};
    assign in4977_2 = {s4946[0],s4951[1]};
    CLA_2 KS_4977(s4977, c4977, in4977_1, in4977_2);
    wire[0:0] s4978, in4978_1, in4978_2;
    wire c4978;
    assign in4978_1 = {s4947[0]};
    assign in4978_2 = {s4948[0]};
    Half_Adder KS_4978(s4978, c4978, in4978_1, in4978_2);
    wire[3:0] s4979, in4979_1, in4979_2;
    wire c4979;
    assign in4979_1 = {s4949[0],s4952[1],s4943[2],pp127[83]};
    assign in4979_2 = {s4950[0],s4953[1],s4944[2],s3424[2]};
    CLA_4 KS_4979(s4979, c4979, in4979_1, in4979_2);
    wire[0:0] s4980, in4980_1, in4980_2;
    wire c4980;
    assign in4980_1 = {s4952[0]};
    assign in4980_2 = {s4953[0]};
    Full_Adder KS_4980(s4980, c4980, in4980_1, in4980_2, s4951[0]);
    wire[3:0] s4981, in4981_1, in4981_2;
    wire c4981;
    assign in4981_1 = {pp86[125],pp85[127],pp86[127],pp87[127]};
    assign in4981_2 = {pp87[124],pp86[126],pp87[126],pp88[126]};
    CLA_4 KS_4981(s4981, c4981, in4981_1, in4981_2);
    wire[3:0] s4982, in4982_1, in4982_2;
    wire c4982;
    assign in4982_1 = {pp88[123],pp87[125],pp88[125],pp89[125]};
    assign in4982_2 = {pp89[122],pp88[124],pp89[124],pp90[124]};
    CLA_4 KS_4982(s4982, c4982, in4982_1, in4982_2);
    wire[3:0] s4983, in4983_1, in4983_2;
    wire c4983;
    assign in4983_1 = {pp90[121],pp89[123],pp90[123],pp91[123]};
    assign in4983_2 = {pp91[120],pp90[122],pp91[122],pp92[122]};
    CLA_4 KS_4983(s4983, c4983, in4983_1, in4983_2);
    wire[3:0] s4984, in4984_1, in4984_2;
    wire c4984;
    assign in4984_1 = {pp92[119],pp91[121],pp92[121],pp93[121]};
    assign in4984_2 = {pp93[118],pp92[120],pp93[120],pp94[120]};
    CLA_4 KS_4984(s4984, c4984, in4984_1, in4984_2);
    wire[3:0] s4985, in4985_1, in4985_2;
    wire c4985;
    assign in4985_1 = {pp94[117],pp93[119],pp94[119],pp95[119]};
    assign in4985_2 = {pp95[116],pp94[118],pp95[118],pp96[118]};
    CLA_4 KS_4985(s4985, c4985, in4985_1, in4985_2);
    wire[3:0] s4986, in4986_1, in4986_2;
    wire c4986;
    assign in4986_1 = {pp96[115],pp95[117],pp96[117],pp97[117]};
    assign in4986_2 = {pp97[114],pp96[116],pp97[116],pp98[116]};
    CLA_4 KS_4986(s4986, c4986, in4986_1, in4986_2);
    wire[3:0] s4987, in4987_1, in4987_2;
    wire c4987;
    assign in4987_1 = {pp98[113],pp97[115],pp98[115],pp99[115]};
    assign in4987_2 = {pp99[112],pp98[114],pp99[114],pp100[114]};
    CLA_4 KS_4987(s4987, c4987, in4987_1, in4987_2);
    wire[3:0] s4988, in4988_1, in4988_2;
    wire c4988;
    assign in4988_1 = {pp100[111],pp99[113],pp100[113],pp101[113]};
    assign in4988_2 = {pp101[110],pp100[112],pp101[112],pp102[112]};
    CLA_4 KS_4988(s4988, c4988, in4988_1, in4988_2);
    wire[3:0] s4989, in4989_1, in4989_2;
    wire c4989;
    assign in4989_1 = {pp102[109],pp101[111],pp102[111],pp103[111]};
    assign in4989_2 = {pp103[108],pp102[110],pp103[110],pp104[110]};
    CLA_4 KS_4989(s4989, c4989, in4989_1, in4989_2);
    wire[3:0] s4990, in4990_1, in4990_2;
    wire c4990;
    assign in4990_1 = {pp104[107],pp103[109],pp104[109],pp105[109]};
    assign in4990_2 = {pp105[106],pp104[108],pp105[108],pp106[108]};
    CLA_4 KS_4990(s4990, c4990, in4990_1, in4990_2);
    wire[3:0] s4991, in4991_1, in4991_2;
    wire c4991;
    assign in4991_1 = {pp106[105],pp105[107],pp106[107],pp107[107]};
    assign in4991_2 = {pp107[104],pp106[106],pp107[106],pp108[106]};
    CLA_4 KS_4991(s4991, c4991, in4991_1, in4991_2);
    wire[3:0] s4992, in4992_1, in4992_2;
    wire c4992;
    assign in4992_1 = {pp108[103],pp107[105],pp108[105],pp109[105]};
    assign in4992_2 = {pp109[102],pp108[104],pp109[104],pp110[104]};
    CLA_4 KS_4992(s4992, c4992, in4992_1, in4992_2);
    wire[3:0] s4993, in4993_1, in4993_2;
    wire c4993;
    assign in4993_1 = {pp110[101],pp109[103],pp110[103],pp111[103]};
    assign in4993_2 = {pp111[100],pp110[102],pp111[102],pp112[102]};
    CLA_4 KS_4993(s4993, c4993, in4993_1, in4993_2);
    wire[3:0] s4994, in4994_1, in4994_2;
    wire c4994;
    assign in4994_1 = {pp112[99],pp111[101],pp112[101],pp113[101]};
    assign in4994_2 = {pp113[98],pp112[100],pp113[100],pp114[100]};
    CLA_4 KS_4994(s4994, c4994, in4994_1, in4994_2);
    wire[3:0] s4995, in4995_1, in4995_2;
    wire c4995;
    assign in4995_1 = {pp114[97],pp113[99],pp114[99],pp115[99]};
    assign in4995_2 = {pp115[96],pp114[98],pp115[98],pp116[98]};
    CLA_4 KS_4995(s4995, c4995, in4995_1, in4995_2);
    wire[2:0] s4996, in4996_1, in4996_2;
    wire c4996;
    assign in4996_1 = {pp116[95],pp115[97],pp116[97]};
    assign in4996_2 = {pp117[94],pp116[96],pp117[96]};
    CLA_3 KS_4996(s4996, c4996, in4996_1, in4996_2);
    wire[1:0] s4997, in4997_1, in4997_2;
    wire c4997;
    assign in4997_1 = {pp118[93],pp117[95]};
    assign in4997_2 = {pp119[92],pp118[94]};
    CLA_2 KS_4997(s4997, c4997, in4997_1, in4997_2);
    wire[3:0] s4998, in4998_1, in4998_2;
    wire c4998;
    assign in4998_1 = {pp120[91],pp119[93],pp118[95],pp117[97]};
    assign in4998_2 = {pp121[90],pp120[92],pp119[94],pp118[96]};
    CLA_4 KS_4998(s4998, c4998, in4998_1, in4998_2);
    wire[0:0] s4999, in4999_1, in4999_2;
    wire c4999;
    assign in4999_1 = {pp122[89]};
    assign in4999_2 = {pp123[88]};
    Half_Adder KS_4999(s4999, c4999, in4999_1, in4999_2);
    wire[1:0] s5000, in5000_1, in5000_2;
    wire c5000;
    assign in5000_1 = {pp124[87],pp121[91]};
    assign in5000_2 = {pp125[86],pp122[90]};
    CLA_2 KS_5000(s5000, c5000, in5000_1, in5000_2);
    wire[0:0] s5001, in5001_1, in5001_2;
    wire c5001;
    assign in5001_1 = {pp126[85]};
    assign in5001_2 = {pp127[84]};
    Half_Adder KS_5001(s5001, c5001, in5001_1, in5001_2);
    wire[2:0] s5002, in5002_1, in5002_2;
    wire c5002;
    assign in5002_1 = {c3424,pp123[89],pp120[93]};
    assign in5002_2 = {s3427[3],pp124[88],pp121[92]};
    CLA_3 KS_5002(s5002, c5002, in5002_1, in5002_2);
    wire[0:0] s5003, in5003_1, in5003_2;
    wire c5003;
    assign in5003_1 = {c4943};
    assign in5003_2 = {c4944};
    Half_Adder KS_5003(s5003, c5003, in5003_1, in5003_2);
    wire[1:0] s5004, in5004_1, in5004_2;
    wire c5004;
    assign in5004_1 = {c4945,pp125[87]};
    assign in5004_2 = {c4946,pp126[86]};
    CLA_2 KS_5004(s5004, c5004, in5004_1, in5004_2);
    wire[0:0] s5005, in5005_1, in5005_2;
    wire c5005;
    assign in5005_1 = {c4947};
    assign in5005_2 = {c4948};
    Half_Adder KS_5005(s5005, c5005, in5005_1, in5005_2);
    wire[3:0] s5006, in5006_1, in5006_2;
    wire c5006;
    assign in5006_1 = {c4949,pp127[85],pp122[91],pp119[95]};
    assign in5006_2 = {c4950,c3427,pp123[90],pp120[94]};
    CLA_4 KS_5006(s5006, c5006, in5006_1, in5006_2);
    wire[0:0] s5007, in5007_1, in5007_2;
    wire c5007;
    assign in5007_1 = {c4951};
    assign in5007_2 = {c4952};
    Half_Adder KS_5007(s5007, c5007, in5007_1, in5007_2);
    wire[1:0] s5008, in5008_1, in5008_2;
    wire c5008;
    assign in5008_1 = {c4953,s4981[1]};
    assign in5008_2 = {c4954,s4982[1]};
    CLA_2 KS_5008(s5008, c5008, in5008_1, in5008_2);
    wire[0:0] s5009, in5009_1, in5009_2;
    wire c5009;
    assign in5009_1 = {c4955};
    assign in5009_2 = {c4956};
    Half_Adder KS_5009(s5009, c5009, in5009_1, in5009_2);
    wire[2:0] s5010, in5010_1, in5010_2;
    wire c5010;
    assign in5010_1 = {c4957,s4983[1],pp124[89]};
    assign in5010_2 = {c4958,s4984[1],pp125[88]};
    CLA_3 KS_5010(s5010, c5010, in5010_1, in5010_2);
    wire[0:0] s5011, in5011_1, in5011_2;
    wire c5011;
    assign in5011_1 = {c4959};
    assign in5011_2 = {c4960};
    Half_Adder KS_5011(s5011, c5011, in5011_1, in5011_2);
    wire[1:0] s5012, in5012_1, in5012_2;
    wire c5012;
    assign in5012_1 = {c4963,s4985[1]};
    assign in5012_2 = {c4971,s4986[1]};
    CLA_2 KS_5012(s5012, c5012, in5012_1, in5012_2);
    wire[0:0] s5013, in5013_1, in5013_2;
    wire c5013;
    assign in5013_1 = {c4979};
    assign in5013_2 = {s4981[0]};
    Half_Adder KS_5013(s5013, c5013, in5013_1, in5013_2);
    wire[3:0] s5014, in5014_1, in5014_2;
    wire c5014;
    assign in5014_1 = {s4982[0],s4987[1],pp126[87],pp121[93]};
    assign in5014_2 = {s4983[0],s4988[1],pp127[86],pp122[92]};
    CLA_4 KS_5014(s5014, c5014, in5014_1, in5014_2);
    wire[0:0] s5015, in5015_1, in5015_2;
    wire c5015;
    assign in5015_1 = {s4984[0]};
    assign in5015_2 = {s4985[0]};
    Half_Adder KS_5015(s5015, c5015, in5015_1, in5015_2);
    wire[1:0] s5016, in5016_1, in5016_2;
    wire c5016;
    assign in5016_1 = {s4986[0],s4989[1]};
    assign in5016_2 = {s4987[0],s4990[1]};
    CLA_2 KS_5016(s5016, c5016, in5016_1, in5016_2);
    wire[0:0] s5017, in5017_1, in5017_2;
    wire c5017;
    assign in5017_1 = {s4989[0]};
    assign in5017_2 = {s4990[0]};
    Full_Adder KS_5017(s5017, c5017, in5017_1, in5017_2, s4988[0]);
    wire[3:0] s5018, in5018_1, in5018_2;
    wire c5018;
    assign in5018_1 = {pp88[127],pp89[127],pp90[127],pp91[127]};
    assign in5018_2 = {pp89[126],pp90[126],pp91[126],pp92[126]};
    CLA_4 KS_5018(s5018, c5018, in5018_1, in5018_2);
    wire[3:0] s5019, in5019_1, in5019_2;
    wire c5019;
    assign in5019_1 = {pp90[125],pp91[125],pp92[125],pp93[125]};
    assign in5019_2 = {pp91[124],pp92[124],pp93[124],pp94[124]};
    CLA_4 KS_5019(s5019, c5019, in5019_1, in5019_2);
    wire[3:0] s5020, in5020_1, in5020_2;
    wire c5020;
    assign in5020_1 = {pp92[123],pp93[123],pp94[123],pp95[123]};
    assign in5020_2 = {pp93[122],pp94[122],pp95[122],pp96[122]};
    CLA_4 KS_5020(s5020, c5020, in5020_1, in5020_2);
    wire[3:0] s5021, in5021_1, in5021_2;
    wire c5021;
    assign in5021_1 = {pp94[121],pp95[121],pp96[121],pp97[121]};
    assign in5021_2 = {pp95[120],pp96[120],pp97[120],pp98[120]};
    CLA_4 KS_5021(s5021, c5021, in5021_1, in5021_2);
    wire[3:0] s5022, in5022_1, in5022_2;
    wire c5022;
    assign in5022_1 = {pp96[119],pp97[119],pp98[119],pp99[119]};
    assign in5022_2 = {pp97[118],pp98[118],pp99[118],pp100[118]};
    CLA_4 KS_5022(s5022, c5022, in5022_1, in5022_2);
    wire[3:0] s5023, in5023_1, in5023_2;
    wire c5023;
    assign in5023_1 = {pp98[117],pp99[117],pp100[117],pp101[117]};
    assign in5023_2 = {pp99[116],pp100[116],pp101[116],pp102[116]};
    CLA_4 KS_5023(s5023, c5023, in5023_1, in5023_2);
    wire[3:0] s5024, in5024_1, in5024_2;
    wire c5024;
    assign in5024_1 = {pp100[115],pp101[115],pp102[115],pp103[115]};
    assign in5024_2 = {pp101[114],pp102[114],pp103[114],pp104[114]};
    CLA_4 KS_5024(s5024, c5024, in5024_1, in5024_2);
    wire[3:0] s5025, in5025_1, in5025_2;
    wire c5025;
    assign in5025_1 = {pp102[113],pp103[113],pp104[113],pp105[113]};
    assign in5025_2 = {pp103[112],pp104[112],pp105[112],pp106[112]};
    CLA_4 KS_5025(s5025, c5025, in5025_1, in5025_2);
    wire[3:0] s5026, in5026_1, in5026_2;
    wire c5026;
    assign in5026_1 = {pp104[111],pp105[111],pp106[111],pp107[111]};
    assign in5026_2 = {pp105[110],pp106[110],pp107[110],pp108[110]};
    CLA_4 KS_5026(s5026, c5026, in5026_1, in5026_2);
    wire[3:0] s5027, in5027_1, in5027_2;
    wire c5027;
    assign in5027_1 = {pp106[109],pp107[109],pp108[109],pp109[109]};
    assign in5027_2 = {pp107[108],pp108[108],pp109[108],pp110[108]};
    CLA_4 KS_5027(s5027, c5027, in5027_1, in5027_2);
    wire[3:0] s5028, in5028_1, in5028_2;
    wire c5028;
    assign in5028_1 = {pp108[107],pp109[107],pp110[107],pp111[107]};
    assign in5028_2 = {pp109[106],pp110[106],pp111[106],pp112[106]};
    CLA_4 KS_5028(s5028, c5028, in5028_1, in5028_2);
    wire[2:0] s5029, in5029_1, in5029_2;
    wire c5029;
    assign in5029_1 = {pp110[105],pp111[105],pp112[105]};
    assign in5029_2 = {pp111[104],pp112[104],pp113[104]};
    CLA_3 KS_5029(s5029, c5029, in5029_1, in5029_2);
    wire[1:0] s5030, in5030_1, in5030_2;
    wire c5030;
    assign in5030_1 = {pp112[103],pp113[103]};
    assign in5030_2 = {pp113[102],pp114[102]};
    CLA_2 KS_5030(s5030, c5030, in5030_1, in5030_2);
    wire[0:0] s5031, in5031_1, in5031_2;
    wire c5031;
    assign in5031_1 = {pp114[101]};
    assign in5031_2 = {pp115[100]};
    Half_Adder KS_5031(s5031, c5031, in5031_1, in5031_2);
    wire[3:0] s5032, in5032_1, in5032_2;
    wire c5032;
    assign in5032_1 = {pp116[99],pp115[101],pp114[103],pp113[105]};
    assign in5032_2 = {pp117[98],pp116[100],pp115[102],pp114[104]};
    CLA_4 KS_5032(s5032, c5032, in5032_1, in5032_2);
    wire[0:0] s5033, in5033_1, in5033_2;
    wire c5033;
    assign in5033_1 = {pp118[97]};
    assign in5033_2 = {pp119[96]};
    Half_Adder KS_5033(s5033, c5033, in5033_1, in5033_2);
    wire[1:0] s5034, in5034_1, in5034_2;
    wire c5034;
    assign in5034_1 = {pp120[95],pp117[99]};
    assign in5034_2 = {pp121[94],pp118[98]};
    CLA_2 KS_5034(s5034, c5034, in5034_1, in5034_2);
    wire[0:0] s5035, in5035_1, in5035_2;
    wire c5035;
    assign in5035_1 = {pp122[93]};
    assign in5035_2 = {pp123[92]};
    Half_Adder KS_5035(s5035, c5035, in5035_1, in5035_2);
    wire[2:0] s5036, in5036_1, in5036_2;
    wire c5036;
    assign in5036_1 = {pp124[91],pp119[97],pp116[101]};
    assign in5036_2 = {pp125[90],pp120[96],pp117[100]};
    CLA_3 KS_5036(s5036, c5036, in5036_1, in5036_2);
    wire[0:0] s5037, in5037_1, in5037_2;
    wire c5037;
    assign in5037_1 = {pp126[89]};
    assign in5037_2 = {pp127[88]};
    Half_Adder KS_5037(s5037, c5037, in5037_1, in5037_2);
    wire[1:0] s5038, in5038_1, in5038_2;
    wire c5038;
    assign in5038_1 = {c4981,pp121[95]};
    assign in5038_2 = {c4982,pp122[94]};
    CLA_2 KS_5038(s5038, c5038, in5038_1, in5038_2);
    wire[0:0] s5039, in5039_1, in5039_2;
    wire c5039;
    assign in5039_1 = {c4983};
    assign in5039_2 = {c4984};
    Half_Adder KS_5039(s5039, c5039, in5039_1, in5039_2);
    wire[3:0] s5040, in5040_1, in5040_2;
    wire c5040;
    assign in5040_1 = {c4985,pp123[93],pp118[99],pp115[103]};
    assign in5040_2 = {c4986,pp124[92],pp119[98],pp116[102]};
    CLA_4 KS_5040(s5040, c5040, in5040_1, in5040_2);
    wire[0:0] s5041, in5041_1, in5041_2;
    wire c5041;
    assign in5041_1 = {c4987};
    assign in5041_2 = {c4988};
    Half_Adder KS_5041(s5041, c5041, in5041_1, in5041_2);
    wire[1:0] s5042, in5042_1, in5042_2;
    wire c5042;
    assign in5042_1 = {c4989,pp125[91]};
    assign in5042_2 = {c4990,pp126[90]};
    CLA_2 KS_5042(s5042, c5042, in5042_1, in5042_2);
    wire[0:0] s5043, in5043_1, in5043_2;
    wire c5043;
    assign in5043_1 = {c4991};
    assign in5043_2 = {c4992};
    Half_Adder KS_5043(s5043, c5043, in5043_1, in5043_2);
    wire[2:0] s5044, in5044_1, in5044_2;
    wire c5044;
    assign in5044_1 = {c4993,pp127[89],pp120[97]};
    assign in5044_2 = {c4994,s5018[1],pp121[96]};
    CLA_3 KS_5044(s5044, c5044, in5044_1, in5044_2);
    wire[0:0] s5045, in5045_1, in5045_2;
    wire c5045;
    assign in5045_1 = {c4995};
    assign in5045_2 = {c4998};
    Half_Adder KS_5045(s5045, c5045, in5045_1, in5045_2);
    wire[1:0] s5046, in5046_1, in5046_2;
    wire c5046;
    assign in5046_1 = {c5006,s5019[1]};
    assign in5046_2 = {c5014,s5020[1]};
    CLA_2 KS_5046(s5046, c5046, in5046_1, in5046_2);
    wire[0:0] s5047, in5047_1, in5047_2;
    wire c5047;
    assign in5047_1 = {s5019[0]};
    assign in5047_2 = {s5020[0]};
    Full_Adder KS_5047(s5047, c5047, in5047_1, in5047_2, s5018[0]);
    wire[3:0] s5048, in5048_1, in5048_2;
    wire c5048;
    assign in5048_1 = {pp92[127],pp93[127],pp94[127],pp95[127]};
    assign in5048_2 = {pp93[126],pp94[126],pp95[126],pp96[126]};
    CLA_4 KS_5048(s5048, c5048, in5048_1, in5048_2);
    wire[3:0] s5049, in5049_1, in5049_2;
    wire c5049;
    assign in5049_1 = {pp94[125],pp95[125],pp96[125],pp97[125]};
    assign in5049_2 = {pp95[124],pp96[124],pp97[124],pp98[124]};
    CLA_4 KS_5049(s5049, c5049, in5049_1, in5049_2);
    wire[3:0] s5050, in5050_1, in5050_2;
    wire c5050;
    assign in5050_1 = {pp96[123],pp97[123],pp98[123],pp99[123]};
    assign in5050_2 = {pp97[122],pp98[122],pp99[122],pp100[122]};
    CLA_4 KS_5050(s5050, c5050, in5050_1, in5050_2);
    wire[3:0] s5051, in5051_1, in5051_2;
    wire c5051;
    assign in5051_1 = {pp98[121],pp99[121],pp100[121],pp101[121]};
    assign in5051_2 = {pp99[120],pp100[120],pp101[120],pp102[120]};
    CLA_4 KS_5051(s5051, c5051, in5051_1, in5051_2);
    wire[3:0] s5052, in5052_1, in5052_2;
    wire c5052;
    assign in5052_1 = {pp100[119],pp101[119],pp102[119],pp103[119]};
    assign in5052_2 = {pp101[118],pp102[118],pp103[118],pp104[118]};
    CLA_4 KS_5052(s5052, c5052, in5052_1, in5052_2);
    wire[3:0] s5053, in5053_1, in5053_2;
    wire c5053;
    assign in5053_1 = {pp102[117],pp103[117],pp104[117],pp105[117]};
    assign in5053_2 = {pp103[116],pp104[116],pp105[116],pp106[116]};
    CLA_4 KS_5053(s5053, c5053, in5053_1, in5053_2);
    wire[3:0] s5054, in5054_1, in5054_2;
    wire c5054;
    assign in5054_1 = {pp104[115],pp105[115],pp106[115],pp107[115]};
    assign in5054_2 = {pp105[114],pp106[114],pp107[114],pp108[114]};
    CLA_4 KS_5054(s5054, c5054, in5054_1, in5054_2);
    wire[2:0] s5055, in5055_1, in5055_2;
    wire c5055;
    assign in5055_1 = {pp106[113],pp107[113],pp108[113]};
    assign in5055_2 = {pp107[112],pp108[112],pp109[112]};
    CLA_3 KS_5055(s5055, c5055, in5055_1, in5055_2);
    wire[1:0] s5056, in5056_1, in5056_2;
    wire c5056;
    assign in5056_1 = {pp108[111],pp109[111]};
    assign in5056_2 = {pp109[110],pp110[110]};
    CLA_2 KS_5056(s5056, c5056, in5056_1, in5056_2);
    wire[0:0] s5057, in5057_1, in5057_2;
    wire c5057;
    assign in5057_1 = {pp110[109]};
    assign in5057_2 = {pp111[108]};
    Half_Adder KS_5057(s5057, c5057, in5057_1, in5057_2);
    wire[3:0] s5058, in5058_1, in5058_2;
    wire c5058;
    assign in5058_1 = {pp112[107],pp111[109],pp110[111],pp109[113]};
    assign in5058_2 = {pp113[106],pp112[108],pp111[110],pp110[112]};
    CLA_4 KS_5058(s5058, c5058, in5058_1, in5058_2);
    wire[0:0] s5059, in5059_1, in5059_2;
    wire c5059;
    assign in5059_1 = {pp114[105]};
    assign in5059_2 = {pp115[104]};
    Half_Adder KS_5059(s5059, c5059, in5059_1, in5059_2);
    wire[1:0] s5060, in5060_1, in5060_2;
    wire c5060;
    assign in5060_1 = {pp116[103],pp113[107]};
    assign in5060_2 = {pp117[102],pp114[106]};
    CLA_2 KS_5060(s5060, c5060, in5060_1, in5060_2);
    wire[0:0] s5061, in5061_1, in5061_2;
    wire c5061;
    assign in5061_1 = {pp118[101]};
    assign in5061_2 = {pp119[100]};
    Half_Adder KS_5061(s5061, c5061, in5061_1, in5061_2);
    wire[2:0] s5062, in5062_1, in5062_2;
    wire c5062;
    assign in5062_1 = {pp120[99],pp115[105],pp112[109]};
    assign in5062_2 = {pp121[98],pp116[104],pp113[108]};
    CLA_3 KS_5062(s5062, c5062, in5062_1, in5062_2);
    wire[0:0] s5063, in5063_1, in5063_2;
    wire c5063;
    assign in5063_1 = {pp122[97]};
    assign in5063_2 = {pp123[96]};
    Half_Adder KS_5063(s5063, c5063, in5063_1, in5063_2);
    wire[1:0] s5064, in5064_1, in5064_2;
    wire c5064;
    assign in5064_1 = {pp124[95],pp117[103]};
    assign in5064_2 = {pp125[94],pp118[102]};
    CLA_2 KS_5064(s5064, c5064, in5064_1, in5064_2);
    wire[0:0] s5065, in5065_1, in5065_2;
    wire c5065;
    assign in5065_1 = {pp126[93]};
    assign in5065_2 = {pp127[92]};
    Half_Adder KS_5065(s5065, c5065, in5065_1, in5065_2);
    wire[3:0] s5066, in5066_1, in5066_2;
    wire c5066;
    assign in5066_1 = {c5018,pp119[101],pp114[107],pp111[111]};
    assign in5066_2 = {c5019,pp120[100],pp115[106],pp112[110]};
    CLA_4 KS_5066(s5066, c5066, in5066_1, in5066_2);
    wire[0:0] s5067, in5067_1, in5067_2;
    wire c5067;
    assign in5067_1 = {c5020};
    assign in5067_2 = {c5021};
    Half_Adder KS_5067(s5067, c5067, in5067_1, in5067_2);
    wire[1:0] s5068, in5068_1, in5068_2;
    wire c5068;
    assign in5068_1 = {c5023,pp121[99]};
    assign in5068_2 = {c5024,pp122[98]};
    CLA_2_c KS_5068(s5068, c5068, in5068_1, in5068_2, c5022);
    wire[3:0] s5069, in5069_1, in5069_2;
    wire c5069;
    assign in5069_1 = {pp96[127],pp97[127],pp98[127],pp99[127]};
    assign in5069_2 = {pp97[126],pp98[126],pp99[126],pp100[126]};
    CLA_4 KS_5069(s5069, c5069, in5069_1, in5069_2);
    wire[3:0] s5070, in5070_1, in5070_2;
    wire c5070;
    assign in5070_1 = {pp98[125],pp99[125],pp100[125],pp101[125]};
    assign in5070_2 = {pp99[124],pp100[124],pp101[124],pp102[124]};
    CLA_4 KS_5070(s5070, c5070, in5070_1, in5070_2);
    wire[3:0] s5071, in5071_1, in5071_2;
    wire c5071;
    assign in5071_1 = {pp100[123],pp101[123],pp102[123],pp103[123]};
    assign in5071_2 = {pp101[122],pp102[122],pp103[122],pp104[122]};
    CLA_4 KS_5071(s5071, c5071, in5071_1, in5071_2);
    wire[2:0] s5072, in5072_1, in5072_2;
    wire c5072;
    assign in5072_1 = {pp102[121],pp103[121],pp104[121]};
    assign in5072_2 = {pp103[120],pp104[120],pp105[120]};
    CLA_3 KS_5072(s5072, c5072, in5072_1, in5072_2);
    wire[1:0] s5073, in5073_1, in5073_2;
    wire c5073;
    assign in5073_1 = {pp104[119],pp105[119]};
    assign in5073_2 = {pp105[118],pp106[118]};
    CLA_2 KS_5073(s5073, c5073, in5073_1, in5073_2);
    wire[0:0] s5074, in5074_1, in5074_2;
    wire c5074;
    assign in5074_1 = {pp106[117]};
    assign in5074_2 = {pp107[116]};
    Half_Adder KS_5074(s5074, c5074, in5074_1, in5074_2);
    wire[3:0] s5075, in5075_1, in5075_2;
    wire c5075;
    assign in5075_1 = {pp108[115],pp107[117],pp106[119],pp105[121]};
    assign in5075_2 = {pp109[114],pp108[116],pp107[118],pp106[120]};
    CLA_4 KS_5075(s5075, c5075, in5075_1, in5075_2);
    wire[0:0] s5076, in5076_1, in5076_2;
    wire c5076;
    assign in5076_1 = {pp110[113]};
    assign in5076_2 = {pp111[112]};
    Half_Adder KS_5076(s5076, c5076, in5076_1, in5076_2);
    wire[1:0] s5077, in5077_1, in5077_2;
    wire c5077;
    assign in5077_1 = {pp112[111],pp109[115]};
    assign in5077_2 = {pp113[110],pp110[114]};
    CLA_2 KS_5077(s5077, c5077, in5077_1, in5077_2);
    wire[0:0] s5078, in5078_1, in5078_2;
    wire c5078;
    assign in5078_1 = {pp114[109]};
    assign in5078_2 = {pp115[108]};
    Half_Adder KS_5078(s5078, c5078, in5078_1, in5078_2);
    wire[2:0] s5079, in5079_1, in5079_2;
    wire c5079;
    assign in5079_1 = {pp116[107],pp111[113],pp108[117]};
    assign in5079_2 = {pp117[106],pp112[112],pp109[116]};
    CLA_3 KS_5079(s5079, c5079, in5079_1, in5079_2);
    wire[0:0] s5080, in5080_1, in5080_2;
    wire c5080;
    assign in5080_1 = {pp118[105]};
    assign in5080_2 = {pp119[104]};
    Half_Adder KS_5080(s5080, c5080, in5080_1, in5080_2);
    wire[1:0] s5081, in5081_1, in5081_2;
    wire c5081;
    assign in5081_1 = {pp121[102],pp113[111]};
    assign in5081_2 = {pp122[101],pp114[110]};
    CLA_2_c KS_5081(s5081, c5081, in5081_1, in5081_2, pp120[103]);
    wire[1:0] s5082, in5082_1, in5082_2;
    wire c5082;
    assign in5082_1 = {pp100[127],pp101[127]};
    assign in5082_2 = {pp101[126],pp102[126]};
    CLA_2 KS_5082(s5082, c5082, in5082_1, in5082_2);
    wire[0:0] s5083, in5083_1, in5083_2;
    wire c5083;
    assign in5083_1 = {pp102[125]};
    assign in5083_2 = {pp103[124]};
    Half_Adder KS_5083(s5083, c5083, in5083_1, in5083_2);
    wire[2:0] s5084, in5084_1, in5084_2;
    wire c5084;
    assign in5084_1 = {pp104[123],pp103[125],pp102[127]};
    assign in5084_2 = {pp105[122],pp104[124],pp103[126]};
    CLA_3 KS_5084(s5084, c5084, in5084_1, in5084_2);
    wire[0:0] s5085, in5085_1, in5085_2;
    wire c5085;
    assign in5085_1 = {pp107[120]};
    assign in5085_2 = {pp108[119]};
    Full_Adder KS_5085(s5085, c5085, in5085_1, in5085_2, pp106[121]);

    /*Stage 4*/
    wire[3:0] s5086, in5086_1, in5086_2;
    wire c5086;
    assign in5086_1 = {pp0[16],pp0[17],pp0[18],pp0[19]};
    assign in5086_2 = {pp1[15],pp1[16],pp1[17],pp1[18]};
    CLA_4 KS_5086(s5086, c5086, in5086_1, in5086_2);
    wire[3:0] s5087, in5087_1, in5087_2;
    wire c5087;
    assign in5087_1 = {pp2[15],pp2[16],pp2[17],pp0[20]};
    assign in5087_2 = {pp3[14],pp3[15],pp3[16],pp1[19]};
    CLA_4 KS_5087(s5087, c5087, in5087_1, in5087_2);
    wire[3:0] s5088, in5088_1, in5088_2;
    wire c5088;
    assign in5088_1 = {pp4[14],pp4[15],pp2[18],pp0[21]};
    assign in5088_2 = {pp5[13],pp5[14],pp3[17],pp1[20]};
    CLA_4 KS_5088(s5088, c5088, in5088_1, in5088_2);
    wire[3:0] s5089, in5089_1, in5089_2;
    wire c5089;
    assign in5089_1 = {pp6[13],pp4[16],pp2[19],pp0[22]};
    assign in5089_2 = {pp7[12],pp5[15],pp3[18],pp1[21]};
    CLA_4 KS_5089(s5089, c5089, in5089_1, in5089_2);
    wire[3:0] s5090, in5090_1, in5090_2;
    wire c5090;
    assign in5090_1 = {pp6[14],pp4[17],pp2[20],pp0[23]};
    assign in5090_2 = {pp7[13],pp5[16],pp3[19],pp1[22]};
    CLA_4 KS_5090(s5090, c5090, in5090_1, in5090_2);
    wire[3:0] s5091, in5091_1, in5091_2;
    wire c5091;
    assign in5091_1 = {pp9[11],pp6[15],pp4[18],pp2[21]};
    assign in5091_2 = {pp10[10],pp7[14],pp5[17],pp3[20]};
    CLA_4_c KS_5091(s5091, c5091, in5091_1, in5091_2, pp8[12]);
    wire[3:0] s5092, in5092_1, in5092_2;
    wire c5092;
    assign in5092_1 = {pp8[13],pp6[16],pp4[19],pp0[24]};
    assign in5092_2 = {pp9[12],pp7[15],pp5[18],pp1[23]};
    CLA_4 KS_5092(s5092, c5092, in5092_1, in5092_2);
    wire[3:0] s5093, in5093_1, in5093_2;
    wire c5093;
    assign in5093_1 = {pp11[10],pp8[14],pp6[17],pp2[22]};
    assign in5093_2 = {pp12[9],pp9[13],pp7[16],pp3[21]};
    CLA_4_c KS_5093(s5093, c5093, in5093_1, in5093_2, pp10[11]);
    wire[3:0] s5094, in5094_1, in5094_2;
    wire c5094;
    assign in5094_1 = {pp10[12],pp8[15],pp4[20],pp0[25]};
    assign in5094_2 = {pp11[11],pp9[14],pp5[19],pp1[24]};
    CLA_4 KS_5094(s5094, c5094, in5094_1, in5094_2);
    wire[3:0] s5095, in5095_1, in5095_2;
    wire c5095;
    assign in5095_1 = {pp13[9],pp10[13],pp6[18],pp2[23]};
    assign in5095_2 = {pp14[8],pp11[12],pp7[17],pp3[22]};
    CLA_4_c KS_5095(s5095, c5095, in5095_1, in5095_2, pp12[10]);
    wire[3:0] s5096, in5096_1, in5096_2;
    wire c5096;
    assign in5096_1 = {pp12[11],pp8[16],pp4[21],pp0[26]};
    assign in5096_2 = {pp13[10],pp9[15],pp5[20],pp1[25]};
    CLA_4 KS_5096(s5096, c5096, in5096_1, in5096_2);
    wire[3:0] s5097, in5097_1, in5097_2;
    wire c5097;
    assign in5097_1 = {pp15[8],pp10[14],pp6[19],pp2[24]};
    assign in5097_2 = {pp16[7],pp11[13],pp7[18],pp3[23]};
    CLA_4_c KS_5097(s5097, c5097, in5097_1, in5097_2, pp14[9]);
    wire[3:0] s5098, in5098_1, in5098_2;
    wire c5098;
    assign in5098_1 = {pp12[12],pp8[17],pp4[22],pp2[25]};
    assign in5098_2 = {pp13[11],pp9[16],pp5[21],pp3[24]};
    CLA_4 KS_5098(s5098, c5098, in5098_1, in5098_2);
    wire[3:0] s5099, in5099_1, in5099_2;
    wire c5099;
    assign in5099_1 = {pp14[10],pp10[15],pp6[20],pp4[23]};
    assign in5099_2 = {pp15[9],pp11[14],pp7[19],pp5[22]};
    CLA_4 KS_5099(s5099, c5099, in5099_1, in5099_2);
    wire[3:0] s5100, in5100_1, in5100_2;
    wire c5100;
    assign in5100_1 = {pp16[8],pp12[13],pp8[18],pp6[21]};
    assign in5100_2 = {pp17[7],pp13[12],pp9[17],pp7[20]};
    CLA_4 KS_5100(s5100, c5100, in5100_1, in5100_2);
    wire[3:0] s5101, in5101_1, in5101_2;
    wire c5101;
    assign in5101_1 = {pp19[5],pp14[11],pp10[16],pp8[19]};
    assign in5101_2 = {pp20[4],pp15[10],pp11[15],pp9[18]};
    CLA_4_c KS_5101(s5101, c5101, in5101_1, in5101_2, pp18[6]);
    wire[3:0] s5102, in5102_1, in5102_2;
    wire c5102;
    assign in5102_1 = {pp16[9],pp12[14],pp10[17],pp4[24]};
    assign in5102_2 = {pp17[8],pp13[13],pp11[16],pp5[23]};
    CLA_4 KS_5102(s5102, c5102, in5102_1, in5102_2);
    wire[3:0] s5103, in5103_1, in5103_2;
    wire c5103;
    assign in5103_1 = {pp18[7],pp14[12],pp12[15],pp6[22]};
    assign in5103_2 = {pp19[6],pp15[11],pp13[14],pp7[21]};
    CLA_4 KS_5103(s5103, c5103, in5103_1, in5103_2);
    wire[3:0] s5104, in5104_1, in5104_2;
    wire c5104;
    assign in5104_1 = {pp21[4],pp16[10],pp14[13],pp8[20]};
    assign in5104_2 = {pp22[3],pp17[9],pp15[12],pp9[19]};
    CLA_4_c KS_5104(s5104, c5104, in5104_1, in5104_2, pp20[5]);
    wire[3:0] s5105, in5105_1, in5105_2;
    wire c5105;
    assign in5105_1 = {pp18[8],pp16[11],pp10[18],pp6[23]};
    assign in5105_2 = {pp19[7],pp17[10],pp11[17],pp7[22]};
    CLA_4 KS_5105(s5105, c5105, in5105_1, in5105_2);
    wire[3:0] s5106, in5106_1, in5106_2;
    wire c5106;
    assign in5106_1 = {pp20[6],pp18[9],pp12[16],pp8[21]};
    assign in5106_2 = {pp21[5],pp19[8],pp13[15],pp9[20]};
    CLA_4 KS_5106(s5106, c5106, in5106_1, in5106_2);
    wire[3:0] s5107, in5107_1, in5107_2;
    wire c5107;
    assign in5107_1 = {pp23[3],pp20[7],pp14[14],pp10[19]};
    assign in5107_2 = {pp24[2],pp21[6],pp15[13],pp11[18]};
    CLA_4_c KS_5107(s5107, c5107, in5107_1, in5107_2, pp22[4]);
    wire[3:0] s5108, in5108_1, in5108_2;
    wire c5108;
    assign in5108_1 = {pp22[5],pp16[12],pp12[17],pp8[22]};
    assign in5108_2 = {pp23[4],pp17[11],pp13[16],pp9[21]};
    CLA_4 KS_5108(s5108, c5108, in5108_1, in5108_2);
    wire[3:0] s5109, in5109_1, in5109_2;
    wire c5109;
    assign in5109_1 = {pp25[2],pp18[10],pp14[15],pp10[20]};
    assign in5109_2 = {pp26[1],pp19[9],pp15[14],pp11[19]};
    CLA_4_c KS_5109(s5109, c5109, in5109_1, in5109_2, pp24[3]);
    wire[3:0] s5110, in5110_1, in5110_2;
    wire c5110;
    assign in5110_1 = {pp20[8],pp16[13],pp12[18],pp11[20]};
    assign in5110_2 = {pp21[7],pp17[12],pp13[17],pp12[19]};
    CLA_4 KS_5110(s5110, c5110, in5110_1, in5110_2);
    wire[3:0] s5111, in5111_1, in5111_2;
    wire c5111;
    assign in5111_1 = {pp22[6],pp18[11],pp14[16],pp13[18]};
    assign in5111_2 = {pp23[5],pp19[10],pp15[15],pp14[17]};
    CLA_4 KS_5111(s5111, c5111, in5111_1, in5111_2);
    wire[3:0] s5112, in5112_1, in5112_2;
    wire c5112;
    assign in5112_1 = {pp24[4],pp20[9],pp16[14],pp15[16]};
    assign in5112_2 = {pp25[3],pp21[8],pp17[13],pp16[15]};
    CLA_4 KS_5112(s5112, c5112, in5112_1, in5112_2);
    wire[3:0] s5113, in5113_1, in5113_2;
    wire c5113;
    assign in5113_1 = {pp26[2],pp22[7],pp18[12],pp17[14]};
    assign in5113_2 = {pp27[1],pp23[6],pp19[11],pp18[13]};
    CLA_4 KS_5113(s5113, c5113, in5113_1, in5113_2);
    wire[3:0] s5114, in5114_1, in5114_2;
    wire c5114;
    assign in5114_1 = {pp28[0],pp24[5],pp20[10],pp19[12]};
    assign in5114_2 = {s3430[1],pp25[4],pp21[9],pp20[11]};
    CLA_4 KS_5114(s5114, c5114, in5114_1, in5114_2);
    wire[3:0] s5115, in5115_1, in5115_2;
    wire c5115;
    assign in5115_1 = {c5098,pp26[3],pp22[8],pp21[10]};
    assign in5115_2 = {c5099,pp27[2],pp23[7],pp22[9]};
    CLA_4_c KS_5115(s5115, c5115, in5115_1, in5115_2, s3431[0]);
    wire[3:0] s5116, in5116_1, in5116_2;
    wire c5116;
    assign in5116_1 = {pp28[1],pp24[6],pp23[8],pp13[19]};
    assign in5116_2 = {pp29[0],pp25[5],pp24[7],pp14[18]};
    CLA_4 KS_5116(s5116, c5116, in5116_1, in5116_2);
    wire[3:0] s5117, in5117_1, in5117_2;
    wire c5117;
    assign in5117_1 = {s3431[1],pp26[4],pp25[6],pp15[17]};
    assign in5117_2 = {s3432[0],pp27[3],pp26[5],pp16[16]};
    CLA_4_c KS_5117(s5117, c5117, in5117_1, in5117_2, s3430[2]);
    wire[3:0] s5118, in5118_1, in5118_2;
    wire c5118;
    assign in5118_1 = {pp28[2],pp27[4],pp17[15],pp15[18]};
    assign in5118_2 = {pp29[1],pp28[3],pp18[14],pp16[17]};
    CLA_4 KS_5118(s5118, c5118, in5118_1, in5118_2);
    wire[3:0] s5119, in5119_1, in5119_2;
    wire c5119;
    assign in5119_1 = {pp30[0],pp29[2],pp19[13],pp17[16]};
    assign in5119_2 = {s3430[3],pp30[1],pp20[12],pp18[15]};
    CLA_4 KS_5119(s5119, c5119, in5119_1, in5119_2);
    wire[3:0] s5120, in5120_1, in5120_2;
    wire c5120;
    assign in5120_1 = {s3432[1],pp31[0],pp21[11],pp19[14]};
    assign in5120_2 = {s3433[0],c3430,pp22[10],pp20[13]};
    CLA_4_c KS_5120(s5120, c5120, in5120_1, in5120_2, s3431[2]);
    wire[3:0] s5121, in5121_1, in5121_2;
    wire c5121;
    assign in5121_1 = {s3432[2],pp23[9],pp21[12],pp17[17]};
    assign in5121_2 = {s3433[1],pp24[8],pp22[11],pp18[16]};
    CLA_4_c KS_5121(s5121, c5121, in5121_1, in5121_2, s3431[3]);
    wire[3:0] s5122, in5122_1, in5122_2;
    wire c5122;
    assign in5122_1 = {pp25[7],pp23[10],pp19[15],pp21[14]};
    assign in5122_2 = {pp26[6],pp24[9],pp20[14],pp22[13]};
    CLA_4 KS_5122(s5122, c5122, in5122_1, in5122_2);
    wire[3:0] s5123, in5123_1, in5123_2;
    wire c5123;
    assign in5123_1 = {pp27[5],pp25[8],pp21[13],pp23[12]};
    assign in5123_2 = {pp28[4],pp26[7],pp22[12],pp24[11]};
    CLA_4 KS_5123(s5123, c5123, in5123_1, in5123_2);
    wire[3:0] s5124, in5124_1, in5124_2;
    wire c5124;
    assign in5124_1 = {pp29[3],pp27[6],pp23[11],pp25[10]};
    assign in5124_2 = {pp30[2],pp28[5],pp24[10],pp26[9]};
    CLA_4 KS_5124(s5124, c5124, in5124_1, in5124_2);
    wire[3:0] s5125, in5125_1, in5125_2;
    wire c5125;
    assign in5125_1 = {pp31[1],pp29[4],pp25[9],pp27[8]};
    assign in5125_2 = {pp32[0],pp30[3],pp26[8],pp28[7]};
    CLA_4 KS_5125(s5125, c5125, in5125_1, in5125_2);
    wire[3:0] s5126, in5126_1, in5126_2;
    wire c5126;
    assign in5126_1 = {c3431,pp31[2],pp27[7],pp29[6]};
    assign in5126_2 = {s3432[3],pp32[1],pp28[6],pp30[5]};
    CLA_4 KS_5126(s5126, c5126, in5126_1, in5126_2);
    wire[3:0] s5127, in5127_1, in5127_2;
    wire c5127;
    assign in5127_1 = {s3433[2],pp33[0],pp29[5],pp31[4]};
    assign in5127_2 = {s3434[1],c3432,pp30[4],pp32[3]};
    CLA_4 KS_5127(s5127, c5127, in5127_1, in5127_2);
    wire[3:0] s5128, in5128_1, in5128_2;
    wire c5128;
    assign in5128_1 = {s3435[1],s3433[3],pp31[3],pp33[2]};
    assign in5128_2 = {s3436[0],s3434[2],pp32[2],pp34[1]};
    CLA_4 KS_5128(s5128, c5128, in5128_1, in5128_2);
    wire[3:0] s5129, in5129_1, in5129_2;
    wire c5129;
    assign in5129_1 = {s3437[0],s3435[2],pp33[1],pp35[0]};
    assign in5129_2 = {c5110,s3436[1],pp34[0],c3434};
    CLA_4 KS_5129(s5129, c5129, in5129_1, in5129_2);
    wire[3:0] s5130, in5130_1, in5130_2;
    wire c5130;
    assign in5130_1 = {c5111,s3437[1],c3433,c3435};
    assign in5130_2 = {c5112,s3438[0],s3434[3],s3436[3]};
    CLA_4 KS_5130(s5130, c5130, in5130_1, in5130_2);
    wire[3:0] s5131, in5131_1, in5131_2;
    wire c5131;
    assign in5131_1 = {c5114,s3439[0],s3435[3],s3437[3]};
    assign in5131_2 = {c5115,c5116,s3436[2],s3438[2]};
    CLA_4_c KS_5131(s5131, c5131, in5131_1, in5131_2, c5113);
    wire[3:0] s5132, in5132_1, in5132_2;
    wire c5132;
    assign in5132_1 = {s3437[2],s3439[2],pp23[13],pp25[12]};
    assign in5132_2 = {s3438[1],s3440[1],pp24[12],pp26[11]};
    CLA_4 KS_5132(s5132, c5132, in5132_1, in5132_2);
    wire[3:0] s5133, in5133_1, in5133_2;
    wire c5133;
    assign in5133_1 = {s3440[0],s3441[1],pp25[11],pp27[10]};
    assign in5133_2 = {s3441[0],s3442[0],pp26[10],pp28[9]};
    CLA_4_c KS_5133(s5133, c5133, in5133_1, in5133_2, s3439[1]);
    wire[3:0] s5134, in5134_1, in5134_2;
    wire c5134;
    assign in5134_1 = {pp27[9],pp29[8],pp27[11],pp33[6]};
    assign in5134_2 = {pp28[8],pp30[7],pp28[10],pp34[5]};
    CLA_4 KS_5134(s5134, c5134, in5134_1, in5134_2);
    wire[3:0] s5135, in5135_1, in5135_2;
    wire c5135;
    assign in5135_1 = {pp29[7],pp31[6],pp29[9],pp35[4]};
    assign in5135_2 = {pp30[6],pp32[5],pp30[8],pp36[3]};
    CLA_4 KS_5135(s5135, c5135, in5135_1, in5135_2);
    wire[3:0] s5136, in5136_1, in5136_2;
    wire c5136;
    assign in5136_1 = {pp31[5],pp33[4],pp31[7],pp37[2]};
    assign in5136_2 = {pp32[4],pp34[3],pp32[6],pp38[1]};
    CLA_4 KS_5136(s5136, c5136, in5136_1, in5136_2);
    wire[3:0] s5137, in5137_1, in5137_2;
    wire c5137;
    assign in5137_1 = {pp33[3],pp35[2],pp33[5],pp39[0]};
    assign in5137_2 = {pp34[2],pp36[1],pp34[4],c3442};
    CLA_4 KS_5137(s5137, c5137, in5137_1, in5137_2);
    wire[3:0] s5138, in5138_1, in5138_2;
    wire c5138;
    assign in5138_1 = {pp35[1],pp37[0],pp35[3],c3443};
    assign in5138_2 = {pp36[0],c3438,pp36[2],c3444};
    CLA_4 KS_5138(s5138, c5138, in5138_1, in5138_2);
    wire[3:0] s5139, in5139_1, in5139_2;
    wire c5139;
    assign in5139_1 = {c3436,c3439,pp37[1],c3445};
    assign in5139_2 = {c3437,s3440[3],pp38[0],s3446[3]};
    CLA_4 KS_5139(s5139, c5139, in5139_1, in5139_2);
    wire[3:0] s5140, in5140_1, in5140_2;
    wire c5140;
    assign in5140_1 = {s3438[3],s3441[3],c3440,s3447[3]};
    assign in5140_2 = {s3439[3],s3442[2],c3441,s3448[3]};
    CLA_4 KS_5140(s5140, c5140, in5140_1, in5140_2);
    wire[3:0] s5141, in5141_1, in5141_2;
    wire c5141;
    assign in5141_1 = {s3440[2],s3443[2],s3442[3],s3449[2]};
    assign in5141_2 = {s3441[2],s3444[2],s3443[3],s3450[2]};
    CLA_4 KS_5141(s5141, c5141, in5141_1, in5141_2);
    wire[3:0] s5142, in5142_1, in5142_2;
    wire c5142;
    assign in5142_1 = {s3442[1],s3445[2],s3444[3],s3451[2]};
    assign in5142_2 = {s3443[1],s3446[1],s3445[3],s3452[1]};
    CLA_4 KS_5142(s5142, c5142, in5142_1, in5142_2);
    wire[3:0] s5143, in5143_1, in5143_2;
    wire c5143;
    assign in5143_1 = {s3444[1],s3447[1],s3446[2],s3453[1]};
    assign in5143_2 = {s3445[1],s3448[1],s3447[2],s3454[1]};
    CLA_4 KS_5143(s5143, c5143, in5143_1, in5143_2);
    wire[0:0] s5144, in5144_1, in5144_2;
    wire c5144;
    assign in5144_1 = {s3446[0]};
    assign in5144_2 = {s3447[0]};
    Half_Adder KS_5144(s5144, c5144, in5144_1, in5144_2);
    wire[3:0] s5145, in5145_1, in5145_2;
    wire c5145;
    assign in5145_1 = {s3448[0],s3449[0],s3448[2],s3455[0]};
    assign in5145_2 = {c5122,s3450[0],s3449[1],s3456[0]};
    CLA_4 KS_5145(s5145, c5145, in5145_1, in5145_2);
    wire[0:0] s5146, in5146_1, in5146_2;
    wire c5146;
    assign in5146_1 = {c5123};
    assign in5146_2 = {c5124};
    Half_Adder KS_5146(s5146, c5146, in5146_1, in5146_2);
    wire[3:0] s5147, in5147_1, in5147_2;
    wire c5147;
    assign in5147_1 = {c5125,s3451[0],s3450[1],s3457[0]};
    assign in5147_2 = {c5126,s5132[3],s3451[1],s3458[0]};
    CLA_4 KS_5147(s5147, c5147, in5147_1, in5147_2);
    wire[0:0] s5148, in5148_1, in5148_2;
    wire c5148;
    assign in5148_1 = {c5127};
    assign in5148_2 = {c5128};
    Half_Adder KS_5148(s5148, c5148, in5148_1, in5148_2);
    wire[2:0] s5149, in5149_1, in5149_2;
    wire c5149;
    assign in5149_1 = {c5129,s5133[3],s3452[0]};
    assign in5149_2 = {c5130,s5134[1],s3453[0]};
    CLA_3 KS_5149(s5149, c5149, in5149_1, in5149_2);
    wire[0:0] s5150, in5150_1, in5150_2;
    wire c5150;
    assign in5150_1 = {c5131};
    assign in5150_2 = {s5132[2]};
    Half_Adder KS_5150(s5150, c5150, in5150_1, in5150_2);
    wire[3:0] s5151, in5151_1, in5151_2;
    wire c5151;
    assign in5151_1 = {s5134[0],s5135[1],s3454[0],s3459[0]};
    assign in5151_2 = {s5135[0],s5136[1],c5132,s3460[0]};
    CLA_4_c KS_5151(s5151, c5151, in5151_1, in5151_2, s5133[2]);
    wire[3:0] s5152, in5152_1, in5152_2;
    wire c5152;
    assign in5152_1 = {pp33[7],pp35[6],pp37[5],c3458};
    assign in5152_2 = {pp34[6],pp36[5],pp38[4],c3459};
    CLA_4 KS_5152(s5152, c5152, in5152_1, in5152_2);
    wire[3:0] s5153, in5153_1, in5153_2;
    wire c5153;
    assign in5153_1 = {pp35[5],pp37[4],pp39[3],c3460};
    assign in5153_2 = {pp36[4],pp38[3],pp40[2],c3461};
    CLA_4 KS_5153(s5153, c5153, in5153_1, in5153_2);
    wire[3:0] s5154, in5154_1, in5154_2;
    wire c5154;
    assign in5154_1 = {pp37[3],pp39[2],pp41[1],s3462[3]};
    assign in5154_2 = {pp38[2],pp40[1],pp42[0],s3463[3]};
    CLA_4 KS_5154(s5154, c5154, in5154_1, in5154_2);
    wire[3:0] s5155, in5155_1, in5155_2;
    wire c5155;
    assign in5155_1 = {pp39[1],pp41[0],c3452,s3464[3]};
    assign in5155_2 = {pp40[0],c3449,c3453,s3465[2]};
    CLA_4 KS_5155(s5155, c5155, in5155_1, in5155_2);
    wire[3:0] s5156, in5156_1, in5156_2;
    wire c5156;
    assign in5156_1 = {c3446,c3450,c3454,s3466[2]};
    assign in5156_2 = {c3447,c3451,s3455[3],s3467[2]};
    CLA_4 KS_5156(s5156, c5156, in5156_1, in5156_2);
    wire[3:0] s5157, in5157_1, in5157_2;
    wire c5157;
    assign in5157_1 = {c3448,s3452[3],s3456[3],s3468[2]};
    assign in5157_2 = {s3449[3],s3453[3],s3457[3],s3469[1]};
    CLA_4 KS_5157(s5157, c5157, in5157_1, in5157_2);
    wire[3:0] s5158, in5158_1, in5158_2;
    wire c5158;
    assign in5158_1 = {s3450[3],s3454[3],s3458[3],s3470[1]};
    assign in5158_2 = {s3451[3],s3455[2],s3459[3],s3471[1]};
    CLA_4 KS_5158(s5158, c5158, in5158_1, in5158_2);
    wire[3:0] s5159, in5159_1, in5159_2;
    wire c5159;
    assign in5159_1 = {s3452[2],s3456[2],s3460[3],s3472[1]};
    assign in5159_2 = {s3453[2],s3457[2],s3461[3],s3473[0]};
    CLA_4 KS_5159(s5159, c5159, in5159_1, in5159_2);
    wire[3:0] s5160, in5160_1, in5160_2;
    wire c5160;
    assign in5160_1 = {s3454[2],s3458[2],s3462[2],s3474[0]};
    assign in5160_2 = {s3455[1],s3459[2],s3463[2],s3475[0]};
    CLA_4 KS_5160(s5160, c5160, in5160_1, in5160_2);
    wire[3:0] s5161, in5161_1, in5161_2;
    wire c5161;
    assign in5161_1 = {s3456[1],s3460[2],s3464[2],s3476[0]};
    assign in5161_2 = {s3457[1],s3461[2],s3465[1],s3477[0]};
    CLA_4 KS_5161(s5161, c5161, in5161_1, in5161_2);
    wire[3:0] s5162, in5162_1, in5162_2;
    wire c5162;
    assign in5162_1 = {s3458[1],s3462[1],s3466[1],s3478[0]};
    assign in5162_2 = {s3459[1],s3463[1],s3467[1],s3479[0]};
    CLA_4 KS_5162(s5162, c5162, in5162_1, in5162_2);
    wire[3:0] s5163, in5163_1, in5163_2;
    wire c5163;
    assign in5163_1 = {s3460[1],s3464[1],s3468[1],s3480[0]};
    assign in5163_2 = {s3461[1],s3465[0],s3469[0],s3481[0]};
    CLA_4 KS_5163(s5163, c5163, in5163_1, in5163_2);
    wire[0:0] s5164, in5164_1, in5164_2;
    wire c5164;
    assign in5164_1 = {s3462[0]};
    assign in5164_2 = {s3463[0]};
    Half_Adder KS_5164(s5164, c5164, in5164_1, in5164_2);
    wire[1:0] s5165, in5165_1, in5165_2;
    wire c5165;
    assign in5165_1 = {s3464[0],s3466[0]};
    assign in5165_2 = {c5134,s3467[0]};
    CLA_2 KS_5165(s5165, c5165, in5165_1, in5165_2);
    wire[0:0] s5166, in5166_1, in5166_2;
    wire c5166;
    assign in5166_1 = {c5135};
    assign in5166_2 = {c5136};
    Half_Adder KS_5166(s5166, c5166, in5166_1, in5166_2);
    wire[2:0] s5167, in5167_1, in5167_2;
    wire c5167;
    assign in5167_1 = {c5137,s3468[0],s3470[0]};
    assign in5167_2 = {c5138,s5152[1],s3471[0]};
    CLA_3 KS_5167(s5167, c5167, in5167_1, in5167_2);
    wire[0:0] s5168, in5168_1, in5168_2;
    wire c5168;
    assign in5168_1 = {c5139};
    assign in5168_2 = {c5140};
    Half_Adder KS_5168(s5168, c5168, in5168_1, in5168_2);
    wire[1:0] s5169, in5169_1, in5169_2;
    wire c5169;
    assign in5169_1 = {c5141,s5153[1]};
    assign in5169_2 = {c5142,s5154[1]};
    CLA_2 KS_5169(s5169, c5169, in5169_1, in5169_2);
    wire[0:0] s5170, in5170_1, in5170_2;
    wire c5170;
    assign in5170_1 = {c5143};
    assign in5170_2 = {c5145};
    Half_Adder KS_5170(s5170, c5170, in5170_1, in5170_2);
    wire[3:0] s5171, in5171_1, in5171_2;
    wire c5171;
    assign in5171_1 = {c5147,s5155[1],s3472[0],s3482[0]};
    assign in5171_2 = {c5151,s5156[1],s5152[2],s3483[0]};
    CLA_4 KS_5171(s5171, c5171, in5171_1, in5171_2);
    wire[0:0] s5172, in5172_1, in5172_2;
    wire c5172;
    assign in5172_1 = {s5152[0]};
    assign in5172_2 = {s5153[0]};
    Half_Adder KS_5172(s5172, c5172, in5172_1, in5172_2);
    wire[1:0] s5173, in5173_1, in5173_2;
    wire c5173;
    assign in5173_1 = {s5154[0],s5157[1]};
    assign in5173_2 = {s5155[0],s5158[1]};
    CLA_2 KS_5173(s5173, c5173, in5173_1, in5173_2);
    wire[0:0] s5174, in5174_1, in5174_2;
    wire c5174;
    assign in5174_1 = {s5157[0]};
    assign in5174_2 = {s5158[0]};
    Full_Adder KS_5174(s5174, c5174, in5174_1, in5174_2, s5156[0]);
    wire[3:0] s5175, in5175_1, in5175_2;
    wire c5175;
    assign in5175_1 = {pp42[2],pp45[0],s1327[1],s3487[2]};
    assign in5175_2 = {pp43[1],s1327[0],s1328[0],s3488[2]};
    CLA_4 KS_5175(s5175, c5175, in5175_1, in5175_2);
    wire[3:0] s5176, in5176_1, in5176_2;
    wire c5176;
    assign in5176_1 = {pp44[0],c3465,c3469,s3489[2]};
    assign in5176_2 = {c3462,c3466,c3470,s3490[1]};
    CLA_4 KS_5176(s5176, c5176, in5176_1, in5176_2);
    wire[3:0] s5177, in5177_1, in5177_2;
    wire c5177;
    assign in5177_1 = {c3463,c3467,c3471,s3491[1]};
    assign in5177_2 = {c3464,c3468,c3472,s3492[1]};
    CLA_4 KS_5177(s5177, c5177, in5177_1, in5177_2);
    wire[3:0] s5178, in5178_1, in5178_2;
    wire c5178;
    assign in5178_1 = {s3465[3],s3469[3],s3473[3],s3493[1]};
    assign in5178_2 = {s3466[3],s3470[3],s3474[3],s3494[0]};
    CLA_4 KS_5178(s5178, c5178, in5178_1, in5178_2);
    wire[3:0] s5179, in5179_1, in5179_2;
    wire c5179;
    assign in5179_1 = {s3467[3],s3471[3],s3475[3],s3495[0]};
    assign in5179_2 = {s3468[3],s3472[3],s3476[3],s3496[0]};
    CLA_4 KS_5179(s5179, c5179, in5179_1, in5179_2);
    wire[3:0] s5180, in5180_1, in5180_2;
    wire c5180;
    assign in5180_1 = {s3469[2],s3473[2],s3477[3],s3497[0]};
    assign in5180_2 = {s3470[2],s3474[2],s3478[3],s3498[0]};
    CLA_4 KS_5180(s5180, c5180, in5180_1, in5180_2);
    wire[3:0] s5181, in5181_1, in5181_2;
    wire c5181;
    assign in5181_1 = {s3471[2],s3475[2],s3479[3],s3499[0]};
    assign in5181_2 = {s3472[2],s3476[2],s3480[3],s3500[0]};
    CLA_4 KS_5181(s5181, c5181, in5181_1, in5181_2);
    wire[3:0] s5182, in5182_1, in5182_2;
    wire c5182;
    assign in5182_1 = {s3473[1],s3477[2],s3481[3],s3501[0]};
    assign in5182_2 = {s3474[1],s3478[2],s3482[3],s3502[0]};
    CLA_4 KS_5182(s5182, c5182, in5182_1, in5182_2);
    wire[3:0] s5183, in5183_1, in5183_2;
    wire c5183;
    assign in5183_1 = {s3475[1],s3479[2],s3483[3],s3503[0]};
    assign in5183_2 = {s3476[1],s3480[2],s3484[3],s3504[0]};
    CLA_4 KS_5183(s5183, c5183, in5183_1, in5183_2);
    wire[3:0] s5184, in5184_1, in5184_2;
    wire c5184;
    assign in5184_1 = {s3477[1],s3481[2],s3485[2],s3505[0]};
    assign in5184_2 = {s3478[1],s3482[2],s3486[1],s3506[0]};
    CLA_4 KS_5184(s5184, c5184, in5184_1, in5184_2);
    wire[3:0] s5185, in5185_1, in5185_2;
    wire c5185;
    assign in5185_1 = {s3479[1],s3483[2],s3487[1],s3507[0]};
    assign in5185_2 = {s3480[1],s3484[2],s3488[1],s3508[0]};
    CLA_4 KS_5185(s5185, c5185, in5185_1, in5185_2);
    wire[3:0] s5186, in5186_1, in5186_2;
    wire c5186;
    assign in5186_1 = {s3481[1],s3485[1],s3489[1],s3509[0]};
    assign in5186_2 = {s3482[1],s3486[0],s3490[0],s3510[0]};
    CLA_4 KS_5186(s5186, c5186, in5186_1, in5186_2);
    wire[0:0] s5187, in5187_1, in5187_2;
    wire c5187;
    assign in5187_1 = {s3483[1]};
    assign in5187_2 = {s3484[1]};
    Half_Adder KS_5187(s5187, c5187, in5187_1, in5187_2);
    wire[1:0] s5188, in5188_1, in5188_2;
    wire c5188;
    assign in5188_1 = {s3485[0],s3487[0]};
    assign in5188_2 = {c5152,s3488[0]};
    CLA_2 KS_5188(s5188, c5188, in5188_1, in5188_2);
    wire[0:0] s5189, in5189_1, in5189_2;
    wire c5189;
    assign in5189_1 = {c5153};
    assign in5189_2 = {c5154};
    Half_Adder KS_5189(s5189, c5189, in5189_1, in5189_2);
    wire[2:0] s5190, in5190_1, in5190_2;
    wire c5190;
    assign in5190_1 = {c5155,s3489[0],s3491[0]};
    assign in5190_2 = {c5156,s5175[1],s3492[0]};
    CLA_3 KS_5190(s5190, c5190, in5190_1, in5190_2);
    wire[0:0] s5191, in5191_1, in5191_2;
    wire c5191;
    assign in5191_1 = {c5157};
    assign in5191_2 = {c5158};
    Half_Adder KS_5191(s5191, c5191, in5191_1, in5191_2);
    wire[1:0] s5192, in5192_1, in5192_2;
    wire c5192;
    assign in5192_1 = {c5159,s5176[1]};
    assign in5192_2 = {c5160,s5177[1]};
    CLA_2 KS_5192(s5192, c5192, in5192_1, in5192_2);
    wire[0:0] s5193, in5193_1, in5193_2;
    wire c5193;
    assign in5193_1 = {c5161};
    assign in5193_2 = {c5162};
    Half_Adder KS_5193(s5193, c5193, in5193_1, in5193_2);
    wire[3:0] s5194, in5194_1, in5194_2;
    wire c5194;
    assign in5194_1 = {c5163,s5178[1],s3493[0],s3511[0]};
    assign in5194_2 = {c5171,s5179[1],s5175[2],s3512[0]};
    CLA_4 KS_5194(s5194, c5194, in5194_1, in5194_2);
    wire[0:0] s5195, in5195_1, in5195_2;
    wire c5195;
    assign in5195_1 = {s5175[0]};
    assign in5195_2 = {s5176[0]};
    Half_Adder KS_5195(s5195, c5195, in5195_1, in5195_2);
    wire[1:0] s5196, in5196_1, in5196_2;
    wire c5196;
    assign in5196_1 = {s5177[0],s5180[1]};
    assign in5196_2 = {s5178[0],s5181[1]};
    CLA_2 KS_5196(s5196, c5196, in5196_1, in5196_2);
    wire[0:0] s5197, in5197_1, in5197_2;
    wire c5197;
    assign in5197_1 = {s5180[0]};
    assign in5197_2 = {s5181[0]};
    Full_Adder KS_5197(s5197, c5197, in5197_1, in5197_2, s5179[0]);
    wire[3:0] s5198, in5198_1, in5198_2;
    wire c5198;
    assign in5198_1 = {s3488[3],s1331[0],s1333[0],s3520[0]};
    assign in5198_2 = {s3489[3],s1332[0],s1334[0],s3521[0]};
    CLA_4 KS_5198(s5198, c5198, in5198_1, in5198_2);
    wire[3:0] s5199, in5199_1, in5199_2;
    wire c5199;
    assign in5199_1 = {s3490[2],c3486,c3490,s3522[0]};
    assign in5199_2 = {s3491[2],c3487,c3491,s3523[0]};
    CLA_4 KS_5199(s5199, c5199, in5199_1, in5199_2);
    wire[3:0] s5200, in5200_1, in5200_2;
    wire c5200;
    assign in5200_1 = {s3492[2],c3488,c3492,s3524[0]};
    assign in5200_2 = {s3493[2],c3489,c3493,s3525[0]};
    CLA_4 KS_5200(s5200, c5200, in5200_1, in5200_2);
    wire[3:0] s5201, in5201_1, in5201_2;
    wire c5201;
    assign in5201_1 = {s3494[1],s3490[3],s3494[3],s3526[0]};
    assign in5201_2 = {s3495[1],s3491[3],s3495[3],s3527[0]};
    CLA_4 KS_5201(s5201, c5201, in5201_1, in5201_2);
    wire[3:0] s5202, in5202_1, in5202_2;
    wire c5202;
    assign in5202_1 = {s3496[1],s3492[3],s3496[3],s3528[0]};
    assign in5202_2 = {s3497[1],s3493[3],s3497[3],s3529[0]};
    CLA_4 KS_5202(s5202, c5202, in5202_1, in5202_2);
    wire[3:0] s5203, in5203_1, in5203_2;
    wire c5203;
    assign in5203_1 = {s3498[1],s3494[2],s3498[3],s3530[0]};
    assign in5203_2 = {s3499[1],s3495[2],s3499[3],s3531[0]};
    CLA_4 KS_5203(s5203, c5203, in5203_1, in5203_2);
    wire[3:0] s5204, in5204_1, in5204_2;
    wire c5204;
    assign in5204_1 = {s3500[1],s3496[2],s3500[3],s3532[0]};
    assign in5204_2 = {s3501[1],s3497[2],s3501[3],s3533[0]};
    CLA_4 KS_5204(s5204, c5204, in5204_1, in5204_2);
    wire[3:0] s5205, in5205_1, in5205_2;
    wire c5205;
    assign in5205_1 = {s3502[1],s3498[2],s3502[3],s3534[0]};
    assign in5205_2 = {s3503[1],s3499[2],s3503[3],s3535[0]};
    CLA_4 KS_5205(s5205, c5205, in5205_1, in5205_2);
    wire[3:0] s5206, in5206_1, in5206_2;
    wire c5206;
    assign in5206_1 = {s3504[1],s3500[2],s3504[3],s3536[0]};
    assign in5206_2 = {s3505[1],s3501[2],s3505[3],s3537[0]};
    CLA_4 KS_5206(s5206, c5206, in5206_1, in5206_2);
    wire[3:0] s5207, in5207_1, in5207_2;
    wire c5207;
    assign in5207_1 = {c3506,s3502[2],s3507[3],s3538[0]};
    assign in5207_2 = {s3507[1],s3503[2],s3509[3],s3539[0]};
    CLA_4 KS_5207(s5207, c5207, in5207_1, in5207_2);
    wire[3:0] s5208, in5208_1, in5208_2;
    wire c5208;
    assign in5208_1 = {c3508,s3504[2],s3511[3],s3540[0]};
    assign in5208_2 = {s3509[1],s3505[2],s3513[3],s3541[0]};
    CLA_4 KS_5208(s5208, c5208, in5208_1, in5208_2);
    wire[3:0] s5209, in5209_1, in5209_2;
    wire c5209;
    assign in5209_1 = {c3510,s3507[2],s3514[1],s3542[0]};
    assign in5209_2 = {s3511[1],s3509[2],s3515[0],s3543[0]};
    CLA_4 KS_5209(s5209, c5209, in5209_1, in5209_2);
    wire[0:0] s5210, in5210_1, in5210_2;
    wire c5210;
    assign in5210_1 = {c3512};
    assign in5210_2 = {s3513[1]};
    Half_Adder KS_5210(s5210, c5210, in5210_1, in5210_2);
    wire[1:0] s5211, in5211_1, in5211_2;
    wire c5211;
    assign in5211_1 = {c5175,s3511[2]};
    assign in5211_2 = {c5176,s3513[2]};
    CLA_2 KS_5211(s5211, c5211, in5211_1, in5211_2);
    wire[0:0] s5212, in5212_1, in5212_2;
    wire c5212;
    assign in5212_1 = {c5177};
    assign in5212_2 = {c5178};
    Half_Adder KS_5212(s5212, c5212, in5212_1, in5212_2);
    wire[2:0] s5213, in5213_1, in5213_2;
    wire c5213;
    assign in5213_1 = {c5179,s3514[0],s3516[0]};
    assign in5213_2 = {c5180,s5198[1],s3517[0]};
    CLA_3 KS_5213(s5213, c5213, in5213_1, in5213_2);
    wire[0:0] s5214, in5214_1, in5214_2;
    wire c5214;
    assign in5214_1 = {c5181};
    assign in5214_2 = {c5182};
    Half_Adder KS_5214(s5214, c5214, in5214_1, in5214_2);
    wire[1:0] s5215, in5215_1, in5215_2;
    wire c5215;
    assign in5215_1 = {c5183,s5199[1]};
    assign in5215_2 = {c5184,s5200[1]};
    CLA_2 KS_5215(s5215, c5215, in5215_1, in5215_2);
    wire[0:0] s5216, in5216_1, in5216_2;
    wire c5216;
    assign in5216_1 = {c5185};
    assign in5216_2 = {c5186};
    Half_Adder KS_5216(s5216, c5216, in5216_1, in5216_2);
    wire[3:0] s5217, in5217_1, in5217_2;
    wire c5217;
    assign in5217_1 = {c5194,s5201[1],s3518[0],s3544[0]};
    assign in5217_2 = {s5198[0],s5202[1],s5198[2],s3545[0]};
    CLA_4 KS_5217(s5217, c5217, in5217_1, in5217_2);
    wire[0:0] s5218, in5218_1, in5218_2;
    wire c5218;
    assign in5218_1 = {s5199[0]};
    assign in5218_2 = {s5200[0]};
    Half_Adder KS_5218(s5218, c5218, in5218_1, in5218_2);
    wire[1:0] s5219, in5219_1, in5219_2;
    wire c5219;
    assign in5219_1 = {s5202[0],s5203[1]};
    assign in5219_2 = {s5203[0],s5204[1]};
    CLA_2_c KS_5219(s5219, c5219, in5219_1, in5219_2, s5201[0]);
    wire[3:0] s5220, in5220_1, in5220_2;
    wire c5220;
    assign in5220_1 = {s3521[1],s1342[0],s1344[0],s3555[0]};
    assign in5220_2 = {s3522[1],c3514,s1345[0],s3556[0]};
    CLA_4 KS_5220(s5220, c5220, in5220_1, in5220_2);
    wire[3:0] s5221, in5221_1, in5221_2;
    wire c5221;
    assign in5221_1 = {s3523[1],s3515[3],c3515,s3557[0]};
    assign in5221_2 = {s3524[1],s3516[3],c3516,s3558[0]};
    CLA_4 KS_5221(s5221, c5221, in5221_1, in5221_2);
    wire[3:0] s5222, in5222_1, in5222_2;
    wire c5222;
    assign in5222_1 = {s3525[1],s3517[3],c3517,s3559[0]};
    assign in5222_2 = {s3526[1],s3518[3],c3518,s3560[0]};
    CLA_4 KS_5222(s5222, c5222, in5222_1, in5222_2);
    wire[3:0] s5223, in5223_1, in5223_2;
    wire c5223;
    assign in5223_1 = {s3527[1],s3519[2],s3519[3],s3561[0]};
    assign in5223_2 = {s3528[1],s3520[2],s3520[3],s3562[0]};
    CLA_4 KS_5223(s5223, c5223, in5223_1, in5223_2);
    wire[3:0] s5224, in5224_1, in5224_2;
    wire c5224;
    assign in5224_1 = {s3529[1],s3521[2],s3521[3],s3563[0]};
    assign in5224_2 = {s3530[1],s3522[2],s3522[3],s3564[0]};
    CLA_4 KS_5224(s5224, c5224, in5224_1, in5224_2);
    wire[3:0] s5225, in5225_1, in5225_2;
    wire c5225;
    assign in5225_1 = {s3531[1],s3523[2],s3523[3],s3565[0]};
    assign in5225_2 = {s3532[1],s3524[2],s3524[3],s3566[0]};
    CLA_4 KS_5225(s5225, c5225, in5225_1, in5225_2);
    wire[3:0] s5226, in5226_1, in5226_2;
    wire c5226;
    assign in5226_1 = {c3533,s3525[2],s3525[3],s3567[0]};
    assign in5226_2 = {s3534[1],s3526[2],s3526[3],s3568[0]};
    CLA_4 KS_5226(s5226, c5226, in5226_1, in5226_2);
    wire[3:0] s5227, in5227_1, in5227_2;
    wire c5227;
    assign in5227_1 = {c3535,s3527[2],s3527[3],s3569[0]};
    assign in5227_2 = {s3536[1],s3528[2],s3528[3],s3570[0]};
    CLA_4 KS_5227(s5227, c5227, in5227_1, in5227_2);
    wire[3:0] s5228, in5228_1, in5228_2;
    wire c5228;
    assign in5228_1 = {c3537,s3529[2],s3529[3],s3571[0]};
    assign in5228_2 = {s3538[1],s3530[2],s3530[3],s3572[0]};
    CLA_4 KS_5228(s5228, c5228, in5228_1, in5228_2);
    wire[3:0] s5229, in5229_1, in5229_2;
    wire c5229;
    assign in5229_1 = {c3539,s3531[2],s3531[3],s3573[0]};
    assign in5229_2 = {s3540[1],s3532[2],s3532[3],s3574[0]};
    CLA_4 KS_5229(s5229, c5229, in5229_1, in5229_2);
    wire[3:0] s5230, in5230_1, in5230_2;
    wire c5230;
    assign in5230_1 = {c3541,s3534[2],s3534[3],s3575[0]};
    assign in5230_2 = {s3542[1],s3536[2],s3536[3],s3576[0]};
    CLA_4 KS_5230(s5230, c5230, in5230_1, in5230_2);
    wire[3:0] s5231, in5231_1, in5231_2;
    wire c5231;
    assign in5231_1 = {c3543,c3538,s3540[3],s3577[0]};
    assign in5231_2 = {s3544[1],s3540[2],s3544[3],s3578[0]};
    CLA_4 KS_5231(s5231, c5231, in5231_1, in5231_2);
    wire[0:0] s5232, in5232_1, in5232_2;
    wire c5232;
    assign in5232_1 = {c3545};
    assign in5232_2 = {s3546[1]};
    Half_Adder KS_5232(s5232, c5232, in5232_1, in5232_2);
    wire[1:0] s5233, in5233_1, in5233_2;
    wire c5233;
    assign in5233_1 = {c5198,c3542};
    assign in5233_2 = {c5199,s3544[2]};
    CLA_2 KS_5233(s5233, c5233, in5233_1, in5233_2);
    wire[0:0] s5234, in5234_1, in5234_2;
    wire c5234;
    assign in5234_1 = {c5200};
    assign in5234_2 = {c5201};
    Half_Adder KS_5234(s5234, c5234, in5234_1, in5234_2);
    wire[2:0] s5235, in5235_1, in5235_2;
    wire c5235;
    assign in5235_1 = {c5202,c3546,s3547[0]};
    assign in5235_2 = {c5203,s5220[1],s3548[0]};
    CLA_3 KS_5235(s5235, c5235, in5235_1, in5235_2);
    wire[0:0] s5236, in5236_1, in5236_2;
    wire c5236;
    assign in5236_1 = {c5204};
    assign in5236_2 = {c5205};
    Half_Adder KS_5236(s5236, c5236, in5236_1, in5236_2);
    wire[1:0] s5237, in5237_1, in5237_2;
    wire c5237;
    assign in5237_1 = {c5206,s5221[1]};
    assign in5237_2 = {c5207,s5222[1]};
    CLA_2 KS_5237(s5237, c5237, in5237_1, in5237_2);
    wire[0:0] s5238, in5238_1, in5238_2;
    wire c5238;
    assign in5238_1 = {c5208};
    assign in5238_2 = {c5209};
    Half_Adder KS_5238(s5238, c5238, in5238_1, in5238_2);
    wire[3:0] s5239, in5239_1, in5239_2;
    wire c5239;
    assign in5239_1 = {c5217,s5223[1],s3549[0],s3579[0]};
    assign in5239_2 = {s5220[0],s5224[1],s5220[2],s3580[0]};
    CLA_4 KS_5239(s5239, c5239, in5239_1, in5239_2);
    wire[0:0] s5240, in5240_1, in5240_2;
    wire c5240;
    assign in5240_1 = {s5221[0]};
    assign in5240_2 = {s5222[0]};
    Half_Adder KS_5240(s5240, c5240, in5240_1, in5240_2);
    wire[1:0] s5241, in5241_1, in5241_2;
    wire c5241;
    assign in5241_1 = {s5224[0],s5225[1]};
    assign in5241_2 = {s5225[0],s5226[1]};
    CLA_2_c KS_5241(s5241, c5241, in5241_1, in5241_2, s5223[0]);
    wire[3:0] s5242, in5242_1, in5242_2;
    wire c5242;
    assign in5242_1 = {s3556[1],s3548[3],s1359[0],s3592[0]};
    assign in5242_2 = {s3557[1],s3549[3],s1360[0],s3593[0]};
    CLA_4 KS_5242(s5242, c5242, in5242_1, in5242_2);
    wire[3:0] s5243, in5243_1, in5243_2;
    wire c5243;
    assign in5243_1 = {s3558[1],s3550[2],s1361[0],s3594[0]};
    assign in5243_2 = {s3559[1],s3551[2],c3547,s3595[0]};
    CLA_4 KS_5243(s5243, c5243, in5243_1, in5243_2);
    wire[3:0] s5244, in5244_1, in5244_2;
    wire c5244;
    assign in5244_1 = {s3560[1],s3552[2],c3548,s3596[0]};
    assign in5244_2 = {s3561[1],s3553[2],c3549,s3597[0]};
    CLA_4 KS_5244(s5244, c5244, in5244_1, in5244_2);
    wire[3:0] s5245, in5245_1, in5245_2;
    wire c5245;
    assign in5245_1 = {s3562[1],s3554[2],s3550[3],s3598[0]};
    assign in5245_2 = {s3563[1],s3555[2],s3551[3],s3599[0]};
    CLA_4 KS_5245(s5245, c5245, in5245_1, in5245_2);
    wire[3:0] s5246, in5246_1, in5246_2;
    wire c5246;
    assign in5246_1 = {s3564[1],s3556[2],s3552[3],s3600[0]};
    assign in5246_2 = {s3565[1],s3557[2],s3553[3],s3601[0]};
    CLA_4 KS_5246(s5246, c5246, in5246_1, in5246_2);
    wire[3:0] s5247, in5247_1, in5247_2;
    wire c5247;
    assign in5247_1 = {c3566,s3558[2],s3554[3],s3602[0]};
    assign in5247_2 = {s3567[1],s3559[2],s3555[3],s3603[0]};
    CLA_4 KS_5247(s5247, c5247, in5247_1, in5247_2);
    wire[3:0] s5248, in5248_1, in5248_2;
    wire c5248;
    assign in5248_1 = {c3568,s3560[2],s3556[3],s3604[0]};
    assign in5248_2 = {s3569[1],s3561[2],s3557[3],s3605[0]};
    CLA_4 KS_5248(s5248, c5248, in5248_1, in5248_2);
    wire[3:0] s5249, in5249_1, in5249_2;
    wire c5249;
    assign in5249_1 = {c3570,s3562[2],s3558[3],s3606[0]};
    assign in5249_2 = {s3571[1],s3563[2],s3559[3],s3607[0]};
    CLA_4 KS_5249(s5249, c5249, in5249_1, in5249_2);
    wire[3:0] s5250, in5250_1, in5250_2;
    wire c5250;
    assign in5250_1 = {c3572,s3564[2],s3560[3],s3608[0]};
    assign in5250_2 = {s3573[1],s3565[2],s3561[3],s3609[0]};
    CLA_4 KS_5250(s5250, c5250, in5250_1, in5250_2);
    wire[3:0] s5251, in5251_1, in5251_2;
    wire c5251;
    assign in5251_1 = {c3574,c3567,s3562[3],s3610[0]};
    assign in5251_2 = {s3575[1],s3569[2],s3563[3],s3611[0]};
    CLA_4 KS_5251(s5251, c5251, in5251_1, in5251_2);
    wire[3:0] s5252, in5252_1, in5252_2;
    wire c5252;
    assign in5252_1 = {c3576,c3571,s3564[3],s3612[0]};
    assign in5252_2 = {s3577[1],s3573[2],s3565[3],s3613[0]};
    CLA_4 KS_5252(s5252, c5252, in5252_1, in5252_2);
    wire[0:0] s5253, in5253_1, in5253_2;
    wire c5253;
    assign in5253_1 = {c3578};
    assign in5253_2 = {s3579[1]};
    Half_Adder KS_5253(s5253, c5253, in5253_1, in5253_2);
    wire[3:0] s5254, in5254_1, in5254_2;
    wire c5254;
    assign in5254_1 = {c3580,c3575,s3569[3],s3614[0]};
    assign in5254_2 = {s3581[1],s3577[2],s3573[3],s3615[0]};
    CLA_4 KS_5254(s5254, c5254, in5254_1, in5254_2);
    wire[0:0] s5255, in5255_1, in5255_2;
    wire c5255;
    assign in5255_1 = {c5220};
    assign in5255_2 = {c5221};
    Half_Adder KS_5255(s5255, c5255, in5255_1, in5255_2);
    wire[1:0] s5256, in5256_1, in5256_2;
    wire c5256;
    assign in5256_1 = {c5222,c3579};
    assign in5256_2 = {c5223,s3581[2]};
    CLA_2 KS_5256(s5256, c5256, in5256_1, in5256_2);
    wire[0:0] s5257, in5257_1, in5257_2;
    wire c5257;
    assign in5257_1 = {c5224};
    assign in5257_2 = {c5225};
    Half_Adder KS_5257(s5257, c5257, in5257_1, in5257_2);
    wire[2:0] s5258, in5258_1, in5258_2;
    wire c5258;
    assign in5258_1 = {c5226,s5242[1],s3577[3]};
    assign in5258_2 = {c5227,s5243[1],s3581[3]};
    CLA_3 KS_5258(s5258, c5258, in5258_1, in5258_2);
    wire[0:0] s5259, in5259_1, in5259_2;
    wire c5259;
    assign in5259_1 = {c5228};
    assign in5259_2 = {c5229};
    Half_Adder KS_5259(s5259, c5259, in5259_1, in5259_2);
    wire[1:0] s5260, in5260_1, in5260_2;
    wire c5260;
    assign in5260_1 = {c5230,s5244[1]};
    assign in5260_2 = {c5231,s5245[1]};
    CLA_2 KS_5260(s5260, c5260, in5260_1, in5260_2);
    wire[0:0] s5261, in5261_1, in5261_2;
    wire c5261;
    assign in5261_1 = {c5239};
    assign in5261_2 = {s5242[0]};
    Half_Adder KS_5261(s5261, c5261, in5261_1, in5261_2);
    wire[3:0] s5262, in5262_1, in5262_2;
    wire c5262;
    assign in5262_1 = {s5243[0],s5246[1],s3582[0],s3616[0]};
    assign in5262_2 = {s5244[0],s5247[1],s5242[2],s3617[0]};
    CLA_4 KS_5262(s5262, c5262, in5262_1, in5262_2);
    wire[0:0] s5263, in5263_1, in5263_2;
    wire c5263;
    assign in5263_1 = {s5246[0]};
    assign in5263_2 = {s5247[0]};
    Full_Adder KS_5263(s5263, c5263, in5263_1, in5263_2, s5245[0]);
    wire[3:0] s5264, in5264_1, in5264_2;
    wire c5264;
    assign in5264_1 = {s3593[1],s3583[2],s1380[1],s3630[0]};
    assign in5264_2 = {s3594[1],s3584[2],s1381[1],s3631[0]};
    CLA_4 KS_5264(s5264, c5264, in5264_1, in5264_2);
    wire[3:0] s5265, in5265_1, in5265_2;
    wire c5265;
    assign in5265_1 = {s3595[1],s3585[2],s1382[0],s3632[0]};
    assign in5265_2 = {s3596[1],s3586[2],c3582,s3633[0]};
    CLA_4 KS_5265(s5265, c5265, in5265_1, in5265_2);
    wire[3:0] s5266, in5266_1, in5266_2;
    wire c5266;
    assign in5266_1 = {s3597[1],s3587[2],s3583[3],s3634[0]};
    assign in5266_2 = {s3598[1],s3588[2],s3584[3],s3635[0]};
    CLA_4 KS_5266(s5266, c5266, in5266_1, in5266_2);
    wire[3:0] s5267, in5267_1, in5267_2;
    wire c5267;
    assign in5267_1 = {s3599[1],s3589[2],s3585[3],s3636[0]};
    assign in5267_2 = {s3600[1],s3590[2],s3586[3],s3637[0]};
    CLA_4 KS_5267(s5267, c5267, in5267_1, in5267_2);
    wire[3:0] s5268, in5268_1, in5268_2;
    wire c5268;
    assign in5268_1 = {c3601,s3591[2],s3587[3],s3638[0]};
    assign in5268_2 = {s3602[1],s3592[2],s3588[3],s3639[0]};
    CLA_4 KS_5268(s5268, c5268, in5268_1, in5268_2);
    wire[3:0] s5269, in5269_1, in5269_2;
    wire c5269;
    assign in5269_1 = {c3603,s3593[2],s3589[3],s3640[0]};
    assign in5269_2 = {s3604[1],s3594[2],s3590[3],s3641[0]};
    CLA_4 KS_5269(s5269, c5269, in5269_1, in5269_2);
    wire[3:0] s5270, in5270_1, in5270_2;
    wire c5270;
    assign in5270_1 = {c3605,s3595[2],s3591[3],s3642[0]};
    assign in5270_2 = {s3606[1],s3596[2],s3592[3],s3643[0]};
    CLA_4 KS_5270(s5270, c5270, in5270_1, in5270_2);
    wire[3:0] s5271, in5271_1, in5271_2;
    wire c5271;
    assign in5271_1 = {c3607,s3597[2],s3593[3],s3644[0]};
    assign in5271_2 = {s3608[1],s3598[2],s3594[3],s3645[0]};
    CLA_4 KS_5271(s5271, c5271, in5271_1, in5271_2);
    wire[3:0] s5272, in5272_1, in5272_2;
    wire c5272;
    assign in5272_1 = {c3609,s3599[2],s3595[3],s3646[0]};
    assign in5272_2 = {s3610[1],s3600[2],s3596[3],s3647[0]};
    CLA_4 KS_5272(s5272, c5272, in5272_1, in5272_2);
    wire[3:0] s5273, in5273_1, in5273_2;
    wire c5273;
    assign in5273_1 = {c3611,c3602,s3597[3],s3648[0]};
    assign in5273_2 = {s3612[1],s3604[2],s3598[3],s3649[0]};
    CLA_4 KS_5273(s5273, c5273, in5273_1, in5273_2);
    wire[3:0] s5274, in5274_1, in5274_2;
    wire c5274;
    assign in5274_1 = {c3613,c3606,s3599[3],s3650[0]};
    assign in5274_2 = {s3614[1],s3608[2],s3600[3],s3651[0]};
    CLA_4 KS_5274(s5274, c5274, in5274_1, in5274_2);
    wire[1:0] s5275, in5275_1, in5275_2;
    wire c5275;
    assign in5275_1 = {c3615,c3610};
    assign in5275_2 = {s3616[1],s3612[2]};
    CLA_2 KS_5275(s5275, c5275, in5275_1, in5275_2);
    wire[0:0] s5276, in5276_1, in5276_2;
    wire c5276;
    assign in5276_1 = {c3617};
    assign in5276_2 = {s3618[1]};
    Half_Adder KS_5276(s5276, c5276, in5276_1, in5276_2);
    wire[3:0] s5277, in5277_1, in5277_2;
    wire c5277;
    assign in5277_1 = {c5242,c3614,s3604[3],s3652[0]};
    assign in5277_2 = {c5243,s3616[2],s3608[3],s3653[0]};
    CLA_4 KS_5277(s5277, c5277, in5277_1, in5277_2);
    wire[0:0] s5278, in5278_1, in5278_2;
    wire c5278;
    assign in5278_1 = {c5244};
    assign in5278_2 = {c5245};
    Half_Adder KS_5278(s5278, c5278, in5278_1, in5278_2);
    wire[1:0] s5279, in5279_1, in5279_2;
    wire c5279;
    assign in5279_1 = {c5246,c3618};
    assign in5279_2 = {c5247,s5264[1]};
    CLA_2 KS_5279(s5279, c5279, in5279_1, in5279_2);
    wire[0:0] s5280, in5280_1, in5280_2;
    wire c5280;
    assign in5280_1 = {c5248};
    assign in5280_2 = {c5249};
    Half_Adder KS_5280(s5280, c5280, in5280_1, in5280_2);
    wire[2:0] s5281, in5281_1, in5281_2;
    wire c5281;
    assign in5281_1 = {c5250,s5265[1],c3612};
    assign in5281_2 = {c5251,s5266[1],s3616[3]};
    CLA_3 KS_5281(s5281, c5281, in5281_1, in5281_2);
    wire[0:0] s5282, in5282_1, in5282_2;
    wire c5282;
    assign in5282_1 = {c5252};
    assign in5282_2 = {c5254};
    Half_Adder KS_5282(s5282, c5282, in5282_1, in5282_2);
    wire[1:0] s5283, in5283_1, in5283_2;
    wire c5283;
    assign in5283_1 = {c5262,s5267[1]};
    assign in5283_2 = {s5264[0],s5268[1]};
    CLA_2 KS_5283(s5283, c5283, in5283_1, in5283_2);
    wire[0:0] s5284, in5284_1, in5284_2;
    wire c5284;
    assign in5284_1 = {s5265[0]};
    assign in5284_2 = {s5266[0]};
    Half_Adder KS_5284(s5284, c5284, in5284_1, in5284_2);
    wire[3:0] s5285, in5285_1, in5285_2;
    wire c5285;
    assign in5285_1 = {s5268[0],s5269[1],s5264[2],s3654[0]};
    assign in5285_2 = {s5269[0],s5270[1],s5265[2],s3655[0]};
    CLA_4_c KS_5285(s5285, c5285, in5285_1, in5285_2, s5267[0]);
    wire[3:0] s5286, in5286_1, in5286_2;
    wire c5286;
    assign in5286_1 = {s3630[1],s3620[2],c1411,s3668[0]};
    assign in5286_2 = {s3631[1],s3621[2],s1412[1],s3669[0]};
    CLA_4 KS_5286(s5286, c5286, in5286_1, in5286_2);
    wire[3:0] s5287, in5287_1, in5287_2;
    wire c5287;
    assign in5287_1 = {s3632[1],s3622[2],c1413,s3670[0]};
    assign in5287_2 = {s3633[1],s3623[2],s3619[3],s3671[0]};
    CLA_4 KS_5287(s5287, c5287, in5287_1, in5287_2);
    wire[3:0] s5288, in5288_1, in5288_2;
    wire c5288;
    assign in5288_1 = {s3634[1],s3624[2],s3620[3],s3672[0]};
    assign in5288_2 = {s3635[1],s3625[2],s3621[3],s3673[0]};
    CLA_4 KS_5288(s5288, c5288, in5288_1, in5288_2);
    wire[3:0] s5289, in5289_1, in5289_2;
    wire c5289;
    assign in5289_1 = {s3636[1],s3626[2],s3622[3],s3674[0]};
    assign in5289_2 = {s3637[1],s3627[2],s3623[3],s3675[0]};
    CLA_4 KS_5289(s5289, c5289, in5289_1, in5289_2);
    wire[3:0] s5290, in5290_1, in5290_2;
    wire c5290;
    assign in5290_1 = {c3638,s3628[2],s3624[3],s3676[0]};
    assign in5290_2 = {s3639[1],s3629[2],s3625[3],s3677[0]};
    CLA_4 KS_5290(s5290, c5290, in5290_1, in5290_2);
    wire[3:0] s5291, in5291_1, in5291_2;
    wire c5291;
    assign in5291_1 = {c3640,s3630[2],s3626[3],s3678[0]};
    assign in5291_2 = {s3641[1],s3631[2],s3627[3],s3679[0]};
    CLA_4 KS_5291(s5291, c5291, in5291_1, in5291_2);
    wire[3:0] s5292, in5292_1, in5292_2;
    wire c5292;
    assign in5292_1 = {c3642,s3632[2],s3628[3],s3680[0]};
    assign in5292_2 = {s3643[1],s3633[2],s3629[3],s3681[0]};
    CLA_4 KS_5292(s5292, c5292, in5292_1, in5292_2);
    wire[3:0] s5293, in5293_1, in5293_2;
    wire c5293;
    assign in5293_1 = {c3644,s3634[2],s3630[3],s3682[0]};
    assign in5293_2 = {s3645[1],s3635[2],s3631[3],s3683[0]};
    CLA_4 KS_5293(s5293, c5293, in5293_1, in5293_2);
    wire[3:0] s5294, in5294_1, in5294_2;
    wire c5294;
    assign in5294_1 = {c3646,s3636[2],s3632[3],s3684[0]};
    assign in5294_2 = {s3647[1],s3637[2],s3633[3],s3685[0]};
    CLA_4 KS_5294(s5294, c5294, in5294_1, in5294_2);
    wire[3:0] s5295, in5295_1, in5295_2;
    wire c5295;
    assign in5295_1 = {c3648,c3639,s3634[3],s3686[0]};
    assign in5295_2 = {s3649[1],s3641[2],s3635[3],s3687[0]};
    CLA_4 KS_5295(s5295, c5295, in5295_1, in5295_2);
    wire[3:0] s5296, in5296_1, in5296_2;
    wire c5296;
    assign in5296_1 = {c3650,c3643,s3636[3],s3688[0]};
    assign in5296_2 = {s3651[1],s3645[2],s3637[3],s3689[0]};
    CLA_4 KS_5296(s5296, c5296, in5296_1, in5296_2);
    wire[1:0] s5297, in5297_1, in5297_2;
    wire c5297;
    assign in5297_1 = {c3652,c3647};
    assign in5297_2 = {s3653[1],s3649[2]};
    CLA_2 KS_5297(s5297, c5297, in5297_1, in5297_2);
    wire[0:0] s5298, in5298_1, in5298_2;
    wire c5298;
    assign in5298_1 = {c3654};
    assign in5298_2 = {s3655[1]};
    Half_Adder KS_5298(s5298, c5298, in5298_1, in5298_2);
    wire[3:0] s5299, in5299_1, in5299_2;
    wire c5299;
    assign in5299_1 = {c3656,c3651,c3641,s3690[0]};
    assign in5299_2 = {c5264,s3653[2],s3645[3],s3691[0]};
    CLA_4 KS_5299(s5299, c5299, in5299_1, in5299_2);
    wire[0:0] s5300, in5300_1, in5300_2;
    wire c5300;
    assign in5300_1 = {c5265};
    assign in5300_2 = {c5266};
    Half_Adder KS_5300(s5300, c5300, in5300_1, in5300_2);
    wire[1:0] s5301, in5301_1, in5301_2;
    wire c5301;
    assign in5301_1 = {c5267,c3655};
    assign in5301_2 = {c5268,s5286[1]};
    CLA_2 KS_5301(s5301, c5301, in5301_1, in5301_2);
    wire[0:0] s5302, in5302_1, in5302_2;
    wire c5302;
    assign in5302_1 = {c5269};
    assign in5302_2 = {c5270};
    Half_Adder KS_5302(s5302, c5302, in5302_1, in5302_2);
    wire[2:0] s5303, in5303_1, in5303_2;
    wire c5303;
    assign in5303_1 = {c5271,s5287[1],c3649};
    assign in5303_2 = {c5272,s5288[1],s3653[3]};
    CLA_3 KS_5303(s5303, c5303, in5303_1, in5303_2);
    wire[0:0] s5304, in5304_1, in5304_2;
    wire c5304;
    assign in5304_1 = {c5273};
    assign in5304_2 = {c5274};
    Half_Adder KS_5304(s5304, c5304, in5304_1, in5304_2);
    wire[1:0] s5305, in5305_1, in5305_2;
    wire c5305;
    assign in5305_1 = {c5277,s5289[1]};
    assign in5305_2 = {c5285,s5290[1]};
    CLA_2 KS_5305(s5305, c5305, in5305_1, in5305_2);
    wire[0:0] s5306, in5306_1, in5306_2;
    wire c5306;
    assign in5306_1 = {s5286[0]};
    assign in5306_2 = {s5287[0]};
    Half_Adder KS_5306(s5306, c5306, in5306_1, in5306_2);
    wire[3:0] s5307, in5307_1, in5307_2;
    wire c5307;
    assign in5307_1 = {s5288[0],s5291[1],s5286[2],s3692[0]};
    assign in5307_2 = {s5289[0],s5292[1],s5287[2],s3693[0]};
    CLA_4 KS_5307(s5307, c5307, in5307_1, in5307_2);
    wire[0:0] s5308, in5308_1, in5308_2;
    wire c5308;
    assign in5308_1 = {s5291[0]};
    assign in5308_2 = {s5292[0]};
    Full_Adder KS_5308(s5308, c5308, in5308_1, in5308_2, s5290[0]);
    wire[3:0] s5309, in5309_1, in5309_2;
    wire c5309;
    assign in5309_1 = {s3668[1],s3658[2],c1451,s3705[0]};
    assign in5309_2 = {s3669[1],s3659[2],s1452[1],s3706[0]};
    CLA_4 KS_5309(s5309, c5309, in5309_1, in5309_2);
    wire[3:0] s5310, in5310_1, in5310_2;
    wire c5310;
    assign in5310_1 = {s3670[1],s3660[2],c1453,s3707[0]};
    assign in5310_2 = {s3671[1],s3661[2],s1454[1],s3708[0]};
    CLA_4 KS_5310(s5310, c5310, in5310_1, in5310_2);
    wire[3:0] s5311, in5311_1, in5311_2;
    wire c5311;
    assign in5311_1 = {s3672[1],s3662[2],s3657[3],s3709[0]};
    assign in5311_2 = {s3673[1],s3663[2],s3658[3],s3710[0]};
    CLA_4 KS_5311(s5311, c5311, in5311_1, in5311_2);
    wire[3:0] s5312, in5312_1, in5312_2;
    wire c5312;
    assign in5312_1 = {s3674[1],s3664[2],s3659[3],s3711[0]};
    assign in5312_2 = {s3675[1],s3665[2],s3660[3],s3712[0]};
    CLA_4 KS_5312(s5312, c5312, in5312_1, in5312_2);
    wire[3:0] s5313, in5313_1, in5313_2;
    wire c5313;
    assign in5313_1 = {c3676,s3666[2],s3661[3],s3713[0]};
    assign in5313_2 = {s3677[1],s3667[2],s3662[3],s3714[0]};
    CLA_4 KS_5313(s5313, c5313, in5313_1, in5313_2);
    wire[3:0] s5314, in5314_1, in5314_2;
    wire c5314;
    assign in5314_1 = {c3678,s3668[2],s3663[3],s3715[0]};
    assign in5314_2 = {s3679[1],s3669[2],s3664[3],s3716[0]};
    CLA_4 KS_5314(s5314, c5314, in5314_1, in5314_2);
    wire[3:0] s5315, in5315_1, in5315_2;
    wire c5315;
    assign in5315_1 = {c3680,s3670[2],s3665[3],s3717[0]};
    assign in5315_2 = {s3681[1],s3671[2],s3666[3],s3718[0]};
    CLA_4 KS_5315(s5315, c5315, in5315_1, in5315_2);
    wire[3:0] s5316, in5316_1, in5316_2;
    wire c5316;
    assign in5316_1 = {c3682,s3672[2],s3667[3],s3719[0]};
    assign in5316_2 = {s3683[1],s3673[2],s3668[3],s3720[0]};
    CLA_4 KS_5316(s5316, c5316, in5316_1, in5316_2);
    wire[3:0] s5317, in5317_1, in5317_2;
    wire c5317;
    assign in5317_1 = {c3684,s3674[2],s3669[3],s3721[0]};
    assign in5317_2 = {s3685[1],s3675[2],s3670[3],s3722[0]};
    CLA_4 KS_5317(s5317, c5317, in5317_1, in5317_2);
    wire[3:0] s5318, in5318_1, in5318_2;
    wire c5318;
    assign in5318_1 = {c3686,c3677,s3671[3],s3723[0]};
    assign in5318_2 = {s3687[1],s3679[2],s3672[3],s3724[0]};
    CLA_4 KS_5318(s5318, c5318, in5318_1, in5318_2);
    wire[3:0] s5319, in5319_1, in5319_2;
    wire c5319;
    assign in5319_1 = {c3688,c3681,s3673[3],s3725[0]};
    assign in5319_2 = {s3689[1],s3683[2],s3674[3],s3726[0]};
    CLA_4 KS_5319(s5319, c5319, in5319_1, in5319_2);
    wire[3:0] s5320, in5320_1, in5320_2;
    wire c5320;
    assign in5320_1 = {c3690,c3685,c3675,s3727[0]};
    assign in5320_2 = {s3691[1],s3687[2],s3679[3],s3728[0]};
    CLA_4 KS_5320(s5320, c5320, in5320_1, in5320_2);
    wire[0:0] s5321, in5321_1, in5321_2;
    wire c5321;
    assign in5321_1 = {c3692};
    assign in5321_2 = {s3693[1]};
    Half_Adder KS_5321(s5321, c5321, in5321_1, in5321_2);
    wire[1:0] s5322, in5322_1, in5322_2;
    wire c5322;
    assign in5322_1 = {c3694,c3689};
    assign in5322_2 = {c5286,s3691[2]};
    CLA_2 KS_5322(s5322, c5322, in5322_1, in5322_2);
    wire[0:0] s5323, in5323_1, in5323_2;
    wire c5323;
    assign in5323_1 = {c5287};
    assign in5323_2 = {c5288};
    Half_Adder KS_5323(s5323, c5323, in5323_1, in5323_2);
    wire[2:0] s5324, in5324_1, in5324_2;
    wire c5324;
    assign in5324_1 = {c5289,c3693,c3683};
    assign in5324_2 = {c5290,s5309[1],s3687[3]};
    CLA_3 KS_5324(s5324, c5324, in5324_1, in5324_2);
    wire[0:0] s5325, in5325_1, in5325_2;
    wire c5325;
    assign in5325_1 = {c5291};
    assign in5325_2 = {c5292};
    Half_Adder KS_5325(s5325, c5325, in5325_1, in5325_2);
    wire[1:0] s5326, in5326_1, in5326_2;
    wire c5326;
    assign in5326_1 = {c5293,s5310[1]};
    assign in5326_2 = {c5294,s5311[1]};
    CLA_2 KS_5326(s5326, c5326, in5326_1, in5326_2);
    wire[0:0] s5327, in5327_1, in5327_2;
    wire c5327;
    assign in5327_1 = {c5295};
    assign in5327_2 = {c5296};
    Half_Adder KS_5327(s5327, c5327, in5327_1, in5327_2);
    wire[3:0] s5328, in5328_1, in5328_2;
    wire c5328;
    assign in5328_1 = {c5299,s5312[1],c3691,s3729[0]};
    assign in5328_2 = {c5307,s5313[1],s5309[2],s3730[0]};
    CLA_4 KS_5328(s5328, c5328, in5328_1, in5328_2);
    wire[0:0] s5329, in5329_1, in5329_2;
    wire c5329;
    assign in5329_1 = {s5309[0]};
    assign in5329_2 = {s5310[0]};
    Half_Adder KS_5329(s5329, c5329, in5329_1, in5329_2);
    wire[1:0] s5330, in5330_1, in5330_2;
    wire c5330;
    assign in5330_1 = {s5311[0],s5314[1]};
    assign in5330_2 = {s5312[0],s5315[1]};
    CLA_2 KS_5330(s5330, c5330, in5330_1, in5330_2);
    wire[0:0] s5331, in5331_1, in5331_2;
    wire c5331;
    assign in5331_1 = {s5314[0]};
    assign in5331_2 = {s5315[0]};
    Full_Adder KS_5331(s5331, c5331, in5331_1, in5331_2, s5313[0]);
    wire[3:0] s5332, in5332_1, in5332_2;
    wire c5332;
    assign in5332_1 = {s3706[1],s3696[2],c1502,s3742[0]};
    assign in5332_2 = {s3707[1],s3697[2],s1503[1],s3743[0]};
    CLA_4 KS_5332(s5332, c5332, in5332_1, in5332_2);
    wire[3:0] s5333, in5333_1, in5333_2;
    wire c5333;
    assign in5333_1 = {s3708[1],s3698[2],c1504,s3744[0]};
    assign in5333_2 = {s3709[1],s3699[2],s1505[1],s3745[0]};
    CLA_4 KS_5333(s5333, c5333, in5333_1, in5333_2);
    wire[3:0] s5334, in5334_1, in5334_2;
    wire c5334;
    assign in5334_1 = {s3710[1],s3700[2],s3695[3],s3746[0]};
    assign in5334_2 = {s3711[1],s3701[2],s3696[3],s3747[0]};
    CLA_4 KS_5334(s5334, c5334, in5334_1, in5334_2);
    wire[3:0] s5335, in5335_1, in5335_2;
    wire c5335;
    assign in5335_1 = {s3712[1],s3702[2],s3697[3],s3748[0]};
    assign in5335_2 = {s3713[1],s3703[2],s3698[3],s3749[0]};
    CLA_4 KS_5335(s5335, c5335, in5335_1, in5335_2);
    wire[3:0] s5336, in5336_1, in5336_2;
    wire c5336;
    assign in5336_1 = {c3714,s3704[2],s3699[3],s3750[0]};
    assign in5336_2 = {s3715[1],s3705[2],s3700[3],s3751[0]};
    CLA_4 KS_5336(s5336, c5336, in5336_1, in5336_2);
    wire[3:0] s5337, in5337_1, in5337_2;
    wire c5337;
    assign in5337_1 = {c3716,s3706[2],s3701[3],s3752[0]};
    assign in5337_2 = {s3717[1],s3707[2],s3702[3],s3753[0]};
    CLA_4 KS_5337(s5337, c5337, in5337_1, in5337_2);
    wire[3:0] s5338, in5338_1, in5338_2;
    wire c5338;
    assign in5338_1 = {c3718,s3708[2],s3703[3],s3754[0]};
    assign in5338_2 = {s3719[1],s3709[2],s3704[3],s3755[0]};
    CLA_4 KS_5338(s5338, c5338, in5338_1, in5338_2);
    wire[3:0] s5339, in5339_1, in5339_2;
    wire c5339;
    assign in5339_1 = {c3720,s3710[2],s3705[3],s3756[0]};
    assign in5339_2 = {s3721[1],s3711[2],s3706[3],s3757[0]};
    CLA_4 KS_5339(s5339, c5339, in5339_1, in5339_2);
    wire[3:0] s5340, in5340_1, in5340_2;
    wire c5340;
    assign in5340_1 = {c3722,s3712[2],s3707[3],s3758[0]};
    assign in5340_2 = {s3723[1],s3713[2],s3708[3],s3759[0]};
    CLA_4 KS_5340(s5340, c5340, in5340_1, in5340_2);
    wire[3:0] s5341, in5341_1, in5341_2;
    wire c5341;
    assign in5341_1 = {c3724,c3715,s3709[3],s3760[0]};
    assign in5341_2 = {s3725[1],s3717[2],s3710[3],s3761[0]};
    CLA_4 KS_5341(s5341, c5341, in5341_1, in5341_2);
    wire[3:0] s5342, in5342_1, in5342_2;
    wire c5342;
    assign in5342_1 = {c3726,c3719,s3711[3],s3762[0]};
    assign in5342_2 = {s3727[1],s3721[2],s3712[3],s3763[0]};
    CLA_4 KS_5342(s5342, c5342, in5342_1, in5342_2);
    wire[3:0] s5343, in5343_1, in5343_2;
    wire c5343;
    assign in5343_1 = {c3728,c3723,c3713,s3764[0]};
    assign in5343_2 = {s3729[1],s3725[2],s3717[3],s3765[0]};
    CLA_4 KS_5343(s5343, c5343, in5343_1, in5343_2);
    wire[0:0] s5344, in5344_1, in5344_2;
    wire c5344;
    assign in5344_1 = {c3730};
    assign in5344_2 = {s3731[1]};
    Half_Adder KS_5344(s5344, c5344, in5344_1, in5344_2);
    wire[1:0] s5345, in5345_1, in5345_2;
    wire c5345;
    assign in5345_1 = {c5309,c3727};
    assign in5345_2 = {c5310,s3729[2]};
    CLA_2 KS_5345(s5345, c5345, in5345_1, in5345_2);
    wire[0:0] s5346, in5346_1, in5346_2;
    wire c5346;
    assign in5346_1 = {c5311};
    assign in5346_2 = {c5312};
    Half_Adder KS_5346(s5346, c5346, in5346_1, in5346_2);
    wire[2:0] s5347, in5347_1, in5347_2;
    wire c5347;
    assign in5347_1 = {c5313,c3731,c3721};
    assign in5347_2 = {c5314,s5332[1],s3725[3]};
    CLA_3 KS_5347(s5347, c5347, in5347_1, in5347_2);
    wire[0:0] s5348, in5348_1, in5348_2;
    wire c5348;
    assign in5348_1 = {c5315};
    assign in5348_2 = {c5316};
    Half_Adder KS_5348(s5348, c5348, in5348_1, in5348_2);
    wire[1:0] s5349, in5349_1, in5349_2;
    wire c5349;
    assign in5349_1 = {c5317,s5333[1]};
    assign in5349_2 = {c5318,s5334[1]};
    CLA_2 KS_5349(s5349, c5349, in5349_1, in5349_2);
    wire[0:0] s5350, in5350_1, in5350_2;
    wire c5350;
    assign in5350_1 = {c5319};
    assign in5350_2 = {c5320};
    Half_Adder KS_5350(s5350, c5350, in5350_1, in5350_2);
    wire[3:0] s5351, in5351_1, in5351_2;
    wire c5351;
    assign in5351_1 = {c5328,s5335[1],c3729,s3766[0]};
    assign in5351_2 = {s5332[0],s5336[1],s5332[2],s3767[0]};
    CLA_4 KS_5351(s5351, c5351, in5351_1, in5351_2);
    wire[0:0] s5352, in5352_1, in5352_2;
    wire c5352;
    assign in5352_1 = {s5333[0]};
    assign in5352_2 = {s5334[0]};
    Half_Adder KS_5352(s5352, c5352, in5352_1, in5352_2);
    wire[1:0] s5353, in5353_1, in5353_2;
    wire c5353;
    assign in5353_1 = {s5336[0],s5337[1]};
    assign in5353_2 = {s5337[0],s5338[1]};
    CLA_2_c KS_5353(s5353, c5353, in5353_1, in5353_2, s5335[0]);
    wire[3:0] s5354, in5354_1, in5354_2;
    wire c5354;
    assign in5354_1 = {s3743[1],s3733[2],c1560,s3779[0]};
    assign in5354_2 = {s3744[1],s3734[2],s1561[1],s3780[0]};
    CLA_4 KS_5354(s5354, c5354, in5354_1, in5354_2);
    wire[3:0] s5355, in5355_1, in5355_2;
    wire c5355;
    assign in5355_1 = {s3745[1],s3735[2],c1562,s3781[0]};
    assign in5355_2 = {s3746[1],s3736[2],s1563[1],s3782[0]};
    CLA_4 KS_5355(s5355, c5355, in5355_1, in5355_2);
    wire[3:0] s5356, in5356_1, in5356_2;
    wire c5356;
    assign in5356_1 = {s3747[1],s3737[2],s3732[3],s3783[0]};
    assign in5356_2 = {s3748[1],s3738[2],s3733[3],s3784[0]};
    CLA_4 KS_5356(s5356, c5356, in5356_1, in5356_2);
    wire[3:0] s5357, in5357_1, in5357_2;
    wire c5357;
    assign in5357_1 = {s3749[1],s3739[2],s3734[3],s3785[0]};
    assign in5357_2 = {s3750[1],s3740[2],s3735[3],s3786[0]};
    CLA_4 KS_5357(s5357, c5357, in5357_1, in5357_2);
    wire[3:0] s5358, in5358_1, in5358_2;
    wire c5358;
    assign in5358_1 = {c3751,s3741[2],s3736[3],s3787[0]};
    assign in5358_2 = {s3752[1],s3742[2],s3737[3],s3788[0]};
    CLA_4 KS_5358(s5358, c5358, in5358_1, in5358_2);
    wire[3:0] s5359, in5359_1, in5359_2;
    wire c5359;
    assign in5359_1 = {c3753,s3743[2],s3738[3],s3789[0]};
    assign in5359_2 = {s3754[1],s3744[2],s3739[3],s3790[0]};
    CLA_4 KS_5359(s5359, c5359, in5359_1, in5359_2);
    wire[3:0] s5360, in5360_1, in5360_2;
    wire c5360;
    assign in5360_1 = {c3755,s3745[2],s3740[3],s3791[0]};
    assign in5360_2 = {s3756[1],s3746[2],s3741[3],s3792[0]};
    CLA_4 KS_5360(s5360, c5360, in5360_1, in5360_2);
    wire[3:0] s5361, in5361_1, in5361_2;
    wire c5361;
    assign in5361_1 = {c3757,s3747[2],s3742[3],s3793[0]};
    assign in5361_2 = {s3758[1],s3748[2],s3743[3],s3794[0]};
    CLA_4 KS_5361(s5361, c5361, in5361_1, in5361_2);
    wire[3:0] s5362, in5362_1, in5362_2;
    wire c5362;
    assign in5362_1 = {c3759,s3749[2],s3744[3],s3795[0]};
    assign in5362_2 = {s3760[1],s3750[2],s3745[3],s3796[0]};
    CLA_4 KS_5362(s5362, c5362, in5362_1, in5362_2);
    wire[3:0] s5363, in5363_1, in5363_2;
    wire c5363;
    assign in5363_1 = {c3761,c3752,s3746[3],s3797[0]};
    assign in5363_2 = {s3762[1],s3754[2],s3747[3],s3798[0]};
    CLA_4 KS_5363(s5363, c5363, in5363_1, in5363_2);
    wire[3:0] s5364, in5364_1, in5364_2;
    wire c5364;
    assign in5364_1 = {c3763,c3756,s3748[3],s3799[0]};
    assign in5364_2 = {s3764[1],s3758[2],s3749[3],s3800[0]};
    CLA_4 KS_5364(s5364, c5364, in5364_1, in5364_2);
    wire[3:0] s5365, in5365_1, in5365_2;
    wire c5365;
    assign in5365_1 = {c3765,c3760,c3750,s3801[0]};
    assign in5365_2 = {s3766[1],s3762[2],s3754[3],s3802[0]};
    CLA_4 KS_5365(s5365, c5365, in5365_1, in5365_2);
    wire[0:0] s5366, in5366_1, in5366_2;
    wire c5366;
    assign in5366_1 = {c3767};
    assign in5366_2 = {s3768[1]};
    Half_Adder KS_5366(s5366, c5366, in5366_1, in5366_2);
    wire[1:0] s5367, in5367_1, in5367_2;
    wire c5367;
    assign in5367_1 = {c5332,c3764};
    assign in5367_2 = {c5333,s3766[2]};
    CLA_2 KS_5367(s5367, c5367, in5367_1, in5367_2);
    wire[0:0] s5368, in5368_1, in5368_2;
    wire c5368;
    assign in5368_1 = {c5334};
    assign in5368_2 = {c5335};
    Half_Adder KS_5368(s5368, c5368, in5368_1, in5368_2);
    wire[2:0] s5369, in5369_1, in5369_2;
    wire c5369;
    assign in5369_1 = {c5336,c3768,c3758};
    assign in5369_2 = {c5337,s5354[1],s3762[3]};
    CLA_3 KS_5369(s5369, c5369, in5369_1, in5369_2);
    wire[0:0] s5370, in5370_1, in5370_2;
    wire c5370;
    assign in5370_1 = {c5338};
    assign in5370_2 = {c5339};
    Half_Adder KS_5370(s5370, c5370, in5370_1, in5370_2);
    wire[1:0] s5371, in5371_1, in5371_2;
    wire c5371;
    assign in5371_1 = {c5340,s5355[1]};
    assign in5371_2 = {c5341,s5356[1]};
    CLA_2 KS_5371(s5371, c5371, in5371_1, in5371_2);
    wire[0:0] s5372, in5372_1, in5372_2;
    wire c5372;
    assign in5372_1 = {c5342};
    assign in5372_2 = {c5343};
    Half_Adder KS_5372(s5372, c5372, in5372_1, in5372_2);
    wire[3:0] s5373, in5373_1, in5373_2;
    wire c5373;
    assign in5373_1 = {c5351,s5357[1],c3766,s3803[0]};
    assign in5373_2 = {s5354[0],s5358[1],s5354[2],s3804[0]};
    CLA_4 KS_5373(s5373, c5373, in5373_1, in5373_2);
    wire[0:0] s5374, in5374_1, in5374_2;
    wire c5374;
    assign in5374_1 = {s5355[0]};
    assign in5374_2 = {s5356[0]};
    Half_Adder KS_5374(s5374, c5374, in5374_1, in5374_2);
    wire[1:0] s5375, in5375_1, in5375_2;
    wire c5375;
    assign in5375_1 = {s5358[0],s5359[1]};
    assign in5375_2 = {s5359[0],s5360[1]};
    CLA_2_c KS_5375(s5375, c5375, in5375_1, in5375_2, s5357[0]);
    wire[3:0] s5376, in5376_1, in5376_2;
    wire c5376;
    assign in5376_1 = {s3780[1],s3770[2],c1618,s3816[0]};
    assign in5376_2 = {s3781[1],s3771[2],s1619[1],s3817[0]};
    CLA_4 KS_5376(s5376, c5376, in5376_1, in5376_2);
    wire[3:0] s5377, in5377_1, in5377_2;
    wire c5377;
    assign in5377_1 = {s3782[1],s3772[2],c1620,s3818[0]};
    assign in5377_2 = {s3783[1],s3773[2],s1621[1],s3819[0]};
    CLA_4 KS_5377(s5377, c5377, in5377_1, in5377_2);
    wire[3:0] s5378, in5378_1, in5378_2;
    wire c5378;
    assign in5378_1 = {s3784[1],s3774[2],s3769[3],s3820[0]};
    assign in5378_2 = {s3785[1],s3775[2],s3770[3],s3821[0]};
    CLA_4 KS_5378(s5378, c5378, in5378_1, in5378_2);
    wire[3:0] s5379, in5379_1, in5379_2;
    wire c5379;
    assign in5379_1 = {s3786[1],s3776[2],s3771[3],s3822[0]};
    assign in5379_2 = {s3787[1],s3777[2],s3772[3],s3823[0]};
    CLA_4 KS_5379(s5379, c5379, in5379_1, in5379_2);
    wire[3:0] s5380, in5380_1, in5380_2;
    wire c5380;
    assign in5380_1 = {c3788,s3778[2],s3773[3],s3824[0]};
    assign in5380_2 = {s3789[1],s3779[2],s3774[3],s3825[0]};
    CLA_4 KS_5380(s5380, c5380, in5380_1, in5380_2);
    wire[3:0] s5381, in5381_1, in5381_2;
    wire c5381;
    assign in5381_1 = {c3790,s3780[2],s3775[3],s3826[0]};
    assign in5381_2 = {s3791[1],s3781[2],s3776[3],s3827[0]};
    CLA_4 KS_5381(s5381, c5381, in5381_1, in5381_2);
    wire[3:0] s5382, in5382_1, in5382_2;
    wire c5382;
    assign in5382_1 = {c3792,s3782[2],s3777[3],s3828[0]};
    assign in5382_2 = {s3793[1],s3783[2],s3778[3],s3829[0]};
    CLA_4 KS_5382(s5382, c5382, in5382_1, in5382_2);
    wire[3:0] s5383, in5383_1, in5383_2;
    wire c5383;
    assign in5383_1 = {c3794,s3784[2],s3779[3],s3830[0]};
    assign in5383_2 = {s3795[1],s3785[2],s3780[3],s3831[0]};
    CLA_4 KS_5383(s5383, c5383, in5383_1, in5383_2);
    wire[3:0] s5384, in5384_1, in5384_2;
    wire c5384;
    assign in5384_1 = {c3796,s3786[2],s3781[3],s3832[0]};
    assign in5384_2 = {s3797[1],s3787[2],s3782[3],s3833[0]};
    CLA_4 KS_5384(s5384, c5384, in5384_1, in5384_2);
    wire[3:0] s5385, in5385_1, in5385_2;
    wire c5385;
    assign in5385_1 = {c3798,c3789,s3783[3],s3834[0]};
    assign in5385_2 = {s3799[1],s3791[2],s3784[3],s3835[0]};
    CLA_4 KS_5385(s5385, c5385, in5385_1, in5385_2);
    wire[3:0] s5386, in5386_1, in5386_2;
    wire c5386;
    assign in5386_1 = {c3800,c3793,s3785[3],s3836[0]};
    assign in5386_2 = {s3801[1],s3795[2],s3786[3],s3837[0]};
    CLA_4 KS_5386(s5386, c5386, in5386_1, in5386_2);
    wire[3:0] s5387, in5387_1, in5387_2;
    wire c5387;
    assign in5387_1 = {c3802,c3797,c3787,s3838[0]};
    assign in5387_2 = {s3803[1],s3799[2],s3791[3],s3839[0]};
    CLA_4 KS_5387(s5387, c5387, in5387_1, in5387_2);
    wire[0:0] s5388, in5388_1, in5388_2;
    wire c5388;
    assign in5388_1 = {c3804};
    assign in5388_2 = {s3805[1]};
    Half_Adder KS_5388(s5388, c5388, in5388_1, in5388_2);
    wire[1:0] s5389, in5389_1, in5389_2;
    wire c5389;
    assign in5389_1 = {c5354,c3801};
    assign in5389_2 = {c5355,s3803[2]};
    CLA_2 KS_5389(s5389, c5389, in5389_1, in5389_2);
    wire[0:0] s5390, in5390_1, in5390_2;
    wire c5390;
    assign in5390_1 = {c5356};
    assign in5390_2 = {c5357};
    Half_Adder KS_5390(s5390, c5390, in5390_1, in5390_2);
    wire[2:0] s5391, in5391_1, in5391_2;
    wire c5391;
    assign in5391_1 = {c5358,c3805,c3795};
    assign in5391_2 = {c5359,s5376[1],s3799[3]};
    CLA_3 KS_5391(s5391, c5391, in5391_1, in5391_2);
    wire[0:0] s5392, in5392_1, in5392_2;
    wire c5392;
    assign in5392_1 = {c5360};
    assign in5392_2 = {c5361};
    Half_Adder KS_5392(s5392, c5392, in5392_1, in5392_2);
    wire[1:0] s5393, in5393_1, in5393_2;
    wire c5393;
    assign in5393_1 = {c5362,s5377[1]};
    assign in5393_2 = {c5363,s5378[1]};
    CLA_2 KS_5393(s5393, c5393, in5393_1, in5393_2);
    wire[0:0] s5394, in5394_1, in5394_2;
    wire c5394;
    assign in5394_1 = {c5364};
    assign in5394_2 = {c5365};
    Half_Adder KS_5394(s5394, c5394, in5394_1, in5394_2);
    wire[3:0] s5395, in5395_1, in5395_2;
    wire c5395;
    assign in5395_1 = {c5373,s5379[1],c3803,s3840[0]};
    assign in5395_2 = {s5376[0],s5380[1],s5376[2],s3841[0]};
    CLA_4 KS_5395(s5395, c5395, in5395_1, in5395_2);
    wire[0:0] s5396, in5396_1, in5396_2;
    wire c5396;
    assign in5396_1 = {s5377[0]};
    assign in5396_2 = {s5378[0]};
    Half_Adder KS_5396(s5396, c5396, in5396_1, in5396_2);
    wire[1:0] s5397, in5397_1, in5397_2;
    wire c5397;
    assign in5397_1 = {s5380[0],s5381[1]};
    assign in5397_2 = {s5381[0],s5382[1]};
    CLA_2_c KS_5397(s5397, c5397, in5397_1, in5397_2, s5379[0]);
    wire[3:0] s5398, in5398_1, in5398_2;
    wire c5398;
    assign in5398_1 = {s3817[1],s3807[2],c1674,s3852[0]};
    assign in5398_2 = {s3818[1],s3808[2],s1675[1],s3853[0]};
    CLA_4 KS_5398(s5398, c5398, in5398_1, in5398_2);
    wire[3:0] s5399, in5399_1, in5399_2;
    wire c5399;
    assign in5399_1 = {s3819[1],s3809[2],c1676,s3854[0]};
    assign in5399_2 = {s3820[1],s3810[2],s1677[1],s3855[0]};
    CLA_4 KS_5399(s5399, c5399, in5399_1, in5399_2);
    wire[3:0] s5400, in5400_1, in5400_2;
    wire c5400;
    assign in5400_1 = {s3821[1],s3811[2],s3806[3],s3856[0]};
    assign in5400_2 = {s3822[1],s3812[2],s3807[3],s3857[0]};
    CLA_4 KS_5400(s5400, c5400, in5400_1, in5400_2);
    wire[3:0] s5401, in5401_1, in5401_2;
    wire c5401;
    assign in5401_1 = {s3823[1],s3813[2],s3808[3],s3858[0]};
    assign in5401_2 = {s3824[1],s3814[2],s3809[3],s3859[0]};
    CLA_4 KS_5401(s5401, c5401, in5401_1, in5401_2);
    wire[3:0] s5402, in5402_1, in5402_2;
    wire c5402;
    assign in5402_1 = {c3825,s3815[2],s3810[3],s3860[0]};
    assign in5402_2 = {s3826[1],s3816[2],s3811[3],s3861[0]};
    CLA_4 KS_5402(s5402, c5402, in5402_1, in5402_2);
    wire[3:0] s5403, in5403_1, in5403_2;
    wire c5403;
    assign in5403_1 = {c3827,s3817[2],s3812[3],s3862[0]};
    assign in5403_2 = {s3828[1],s3818[2],s3813[3],s3863[0]};
    CLA_4 KS_5403(s5403, c5403, in5403_1, in5403_2);
    wire[3:0] s5404, in5404_1, in5404_2;
    wire c5404;
    assign in5404_1 = {c3829,s3819[2],s3814[3],s3864[0]};
    assign in5404_2 = {s3830[1],s3820[2],s3815[3],s3865[0]};
    CLA_4 KS_5404(s5404, c5404, in5404_1, in5404_2);
    wire[3:0] s5405, in5405_1, in5405_2;
    wire c5405;
    assign in5405_1 = {c3831,s3821[2],s3816[3],s3866[0]};
    assign in5405_2 = {s3832[1],s3822[2],s3817[3],s3867[0]};
    CLA_4 KS_5405(s5405, c5405, in5405_1, in5405_2);
    wire[3:0] s5406, in5406_1, in5406_2;
    wire c5406;
    assign in5406_1 = {c3833,s3823[2],s3818[3],s3868[0]};
    assign in5406_2 = {s3834[1],s3824[2],s3819[3],s3869[0]};
    CLA_4 KS_5406(s5406, c5406, in5406_1, in5406_2);
    wire[3:0] s5407, in5407_1, in5407_2;
    wire c5407;
    assign in5407_1 = {c3835,c3826,s3820[3],s3870[0]};
    assign in5407_2 = {s3836[1],s3828[2],s3821[3],s3871[0]};
    CLA_4 KS_5407(s5407, c5407, in5407_1, in5407_2);
    wire[3:0] s5408, in5408_1, in5408_2;
    wire c5408;
    assign in5408_1 = {c3837,c3830,s3822[3],s3872[0]};
    assign in5408_2 = {s3838[1],s3832[2],s3823[3],s3873[0]};
    CLA_4 KS_5408(s5408, c5408, in5408_1, in5408_2);
    wire[3:0] s5409, in5409_1, in5409_2;
    wire c5409;
    assign in5409_1 = {c3839,c3834,c3824,s3874[0]};
    assign in5409_2 = {s3840[1],s3836[2],s3828[3],s3875[0]};
    CLA_4 KS_5409(s5409, c5409, in5409_1, in5409_2);
    wire[0:0] s5410, in5410_1, in5410_2;
    wire c5410;
    assign in5410_1 = {c3841};
    assign in5410_2 = {s3842[1]};
    Half_Adder KS_5410(s5410, c5410, in5410_1, in5410_2);
    wire[1:0] s5411, in5411_1, in5411_2;
    wire c5411;
    assign in5411_1 = {c5376,c3838};
    assign in5411_2 = {c5377,s3840[2]};
    CLA_2 KS_5411(s5411, c5411, in5411_1, in5411_2);
    wire[0:0] s5412, in5412_1, in5412_2;
    wire c5412;
    assign in5412_1 = {c5378};
    assign in5412_2 = {c5379};
    Half_Adder KS_5412(s5412, c5412, in5412_1, in5412_2);
    wire[2:0] s5413, in5413_1, in5413_2;
    wire c5413;
    assign in5413_1 = {c5380,c3842,c3832};
    assign in5413_2 = {c5381,s5398[1],s3836[3]};
    CLA_3 KS_5413(s5413, c5413, in5413_1, in5413_2);
    wire[0:0] s5414, in5414_1, in5414_2;
    wire c5414;
    assign in5414_1 = {c5382};
    assign in5414_2 = {c5383};
    Half_Adder KS_5414(s5414, c5414, in5414_1, in5414_2);
    wire[1:0] s5415, in5415_1, in5415_2;
    wire c5415;
    assign in5415_1 = {c5384,s5399[1]};
    assign in5415_2 = {c5385,s5400[1]};
    CLA_2 KS_5415(s5415, c5415, in5415_1, in5415_2);
    wire[0:0] s5416, in5416_1, in5416_2;
    wire c5416;
    assign in5416_1 = {c5386};
    assign in5416_2 = {c5387};
    Half_Adder KS_5416(s5416, c5416, in5416_1, in5416_2);
    wire[3:0] s5417, in5417_1, in5417_2;
    wire c5417;
    assign in5417_1 = {c5395,s5401[1],c3840,s3876[0]};
    assign in5417_2 = {s5398[0],s5402[1],s5398[2],s3877[0]};
    CLA_4 KS_5417(s5417, c5417, in5417_1, in5417_2);
    wire[0:0] s5418, in5418_1, in5418_2;
    wire c5418;
    assign in5418_1 = {s5399[0]};
    assign in5418_2 = {s5400[0]};
    Half_Adder KS_5418(s5418, c5418, in5418_1, in5418_2);
    wire[1:0] s5419, in5419_1, in5419_2;
    wire c5419;
    assign in5419_1 = {s5402[0],s5403[1]};
    assign in5419_2 = {s5403[0],s5404[1]};
    CLA_2_c KS_5419(s5419, c5419, in5419_1, in5419_2, s5401[0]);
    wire[3:0] s5420, in5420_1, in5420_2;
    wire c5420;
    assign in5420_1 = {s3852[1],s3844[2],c1726,s3888[0]};
    assign in5420_2 = {s3853[1],s3845[2],s1727[1],s3889[0]};
    CLA_4 KS_5420(s5420, c5420, in5420_1, in5420_2);
    wire[3:0] s5421, in5421_1, in5421_2;
    wire c5421;
    assign in5421_1 = {s3854[1],s3846[2],c1728,s3890[0]};
    assign in5421_2 = {s3855[1],s3847[2],s1729[1],s3891[0]};
    CLA_4 KS_5421(s5421, c5421, in5421_1, in5421_2);
    wire[3:0] s5422, in5422_1, in5422_2;
    wire c5422;
    assign in5422_1 = {s3856[1],s3848[2],s3843[3],s3892[0]};
    assign in5422_2 = {s3857[1],s3849[2],s3844[3],s3893[0]};
    CLA_4 KS_5422(s5422, c5422, in5422_1, in5422_2);
    wire[3:0] s5423, in5423_1, in5423_2;
    wire c5423;
    assign in5423_1 = {s3858[1],s3850[2],s3845[3],s3894[0]};
    assign in5423_2 = {s3859[1],s3851[2],s3846[3],s3895[0]};
    CLA_4 KS_5423(s5423, c5423, in5423_1, in5423_2);
    wire[3:0] s5424, in5424_1, in5424_2;
    wire c5424;
    assign in5424_1 = {s3860[1],s3852[2],s3847[3],s3896[0]};
    assign in5424_2 = {s3861[1],s3853[2],s3848[3],s3897[0]};
    CLA_4 KS_5424(s5424, c5424, in5424_1, in5424_2);
    wire[3:0] s5425, in5425_1, in5425_2;
    wire c5425;
    assign in5425_1 = {c3862,s3854[2],s3849[3],s3898[0]};
    assign in5425_2 = {s3863[1],s3855[2],s3850[3],s3899[0]};
    CLA_4 KS_5425(s5425, c5425, in5425_1, in5425_2);
    wire[3:0] s5426, in5426_1, in5426_2;
    wire c5426;
    assign in5426_1 = {c3864,s3856[2],s3851[3],s3900[0]};
    assign in5426_2 = {s3865[1],s3857[2],s3852[3],s3901[0]};
    CLA_4 KS_5426(s5426, c5426, in5426_1, in5426_2);
    wire[3:0] s5427, in5427_1, in5427_2;
    wire c5427;
    assign in5427_1 = {c3866,s3858[2],s3853[3],s3902[0]};
    assign in5427_2 = {s3867[1],s3859[2],s3854[3],s3903[0]};
    CLA_4 KS_5427(s5427, c5427, in5427_1, in5427_2);
    wire[3:0] s5428, in5428_1, in5428_2;
    wire c5428;
    assign in5428_1 = {c3868,s3860[2],s3855[3],s3904[0]};
    assign in5428_2 = {s3869[1],s3861[2],s3856[3],s3905[0]};
    CLA_4 KS_5428(s5428, c5428, in5428_1, in5428_2);
    wire[3:0] s5429, in5429_1, in5429_2;
    wire c5429;
    assign in5429_1 = {c3870,c3863,s3857[3],s3906[0]};
    assign in5429_2 = {s3871[1],s3865[2],s3858[3],s3907[0]};
    CLA_4 KS_5429(s5429, c5429, in5429_1, in5429_2);
    wire[3:0] s5430, in5430_1, in5430_2;
    wire c5430;
    assign in5430_1 = {c3872,c3867,s3859[3],s3908[0]};
    assign in5430_2 = {s3873[1],s3869[2],s3860[3],s3909[0]};
    CLA_4 KS_5430(s5430, c5430, in5430_1, in5430_2);
    wire[0:0] s5431, in5431_1, in5431_2;
    wire c5431;
    assign in5431_1 = {c3874};
    assign in5431_2 = {s3875[1]};
    Half_Adder KS_5431(s5431, c5431, in5431_1, in5431_2);
    wire[3:0] s5432, in5432_1, in5432_2;
    wire c5432;
    assign in5432_1 = {c3876,c3871,c3861,s3910[0]};
    assign in5432_2 = {s3877[1],s3873[2],s3865[3],s3911[0]};
    CLA_4 KS_5432(s5432, c5432, in5432_1, in5432_2);
    wire[0:0] s5433, in5433_1, in5433_2;
    wire c5433;
    assign in5433_1 = {c3878};
    assign in5433_2 = {c5398};
    Half_Adder KS_5433(s5433, c5433, in5433_1, in5433_2);
    wire[1:0] s5434, in5434_1, in5434_2;
    wire c5434;
    assign in5434_1 = {c5399,c3875};
    assign in5434_2 = {c5400,s3877[2]};
    CLA_2 KS_5434(s5434, c5434, in5434_1, in5434_2);
    wire[0:0] s5435, in5435_1, in5435_2;
    wire c5435;
    assign in5435_1 = {c5401};
    assign in5435_2 = {c5402};
    Half_Adder KS_5435(s5435, c5435, in5435_1, in5435_2);
    wire[2:0] s5436, in5436_1, in5436_2;
    wire c5436;
    assign in5436_1 = {c5403,s5420[1],c3869};
    assign in5436_2 = {c5404,s5421[1],s3873[3]};
    CLA_3 KS_5436(s5436, c5436, in5436_1, in5436_2);
    wire[0:0] s5437, in5437_1, in5437_2;
    wire c5437;
    assign in5437_1 = {c5405};
    assign in5437_2 = {c5406};
    Half_Adder KS_5437(s5437, c5437, in5437_1, in5437_2);
    wire[1:0] s5438, in5438_1, in5438_2;
    wire c5438;
    assign in5438_1 = {c5407,s5422[1]};
    assign in5438_2 = {c5408,s5423[1]};
    CLA_2 KS_5438(s5438, c5438, in5438_1, in5438_2);
    wire[0:0] s5439, in5439_1, in5439_2;
    wire c5439;
    assign in5439_1 = {c5409};
    assign in5439_2 = {c5417};
    Half_Adder KS_5439(s5439, c5439, in5439_1, in5439_2);
    wire[3:0] s5440, in5440_1, in5440_2;
    wire c5440;
    assign in5440_1 = {s5420[0],s5424[1],c3877,s3912[0]};
    assign in5440_2 = {s5421[0],s5425[1],s5420[2],s3913[0]};
    CLA_4 KS_5440(s5440, c5440, in5440_1, in5440_2);
    wire[0:0] s5441, in5441_1, in5441_2;
    wire c5441;
    assign in5441_1 = {s5422[0]};
    assign in5441_2 = {s5423[0]};
    Half_Adder KS_5441(s5441, c5441, in5441_1, in5441_2);
    wire[1:0] s5442, in5442_1, in5442_2;
    wire c5442;
    assign in5442_1 = {s5425[0],s5426[1]};
    assign in5442_2 = {s5426[0],s5427[1]};
    CLA_2_c KS_5442(s5442, c5442, in5442_1, in5442_2, s5424[0]);
    wire[3:0] s5443, in5443_1, in5443_2;
    wire c5443;
    assign in5443_1 = {s3888[1],s3880[2],c1770,s3926[0]};
    assign in5443_2 = {s3889[1],s3881[2],s1771[1],s3927[0]};
    CLA_4 KS_5443(s5443, c5443, in5443_1, in5443_2);
    wire[3:0] s5444, in5444_1, in5444_2;
    wire c5444;
    assign in5444_1 = {s3890[1],s3882[2],c1772,s3928[0]};
    assign in5444_2 = {s3891[1],s3883[2],s3879[3],s3929[0]};
    CLA_4 KS_5444(s5444, c5444, in5444_1, in5444_2);
    wire[3:0] s5445, in5445_1, in5445_2;
    wire c5445;
    assign in5445_1 = {s3892[1],s3884[2],s3880[3],s3930[0]};
    assign in5445_2 = {s3893[1],s3885[2],s3881[3],s3931[0]};
    CLA_4 KS_5445(s5445, c5445, in5445_1, in5445_2);
    wire[3:0] s5446, in5446_1, in5446_2;
    wire c5446;
    assign in5446_1 = {s3894[1],s3886[2],s3882[3],s3932[0]};
    assign in5446_2 = {s3895[1],s3887[2],s3883[3],s3933[0]};
    CLA_4 KS_5446(s5446, c5446, in5446_1, in5446_2);
    wire[3:0] s5447, in5447_1, in5447_2;
    wire c5447;
    assign in5447_1 = {s3896[1],s3888[2],s3884[3],s3934[0]};
    assign in5447_2 = {s3897[1],s3889[2],s3885[3],s3935[0]};
    CLA_4 KS_5447(s5447, c5447, in5447_1, in5447_2);
    wire[3:0] s5448, in5448_1, in5448_2;
    wire c5448;
    assign in5448_1 = {c3898,s3890[2],s3886[3],s3936[0]};
    assign in5448_2 = {s3899[1],s3891[2],s3887[3],s3937[0]};
    CLA_4 KS_5448(s5448, c5448, in5448_1, in5448_2);
    wire[3:0] s5449, in5449_1, in5449_2;
    wire c5449;
    assign in5449_1 = {c3900,s3892[2],s3888[3],s3938[0]};
    assign in5449_2 = {s3901[1],s3893[2],s3889[3],s3939[0]};
    CLA_4 KS_5449(s5449, c5449, in5449_1, in5449_2);
    wire[3:0] s5450, in5450_1, in5450_2;
    wire c5450;
    assign in5450_1 = {c3902,s3894[2],s3890[3],s3940[0]};
    assign in5450_2 = {s3903[1],s3895[2],s3891[3],s3941[0]};
    CLA_4 KS_5450(s5450, c5450, in5450_1, in5450_2);
    wire[3:0] s5451, in5451_1, in5451_2;
    wire c5451;
    assign in5451_1 = {c3904,s3896[2],s3892[3],s3942[0]};
    assign in5451_2 = {s3905[1],s3897[2],s3893[3],s3943[0]};
    CLA_4 KS_5451(s5451, c5451, in5451_1, in5451_2);
    wire[3:0] s5452, in5452_1, in5452_2;
    wire c5452;
    assign in5452_1 = {c3906,c3899,s3894[3],s3944[0]};
    assign in5452_2 = {s3907[1],s3901[2],s3895[3],s3945[0]};
    CLA_4 KS_5452(s5452, c5452, in5452_1, in5452_2);
    wire[3:0] s5453, in5453_1, in5453_2;
    wire c5453;
    assign in5453_1 = {c3908,c3903,s3896[3],s3946[0]};
    assign in5453_2 = {s3909[1],s3905[2],s3897[3],s3947[0]};
    CLA_4 KS_5453(s5453, c5453, in5453_1, in5453_2);
    wire[0:0] s5454, in5454_1, in5454_2;
    wire c5454;
    assign in5454_1 = {c3910};
    assign in5454_2 = {s3911[1]};
    Half_Adder KS_5454(s5454, c5454, in5454_1, in5454_2);
    wire[1:0] s5455, in5455_1, in5455_2;
    wire c5455;
    assign in5455_1 = {c3912,c3907};
    assign in5455_2 = {s3913[1],s3909[2]};
    CLA_2 KS_5455(s5455, c5455, in5455_1, in5455_2);
    wire[0:0] s5456, in5456_1, in5456_2;
    wire c5456;
    assign in5456_1 = {c3914};
    assign in5456_2 = {c5420};
    Half_Adder KS_5456(s5456, c5456, in5456_1, in5456_2);
    wire[3:0] s5457, in5457_1, in5457_2;
    wire c5457;
    assign in5457_1 = {c5421,c3911,c3901,s3948[0]};
    assign in5457_2 = {c5422,s3913[2],s3905[3],s3949[0]};
    CLA_4 KS_5457(s5457, c5457, in5457_1, in5457_2);
    wire[0:0] s5458, in5458_1, in5458_2;
    wire c5458;
    assign in5458_1 = {c5423};
    assign in5458_2 = {c5424};
    Half_Adder KS_5458(s5458, c5458, in5458_1, in5458_2);
    wire[1:0] s5459, in5459_1, in5459_2;
    wire c5459;
    assign in5459_1 = {c5425,s5443[1]};
    assign in5459_2 = {c5426,s5444[1]};
    CLA_2 KS_5459(s5459, c5459, in5459_1, in5459_2);
    wire[0:0] s5460, in5460_1, in5460_2;
    wire c5460;
    assign in5460_1 = {c5427};
    assign in5460_2 = {c5428};
    Half_Adder KS_5460(s5460, c5460, in5460_1, in5460_2);
    wire[2:0] s5461, in5461_1, in5461_2;
    wire c5461;
    assign in5461_1 = {c5429,s5445[1],c3909};
    assign in5461_2 = {c5430,s5446[1],s3913[3]};
    CLA_3 KS_5461(s5461, c5461, in5461_1, in5461_2);
    wire[0:0] s5462, in5462_1, in5462_2;
    wire c5462;
    assign in5462_1 = {c5432};
    assign in5462_2 = {c5440};
    Half_Adder KS_5462(s5462, c5462, in5462_1, in5462_2);
    wire[1:0] s5463, in5463_1, in5463_2;
    wire c5463;
    assign in5463_1 = {s5443[0],s5447[1]};
    assign in5463_2 = {s5444[0],s5448[1]};
    CLA_2 KS_5463(s5463, c5463, in5463_1, in5463_2);
    wire[0:0] s5464, in5464_1, in5464_2;
    wire c5464;
    assign in5464_1 = {s5445[0]};
    assign in5464_2 = {s5446[0]};
    Half_Adder KS_5464(s5464, c5464, in5464_1, in5464_2);
    wire[3:0] s5465, in5465_1, in5465_2;
    wire c5465;
    assign in5465_1 = {s5448[0],s5449[1],s5443[2],s3950[0]};
    assign in5465_2 = {s5449[0],s5450[1],s5444[2],s3951[0]};
    CLA_4_c KS_5465(s5465, c5465, in5465_1, in5465_2, s5447[0]);
    wire[3:0] s5466, in5466_1, in5466_2;
    wire c5466;
    assign in5466_1 = {s3926[1],s3917[2],c1830,s3962[0]};
    assign in5466_2 = {s3927[1],s3918[2],s1832[2],s3963[0]};
    CLA_4 KS_5466(s5466, c5466, in5466_1, in5466_2);
    wire[3:0] s5467, in5467_1, in5467_2;
    wire c5467;
    assign in5467_1 = {s3928[1],s3919[2],c1834,s3964[0]};
    assign in5467_2 = {s3929[1],s3920[2],s1836[2],s3965[0]};
    CLA_4 KS_5467(s5467, c5467, in5467_1, in5467_2);
    wire[3:0] s5468, in5468_1, in5468_2;
    wire c5468;
    assign in5468_1 = {s3930[1],s3921[2],s3915[3],s3966[0]};
    assign in5468_2 = {s3931[1],s3922[2],s3916[3],s3967[0]};
    CLA_4 KS_5468(s5468, c5468, in5468_1, in5468_2);
    wire[3:0] s5469, in5469_1, in5469_2;
    wire c5469;
    assign in5469_1 = {s3932[1],s3923[2],s3917[3],s3968[0]};
    assign in5469_2 = {s3933[1],s3924[2],s3918[3],s3969[0]};
    CLA_4 KS_5469(s5469, c5469, in5469_1, in5469_2);
    wire[3:0] s5470, in5470_1, in5470_2;
    wire c5470;
    assign in5470_1 = {c3934,s3925[2],s3919[3],s3970[0]};
    assign in5470_2 = {s3935[1],s3926[2],s3920[3],s3971[0]};
    CLA_4 KS_5470(s5470, c5470, in5470_1, in5470_2);
    wire[3:0] s5471, in5471_1, in5471_2;
    wire c5471;
    assign in5471_1 = {c3936,s3927[2],s3921[3],s3972[0]};
    assign in5471_2 = {s3937[1],s3928[2],s3922[3],s3973[0]};
    CLA_4 KS_5471(s5471, c5471, in5471_1, in5471_2);
    wire[3:0] s5472, in5472_1, in5472_2;
    wire c5472;
    assign in5472_1 = {c3938,s3929[2],s3923[3],s3974[0]};
    assign in5472_2 = {s3939[1],s3930[2],s3924[3],s3975[0]};
    CLA_4 KS_5472(s5472, c5472, in5472_1, in5472_2);
    wire[3:0] s5473, in5473_1, in5473_2;
    wire c5473;
    assign in5473_1 = {c3940,s3931[2],s3925[3],s3976[0]};
    assign in5473_2 = {s3941[1],s3932[2],s3926[3],s3977[0]};
    CLA_4 KS_5473(s5473, c5473, in5473_1, in5473_2);
    wire[3:0] s5474, in5474_1, in5474_2;
    wire c5474;
    assign in5474_1 = {c3942,c3933,s3927[3],s3978[0]};
    assign in5474_2 = {s3943[1],s3935[2],s3928[3],s3979[0]};
    CLA_4 KS_5474(s5474, c5474, in5474_1, in5474_2);
    wire[3:0] s5475, in5475_1, in5475_2;
    wire c5475;
    assign in5475_1 = {c3944,c3937,s3929[3],s3980[0]};
    assign in5475_2 = {s3945[1],s3939[2],s3930[3],s3981[0]};
    CLA_4 KS_5475(s5475, c5475, in5475_1, in5475_2);
    wire[3:0] s5476, in5476_1, in5476_2;
    wire c5476;
    assign in5476_1 = {c3946,c3941,s3931[3],s3982[0]};
    assign in5476_2 = {s3947[1],s3943[2],s3932[3],s3983[0]};
    CLA_4 KS_5476(s5476, c5476, in5476_1, in5476_2);
    wire[0:0] s5477, in5477_1, in5477_2;
    wire c5477;
    assign in5477_1 = {c3948};
    assign in5477_2 = {s3949[1]};
    Half_Adder KS_5477(s5477, c5477, in5477_1, in5477_2);
    wire[3:0] s5478, in5478_1, in5478_2;
    wire c5478;
    assign in5478_1 = {c3950,c3945,c3935,s3984[0]};
    assign in5478_2 = {s3951[1],s3947[2],s3939[3],s3985[0]};
    CLA_4 KS_5478(s5478, c5478, in5478_1, in5478_2);
    wire[0:0] s5479, in5479_1, in5479_2;
    wire c5479;
    assign in5479_1 = {c3952};
    assign in5479_2 = {c5443};
    Half_Adder KS_5479(s5479, c5479, in5479_1, in5479_2);
    wire[1:0] s5480, in5480_1, in5480_2;
    wire c5480;
    assign in5480_1 = {c5444,c3949};
    assign in5480_2 = {c5445,s3951[2]};
    CLA_2 KS_5480(s5480, c5480, in5480_1, in5480_2);
    wire[0:0] s5481, in5481_1, in5481_2;
    wire c5481;
    assign in5481_1 = {c5446};
    assign in5481_2 = {c5447};
    Half_Adder KS_5481(s5481, c5481, in5481_1, in5481_2);
    wire[2:0] s5482, in5482_1, in5482_2;
    wire c5482;
    assign in5482_1 = {c5448,s5466[1],c3943};
    assign in5482_2 = {c5449,s5467[1],s3947[3]};
    CLA_3 KS_5482(s5482, c5482, in5482_1, in5482_2);
    wire[0:0] s5483, in5483_1, in5483_2;
    wire c5483;
    assign in5483_1 = {c5450};
    assign in5483_2 = {c5451};
    Half_Adder KS_5483(s5483, c5483, in5483_1, in5483_2);
    wire[1:0] s5484, in5484_1, in5484_2;
    wire c5484;
    assign in5484_1 = {c5452,s5468[1]};
    assign in5484_2 = {c5453,s5469[1]};
    CLA_2 KS_5484(s5484, c5484, in5484_1, in5484_2);
    wire[0:0] s5485, in5485_1, in5485_2;
    wire c5485;
    assign in5485_1 = {c5457};
    assign in5485_2 = {c5465};
    Half_Adder KS_5485(s5485, c5485, in5485_1, in5485_2);
    wire[3:0] s5486, in5486_1, in5486_2;
    wire c5486;
    assign in5486_1 = {s5466[0],s5470[1],c3951,s3986[0]};
    assign in5486_2 = {s5467[0],s5471[1],s5466[2],s3987[0]};
    CLA_4 KS_5486(s5486, c5486, in5486_1, in5486_2);
    wire[0:0] s5487, in5487_1, in5487_2;
    wire c5487;
    assign in5487_1 = {s5468[0]};
    assign in5487_2 = {s5469[0]};
    Half_Adder KS_5487(s5487, c5487, in5487_1, in5487_2);
    wire[1:0] s5488, in5488_1, in5488_2;
    wire c5488;
    assign in5488_1 = {s5471[0],s5472[1]};
    assign in5488_2 = {s5472[0],s5473[1]};
    CLA_2_c KS_5488(s5488, c5488, in5488_1, in5488_2, s5470[0]);
    wire[3:0] s5489, in5489_1, in5489_2;
    wire c5489;
    assign in5489_1 = {s3962[1],s3954[2],c1895,s3998[0]};
    assign in5489_2 = {s3963[1],s3955[2],s1897[2],s3999[0]};
    CLA_4 KS_5489(s5489, c5489, in5489_1, in5489_2);
    wire[3:0] s5490, in5490_1, in5490_2;
    wire c5490;
    assign in5490_1 = {s3964[1],s3956[2],c1899,s4000[0]};
    assign in5490_2 = {s3965[1],s3957[2],s1901[2],s4001[0]};
    CLA_4 KS_5490(s5490, c5490, in5490_1, in5490_2);
    wire[3:0] s5491, in5491_1, in5491_2;
    wire c5491;
    assign in5491_1 = {s3966[1],s3958[2],s3953[3],s4002[0]};
    assign in5491_2 = {s3967[1],s3959[2],s3954[3],s4003[0]};
    CLA_4 KS_5491(s5491, c5491, in5491_1, in5491_2);
    wire[3:0] s5492, in5492_1, in5492_2;
    wire c5492;
    assign in5492_1 = {s3968[1],s3960[2],s3955[3],s4004[0]};
    assign in5492_2 = {s3969[1],s3961[2],s3956[3],s4005[0]};
    CLA_4 KS_5492(s5492, c5492, in5492_1, in5492_2);
    wire[3:0] s5493, in5493_1, in5493_2;
    wire c5493;
    assign in5493_1 = {s3970[1],s3962[2],s3957[3],s4006[0]};
    assign in5493_2 = {s3971[1],s3963[2],s3958[3],s4007[0]};
    CLA_4 KS_5493(s5493, c5493, in5493_1, in5493_2);
    wire[3:0] s5494, in5494_1, in5494_2;
    wire c5494;
    assign in5494_1 = {c3972,s3964[2],s3959[3],s4008[0]};
    assign in5494_2 = {s3973[1],s3965[2],s3960[3],s4009[0]};
    CLA_4 KS_5494(s5494, c5494, in5494_1, in5494_2);
    wire[3:0] s5495, in5495_1, in5495_2;
    wire c5495;
    assign in5495_1 = {c3974,s3966[2],s3961[3],s4010[0]};
    assign in5495_2 = {s3975[1],s3967[2],s3962[3],s4011[0]};
    CLA_4 KS_5495(s5495, c5495, in5495_1, in5495_2);
    wire[3:0] s5496, in5496_1, in5496_2;
    wire c5496;
    assign in5496_1 = {c3976,s3968[2],s3963[3],s4012[0]};
    assign in5496_2 = {s3977[1],s3969[2],s3964[3],s4013[0]};
    CLA_4 KS_5496(s5496, c5496, in5496_1, in5496_2);
    wire[3:0] s5497, in5497_1, in5497_2;
    wire c5497;
    assign in5497_1 = {c3978,s3970[2],s3965[3],s4014[0]};
    assign in5497_2 = {s3979[1],s3971[2],s3966[3],s4015[0]};
    CLA_4 KS_5497(s5497, c5497, in5497_1, in5497_2);
    wire[3:0] s5498, in5498_1, in5498_2;
    wire c5498;
    assign in5498_1 = {c3980,c3973,s3967[3],s4016[0]};
    assign in5498_2 = {s3981[1],s3975[2],s3968[3],s4017[0]};
    CLA_4 KS_5498(s5498, c5498, in5498_1, in5498_2);
    wire[3:0] s5499, in5499_1, in5499_2;
    wire c5499;
    assign in5499_1 = {c3982,c3977,s3969[3],s4018[0]};
    assign in5499_2 = {s3983[1],s3979[2],s3970[3],s4019[0]};
    CLA_4 KS_5499(s5499, c5499, in5499_1, in5499_2);
    wire[0:0] s5500, in5500_1, in5500_2;
    wire c5500;
    assign in5500_1 = {c3984};
    assign in5500_2 = {s3985[1]};
    Half_Adder KS_5500(s5500, c5500, in5500_1, in5500_2);
    wire[3:0] s5501, in5501_1, in5501_2;
    wire c5501;
    assign in5501_1 = {c3986,c3981,c3971,s4020[0]};
    assign in5501_2 = {s3987[1],s3983[2],s3975[3],s4021[0]};
    CLA_4 KS_5501(s5501, c5501, in5501_1, in5501_2);
    wire[0:0] s5502, in5502_1, in5502_2;
    wire c5502;
    assign in5502_1 = {c3988};
    assign in5502_2 = {c5466};
    Half_Adder KS_5502(s5502, c5502, in5502_1, in5502_2);
    wire[1:0] s5503, in5503_1, in5503_2;
    wire c5503;
    assign in5503_1 = {c5467,c3985};
    assign in5503_2 = {c5468,s3987[2]};
    CLA_2 KS_5503(s5503, c5503, in5503_1, in5503_2);
    wire[0:0] s5504, in5504_1, in5504_2;
    wire c5504;
    assign in5504_1 = {c5469};
    assign in5504_2 = {c5470};
    Half_Adder KS_5504(s5504, c5504, in5504_1, in5504_2);
    wire[2:0] s5505, in5505_1, in5505_2;
    wire c5505;
    assign in5505_1 = {c5471,s5489[1],c3979};
    assign in5505_2 = {c5472,s5490[1],s3983[3]};
    CLA_3 KS_5505(s5505, c5505, in5505_1, in5505_2);
    wire[0:0] s5506, in5506_1, in5506_2;
    wire c5506;
    assign in5506_1 = {c5473};
    assign in5506_2 = {c5474};
    Half_Adder KS_5506(s5506, c5506, in5506_1, in5506_2);
    wire[1:0] s5507, in5507_1, in5507_2;
    wire c5507;
    assign in5507_1 = {c5475,s5491[1]};
    assign in5507_2 = {c5476,s5492[1]};
    CLA_2 KS_5507(s5507, c5507, in5507_1, in5507_2);
    wire[0:0] s5508, in5508_1, in5508_2;
    wire c5508;
    assign in5508_1 = {c5478};
    assign in5508_2 = {c5486};
    Half_Adder KS_5508(s5508, c5508, in5508_1, in5508_2);
    wire[3:0] s5509, in5509_1, in5509_2;
    wire c5509;
    assign in5509_1 = {s5489[0],s5493[1],c3987,s4022[0]};
    assign in5509_2 = {s5490[0],s5494[1],s5489[2],s4023[0]};
    CLA_4 KS_5509(s5509, c5509, in5509_1, in5509_2);
    wire[0:0] s5510, in5510_1, in5510_2;
    wire c5510;
    assign in5510_1 = {s5491[0]};
    assign in5510_2 = {s5492[0]};
    Half_Adder KS_5510(s5510, c5510, in5510_1, in5510_2);
    wire[1:0] s5511, in5511_1, in5511_2;
    wire c5511;
    assign in5511_1 = {s5494[0],s5495[1]};
    assign in5511_2 = {s5495[0],s5496[1]};
    CLA_2_c KS_5511(s5511, c5511, in5511_1, in5511_2, s5493[0]);
    wire[3:0] s5512, in5512_1, in5512_2;
    wire c5512;
    assign in5512_1 = {s3998[1],s3990[2],c1961,s4034[0]};
    assign in5512_2 = {s3999[1],s3991[2],s1963[2],s4035[0]};
    CLA_4 KS_5512(s5512, c5512, in5512_1, in5512_2);
    wire[3:0] s5513, in5513_1, in5513_2;
    wire c5513;
    assign in5513_1 = {s4000[1],s3992[2],c1965,s4036[0]};
    assign in5513_2 = {s4001[1],s3993[2],s1967[2],s4037[0]};
    CLA_4 KS_5513(s5513, c5513, in5513_1, in5513_2);
    wire[3:0] s5514, in5514_1, in5514_2;
    wire c5514;
    assign in5514_1 = {s4002[1],s3994[2],s3989[3],s4038[0]};
    assign in5514_2 = {s4003[1],s3995[2],s3990[3],s4039[0]};
    CLA_4 KS_5514(s5514, c5514, in5514_1, in5514_2);
    wire[3:0] s5515, in5515_1, in5515_2;
    wire c5515;
    assign in5515_1 = {s4004[1],s3996[2],s3991[3],s4040[0]};
    assign in5515_2 = {s4005[1],s3997[2],s3992[3],s4041[0]};
    CLA_4 KS_5515(s5515, c5515, in5515_1, in5515_2);
    wire[3:0] s5516, in5516_1, in5516_2;
    wire c5516;
    assign in5516_1 = {s4006[1],s3998[2],s3993[3],s4042[0]};
    assign in5516_2 = {s4007[1],s3999[2],s3994[3],s4043[0]};
    CLA_4 KS_5516(s5516, c5516, in5516_1, in5516_2);
    wire[3:0] s5517, in5517_1, in5517_2;
    wire c5517;
    assign in5517_1 = {c4008,s4000[2],s3995[3],s4044[0]};
    assign in5517_2 = {s4009[1],s4001[2],s3996[3],s4045[0]};
    CLA_4 KS_5517(s5517, c5517, in5517_1, in5517_2);
    wire[3:0] s5518, in5518_1, in5518_2;
    wire c5518;
    assign in5518_1 = {c4010,s4002[2],s3997[3],s4046[0]};
    assign in5518_2 = {s4011[1],s4003[2],s3998[3],s4047[0]};
    CLA_4 KS_5518(s5518, c5518, in5518_1, in5518_2);
    wire[3:0] s5519, in5519_1, in5519_2;
    wire c5519;
    assign in5519_1 = {c4012,s4004[2],s3999[3],s4048[0]};
    assign in5519_2 = {s4013[1],s4005[2],s4000[3],s4049[0]};
    CLA_4 KS_5519(s5519, c5519, in5519_1, in5519_2);
    wire[3:0] s5520, in5520_1, in5520_2;
    wire c5520;
    assign in5520_1 = {c4014,s4006[2],s4001[3],s4050[0]};
    assign in5520_2 = {s4015[1],s4007[2],s4002[3],s4051[0]};
    CLA_4 KS_5520(s5520, c5520, in5520_1, in5520_2);
    wire[3:0] s5521, in5521_1, in5521_2;
    wire c5521;
    assign in5521_1 = {c4016,c4009,s4003[3],s4052[0]};
    assign in5521_2 = {s4017[1],s4011[2],s4004[3],s4053[0]};
    CLA_4 KS_5521(s5521, c5521, in5521_1, in5521_2);
    wire[3:0] s5522, in5522_1, in5522_2;
    wire c5522;
    assign in5522_1 = {c4018,c4013,s4005[3],s4054[0]};
    assign in5522_2 = {s4019[1],s4015[2],s4006[3],s4055[0]};
    CLA_4 KS_5522(s5522, c5522, in5522_1, in5522_2);
    wire[0:0] s5523, in5523_1, in5523_2;
    wire c5523;
    assign in5523_1 = {c4020};
    assign in5523_2 = {s4021[1]};
    Half_Adder KS_5523(s5523, c5523, in5523_1, in5523_2);
    wire[3:0] s5524, in5524_1, in5524_2;
    wire c5524;
    assign in5524_1 = {c4022,c4017,c4007,s4056[0]};
    assign in5524_2 = {s4023[1],s4019[2],s4011[3],s4057[0]};
    CLA_4 KS_5524(s5524, c5524, in5524_1, in5524_2);
    wire[0:0] s5525, in5525_1, in5525_2;
    wire c5525;
    assign in5525_1 = {c4024};
    assign in5525_2 = {c5489};
    Half_Adder KS_5525(s5525, c5525, in5525_1, in5525_2);
    wire[1:0] s5526, in5526_1, in5526_2;
    wire c5526;
    assign in5526_1 = {c5490,c4021};
    assign in5526_2 = {c5491,s4023[2]};
    CLA_2 KS_5526(s5526, c5526, in5526_1, in5526_2);
    wire[0:0] s5527, in5527_1, in5527_2;
    wire c5527;
    assign in5527_1 = {c5492};
    assign in5527_2 = {c5493};
    Half_Adder KS_5527(s5527, c5527, in5527_1, in5527_2);
    wire[2:0] s5528, in5528_1, in5528_2;
    wire c5528;
    assign in5528_1 = {c5494,s5512[1],c4015};
    assign in5528_2 = {c5495,s5513[1],s4019[3]};
    CLA_3 KS_5528(s5528, c5528, in5528_1, in5528_2);
    wire[0:0] s5529, in5529_1, in5529_2;
    wire c5529;
    assign in5529_1 = {c5496};
    assign in5529_2 = {c5497};
    Half_Adder KS_5529(s5529, c5529, in5529_1, in5529_2);
    wire[1:0] s5530, in5530_1, in5530_2;
    wire c5530;
    assign in5530_1 = {c5498,s5514[1]};
    assign in5530_2 = {c5499,s5515[1]};
    CLA_2 KS_5530(s5530, c5530, in5530_1, in5530_2);
    wire[0:0] s5531, in5531_1, in5531_2;
    wire c5531;
    assign in5531_1 = {c5501};
    assign in5531_2 = {c5509};
    Half_Adder KS_5531(s5531, c5531, in5531_1, in5531_2);
    wire[3:0] s5532, in5532_1, in5532_2;
    wire c5532;
    assign in5532_1 = {s5512[0],s5516[1],c4023,s4058[0]};
    assign in5532_2 = {s5513[0],s5517[1],s5512[2],s4059[0]};
    CLA_4 KS_5532(s5532, c5532, in5532_1, in5532_2);
    wire[0:0] s5533, in5533_1, in5533_2;
    wire c5533;
    assign in5533_1 = {s5514[0]};
    assign in5533_2 = {s5515[0]};
    Half_Adder KS_5533(s5533, c5533, in5533_1, in5533_2);
    wire[1:0] s5534, in5534_1, in5534_2;
    wire c5534;
    assign in5534_1 = {s5517[0],s5518[1]};
    assign in5534_2 = {s5518[0],s5519[1]};
    CLA_2_c KS_5534(s5534, c5534, in5534_1, in5534_2, s5516[0]);
    wire[3:0] s5535, in5535_1, in5535_2;
    wire c5535;
    assign in5535_1 = {s4034[1],s4025[2],c2026,s4070[0]};
    assign in5535_2 = {s4035[1],s4026[2],s2028[2],s4071[0]};
    CLA_4 KS_5535(s5535, c5535, in5535_1, in5535_2);
    wire[3:0] s5536, in5536_1, in5536_2;
    wire c5536;
    assign in5536_1 = {s4036[1],s4027[2],c2030,s4072[0]};
    assign in5536_2 = {s4037[1],s4028[2],s2032[2],s4073[0]};
    CLA_4 KS_5536(s5536, c5536, in5536_1, in5536_2);
    wire[3:0] s5537, in5537_1, in5537_2;
    wire c5537;
    assign in5537_1 = {s4038[1],s4029[2],c2034,s4074[0]};
    assign in5537_2 = {s4039[1],s4030[2],s4025[3],s4075[0]};
    CLA_4 KS_5537(s5537, c5537, in5537_1, in5537_2);
    wire[3:0] s5538, in5538_1, in5538_2;
    wire c5538;
    assign in5538_1 = {s4040[1],s4031[2],s4026[3],s4076[0]};
    assign in5538_2 = {s4041[1],s4032[2],s4027[3],s4077[0]};
    CLA_4 KS_5538(s5538, c5538, in5538_1, in5538_2);
    wire[3:0] s5539, in5539_1, in5539_2;
    wire c5539;
    assign in5539_1 = {s4042[1],s4033[2],s4028[3],s4078[0]};
    assign in5539_2 = {s4043[1],s4034[2],s4029[3],s4079[0]};
    CLA_4 KS_5539(s5539, c5539, in5539_1, in5539_2);
    wire[3:0] s5540, in5540_1, in5540_2;
    wire c5540;
    assign in5540_1 = {c4044,s4035[2],s4030[3],s4080[0]};
    assign in5540_2 = {s4045[1],s4036[2],s4031[3],s4081[0]};
    CLA_4 KS_5540(s5540, c5540, in5540_1, in5540_2);
    wire[3:0] s5541, in5541_1, in5541_2;
    wire c5541;
    assign in5541_1 = {c4046,s4037[2],s4032[3],s4082[0]};
    assign in5541_2 = {s4047[1],s4038[2],s4033[3],s4083[0]};
    CLA_4 KS_5541(s5541, c5541, in5541_1, in5541_2);
    wire[3:0] s5542, in5542_1, in5542_2;
    wire c5542;
    assign in5542_1 = {c4048,s4039[2],s4034[3],s4084[0]};
    assign in5542_2 = {s4049[1],s4040[2],s4035[3],s4085[0]};
    CLA_4 KS_5542(s5542, c5542, in5542_1, in5542_2);
    wire[3:0] s5543, in5543_1, in5543_2;
    wire c5543;
    assign in5543_1 = {c4050,s4041[2],s4036[3],s4086[0]};
    assign in5543_2 = {s4051[1],s4042[2],s4037[3],s4087[0]};
    CLA_4 KS_5543(s5543, c5543, in5543_1, in5543_2);
    wire[3:0] s5544, in5544_1, in5544_2;
    wire c5544;
    assign in5544_1 = {c4052,c4043,s4038[3],s4088[0]};
    assign in5544_2 = {s4053[1],s4045[2],s4039[3],s4089[0]};
    CLA_4 KS_5544(s5544, c5544, in5544_1, in5544_2);
    wire[3:0] s5545, in5545_1, in5545_2;
    wire c5545;
    assign in5545_1 = {c4054,c4047,s4040[3],s4090[0]};
    assign in5545_2 = {s4055[1],s4049[2],s4041[3],s4091[0]};
    CLA_4 KS_5545(s5545, c5545, in5545_1, in5545_2);
    wire[3:0] s5546, in5546_1, in5546_2;
    wire c5546;
    assign in5546_1 = {c4056,c4051,s4042[3],s4092[0]};
    assign in5546_2 = {s4057[1],s4053[2],s4045[3],s4093[0]};
    CLA_4 KS_5546(s5546, c5546, in5546_1, in5546_2);
    wire[0:0] s5547, in5547_1, in5547_2;
    wire c5547;
    assign in5547_1 = {c4058};
    assign in5547_2 = {s4059[1]};
    Half_Adder KS_5547(s5547, c5547, in5547_1, in5547_2);
    wire[1:0] s5548, in5548_1, in5548_2;
    wire c5548;
    assign in5548_1 = {c4060,c4055};
    assign in5548_2 = {c5512,s4057[2]};
    CLA_2 KS_5548(s5548, c5548, in5548_1, in5548_2);
    wire[0:0] s5549, in5549_1, in5549_2;
    wire c5549;
    assign in5549_1 = {c5513};
    assign in5549_2 = {c5514};
    Half_Adder KS_5549(s5549, c5549, in5549_1, in5549_2);
    wire[2:0] s5550, in5550_1, in5550_2;
    wire c5550;
    assign in5550_1 = {c5515,c4059,c4049};
    assign in5550_2 = {c5516,s5535[1],s4053[3]};
    CLA_3 KS_5550(s5550, c5550, in5550_1, in5550_2);
    wire[0:0] s5551, in5551_1, in5551_2;
    wire c5551;
    assign in5551_1 = {c5517};
    assign in5551_2 = {c5518};
    Half_Adder KS_5551(s5551, c5551, in5551_1, in5551_2);
    wire[1:0] s5552, in5552_1, in5552_2;
    wire c5552;
    assign in5552_1 = {c5519,s5536[1]};
    assign in5552_2 = {c5520,s5537[1]};
    CLA_2 KS_5552(s5552, c5552, in5552_1, in5552_2);
    wire[0:0] s5553, in5553_1, in5553_2;
    wire c5553;
    assign in5553_1 = {c5521};
    assign in5553_2 = {c5522};
    Half_Adder KS_5553(s5553, c5553, in5553_1, in5553_2);
    wire[3:0] s5554, in5554_1, in5554_2;
    wire c5554;
    assign in5554_1 = {c5524,s5538[1],c4057,s4094[0]};
    assign in5554_2 = {c5532,s5539[1],s5535[2],s4095[0]};
    CLA_4 KS_5554(s5554, c5554, in5554_1, in5554_2);
    wire[0:0] s5555, in5555_1, in5555_2;
    wire c5555;
    assign in5555_1 = {s5535[0]};
    assign in5555_2 = {s5536[0]};
    Half_Adder KS_5555(s5555, c5555, in5555_1, in5555_2);
    wire[1:0] s5556, in5556_1, in5556_2;
    wire c5556;
    assign in5556_1 = {s5537[0],s5540[1]};
    assign in5556_2 = {s5538[0],s5541[1]};
    CLA_2 KS_5556(s5556, c5556, in5556_1, in5556_2);
    wire[0:0] s5557, in5557_1, in5557_2;
    wire c5557;
    assign in5557_1 = {s5540[0]};
    assign in5557_2 = {s5541[0]};
    Full_Adder KS_5557(s5557, c5557, in5557_1, in5557_2, s5539[0]);
    wire[3:0] s5558, in5558_1, in5558_2;
    wire c5558;
    assign in5558_1 = {s4070[1],s4061[2],c2094,s4106[0]};
    assign in5558_2 = {s4071[1],s4062[2],s2096[2],s4107[0]};
    CLA_4 KS_5558(s5558, c5558, in5558_1, in5558_2);
    wire[3:0] s5559, in5559_1, in5559_2;
    wire c5559;
    assign in5559_1 = {s4072[1],s4063[2],c2098,s4108[0]};
    assign in5559_2 = {s4073[1],s4064[2],s2100[2],s4109[0]};
    CLA_4 KS_5559(s5559, c5559, in5559_1, in5559_2);
    wire[3:0] s5560, in5560_1, in5560_2;
    wire c5560;
    assign in5560_1 = {s4074[1],s4065[2],s4061[3],s4110[0]};
    assign in5560_2 = {s4075[1],s4066[2],s4062[3],s4111[0]};
    CLA_4 KS_5560(s5560, c5560, in5560_1, in5560_2);
    wire[3:0] s5561, in5561_1, in5561_2;
    wire c5561;
    assign in5561_1 = {s4076[1],s4067[2],s4063[3],s4112[0]};
    assign in5561_2 = {s4077[1],s4068[2],s4064[3],s4113[0]};
    CLA_4 KS_5561(s5561, c5561, in5561_1, in5561_2);
    wire[3:0] s5562, in5562_1, in5562_2;
    wire c5562;
    assign in5562_1 = {s4078[1],s4069[2],s4065[3],s4114[0]};
    assign in5562_2 = {s4079[1],s4070[2],s4066[3],s4115[0]};
    CLA_4 KS_5562(s5562, c5562, in5562_1, in5562_2);
    wire[3:0] s5563, in5563_1, in5563_2;
    wire c5563;
    assign in5563_1 = {c4080,s4071[2],s4067[3],s4116[0]};
    assign in5563_2 = {s4081[1],s4072[2],s4068[3],s4117[0]};
    CLA_4 KS_5563(s5563, c5563, in5563_1, in5563_2);
    wire[3:0] s5564, in5564_1, in5564_2;
    wire c5564;
    assign in5564_1 = {c4082,s4073[2],s4069[3],s4118[0]};
    assign in5564_2 = {s4083[1],s4074[2],s4070[3],s4119[0]};
    CLA_4 KS_5564(s5564, c5564, in5564_1, in5564_2);
    wire[3:0] s5565, in5565_1, in5565_2;
    wire c5565;
    assign in5565_1 = {c4084,s4075[2],s4071[3],s4120[0]};
    assign in5565_2 = {s4085[1],s4076[2],s4072[3],s4121[0]};
    CLA_4 KS_5565(s5565, c5565, in5565_1, in5565_2);
    wire[3:0] s5566, in5566_1, in5566_2;
    wire c5566;
    assign in5566_1 = {c4086,s4077[2],s4073[3],s4122[0]};
    assign in5566_2 = {s4087[1],s4078[2],s4074[3],s4123[0]};
    CLA_4 KS_5566(s5566, c5566, in5566_1, in5566_2);
    wire[3:0] s5567, in5567_1, in5567_2;
    wire c5567;
    assign in5567_1 = {c4088,c4079,s4075[3],s4124[0]};
    assign in5567_2 = {s4089[1],s4081[2],s4076[3],s4125[0]};
    CLA_4 KS_5567(s5567, c5567, in5567_1, in5567_2);
    wire[3:0] s5568, in5568_1, in5568_2;
    wire c5568;
    assign in5568_1 = {c4090,c4083,s4077[3],s4126[0]};
    assign in5568_2 = {s4091[1],s4085[2],s4078[3],s4127[0]};
    CLA_4 KS_5568(s5568, c5568, in5568_1, in5568_2);
    wire[1:0] s5569, in5569_1, in5569_2;
    wire c5569;
    assign in5569_1 = {c4092,c4087};
    assign in5569_2 = {s4093[1],s4089[2]};
    CLA_2 KS_5569(s5569, c5569, in5569_1, in5569_2);
    wire[0:0] s5570, in5570_1, in5570_2;
    wire c5570;
    assign in5570_1 = {c4094};
    assign in5570_2 = {s4095[1]};
    Half_Adder KS_5570(s5570, c5570, in5570_1, in5570_2);
    wire[3:0] s5571, in5571_1, in5571_2;
    wire c5571;
    assign in5571_1 = {c4096,c4091,c4081,s4128[0]};
    assign in5571_2 = {c5535,s4093[2],s4085[3],s4129[0]};
    CLA_4 KS_5571(s5571, c5571, in5571_1, in5571_2);
    wire[0:0] s5572, in5572_1, in5572_2;
    wire c5572;
    assign in5572_1 = {c5536};
    assign in5572_2 = {c5537};
    Half_Adder KS_5572(s5572, c5572, in5572_1, in5572_2);
    wire[1:0] s5573, in5573_1, in5573_2;
    wire c5573;
    assign in5573_1 = {c5538,c4095};
    assign in5573_2 = {c5539,s5558[1]};
    CLA_2 KS_5573(s5573, c5573, in5573_1, in5573_2);
    wire[0:0] s5574, in5574_1, in5574_2;
    wire c5574;
    assign in5574_1 = {c5540};
    assign in5574_2 = {c5541};
    Half_Adder KS_5574(s5574, c5574, in5574_1, in5574_2);
    wire[2:0] s5575, in5575_1, in5575_2;
    wire c5575;
    assign in5575_1 = {c5542,s5559[1],c4089};
    assign in5575_2 = {c5543,s5560[1],s4093[3]};
    CLA_3 KS_5575(s5575, c5575, in5575_1, in5575_2);
    wire[0:0] s5576, in5576_1, in5576_2;
    wire c5576;
    assign in5576_1 = {c5544};
    assign in5576_2 = {c5545};
    Half_Adder KS_5576(s5576, c5576, in5576_1, in5576_2);
    wire[1:0] s5577, in5577_1, in5577_2;
    wire c5577;
    assign in5577_1 = {c5546,s5561[1]};
    assign in5577_2 = {c5554,s5562[1]};
    CLA_2 KS_5577(s5577, c5577, in5577_1, in5577_2);
    wire[0:0] s5578, in5578_1, in5578_2;
    wire c5578;
    assign in5578_1 = {s5558[0]};
    assign in5578_2 = {s5559[0]};
    Half_Adder KS_5578(s5578, c5578, in5578_1, in5578_2);
    wire[3:0] s5579, in5579_1, in5579_2;
    wire c5579;
    assign in5579_1 = {s5560[0],s5563[1],s5558[2],s4130[0]};
    assign in5579_2 = {s5561[0],s5564[1],s5559[2],s4131[0]};
    CLA_4 KS_5579(s5579, c5579, in5579_1, in5579_2);
    wire[0:0] s5580, in5580_1, in5580_2;
    wire c5580;
    assign in5580_1 = {s5563[0]};
    assign in5580_2 = {s5564[0]};
    Full_Adder KS_5580(s5580, c5580, in5580_1, in5580_2, s5562[0]);
    wire[3:0] s5581, in5581_1, in5581_2;
    wire c5581;
    assign in5581_1 = {s4106[1],s4097[2],c2160,s4142[0]};
    assign in5581_2 = {s4107[1],s4098[2],s2162[2],s4143[0]};
    CLA_4 KS_5581(s5581, c5581, in5581_1, in5581_2);
    wire[3:0] s5582, in5582_1, in5582_2;
    wire c5582;
    assign in5582_1 = {s4108[1],s4099[2],c2164,s4144[0]};
    assign in5582_2 = {s4109[1],s4100[2],s2166[2],s4145[0]};
    CLA_4 KS_5582(s5582, c5582, in5582_1, in5582_2);
    wire[3:0] s5583, in5583_1, in5583_2;
    wire c5583;
    assign in5583_1 = {s4110[1],s4101[2],s4097[3],s4146[0]};
    assign in5583_2 = {s4111[1],s4102[2],s4098[3],s4147[0]};
    CLA_4 KS_5583(s5583, c5583, in5583_1, in5583_2);
    wire[3:0] s5584, in5584_1, in5584_2;
    wire c5584;
    assign in5584_1 = {s4112[1],s4103[2],s4099[3],s4148[0]};
    assign in5584_2 = {s4113[1],s4104[2],s4100[3],s4149[0]};
    CLA_4 KS_5584(s5584, c5584, in5584_1, in5584_2);
    wire[3:0] s5585, in5585_1, in5585_2;
    wire c5585;
    assign in5585_1 = {s4114[1],s4105[2],s4101[3],s4150[0]};
    assign in5585_2 = {s4115[1],s4106[2],s4102[3],s4151[0]};
    CLA_4 KS_5585(s5585, c5585, in5585_1, in5585_2);
    wire[3:0] s5586, in5586_1, in5586_2;
    wire c5586;
    assign in5586_1 = {c4116,s4107[2],s4103[3],s4152[0]};
    assign in5586_2 = {s4117[1],s4108[2],s4104[3],s4153[0]};
    CLA_4 KS_5586(s5586, c5586, in5586_1, in5586_2);
    wire[3:0] s5587, in5587_1, in5587_2;
    wire c5587;
    assign in5587_1 = {c4118,s4109[2],s4105[3],s4154[0]};
    assign in5587_2 = {s4119[1],s4110[2],s4106[3],s4155[0]};
    CLA_4 KS_5587(s5587, c5587, in5587_1, in5587_2);
    wire[3:0] s5588, in5588_1, in5588_2;
    wire c5588;
    assign in5588_1 = {c4120,s4111[2],s4107[3],s4156[0]};
    assign in5588_2 = {s4121[1],s4112[2],s4108[3],s4157[0]};
    CLA_4 KS_5588(s5588, c5588, in5588_1, in5588_2);
    wire[3:0] s5589, in5589_1, in5589_2;
    wire c5589;
    assign in5589_1 = {c4122,s4113[2],s4109[3],s4158[0]};
    assign in5589_2 = {s4123[1],s4114[2],s4110[3],s4159[0]};
    CLA_4 KS_5589(s5589, c5589, in5589_1, in5589_2);
    wire[3:0] s5590, in5590_1, in5590_2;
    wire c5590;
    assign in5590_1 = {c4124,c4115,s4111[3],s4160[0]};
    assign in5590_2 = {s4125[1],s4117[2],s4112[3],s4161[0]};
    CLA_4 KS_5590(s5590, c5590, in5590_1, in5590_2);
    wire[3:0] s5591, in5591_1, in5591_2;
    wire c5591;
    assign in5591_1 = {c4126,c4119,s4113[3],s4162[0]};
    assign in5591_2 = {s4127[1],s4121[2],s4114[3],s4163[0]};
    CLA_4 KS_5591(s5591, c5591, in5591_1, in5591_2);
    wire[1:0] s5592, in5592_1, in5592_2;
    wire c5592;
    assign in5592_1 = {c4128,c4123};
    assign in5592_2 = {s4129[1],s4125[2]};
    CLA_2 KS_5592(s5592, c5592, in5592_1, in5592_2);
    wire[0:0] s5593, in5593_1, in5593_2;
    wire c5593;
    assign in5593_1 = {c4130};
    assign in5593_2 = {s4131[1]};
    Half_Adder KS_5593(s5593, c5593, in5593_1, in5593_2);
    wire[3:0] s5594, in5594_1, in5594_2;
    wire c5594;
    assign in5594_1 = {c4132,c4127,c4117,s4164[0]};
    assign in5594_2 = {c5558,s4129[2],s4121[3],s4165[0]};
    CLA_4 KS_5594(s5594, c5594, in5594_1, in5594_2);
    wire[0:0] s5595, in5595_1, in5595_2;
    wire c5595;
    assign in5595_1 = {c5559};
    assign in5595_2 = {c5560};
    Half_Adder KS_5595(s5595, c5595, in5595_1, in5595_2);
    wire[1:0] s5596, in5596_1, in5596_2;
    wire c5596;
    assign in5596_1 = {c5561,c4131};
    assign in5596_2 = {c5562,s5581[1]};
    CLA_2 KS_5596(s5596, c5596, in5596_1, in5596_2);
    wire[0:0] s5597, in5597_1, in5597_2;
    wire c5597;
    assign in5597_1 = {c5563};
    assign in5597_2 = {c5564};
    Half_Adder KS_5597(s5597, c5597, in5597_1, in5597_2);
    wire[2:0] s5598, in5598_1, in5598_2;
    wire c5598;
    assign in5598_1 = {c5565,s5582[1],c4125};
    assign in5598_2 = {c5566,s5583[1],s4129[3]};
    CLA_3 KS_5598(s5598, c5598, in5598_1, in5598_2);
    wire[0:0] s5599, in5599_1, in5599_2;
    wire c5599;
    assign in5599_1 = {c5567};
    assign in5599_2 = {c5568};
    Half_Adder KS_5599(s5599, c5599, in5599_1, in5599_2);
    wire[1:0] s5600, in5600_1, in5600_2;
    wire c5600;
    assign in5600_1 = {c5571,s5584[1]};
    assign in5600_2 = {c5579,s5585[1]};
    CLA_2 KS_5600(s5600, c5600, in5600_1, in5600_2);
    wire[0:0] s5601, in5601_1, in5601_2;
    wire c5601;
    assign in5601_1 = {s5581[0]};
    assign in5601_2 = {s5582[0]};
    Half_Adder KS_5601(s5601, c5601, in5601_1, in5601_2);
    wire[3:0] s5602, in5602_1, in5602_2;
    wire c5602;
    assign in5602_1 = {s5583[0],s5586[1],s5581[2],s4166[0]};
    assign in5602_2 = {s5584[0],s5587[1],s5582[2],s4167[0]};
    CLA_4 KS_5602(s5602, c5602, in5602_1, in5602_2);
    wire[0:0] s5603, in5603_1, in5603_2;
    wire c5603;
    assign in5603_1 = {s5586[0]};
    assign in5603_2 = {s5587[0]};
    Full_Adder KS_5603(s5603, c5603, in5603_1, in5603_2, s5585[0]);
    wire[3:0] s5604, in5604_1, in5604_2;
    wire c5604;
    assign in5604_1 = {s4142[1],s4134[2],c2227,s4180[0]};
    assign in5604_2 = {s4143[1],s4135[2],s2229[2],s4181[0]};
    CLA_4 KS_5604(s5604, c5604, in5604_1, in5604_2);
    wire[3:0] s5605, in5605_1, in5605_2;
    wire c5605;
    assign in5605_1 = {s4144[1],s4136[2],c2231,s4182[0]};
    assign in5605_2 = {s4145[1],s4137[2],s4133[3],s4183[0]};
    CLA_4 KS_5605(s5605, c5605, in5605_1, in5605_2);
    wire[3:0] s5606, in5606_1, in5606_2;
    wire c5606;
    assign in5606_1 = {s4146[1],s4138[2],s4134[3],s4184[0]};
    assign in5606_2 = {s4147[1],s4139[2],s4135[3],s4185[0]};
    CLA_4 KS_5606(s5606, c5606, in5606_1, in5606_2);
    wire[3:0] s5607, in5607_1, in5607_2;
    wire c5607;
    assign in5607_1 = {s4148[1],s4140[2],s4136[3],s4186[0]};
    assign in5607_2 = {s4149[1],s4141[2],s4137[3],s4187[0]};
    CLA_4 KS_5607(s5607, c5607, in5607_1, in5607_2);
    wire[3:0] s5608, in5608_1, in5608_2;
    wire c5608;
    assign in5608_1 = {s4150[1],s4142[2],s4138[3],s4188[0]};
    assign in5608_2 = {s4151[1],s4143[2],s4139[3],s4189[0]};
    CLA_4 KS_5608(s5608, c5608, in5608_1, in5608_2);
    wire[3:0] s5609, in5609_1, in5609_2;
    wire c5609;
    assign in5609_1 = {c4152,s4144[2],s4140[3],s4190[0]};
    assign in5609_2 = {s4153[1],s4145[2],s4141[3],s4191[0]};
    CLA_4 KS_5609(s5609, c5609, in5609_1, in5609_2);
    wire[3:0] s5610, in5610_1, in5610_2;
    wire c5610;
    assign in5610_1 = {c4154,s4146[2],s4142[3],s4192[0]};
    assign in5610_2 = {s4155[1],s4147[2],s4143[3],s4193[0]};
    CLA_4 KS_5610(s5610, c5610, in5610_1, in5610_2);
    wire[3:0] s5611, in5611_1, in5611_2;
    wire c5611;
    assign in5611_1 = {c4156,s4148[2],s4144[3],s4194[0]};
    assign in5611_2 = {s4157[1],s4149[2],s4145[3],s4195[0]};
    CLA_4 KS_5611(s5611, c5611, in5611_1, in5611_2);
    wire[3:0] s5612, in5612_1, in5612_2;
    wire c5612;
    assign in5612_1 = {c4158,s4150[2],s4146[3],s4196[0]};
    assign in5612_2 = {s4159[1],s4151[2],s4147[3],s4197[0]};
    CLA_4 KS_5612(s5612, c5612, in5612_1, in5612_2);
    wire[3:0] s5613, in5613_1, in5613_2;
    wire c5613;
    assign in5613_1 = {c4160,c4153,s4148[3],s4198[0]};
    assign in5613_2 = {s4161[1],s4155[2],s4149[3],s4199[0]};
    CLA_4 KS_5613(s5613, c5613, in5613_1, in5613_2);
    wire[3:0] s5614, in5614_1, in5614_2;
    wire c5614;
    assign in5614_1 = {c4162,c4157,s4150[3],s4200[0]};
    assign in5614_2 = {s4163[1],s4159[2],s4151[3],s4201[0]};
    CLA_4 KS_5614(s5614, c5614, in5614_1, in5614_2);
    wire[0:0] s5615, in5615_1, in5615_2;
    wire c5615;
    assign in5615_1 = {c4164};
    assign in5615_2 = {s4165[1]};
    Half_Adder KS_5615(s5615, c5615, in5615_1, in5615_2);
    wire[1:0] s5616, in5616_1, in5616_2;
    wire c5616;
    assign in5616_1 = {c4166,c4161};
    assign in5616_2 = {s4167[1],s4163[2]};
    CLA_2 KS_5616(s5616, c5616, in5616_1, in5616_2);
    wire[0:0] s5617, in5617_1, in5617_2;
    wire c5617;
    assign in5617_1 = {c4168};
    assign in5617_2 = {c5581};
    Half_Adder KS_5617(s5617, c5617, in5617_1, in5617_2);
    wire[3:0] s5618, in5618_1, in5618_2;
    wire c5618;
    assign in5618_1 = {c5582,c4165,c4155,s4202[0]};
    assign in5618_2 = {c5583,s4167[2],s4159[3],s4203[0]};
    CLA_4 KS_5618(s5618, c5618, in5618_1, in5618_2);
    wire[0:0] s5619, in5619_1, in5619_2;
    wire c5619;
    assign in5619_1 = {c5584};
    assign in5619_2 = {c5585};
    Half_Adder KS_5619(s5619, c5619, in5619_1, in5619_2);
    wire[1:0] s5620, in5620_1, in5620_2;
    wire c5620;
    assign in5620_1 = {c5586,s5604[1]};
    assign in5620_2 = {c5587,s5605[1]};
    CLA_2 KS_5620(s5620, c5620, in5620_1, in5620_2);
    wire[0:0] s5621, in5621_1, in5621_2;
    wire c5621;
    assign in5621_1 = {c5588};
    assign in5621_2 = {c5589};
    Half_Adder KS_5621(s5621, c5621, in5621_1, in5621_2);
    wire[2:0] s5622, in5622_1, in5622_2;
    wire c5622;
    assign in5622_1 = {c5590,s5606[1],c4163};
    assign in5622_2 = {c5591,s5607[1],s4167[3]};
    CLA_3 KS_5622(s5622, c5622, in5622_1, in5622_2);
    wire[0:0] s5623, in5623_1, in5623_2;
    wire c5623;
    assign in5623_1 = {c5594};
    assign in5623_2 = {c5602};
    Half_Adder KS_5623(s5623, c5623, in5623_1, in5623_2);
    wire[1:0] s5624, in5624_1, in5624_2;
    wire c5624;
    assign in5624_1 = {s5604[0],s5608[1]};
    assign in5624_2 = {s5605[0],s5609[1]};
    CLA_2 KS_5624(s5624, c5624, in5624_1, in5624_2);
    wire[0:0] s5625, in5625_1, in5625_2;
    wire c5625;
    assign in5625_1 = {s5606[0]};
    assign in5625_2 = {s5607[0]};
    Half_Adder KS_5625(s5625, c5625, in5625_1, in5625_2);
    wire[3:0] s5626, in5626_1, in5626_2;
    wire c5626;
    assign in5626_1 = {s5609[0],s5610[1],s5604[2],s4204[0]};
    assign in5626_2 = {s5610[0],s5611[1],s5605[2],s4205[0]};
    CLA_4_c KS_5626(s5626, c5626, in5626_1, in5626_2, s5608[0]);
    wire[3:0] s5627, in5627_1, in5627_2;
    wire c5627;
    assign in5627_1 = {s4180[1],s4171[2],c2292,s4218[0]};
    assign in5627_2 = {s4181[1],s4172[2],s2294[2],s4219[0]};
    CLA_4 KS_5627(s5627, c5627, in5627_1, in5627_2);
    wire[3:0] s5628, in5628_1, in5628_2;
    wire c5628;
    assign in5628_1 = {s4182[1],s4173[2],c2296,s4220[0]};
    assign in5628_2 = {s4183[1],s4174[2],s4169[3],s4221[0]};
    CLA_4 KS_5628(s5628, c5628, in5628_1, in5628_2);
    wire[3:0] s5629, in5629_1, in5629_2;
    wire c5629;
    assign in5629_1 = {s4184[1],s4175[2],s4170[3],s4222[0]};
    assign in5629_2 = {s4185[1],s4176[2],s4171[3],s4223[0]};
    CLA_4 KS_5629(s5629, c5629, in5629_1, in5629_2);
    wire[3:0] s5630, in5630_1, in5630_2;
    wire c5630;
    assign in5630_1 = {s4186[1],s4177[2],s4172[3],s4224[0]};
    assign in5630_2 = {s4187[1],s4178[2],s4173[3],s4225[0]};
    CLA_4 KS_5630(s5630, c5630, in5630_1, in5630_2);
    wire[3:0] s5631, in5631_1, in5631_2;
    wire c5631;
    assign in5631_1 = {c4188,s4179[2],s4174[3],s4226[0]};
    assign in5631_2 = {s4189[1],s4180[2],s4175[3],s4227[0]};
    CLA_4 KS_5631(s5631, c5631, in5631_1, in5631_2);
    wire[3:0] s5632, in5632_1, in5632_2;
    wire c5632;
    assign in5632_1 = {c4190,s4181[2],s4176[3],s4228[0]};
    assign in5632_2 = {s4191[1],s4182[2],s4177[3],s4229[0]};
    CLA_4 KS_5632(s5632, c5632, in5632_1, in5632_2);
    wire[3:0] s5633, in5633_1, in5633_2;
    wire c5633;
    assign in5633_1 = {c4192,s4183[2],s4178[3],s4230[0]};
    assign in5633_2 = {s4193[1],s4184[2],s4179[3],s4231[0]};
    CLA_4 KS_5633(s5633, c5633, in5633_1, in5633_2);
    wire[3:0] s5634, in5634_1, in5634_2;
    wire c5634;
    assign in5634_1 = {c4194,s4185[2],s4180[3],s4232[0]};
    assign in5634_2 = {s4195[1],s4186[2],s4181[3],s4233[0]};
    CLA_4 KS_5634(s5634, c5634, in5634_1, in5634_2);
    wire[3:0] s5635, in5635_1, in5635_2;
    wire c5635;
    assign in5635_1 = {c4196,c4187,s4182[3],s4234[0]};
    assign in5635_2 = {s4197[1],s4189[2],s4183[3],s4235[0]};
    CLA_4 KS_5635(s5635, c5635, in5635_1, in5635_2);
    wire[3:0] s5636, in5636_1, in5636_2;
    wire c5636;
    assign in5636_1 = {c4198,c4191,s4184[3],s4236[0]};
    assign in5636_2 = {s4199[1],s4193[2],s4185[3],s4237[0]};
    CLA_4 KS_5636(s5636, c5636, in5636_1, in5636_2);
    wire[3:0] s5637, in5637_1, in5637_2;
    wire c5637;
    assign in5637_1 = {c4200,c4195,s4186[3],s4238[0]};
    assign in5637_2 = {s4201[1],s4197[2],s4189[3],s4239[0]};
    CLA_4 KS_5637(s5637, c5637, in5637_1, in5637_2);
    wire[0:0] s5638, in5638_1, in5638_2;
    wire c5638;
    assign in5638_1 = {c4202};
    assign in5638_2 = {s4203[1]};
    Half_Adder KS_5638(s5638, c5638, in5638_1, in5638_2);
    wire[1:0] s5639, in5639_1, in5639_2;
    wire c5639;
    assign in5639_1 = {c4204,c4199};
    assign in5639_2 = {s4205[1],s4201[2]};
    CLA_2 KS_5639(s5639, c5639, in5639_1, in5639_2);
    wire[0:0] s5640, in5640_1, in5640_2;
    wire c5640;
    assign in5640_1 = {c4206};
    assign in5640_2 = {c5604};
    Half_Adder KS_5640(s5640, c5640, in5640_1, in5640_2);
    wire[3:0] s5641, in5641_1, in5641_2;
    wire c5641;
    assign in5641_1 = {c5605,c4203,c4193,s4240[0]};
    assign in5641_2 = {c5606,s4205[2],s4197[3],s4241[0]};
    CLA_4 KS_5641(s5641, c5641, in5641_1, in5641_2);
    wire[0:0] s5642, in5642_1, in5642_2;
    wire c5642;
    assign in5642_1 = {c5607};
    assign in5642_2 = {c5608};
    Half_Adder KS_5642(s5642, c5642, in5642_1, in5642_2);
    wire[1:0] s5643, in5643_1, in5643_2;
    wire c5643;
    assign in5643_1 = {c5609,s5627[1]};
    assign in5643_2 = {c5610,s5628[1]};
    CLA_2 KS_5643(s5643, c5643, in5643_1, in5643_2);
    wire[0:0] s5644, in5644_1, in5644_2;
    wire c5644;
    assign in5644_1 = {c5611};
    assign in5644_2 = {c5612};
    Half_Adder KS_5644(s5644, c5644, in5644_1, in5644_2);
    wire[2:0] s5645, in5645_1, in5645_2;
    wire c5645;
    assign in5645_1 = {c5613,s5629[1],c4201};
    assign in5645_2 = {c5614,s5630[1],s4205[3]};
    CLA_3 KS_5645(s5645, c5645, in5645_1, in5645_2);
    wire[0:0] s5646, in5646_1, in5646_2;
    wire c5646;
    assign in5646_1 = {c5618};
    assign in5646_2 = {c5626};
    Half_Adder KS_5646(s5646, c5646, in5646_1, in5646_2);
    wire[1:0] s5647, in5647_1, in5647_2;
    wire c5647;
    assign in5647_1 = {s5627[0],s5631[1]};
    assign in5647_2 = {s5628[0],s5632[1]};
    CLA_2 KS_5647(s5647, c5647, in5647_1, in5647_2);
    wire[0:0] s5648, in5648_1, in5648_2;
    wire c5648;
    assign in5648_1 = {s5629[0]};
    assign in5648_2 = {s5630[0]};
    Half_Adder KS_5648(s5648, c5648, in5648_1, in5648_2);
    wire[3:0] s5649, in5649_1, in5649_2;
    wire c5649;
    assign in5649_1 = {s5632[0],s5633[1],s5627[2],s4242[0]};
    assign in5649_2 = {s5633[0],s5634[1],s5628[2],s4243[0]};
    CLA_4_c KS_5649(s5649, c5649, in5649_1, in5649_2, s5631[0]);
    wire[3:0] s5650, in5650_1, in5650_2;
    wire c5650;
    assign in5650_1 = {s4218[1],s4209[2],c2354,s4254[0]};
    assign in5650_2 = {s4219[1],s4210[2],s2356[2],s4255[0]};
    CLA_4 KS_5650(s5650, c5650, in5650_1, in5650_2);
    wire[3:0] s5651, in5651_1, in5651_2;
    wire c5651;
    assign in5651_1 = {s4220[1],s4211[2],c2358,s4256[0]};
    assign in5651_2 = {s4221[1],s4212[2],s2360[2],s4257[0]};
    CLA_4 KS_5651(s5651, c5651, in5651_1, in5651_2);
    wire[3:0] s5652, in5652_1, in5652_2;
    wire c5652;
    assign in5652_1 = {s4222[1],s4213[2],s4207[3],s4258[0]};
    assign in5652_2 = {s4223[1],s4214[2],s4208[3],s4259[0]};
    CLA_4 KS_5652(s5652, c5652, in5652_1, in5652_2);
    wire[3:0] s5653, in5653_1, in5653_2;
    wire c5653;
    assign in5653_1 = {s4224[1],s4215[2],s4209[3],s4260[0]};
    assign in5653_2 = {s4225[1],s4216[2],s4210[3],s4261[0]};
    CLA_4 KS_5653(s5653, c5653, in5653_1, in5653_2);
    wire[3:0] s5654, in5654_1, in5654_2;
    wire c5654;
    assign in5654_1 = {c4226,s4217[2],s4211[3],s4262[0]};
    assign in5654_2 = {s4227[1],s4218[2],s4212[3],s4263[0]};
    CLA_4 KS_5654(s5654, c5654, in5654_1, in5654_2);
    wire[3:0] s5655, in5655_1, in5655_2;
    wire c5655;
    assign in5655_1 = {c4228,s4219[2],s4213[3],s4264[0]};
    assign in5655_2 = {s4229[1],s4220[2],s4214[3],s4265[0]};
    CLA_4 KS_5655(s5655, c5655, in5655_1, in5655_2);
    wire[3:0] s5656, in5656_1, in5656_2;
    wire c5656;
    assign in5656_1 = {c4230,s4221[2],s4215[3],s4266[0]};
    assign in5656_2 = {s4231[1],s4222[2],s4216[3],s4267[0]};
    CLA_4 KS_5656(s5656, c5656, in5656_1, in5656_2);
    wire[3:0] s5657, in5657_1, in5657_2;
    wire c5657;
    assign in5657_1 = {c4232,s4223[2],s4217[3],s4268[0]};
    assign in5657_2 = {s4233[1],s4224[2],s4218[3],s4269[0]};
    CLA_4 KS_5657(s5657, c5657, in5657_1, in5657_2);
    wire[3:0] s5658, in5658_1, in5658_2;
    wire c5658;
    assign in5658_1 = {c4234,c4225,s4219[3],s4270[0]};
    assign in5658_2 = {s4235[1],s4227[2],s4220[3],s4271[0]};
    CLA_4 KS_5658(s5658, c5658, in5658_1, in5658_2);
    wire[3:0] s5659, in5659_1, in5659_2;
    wire c5659;
    assign in5659_1 = {c4236,c4229,s4221[3],s4272[0]};
    assign in5659_2 = {s4237[1],s4231[2],s4222[3],s4273[0]};
    CLA_4 KS_5659(s5659, c5659, in5659_1, in5659_2);
    wire[3:0] s5660, in5660_1, in5660_2;
    wire c5660;
    assign in5660_1 = {c4238,c4233,s4223[3],s4274[0]};
    assign in5660_2 = {s4239[1],s4235[2],s4224[3],s4275[0]};
    CLA_4 KS_5660(s5660, c5660, in5660_1, in5660_2);
    wire[0:0] s5661, in5661_1, in5661_2;
    wire c5661;
    assign in5661_1 = {c4240};
    assign in5661_2 = {s4241[1]};
    Half_Adder KS_5661(s5661, c5661, in5661_1, in5661_2);
    wire[3:0] s5662, in5662_1, in5662_2;
    wire c5662;
    assign in5662_1 = {c4242,c4237,c4227,s4276[0]};
    assign in5662_2 = {s4243[1],s4239[2],s4231[3],s4277[0]};
    CLA_4 KS_5662(s5662, c5662, in5662_1, in5662_2);
    wire[0:0] s5663, in5663_1, in5663_2;
    wire c5663;
    assign in5663_1 = {c4244};
    assign in5663_2 = {c5627};
    Half_Adder KS_5663(s5663, c5663, in5663_1, in5663_2);
    wire[1:0] s5664, in5664_1, in5664_2;
    wire c5664;
    assign in5664_1 = {c5628,c4241};
    assign in5664_2 = {c5629,s4243[2]};
    CLA_2 KS_5664(s5664, c5664, in5664_1, in5664_2);
    wire[0:0] s5665, in5665_1, in5665_2;
    wire c5665;
    assign in5665_1 = {c5630};
    assign in5665_2 = {c5631};
    Half_Adder KS_5665(s5665, c5665, in5665_1, in5665_2);
    wire[2:0] s5666, in5666_1, in5666_2;
    wire c5666;
    assign in5666_1 = {c5632,s5650[1],c4235};
    assign in5666_2 = {c5633,s5651[1],s4239[3]};
    CLA_3 KS_5666(s5666, c5666, in5666_1, in5666_2);
    wire[0:0] s5667, in5667_1, in5667_2;
    wire c5667;
    assign in5667_1 = {c5634};
    assign in5667_2 = {c5635};
    Half_Adder KS_5667(s5667, c5667, in5667_1, in5667_2);
    wire[1:0] s5668, in5668_1, in5668_2;
    wire c5668;
    assign in5668_1 = {c5636,s5652[1]};
    assign in5668_2 = {c5637,s5653[1]};
    CLA_2 KS_5668(s5668, c5668, in5668_1, in5668_2);
    wire[0:0] s5669, in5669_1, in5669_2;
    wire c5669;
    assign in5669_1 = {c5641};
    assign in5669_2 = {c5649};
    Half_Adder KS_5669(s5669, c5669, in5669_1, in5669_2);
    wire[3:0] s5670, in5670_1, in5670_2;
    wire c5670;
    assign in5670_1 = {s5650[0],s5654[1],c4243,s4278[0]};
    assign in5670_2 = {s5651[0],s5655[1],s5650[2],s4279[0]};
    CLA_4 KS_5670(s5670, c5670, in5670_1, in5670_2);
    wire[0:0] s5671, in5671_1, in5671_2;
    wire c5671;
    assign in5671_1 = {s5652[0]};
    assign in5671_2 = {s5653[0]};
    Half_Adder KS_5671(s5671, c5671, in5671_1, in5671_2);
    wire[1:0] s5672, in5672_1, in5672_2;
    wire c5672;
    assign in5672_1 = {s5655[0],s5656[1]};
    assign in5672_2 = {s5656[0],s5657[1]};
    CLA_2_c KS_5672(s5672, c5672, in5672_1, in5672_2, s5654[0]);
    wire[3:0] s5673, in5673_1, in5673_2;
    wire c5673;
    assign in5673_1 = {s4254[1],s4246[2],c2418,s4290[0]};
    assign in5673_2 = {s4255[1],s4247[2],s2420[2],s4291[0]};
    CLA_4 KS_5673(s5673, c5673, in5673_1, in5673_2);
    wire[3:0] s5674, in5674_1, in5674_2;
    wire c5674;
    assign in5674_1 = {s4256[1],s4248[2],c2422,s4292[0]};
    assign in5674_2 = {s4257[1],s4249[2],s2424[2],s4293[0]};
    CLA_4 KS_5674(s5674, c5674, in5674_1, in5674_2);
    wire[3:0] s5675, in5675_1, in5675_2;
    wire c5675;
    assign in5675_1 = {s4258[1],s4250[2],s4245[3],s4294[0]};
    assign in5675_2 = {s4259[1],s4251[2],s4246[3],s4295[0]};
    CLA_4 KS_5675(s5675, c5675, in5675_1, in5675_2);
    wire[3:0] s5676, in5676_1, in5676_2;
    wire c5676;
    assign in5676_1 = {s4260[1],s4252[2],s4247[3],s4296[0]};
    assign in5676_2 = {s4261[1],s4253[2],s4248[3],s4297[0]};
    CLA_4 KS_5676(s5676, c5676, in5676_1, in5676_2);
    wire[3:0] s5677, in5677_1, in5677_2;
    wire c5677;
    assign in5677_1 = {s4262[1],s4254[2],s4249[3],s4298[0]};
    assign in5677_2 = {s4263[1],s4255[2],s4250[3],s4299[0]};
    CLA_4 KS_5677(s5677, c5677, in5677_1, in5677_2);
    wire[3:0] s5678, in5678_1, in5678_2;
    wire c5678;
    assign in5678_1 = {c4264,s4256[2],s4251[3],s4300[0]};
    assign in5678_2 = {s4265[1],s4257[2],s4252[3],s4301[0]};
    CLA_4 KS_5678(s5678, c5678, in5678_1, in5678_2);
    wire[3:0] s5679, in5679_1, in5679_2;
    wire c5679;
    assign in5679_1 = {c4266,s4258[2],s4253[3],s4302[0]};
    assign in5679_2 = {s4267[1],s4259[2],s4254[3],s4303[0]};
    CLA_4 KS_5679(s5679, c5679, in5679_1, in5679_2);
    wire[3:0] s5680, in5680_1, in5680_2;
    wire c5680;
    assign in5680_1 = {c4268,s4260[2],s4255[3],s4304[0]};
    assign in5680_2 = {s4269[1],s4261[2],s4256[3],s4305[0]};
    CLA_4 KS_5680(s5680, c5680, in5680_1, in5680_2);
    wire[3:0] s5681, in5681_1, in5681_2;
    wire c5681;
    assign in5681_1 = {c4270,s4262[2],s4257[3],s4306[0]};
    assign in5681_2 = {s4271[1],s4263[2],s4258[3],s4307[0]};
    CLA_4 KS_5681(s5681, c5681, in5681_1, in5681_2);
    wire[3:0] s5682, in5682_1, in5682_2;
    wire c5682;
    assign in5682_1 = {c4272,c4265,s4259[3],s4308[0]};
    assign in5682_2 = {s4273[1],s4267[2],s4260[3],s4309[0]};
    CLA_4 KS_5682(s5682, c5682, in5682_1, in5682_2);
    wire[3:0] s5683, in5683_1, in5683_2;
    wire c5683;
    assign in5683_1 = {c4274,c4269,s4261[3],s4310[0]};
    assign in5683_2 = {s4275[1],s4271[2],s4262[3],s4311[0]};
    CLA_4 KS_5683(s5683, c5683, in5683_1, in5683_2);
    wire[0:0] s5684, in5684_1, in5684_2;
    wire c5684;
    assign in5684_1 = {c4276};
    assign in5684_2 = {s4277[1]};
    Half_Adder KS_5684(s5684, c5684, in5684_1, in5684_2);
    wire[3:0] s5685, in5685_1, in5685_2;
    wire c5685;
    assign in5685_1 = {c4278,c4273,c4263,s4312[0]};
    assign in5685_2 = {s4279[1],s4275[2],s4267[3],s4313[0]};
    CLA_4 KS_5685(s5685, c5685, in5685_1, in5685_2);
    wire[0:0] s5686, in5686_1, in5686_2;
    wire c5686;
    assign in5686_1 = {c4280};
    assign in5686_2 = {c5650};
    Half_Adder KS_5686(s5686, c5686, in5686_1, in5686_2);
    wire[1:0] s5687, in5687_1, in5687_2;
    wire c5687;
    assign in5687_1 = {c5651,c4277};
    assign in5687_2 = {c5652,s4279[2]};
    CLA_2 KS_5687(s5687, c5687, in5687_1, in5687_2);
    wire[0:0] s5688, in5688_1, in5688_2;
    wire c5688;
    assign in5688_1 = {c5653};
    assign in5688_2 = {c5654};
    Half_Adder KS_5688(s5688, c5688, in5688_1, in5688_2);
    wire[2:0] s5689, in5689_1, in5689_2;
    wire c5689;
    assign in5689_1 = {c5655,s5673[1],c4271};
    assign in5689_2 = {c5656,s5674[1],s4275[3]};
    CLA_3 KS_5689(s5689, c5689, in5689_1, in5689_2);
    wire[0:0] s5690, in5690_1, in5690_2;
    wire c5690;
    assign in5690_1 = {c5657};
    assign in5690_2 = {c5658};
    Half_Adder KS_5690(s5690, c5690, in5690_1, in5690_2);
    wire[1:0] s5691, in5691_1, in5691_2;
    wire c5691;
    assign in5691_1 = {c5659,s5675[1]};
    assign in5691_2 = {c5660,s5676[1]};
    CLA_2 KS_5691(s5691, c5691, in5691_1, in5691_2);
    wire[0:0] s5692, in5692_1, in5692_2;
    wire c5692;
    assign in5692_1 = {c5662};
    assign in5692_2 = {c5670};
    Half_Adder KS_5692(s5692, c5692, in5692_1, in5692_2);
    wire[3:0] s5693, in5693_1, in5693_2;
    wire c5693;
    assign in5693_1 = {s5673[0],s5677[1],c4279,s4314[0]};
    assign in5693_2 = {s5674[0],s5678[1],s5673[2],s4315[0]};
    CLA_4 KS_5693(s5693, c5693, in5693_1, in5693_2);
    wire[0:0] s5694, in5694_1, in5694_2;
    wire c5694;
    assign in5694_1 = {s5675[0]};
    assign in5694_2 = {s5676[0]};
    Half_Adder KS_5694(s5694, c5694, in5694_1, in5694_2);
    wire[1:0] s5695, in5695_1, in5695_2;
    wire c5695;
    assign in5695_1 = {s5678[0],s5679[1]};
    assign in5695_2 = {s5679[0],s5680[1]};
    CLA_2_c KS_5695(s5695, c5695, in5695_1, in5695_2, s5677[0]);
    wire[3:0] s5696, in5696_1, in5696_2;
    wire c5696;
    assign in5696_1 = {s4290[1],s4282[2],c2485,s4328[0]};
    assign in5696_2 = {s4291[1],s4283[2],s2487[2],s4329[0]};
    CLA_4 KS_5696(s5696, c5696, in5696_1, in5696_2);
    wire[3:0] s5697, in5697_1, in5697_2;
    wire c5697;
    assign in5697_1 = {s4292[1],s4284[2],c2489,s4330[0]};
    assign in5697_2 = {s4293[1],s4285[2],s4281[3],s4331[0]};
    CLA_4 KS_5697(s5697, c5697, in5697_1, in5697_2);
    wire[3:0] s5698, in5698_1, in5698_2;
    wire c5698;
    assign in5698_1 = {s4294[1],s4286[2],s4282[3],s4332[0]};
    assign in5698_2 = {s4295[1],s4287[2],s4283[3],s4333[0]};
    CLA_4 KS_5698(s5698, c5698, in5698_1, in5698_2);
    wire[3:0] s5699, in5699_1, in5699_2;
    wire c5699;
    assign in5699_1 = {s4296[1],s4288[2],s4284[3],s4334[0]};
    assign in5699_2 = {s4297[1],s4289[2],s4285[3],s4335[0]};
    CLA_4 KS_5699(s5699, c5699, in5699_1, in5699_2);
    wire[3:0] s5700, in5700_1, in5700_2;
    wire c5700;
    assign in5700_1 = {s4298[1],s4290[2],s4286[3],s4336[0]};
    assign in5700_2 = {s4299[1],s4291[2],s4287[3],s4337[0]};
    CLA_4 KS_5700(s5700, c5700, in5700_1, in5700_2);
    wire[3:0] s5701, in5701_1, in5701_2;
    wire c5701;
    assign in5701_1 = {c4300,s4292[2],s4288[3],s4338[0]};
    assign in5701_2 = {s4301[1],s4293[2],s4289[3],s4339[0]};
    CLA_4 KS_5701(s5701, c5701, in5701_1, in5701_2);
    wire[3:0] s5702, in5702_1, in5702_2;
    wire c5702;
    assign in5702_1 = {c4302,s4294[2],s4290[3],s4340[0]};
    assign in5702_2 = {s4303[1],s4295[2],s4291[3],s4341[0]};
    CLA_4 KS_5702(s5702, c5702, in5702_1, in5702_2);
    wire[3:0] s5703, in5703_1, in5703_2;
    wire c5703;
    assign in5703_1 = {c4304,s4296[2],s4292[3],s4342[0]};
    assign in5703_2 = {s4305[1],s4297[2],s4293[3],s4343[0]};
    CLA_4 KS_5703(s5703, c5703, in5703_1, in5703_2);
    wire[3:0] s5704, in5704_1, in5704_2;
    wire c5704;
    assign in5704_1 = {c4306,s4298[2],s4294[3],s4344[0]};
    assign in5704_2 = {s4307[1],s4299[2],s4295[3],s4345[0]};
    CLA_4 KS_5704(s5704, c5704, in5704_1, in5704_2);
    wire[3:0] s5705, in5705_1, in5705_2;
    wire c5705;
    assign in5705_1 = {c4308,c4301,s4296[3],s4346[0]};
    assign in5705_2 = {s4309[1],s4303[2],s4297[3],s4347[0]};
    CLA_4 KS_5705(s5705, c5705, in5705_1, in5705_2);
    wire[3:0] s5706, in5706_1, in5706_2;
    wire c5706;
    assign in5706_1 = {c4310,c4305,s4298[3],s4348[0]};
    assign in5706_2 = {s4311[1],s4307[2],s4299[3],s4349[0]};
    CLA_4 KS_5706(s5706, c5706, in5706_1, in5706_2);
    wire[0:0] s5707, in5707_1, in5707_2;
    wire c5707;
    assign in5707_1 = {c4312};
    assign in5707_2 = {s4313[1]};
    Half_Adder KS_5707(s5707, c5707, in5707_1, in5707_2);
    wire[1:0] s5708, in5708_1, in5708_2;
    wire c5708;
    assign in5708_1 = {c4314,c4309};
    assign in5708_2 = {s4315[1],s4311[2]};
    CLA_2 KS_5708(s5708, c5708, in5708_1, in5708_2);
    wire[0:0] s5709, in5709_1, in5709_2;
    wire c5709;
    assign in5709_1 = {c4316};
    assign in5709_2 = {c5673};
    Half_Adder KS_5709(s5709, c5709, in5709_1, in5709_2);
    wire[3:0] s5710, in5710_1, in5710_2;
    wire c5710;
    assign in5710_1 = {c5674,c4313,c4303,s4350[0]};
    assign in5710_2 = {c5675,s4315[2],s4307[3],s4351[0]};
    CLA_4 KS_5710(s5710, c5710, in5710_1, in5710_2);
    wire[0:0] s5711, in5711_1, in5711_2;
    wire c5711;
    assign in5711_1 = {c5676};
    assign in5711_2 = {c5677};
    Half_Adder KS_5711(s5711, c5711, in5711_1, in5711_2);
    wire[1:0] s5712, in5712_1, in5712_2;
    wire c5712;
    assign in5712_1 = {c5678,s5696[1]};
    assign in5712_2 = {c5679,s5697[1]};
    CLA_2 KS_5712(s5712, c5712, in5712_1, in5712_2);
    wire[0:0] s5713, in5713_1, in5713_2;
    wire c5713;
    assign in5713_1 = {c5680};
    assign in5713_2 = {c5681};
    Half_Adder KS_5713(s5713, c5713, in5713_1, in5713_2);
    wire[2:0] s5714, in5714_1, in5714_2;
    wire c5714;
    assign in5714_1 = {c5682,s5698[1],c4311};
    assign in5714_2 = {c5683,s5699[1],s4315[3]};
    CLA_3 KS_5714(s5714, c5714, in5714_1, in5714_2);
    wire[0:0] s5715, in5715_1, in5715_2;
    wire c5715;
    assign in5715_1 = {c5685};
    assign in5715_2 = {c5693};
    Half_Adder KS_5715(s5715, c5715, in5715_1, in5715_2);
    wire[1:0] s5716, in5716_1, in5716_2;
    wire c5716;
    assign in5716_1 = {s5696[0],s5700[1]};
    assign in5716_2 = {s5697[0],s5701[1]};
    CLA_2 KS_5716(s5716, c5716, in5716_1, in5716_2);
    wire[0:0] s5717, in5717_1, in5717_2;
    wire c5717;
    assign in5717_1 = {s5698[0]};
    assign in5717_2 = {s5699[0]};
    Half_Adder KS_5717(s5717, c5717, in5717_1, in5717_2);
    wire[3:0] s5718, in5718_1, in5718_2;
    wire c5718;
    assign in5718_1 = {s5701[0],s5702[1],s5696[2],s4352[0]};
    assign in5718_2 = {s5702[0],s5703[1],s5697[2],s4353[0]};
    CLA_4_c KS_5718(s5718, c5718, in5718_1, in5718_2, s5700[0]);
    wire[3:0] s5719, in5719_1, in5719_2;
    wire c5719;
    assign in5719_1 = {s4328[1],s4319[2],c2548,s4364[0]};
    assign in5719_2 = {s4329[1],s4320[2],s2550[2],s4365[0]};
    CLA_4 KS_5719(s5719, c5719, in5719_1, in5719_2);
    wire[3:0] s5720, in5720_1, in5720_2;
    wire c5720;
    assign in5720_1 = {s4330[1],s4321[2],c2552,s4366[0]};
    assign in5720_2 = {s4331[1],s4322[2],s2554[2],s4367[0]};
    CLA_4 KS_5720(s5720, c5720, in5720_1, in5720_2);
    wire[3:0] s5721, in5721_1, in5721_2;
    wire c5721;
    assign in5721_1 = {s4332[1],s4323[2],s4317[3],s4368[0]};
    assign in5721_2 = {s4333[1],s4324[2],s4318[3],s4369[0]};
    CLA_4 KS_5721(s5721, c5721, in5721_1, in5721_2);
    wire[3:0] s5722, in5722_1, in5722_2;
    wire c5722;
    assign in5722_1 = {s4334[1],s4325[2],s4319[3],s4370[0]};
    assign in5722_2 = {s4335[1],s4326[2],s4320[3],s4371[0]};
    CLA_4 KS_5722(s5722, c5722, in5722_1, in5722_2);
    wire[3:0] s5723, in5723_1, in5723_2;
    wire c5723;
    assign in5723_1 = {c4336,s4327[2],s4321[3],s4372[0]};
    assign in5723_2 = {s4337[1],s4328[2],s4322[3],s4373[0]};
    CLA_4 KS_5723(s5723, c5723, in5723_1, in5723_2);
    wire[3:0] s5724, in5724_1, in5724_2;
    wire c5724;
    assign in5724_1 = {c4338,s4329[2],s4323[3],s4374[0]};
    assign in5724_2 = {s4339[1],s4330[2],s4324[3],s4375[0]};
    CLA_4 KS_5724(s5724, c5724, in5724_1, in5724_2);
    wire[3:0] s5725, in5725_1, in5725_2;
    wire c5725;
    assign in5725_1 = {c4340,s4331[2],s4325[3],s4376[0]};
    assign in5725_2 = {s4341[1],s4332[2],s4326[3],s4377[0]};
    CLA_4 KS_5725(s5725, c5725, in5725_1, in5725_2);
    wire[3:0] s5726, in5726_1, in5726_2;
    wire c5726;
    assign in5726_1 = {c4342,s4333[2],s4327[3],s4378[0]};
    assign in5726_2 = {s4343[1],s4334[2],s4328[3],s4379[0]};
    CLA_4 KS_5726(s5726, c5726, in5726_1, in5726_2);
    wire[3:0] s5727, in5727_1, in5727_2;
    wire c5727;
    assign in5727_1 = {c4344,c4335,s4329[3],s4380[0]};
    assign in5727_2 = {s4345[1],s4337[2],s4330[3],s4381[0]};
    CLA_4 KS_5727(s5727, c5727, in5727_1, in5727_2);
    wire[3:0] s5728, in5728_1, in5728_2;
    wire c5728;
    assign in5728_1 = {c4346,c4339,s4331[3],s4382[0]};
    assign in5728_2 = {s4347[1],s4341[2],s4332[3],s4383[0]};
    CLA_4 KS_5728(s5728, c5728, in5728_1, in5728_2);
    wire[3:0] s5729, in5729_1, in5729_2;
    wire c5729;
    assign in5729_1 = {c4348,c4343,s4333[3],s4384[0]};
    assign in5729_2 = {s4349[1],s4345[2],s4334[3],s4385[0]};
    CLA_4 KS_5729(s5729, c5729, in5729_1, in5729_2);
    wire[0:0] s5730, in5730_1, in5730_2;
    wire c5730;
    assign in5730_1 = {c4350};
    assign in5730_2 = {s4351[1]};
    Half_Adder KS_5730(s5730, c5730, in5730_1, in5730_2);
    wire[3:0] s5731, in5731_1, in5731_2;
    wire c5731;
    assign in5731_1 = {c4352,c4347,c4337,s4386[0]};
    assign in5731_2 = {s4353[1],s4349[2],s4341[3],s4387[0]};
    CLA_4 KS_5731(s5731, c5731, in5731_1, in5731_2);
    wire[0:0] s5732, in5732_1, in5732_2;
    wire c5732;
    assign in5732_1 = {c4354};
    assign in5732_2 = {c5696};
    Half_Adder KS_5732(s5732, c5732, in5732_1, in5732_2);
    wire[1:0] s5733, in5733_1, in5733_2;
    wire c5733;
    assign in5733_1 = {c5697,c4351};
    assign in5733_2 = {c5698,s4353[2]};
    CLA_2 KS_5733(s5733, c5733, in5733_1, in5733_2);
    wire[0:0] s5734, in5734_1, in5734_2;
    wire c5734;
    assign in5734_1 = {c5699};
    assign in5734_2 = {c5700};
    Half_Adder KS_5734(s5734, c5734, in5734_1, in5734_2);
    wire[2:0] s5735, in5735_1, in5735_2;
    wire c5735;
    assign in5735_1 = {c5701,s5719[1],c4345};
    assign in5735_2 = {c5702,s5720[1],s4349[3]};
    CLA_3 KS_5735(s5735, c5735, in5735_1, in5735_2);
    wire[0:0] s5736, in5736_1, in5736_2;
    wire c5736;
    assign in5736_1 = {c5703};
    assign in5736_2 = {c5704};
    Half_Adder KS_5736(s5736, c5736, in5736_1, in5736_2);
    wire[1:0] s5737, in5737_1, in5737_2;
    wire c5737;
    assign in5737_1 = {c5705,s5721[1]};
    assign in5737_2 = {c5706,s5722[1]};
    CLA_2 KS_5737(s5737, c5737, in5737_1, in5737_2);
    wire[0:0] s5738, in5738_1, in5738_2;
    wire c5738;
    assign in5738_1 = {c5710};
    assign in5738_2 = {c5718};
    Half_Adder KS_5738(s5738, c5738, in5738_1, in5738_2);
    wire[3:0] s5739, in5739_1, in5739_2;
    wire c5739;
    assign in5739_1 = {s5719[0],s5723[1],c4353,s4388[0]};
    assign in5739_2 = {s5720[0],s5724[1],s5719[2],s4389[0]};
    CLA_4 KS_5739(s5739, c5739, in5739_1, in5739_2);
    wire[0:0] s5740, in5740_1, in5740_2;
    wire c5740;
    assign in5740_1 = {s5721[0]};
    assign in5740_2 = {s5722[0]};
    Half_Adder KS_5740(s5740, c5740, in5740_1, in5740_2);
    wire[1:0] s5741, in5741_1, in5741_2;
    wire c5741;
    assign in5741_1 = {s5724[0],s5725[1]};
    assign in5741_2 = {s5725[0],s5726[1]};
    CLA_2_c KS_5741(s5741, c5741, in5741_1, in5741_2, s5723[0]);
    wire[3:0] s5742, in5742_1, in5742_2;
    wire c5742;
    assign in5742_1 = {s4364[1],s4356[2],c2615,s4402[0]};
    assign in5742_2 = {s4365[1],s4357[2],s2617[2],s4403[0]};
    CLA_4 KS_5742(s5742, c5742, in5742_1, in5742_2);
    wire[3:0] s5743, in5743_1, in5743_2;
    wire c5743;
    assign in5743_1 = {s4366[1],s4358[2],c2619,s4404[0]};
    assign in5743_2 = {s4367[1],s4359[2],s4355[3],s4405[0]};
    CLA_4 KS_5743(s5743, c5743, in5743_1, in5743_2);
    wire[3:0] s5744, in5744_1, in5744_2;
    wire c5744;
    assign in5744_1 = {s4368[1],s4360[2],s4356[3],s4406[0]};
    assign in5744_2 = {s4369[1],s4361[2],s4357[3],s4407[0]};
    CLA_4 KS_5744(s5744, c5744, in5744_1, in5744_2);
    wire[3:0] s5745, in5745_1, in5745_2;
    wire c5745;
    assign in5745_1 = {s4370[1],s4362[2],s4358[3],s4408[0]};
    assign in5745_2 = {s4371[1],s4363[2],s4359[3],s4409[0]};
    CLA_4 KS_5745(s5745, c5745, in5745_1, in5745_2);
    wire[3:0] s5746, in5746_1, in5746_2;
    wire c5746;
    assign in5746_1 = {s4372[1],s4364[2],s4360[3],s4410[0]};
    assign in5746_2 = {s4373[1],s4365[2],s4361[3],s4411[0]};
    CLA_4 KS_5746(s5746, c5746, in5746_1, in5746_2);
    wire[3:0] s5747, in5747_1, in5747_2;
    wire c5747;
    assign in5747_1 = {c4374,s4366[2],s4362[3],s4412[0]};
    assign in5747_2 = {s4375[1],s4367[2],s4363[3],s4413[0]};
    CLA_4 KS_5747(s5747, c5747, in5747_1, in5747_2);
    wire[3:0] s5748, in5748_1, in5748_2;
    wire c5748;
    assign in5748_1 = {c4376,s4368[2],s4364[3],s4414[0]};
    assign in5748_2 = {s4377[1],s4369[2],s4365[3],s4415[0]};
    CLA_4 KS_5748(s5748, c5748, in5748_1, in5748_2);
    wire[3:0] s5749, in5749_1, in5749_2;
    wire c5749;
    assign in5749_1 = {c4378,s4370[2],s4366[3],s4416[0]};
    assign in5749_2 = {s4379[1],s4371[2],s4367[3],s4417[0]};
    CLA_4 KS_5749(s5749, c5749, in5749_1, in5749_2);
    wire[3:0] s5750, in5750_1, in5750_2;
    wire c5750;
    assign in5750_1 = {c4380,s4372[2],s4368[3],s4418[0]};
    assign in5750_2 = {s4381[1],s4373[2],s4369[3],s4419[0]};
    CLA_4 KS_5750(s5750, c5750, in5750_1, in5750_2);
    wire[3:0] s5751, in5751_1, in5751_2;
    wire c5751;
    assign in5751_1 = {c4382,c4375,s4370[3],s4420[0]};
    assign in5751_2 = {s4383[1],s4377[2],s4371[3],s4421[0]};
    CLA_4 KS_5751(s5751, c5751, in5751_1, in5751_2);
    wire[3:0] s5752, in5752_1, in5752_2;
    wire c5752;
    assign in5752_1 = {c4384,c4379,s4372[3],s4422[0]};
    assign in5752_2 = {s4385[1],s4381[2],s4373[3],s4423[0]};
    CLA_4 KS_5752(s5752, c5752, in5752_1, in5752_2);
    wire[0:0] s5753, in5753_1, in5753_2;
    wire c5753;
    assign in5753_1 = {c4386};
    assign in5753_2 = {s4387[1]};
    Half_Adder KS_5753(s5753, c5753, in5753_1, in5753_2);
    wire[1:0] s5754, in5754_1, in5754_2;
    wire c5754;
    assign in5754_1 = {c4388,c4383};
    assign in5754_2 = {s4389[1],s4385[2]};
    CLA_2 KS_5754(s5754, c5754, in5754_1, in5754_2);
    wire[0:0] s5755, in5755_1, in5755_2;
    wire c5755;
    assign in5755_1 = {c4390};
    assign in5755_2 = {c5719};
    Half_Adder KS_5755(s5755, c5755, in5755_1, in5755_2);
    wire[3:0] s5756, in5756_1, in5756_2;
    wire c5756;
    assign in5756_1 = {c5720,c4387,c4377,s4424[0]};
    assign in5756_2 = {c5721,s4389[2],s4381[3],s4425[0]};
    CLA_4 KS_5756(s5756, c5756, in5756_1, in5756_2);
    wire[0:0] s5757, in5757_1, in5757_2;
    wire c5757;
    assign in5757_1 = {c5722};
    assign in5757_2 = {c5723};
    Half_Adder KS_5757(s5757, c5757, in5757_1, in5757_2);
    wire[1:0] s5758, in5758_1, in5758_2;
    wire c5758;
    assign in5758_1 = {c5724,s5742[1]};
    assign in5758_2 = {c5725,s5743[1]};
    CLA_2 KS_5758(s5758, c5758, in5758_1, in5758_2);
    wire[0:0] s5759, in5759_1, in5759_2;
    wire c5759;
    assign in5759_1 = {c5726};
    assign in5759_2 = {c5727};
    Half_Adder KS_5759(s5759, c5759, in5759_1, in5759_2);
    wire[2:0] s5760, in5760_1, in5760_2;
    wire c5760;
    assign in5760_1 = {c5728,s5744[1],c4385};
    assign in5760_2 = {c5729,s5745[1],s4389[3]};
    CLA_3 KS_5760(s5760, c5760, in5760_1, in5760_2);
    wire[0:0] s5761, in5761_1, in5761_2;
    wire c5761;
    assign in5761_1 = {c5731};
    assign in5761_2 = {c5739};
    Half_Adder KS_5761(s5761, c5761, in5761_1, in5761_2);
    wire[1:0] s5762, in5762_1, in5762_2;
    wire c5762;
    assign in5762_1 = {s5742[0],s5746[1]};
    assign in5762_2 = {s5743[0],s5747[1]};
    CLA_2 KS_5762(s5762, c5762, in5762_1, in5762_2);
    wire[0:0] s5763, in5763_1, in5763_2;
    wire c5763;
    assign in5763_1 = {s5744[0]};
    assign in5763_2 = {s5745[0]};
    Half_Adder KS_5763(s5763, c5763, in5763_1, in5763_2);
    wire[3:0] s5764, in5764_1, in5764_2;
    wire c5764;
    assign in5764_1 = {s5747[0],s5748[1],s5742[2],s4426[0]};
    assign in5764_2 = {s5748[0],s5749[1],s5743[2],s4427[0]};
    CLA_4_c KS_5764(s5764, c5764, in5764_1, in5764_2, s5746[0]);
    wire[3:0] s5765, in5765_1, in5765_2;
    wire c5765;
    assign in5765_1 = {s4402[1],s4393[2],c2679,s4438[0]};
    assign in5765_2 = {s4403[1],s4394[2],s2681[2],s4439[0]};
    CLA_4 KS_5765(s5765, c5765, in5765_1, in5765_2);
    wire[3:0] s5766, in5766_1, in5766_2;
    wire c5766;
    assign in5766_1 = {s4404[1],s4395[2],c2683,s4440[0]};
    assign in5766_2 = {s4405[1],s4396[2],s2685[2],s4441[0]};
    CLA_4 KS_5766(s5766, c5766, in5766_1, in5766_2);
    wire[3:0] s5767, in5767_1, in5767_2;
    wire c5767;
    assign in5767_1 = {s4406[1],s4397[2],s4391[3],s4442[0]};
    assign in5767_2 = {s4407[1],s4398[2],s4392[3],s4443[0]};
    CLA_4 KS_5767(s5767, c5767, in5767_1, in5767_2);
    wire[3:0] s5768, in5768_1, in5768_2;
    wire c5768;
    assign in5768_1 = {s4408[1],s4399[2],s4393[3],s4444[0]};
    assign in5768_2 = {s4409[1],s4400[2],s4394[3],s4445[0]};
    CLA_4 KS_5768(s5768, c5768, in5768_1, in5768_2);
    wire[3:0] s5769, in5769_1, in5769_2;
    wire c5769;
    assign in5769_1 = {c4410,s4401[2],s4395[3],s4446[0]};
    assign in5769_2 = {s4411[1],s4402[2],s4396[3],s4447[0]};
    CLA_4 KS_5769(s5769, c5769, in5769_1, in5769_2);
    wire[3:0] s5770, in5770_1, in5770_2;
    wire c5770;
    assign in5770_1 = {c4412,s4403[2],s4397[3],s4448[0]};
    assign in5770_2 = {s4413[1],s4404[2],s4398[3],s4449[0]};
    CLA_4 KS_5770(s5770, c5770, in5770_1, in5770_2);
    wire[3:0] s5771, in5771_1, in5771_2;
    wire c5771;
    assign in5771_1 = {c4414,s4405[2],s4399[3],s4450[0]};
    assign in5771_2 = {s4415[1],s4406[2],s4400[3],s4451[0]};
    CLA_4 KS_5771(s5771, c5771, in5771_1, in5771_2);
    wire[3:0] s5772, in5772_1, in5772_2;
    wire c5772;
    assign in5772_1 = {c4416,s4407[2],s4401[3],s4452[0]};
    assign in5772_2 = {s4417[1],s4408[2],s4402[3],s4453[0]};
    CLA_4 KS_5772(s5772, c5772, in5772_1, in5772_2);
    wire[3:0] s5773, in5773_1, in5773_2;
    wire c5773;
    assign in5773_1 = {c4418,c4409,s4403[3],s4454[0]};
    assign in5773_2 = {s4419[1],s4411[2],s4404[3],s4455[0]};
    CLA_4 KS_5773(s5773, c5773, in5773_1, in5773_2);
    wire[3:0] s5774, in5774_1, in5774_2;
    wire c5774;
    assign in5774_1 = {c4420,c4413,s4405[3],s4456[0]};
    assign in5774_2 = {s4421[1],s4415[2],s4406[3],s4457[0]};
    CLA_4 KS_5774(s5774, c5774, in5774_1, in5774_2);
    wire[3:0] s5775, in5775_1, in5775_2;
    wire c5775;
    assign in5775_1 = {c4422,c4417,s4407[3],s4458[0]};
    assign in5775_2 = {s4423[1],s4419[2],s4408[3],s4459[0]};
    CLA_4 KS_5775(s5775, c5775, in5775_1, in5775_2);
    wire[0:0] s5776, in5776_1, in5776_2;
    wire c5776;
    assign in5776_1 = {c4424};
    assign in5776_2 = {s4425[1]};
    Half_Adder KS_5776(s5776, c5776, in5776_1, in5776_2);
    wire[3:0] s5777, in5777_1, in5777_2;
    wire c5777;
    assign in5777_1 = {c4426,c4421,c4411,s4460[0]};
    assign in5777_2 = {s4427[1],s4423[2],s4415[3],s4461[0]};
    CLA_4 KS_5777(s5777, c5777, in5777_1, in5777_2);
    wire[0:0] s5778, in5778_1, in5778_2;
    wire c5778;
    assign in5778_1 = {c4428};
    assign in5778_2 = {c5742};
    Half_Adder KS_5778(s5778, c5778, in5778_1, in5778_2);
    wire[1:0] s5779, in5779_1, in5779_2;
    wire c5779;
    assign in5779_1 = {c5743,c4425};
    assign in5779_2 = {c5744,s4427[2]};
    CLA_2 KS_5779(s5779, c5779, in5779_1, in5779_2);
    wire[0:0] s5780, in5780_1, in5780_2;
    wire c5780;
    assign in5780_1 = {c5745};
    assign in5780_2 = {c5746};
    Half_Adder KS_5780(s5780, c5780, in5780_1, in5780_2);
    wire[2:0] s5781, in5781_1, in5781_2;
    wire c5781;
    assign in5781_1 = {c5747,s5765[1],c4419};
    assign in5781_2 = {c5748,s5766[1],s4423[3]};
    CLA_3 KS_5781(s5781, c5781, in5781_1, in5781_2);
    wire[0:0] s5782, in5782_1, in5782_2;
    wire c5782;
    assign in5782_1 = {c5749};
    assign in5782_2 = {c5750};
    Half_Adder KS_5782(s5782, c5782, in5782_1, in5782_2);
    wire[1:0] s5783, in5783_1, in5783_2;
    wire c5783;
    assign in5783_1 = {c5751,s5767[1]};
    assign in5783_2 = {c5752,s5768[1]};
    CLA_2 KS_5783(s5783, c5783, in5783_1, in5783_2);
    wire[0:0] s5784, in5784_1, in5784_2;
    wire c5784;
    assign in5784_1 = {c5756};
    assign in5784_2 = {c5764};
    Half_Adder KS_5784(s5784, c5784, in5784_1, in5784_2);
    wire[3:0] s5785, in5785_1, in5785_2;
    wire c5785;
    assign in5785_1 = {s5765[0],s5769[1],c4427,s4462[0]};
    assign in5785_2 = {s5766[0],s5770[1],s5765[2],s4463[0]};
    CLA_4 KS_5785(s5785, c5785, in5785_1, in5785_2);
    wire[0:0] s5786, in5786_1, in5786_2;
    wire c5786;
    assign in5786_1 = {s5767[0]};
    assign in5786_2 = {s5768[0]};
    Half_Adder KS_5786(s5786, c5786, in5786_1, in5786_2);
    wire[1:0] s5787, in5787_1, in5787_2;
    wire c5787;
    assign in5787_1 = {s5770[0],s5771[1]};
    assign in5787_2 = {s5771[0],s5772[1]};
    CLA_2_c KS_5787(s5787, c5787, in5787_1, in5787_2, s5769[0]);
    wire[3:0] s5788, in5788_1, in5788_2;
    wire c5788;
    assign in5788_1 = {s4438[1],s4429[2],c2742,s4475[0]};
    assign in5788_2 = {s4439[1],s4430[2],s2744[2],s4476[0]};
    CLA_4 KS_5788(s5788, c5788, in5788_1, in5788_2);
    wire[3:0] s5789, in5789_1, in5789_2;
    wire c5789;
    assign in5789_1 = {s4440[1],s4431[2],c2746,s4477[0]};
    assign in5789_2 = {s4441[1],s4432[2],s2748[2],s4478[0]};
    CLA_4 KS_5789(s5789, c5789, in5789_1, in5789_2);
    wire[3:0] s5790, in5790_1, in5790_2;
    wire c5790;
    assign in5790_1 = {s4442[1],s4433[2],c2750,s4479[0]};
    assign in5790_2 = {s4443[1],s4434[2],s4429[3],s4480[0]};
    CLA_4 KS_5790(s5790, c5790, in5790_1, in5790_2);
    wire[3:0] s5791, in5791_1, in5791_2;
    wire c5791;
    assign in5791_1 = {s4444[1],s4435[2],s4430[3],s4481[0]};
    assign in5791_2 = {s4445[1],s4436[2],s4431[3],s4482[0]};
    CLA_4 KS_5791(s5791, c5791, in5791_1, in5791_2);
    wire[3:0] s5792, in5792_1, in5792_2;
    wire c5792;
    assign in5792_1 = {s4446[1],s4437[2],s4432[3],s4483[0]};
    assign in5792_2 = {s4447[1],s4438[2],s4433[3],s4484[0]};
    CLA_4 KS_5792(s5792, c5792, in5792_1, in5792_2);
    wire[3:0] s5793, in5793_1, in5793_2;
    wire c5793;
    assign in5793_1 = {c4448,s4439[2],s4434[3],s4485[0]};
    assign in5793_2 = {s4449[1],s4440[2],s4435[3],s4486[0]};
    CLA_4 KS_5793(s5793, c5793, in5793_1, in5793_2);
    wire[3:0] s5794, in5794_1, in5794_2;
    wire c5794;
    assign in5794_1 = {c4450,s4441[2],s4436[3],s4487[0]};
    assign in5794_2 = {s4451[1],s4442[2],s4437[3],s4488[0]};
    CLA_4 KS_5794(s5794, c5794, in5794_1, in5794_2);
    wire[3:0] s5795, in5795_1, in5795_2;
    wire c5795;
    assign in5795_1 = {c4452,s4443[2],s4438[3],s4489[0]};
    assign in5795_2 = {s4453[1],s4444[2],s4439[3],s4490[0]};
    CLA_4 KS_5795(s5795, c5795, in5795_1, in5795_2);
    wire[3:0] s5796, in5796_1, in5796_2;
    wire c5796;
    assign in5796_1 = {c4454,s4445[2],s4440[3],s4491[0]};
    assign in5796_2 = {s4455[1],s4446[2],s4441[3],s4492[0]};
    CLA_4 KS_5796(s5796, c5796, in5796_1, in5796_2);
    wire[3:0] s5797, in5797_1, in5797_2;
    wire c5797;
    assign in5797_1 = {c4456,c4447,s4442[3],s4493[0]};
    assign in5797_2 = {s4457[1],s4449[2],s4443[3],s4494[0]};
    CLA_4 KS_5797(s5797, c5797, in5797_1, in5797_2);
    wire[3:0] s5798, in5798_1, in5798_2;
    wire c5798;
    assign in5798_1 = {c4458,c4451,s4444[3],s4495[0]};
    assign in5798_2 = {s4459[1],s4453[2],s4445[3],s4496[0]};
    CLA_4 KS_5798(s5798, c5798, in5798_1, in5798_2);
    wire[3:0] s5799, in5799_1, in5799_2;
    wire c5799;
    assign in5799_1 = {c4460,c4455,s4446[3],s4497[0]};
    assign in5799_2 = {s4461[1],s4457[2],s4449[3],s4498[0]};
    CLA_4 KS_5799(s5799, c5799, in5799_1, in5799_2);
    wire[0:0] s5800, in5800_1, in5800_2;
    wire c5800;
    assign in5800_1 = {c4462};
    assign in5800_2 = {s4463[1]};
    Half_Adder KS_5800(s5800, c5800, in5800_1, in5800_2);
    wire[1:0] s5801, in5801_1, in5801_2;
    wire c5801;
    assign in5801_1 = {c4464,c4459};
    assign in5801_2 = {c5765,s4461[2]};
    CLA_2 KS_5801(s5801, c5801, in5801_1, in5801_2);
    wire[0:0] s5802, in5802_1, in5802_2;
    wire c5802;
    assign in5802_1 = {c5766};
    assign in5802_2 = {c5767};
    Half_Adder KS_5802(s5802, c5802, in5802_1, in5802_2);
    wire[2:0] s5803, in5803_1, in5803_2;
    wire c5803;
    assign in5803_1 = {c5768,c4463,c4453};
    assign in5803_2 = {c5769,s5788[1],s4457[3]};
    CLA_3 KS_5803(s5803, c5803, in5803_1, in5803_2);
    wire[0:0] s5804, in5804_1, in5804_2;
    wire c5804;
    assign in5804_1 = {c5770};
    assign in5804_2 = {c5771};
    Half_Adder KS_5804(s5804, c5804, in5804_1, in5804_2);
    wire[1:0] s5805, in5805_1, in5805_2;
    wire c5805;
    assign in5805_1 = {c5772,s5789[1]};
    assign in5805_2 = {c5773,s5790[1]};
    CLA_2 KS_5805(s5805, c5805, in5805_1, in5805_2);
    wire[0:0] s5806, in5806_1, in5806_2;
    wire c5806;
    assign in5806_1 = {c5774};
    assign in5806_2 = {c5775};
    Half_Adder KS_5806(s5806, c5806, in5806_1, in5806_2);
    wire[3:0] s5807, in5807_1, in5807_2;
    wire c5807;
    assign in5807_1 = {c5777,s5791[1],c4461,s4499[0]};
    assign in5807_2 = {c5785,s5792[1],s5788[2],s4500[0]};
    CLA_4 KS_5807(s5807, c5807, in5807_1, in5807_2);
    wire[0:0] s5808, in5808_1, in5808_2;
    wire c5808;
    assign in5808_1 = {s5788[0]};
    assign in5808_2 = {s5789[0]};
    Half_Adder KS_5808(s5808, c5808, in5808_1, in5808_2);
    wire[1:0] s5809, in5809_1, in5809_2;
    wire c5809;
    assign in5809_1 = {s5790[0],s5793[1]};
    assign in5809_2 = {s5791[0],s5794[1]};
    CLA_2 KS_5809(s5809, c5809, in5809_1, in5809_2);
    wire[0:0] s5810, in5810_1, in5810_2;
    wire c5810;
    assign in5810_1 = {s5793[0]};
    assign in5810_2 = {s5794[0]};
    Full_Adder KS_5810(s5810, c5810, in5810_1, in5810_2, s5792[0]);
    wire[3:0] s5811, in5811_1, in5811_2;
    wire c5811;
    assign in5811_1 = {s4476[1],s4466[2],c2809,s4513[0]};
    assign in5811_2 = {s4477[1],s4467[2],s2811[2],s4514[0]};
    CLA_4 KS_5811(s5811, c5811, in5811_1, in5811_2);
    wire[3:0] s5812, in5812_1, in5812_2;
    wire c5812;
    assign in5812_1 = {s4478[1],s4468[2],c2813,s4515[0]};
    assign in5812_2 = {s4479[1],s4469[2],s4465[3],s4516[0]};
    CLA_4 KS_5812(s5812, c5812, in5812_1, in5812_2);
    wire[3:0] s5813, in5813_1, in5813_2;
    wire c5813;
    assign in5813_1 = {s4480[1],s4470[2],s4466[3],s4517[0]};
    assign in5813_2 = {s4481[1],s4471[2],s4467[3],s4518[0]};
    CLA_4 KS_5813(s5813, c5813, in5813_1, in5813_2);
    wire[3:0] s5814, in5814_1, in5814_2;
    wire c5814;
    assign in5814_1 = {s4482[1],s4472[2],s4468[3],s4519[0]};
    assign in5814_2 = {s4483[1],s4473[2],s4469[3],s4520[0]};
    CLA_4 KS_5814(s5814, c5814, in5814_1, in5814_2);
    wire[3:0] s5815, in5815_1, in5815_2;
    wire c5815;
    assign in5815_1 = {c4484,s4474[2],s4470[3],s4521[0]};
    assign in5815_2 = {s4485[1],s4475[2],s4471[3],s4522[0]};
    CLA_4 KS_5815(s5815, c5815, in5815_1, in5815_2);
    wire[3:0] s5816, in5816_1, in5816_2;
    wire c5816;
    assign in5816_1 = {c4486,s4476[2],s4472[3],s4523[0]};
    assign in5816_2 = {s4487[1],s4477[2],s4473[3],s4524[0]};
    CLA_4 KS_5816(s5816, c5816, in5816_1, in5816_2);
    wire[3:0] s5817, in5817_1, in5817_2;
    wire c5817;
    assign in5817_1 = {c4488,s4478[2],s4474[3],s4525[0]};
    assign in5817_2 = {s4489[1],s4479[2],s4475[3],s4526[0]};
    CLA_4 KS_5817(s5817, c5817, in5817_1, in5817_2);
    wire[3:0] s5818, in5818_1, in5818_2;
    wire c5818;
    assign in5818_1 = {c4490,s4480[2],s4476[3],s4527[0]};
    assign in5818_2 = {s4491[1],s4481[2],s4477[3],s4528[0]};
    CLA_4 KS_5818(s5818, c5818, in5818_1, in5818_2);
    wire[3:0] s5819, in5819_1, in5819_2;
    wire c5819;
    assign in5819_1 = {c4492,s4482[2],s4478[3],s4529[0]};
    assign in5819_2 = {s4493[1],s4483[2],s4479[3],s4530[0]};
    CLA_4 KS_5819(s5819, c5819, in5819_1, in5819_2);
    wire[3:0] s5820, in5820_1, in5820_2;
    wire c5820;
    assign in5820_1 = {c4494,c4485,s4480[3],s4531[0]};
    assign in5820_2 = {s4495[1],s4487[2],s4481[3],s4532[0]};
    CLA_4 KS_5820(s5820, c5820, in5820_1, in5820_2);
    wire[3:0] s5821, in5821_1, in5821_2;
    wire c5821;
    assign in5821_1 = {c4496,c4489,s4482[3],s4533[0]};
    assign in5821_2 = {s4497[1],s4491[2],s4483[3],s4534[0]};
    CLA_4 KS_5821(s5821, c5821, in5821_1, in5821_2);
    wire[1:0] s5822, in5822_1, in5822_2;
    wire c5822;
    assign in5822_1 = {c4498,c4493};
    assign in5822_2 = {s4499[1],s4495[2]};
    CLA_2 KS_5822(s5822, c5822, in5822_1, in5822_2);
    wire[0:0] s5823, in5823_1, in5823_2;
    wire c5823;
    assign in5823_1 = {c4500};
    assign in5823_2 = {s4501[1]};
    Half_Adder KS_5823(s5823, c5823, in5823_1, in5823_2);
    wire[3:0] s5824, in5824_1, in5824_2;
    wire c5824;
    assign in5824_1 = {c5788,c4497,c4487,s4535[0]};
    assign in5824_2 = {c5789,s4499[2],s4491[3],s4536[0]};
    CLA_4 KS_5824(s5824, c5824, in5824_1, in5824_2);
    wire[0:0] s5825, in5825_1, in5825_2;
    wire c5825;
    assign in5825_1 = {c5790};
    assign in5825_2 = {c5791};
    Half_Adder KS_5825(s5825, c5825, in5825_1, in5825_2);
    wire[1:0] s5826, in5826_1, in5826_2;
    wire c5826;
    assign in5826_1 = {c5792,c4501};
    assign in5826_2 = {c5793,s5811[1]};
    CLA_2 KS_5826(s5826, c5826, in5826_1, in5826_2);
    wire[0:0] s5827, in5827_1, in5827_2;
    wire c5827;
    assign in5827_1 = {c5794};
    assign in5827_2 = {c5795};
    Half_Adder KS_5827(s5827, c5827, in5827_1, in5827_2);
    wire[2:0] s5828, in5828_1, in5828_2;
    wire c5828;
    assign in5828_1 = {c5796,s5812[1],c4495};
    assign in5828_2 = {c5797,s5813[1],s4499[3]};
    CLA_3 KS_5828(s5828, c5828, in5828_1, in5828_2);
    wire[0:0] s5829, in5829_1, in5829_2;
    wire c5829;
    assign in5829_1 = {c5798};
    assign in5829_2 = {c5799};
    Half_Adder KS_5829(s5829, c5829, in5829_1, in5829_2);
    wire[1:0] s5830, in5830_1, in5830_2;
    wire c5830;
    assign in5830_1 = {c5807,s5814[1]};
    assign in5830_2 = {s5811[0],s5815[1]};
    CLA_2 KS_5830(s5830, c5830, in5830_1, in5830_2);
    wire[0:0] s5831, in5831_1, in5831_2;
    wire c5831;
    assign in5831_1 = {s5812[0]};
    assign in5831_2 = {s5813[0]};
    Half_Adder KS_5831(s5831, c5831, in5831_1, in5831_2);
    wire[3:0] s5832, in5832_1, in5832_2;
    wire c5832;
    assign in5832_1 = {s5815[0],s5816[1],s5811[2],s4537[0]};
    assign in5832_2 = {s5816[0],s5817[1],s5812[2],s4538[0]};
    CLA_4_c KS_5832(s5832, c5832, in5832_1, in5832_2, s5814[0]);
    wire[3:0] s5833, in5833_1, in5833_2;
    wire c5833;
    assign in5833_1 = {s4513[1],s4503[2],c2872,s4549[0]};
    assign in5833_2 = {s4514[1],s4504[2],s2874[2],s4550[0]};
    CLA_4 KS_5833(s5833, c5833, in5833_1, in5833_2);
    wire[3:0] s5834, in5834_1, in5834_2;
    wire c5834;
    assign in5834_1 = {s4515[1],s4505[2],c2876,s4551[0]};
    assign in5834_2 = {s4516[1],s4506[2],s2878[2],s4552[0]};
    CLA_4 KS_5834(s5834, c5834, in5834_1, in5834_2);
    wire[3:0] s5835, in5835_1, in5835_2;
    wire c5835;
    assign in5835_1 = {s4517[1],s4507[2],s4502[3],s4553[0]};
    assign in5835_2 = {s4518[1],s4508[2],s4503[3],s4554[0]};
    CLA_4 KS_5835(s5835, c5835, in5835_1, in5835_2);
    wire[3:0] s5836, in5836_1, in5836_2;
    wire c5836;
    assign in5836_1 = {s4519[1],s4509[2],s4504[3],s4555[0]};
    assign in5836_2 = {s4520[1],s4510[2],s4505[3],s4556[0]};
    CLA_4 KS_5836(s5836, c5836, in5836_1, in5836_2);
    wire[3:0] s5837, in5837_1, in5837_2;
    wire c5837;
    assign in5837_1 = {c4521,s4511[2],s4506[3],s4557[0]};
    assign in5837_2 = {s4522[1],s4512[2],s4507[3],s4558[0]};
    CLA_4 KS_5837(s5837, c5837, in5837_1, in5837_2);
    wire[3:0] s5838, in5838_1, in5838_2;
    wire c5838;
    assign in5838_1 = {c4523,s4513[2],s4508[3],s4559[0]};
    assign in5838_2 = {s4524[1],s4514[2],s4509[3],s4560[0]};
    CLA_4 KS_5838(s5838, c5838, in5838_1, in5838_2);
    wire[3:0] s5839, in5839_1, in5839_2;
    wire c5839;
    assign in5839_1 = {c4525,s4515[2],s4510[3],s4561[0]};
    assign in5839_2 = {s4526[1],s4516[2],s4511[3],s4562[0]};
    CLA_4 KS_5839(s5839, c5839, in5839_1, in5839_2);
    wire[3:0] s5840, in5840_1, in5840_2;
    wire c5840;
    assign in5840_1 = {c4527,s4517[2],s4512[3],s4563[0]};
    assign in5840_2 = {s4528[1],s4518[2],s4513[3],s4564[0]};
    CLA_4 KS_5840(s5840, c5840, in5840_1, in5840_2);
    wire[3:0] s5841, in5841_1, in5841_2;
    wire c5841;
    assign in5841_1 = {c4529,s4519[2],s4514[3],s4565[0]};
    assign in5841_2 = {s4530[1],s4520[2],s4515[3],s4566[0]};
    CLA_4 KS_5841(s5841, c5841, in5841_1, in5841_2);
    wire[3:0] s5842, in5842_1, in5842_2;
    wire c5842;
    assign in5842_1 = {c4531,c4522,s4516[3],s4567[0]};
    assign in5842_2 = {s4532[1],s4524[2],s4517[3],s4568[0]};
    CLA_4 KS_5842(s5842, c5842, in5842_1, in5842_2);
    wire[3:0] s5843, in5843_1, in5843_2;
    wire c5843;
    assign in5843_1 = {c4533,c4526,s4518[3],s4569[0]};
    assign in5843_2 = {s4534[1],s4528[2],s4519[3],s4570[0]};
    CLA_4 KS_5843(s5843, c5843, in5843_1, in5843_2);
    wire[3:0] s5844, in5844_1, in5844_2;
    wire c5844;
    assign in5844_1 = {c4535,c4530,c4520,s4571[0]};
    assign in5844_2 = {s4536[1],s4532[2],s4524[3],s4572[0]};
    CLA_4 KS_5844(s5844, c5844, in5844_1, in5844_2);
    wire[0:0] s5845, in5845_1, in5845_2;
    wire c5845;
    assign in5845_1 = {c4537};
    assign in5845_2 = {s4538[1]};
    Half_Adder KS_5845(s5845, c5845, in5845_1, in5845_2);
    wire[1:0] s5846, in5846_1, in5846_2;
    wire c5846;
    assign in5846_1 = {c4539,c4534};
    assign in5846_2 = {c5811,s4536[2]};
    CLA_2 KS_5846(s5846, c5846, in5846_1, in5846_2);
    wire[0:0] s5847, in5847_1, in5847_2;
    wire c5847;
    assign in5847_1 = {c5812};
    assign in5847_2 = {c5813};
    Half_Adder KS_5847(s5847, c5847, in5847_1, in5847_2);
    wire[2:0] s5848, in5848_1, in5848_2;
    wire c5848;
    assign in5848_1 = {c5814,c4538,c4528};
    assign in5848_2 = {c5815,s5833[1],s4532[3]};
    CLA_3 KS_5848(s5848, c5848, in5848_1, in5848_2);
    wire[0:0] s5849, in5849_1, in5849_2;
    wire c5849;
    assign in5849_1 = {c5816};
    assign in5849_2 = {c5817};
    Half_Adder KS_5849(s5849, c5849, in5849_1, in5849_2);
    wire[1:0] s5850, in5850_1, in5850_2;
    wire c5850;
    assign in5850_1 = {c5818,s5834[1]};
    assign in5850_2 = {c5819,s5835[1]};
    CLA_2 KS_5850(s5850, c5850, in5850_1, in5850_2);
    wire[0:0] s5851, in5851_1, in5851_2;
    wire c5851;
    assign in5851_1 = {c5820};
    assign in5851_2 = {c5821};
    Half_Adder KS_5851(s5851, c5851, in5851_1, in5851_2);
    wire[3:0] s5852, in5852_1, in5852_2;
    wire c5852;
    assign in5852_1 = {c5824,s5836[1],c4536,s4573[0]};
    assign in5852_2 = {c5832,s5837[1],s5833[2],s4574[0]};
    CLA_4 KS_5852(s5852, c5852, in5852_1, in5852_2);
    wire[0:0] s5853, in5853_1, in5853_2;
    wire c5853;
    assign in5853_1 = {s5833[0]};
    assign in5853_2 = {s5834[0]};
    Half_Adder KS_5853(s5853, c5853, in5853_1, in5853_2);
    wire[1:0] s5854, in5854_1, in5854_2;
    wire c5854;
    assign in5854_1 = {s5835[0],s5838[1]};
    assign in5854_2 = {s5836[0],s5839[1]};
    CLA_2 KS_5854(s5854, c5854, in5854_1, in5854_2);
    wire[0:0] s5855, in5855_1, in5855_2;
    wire c5855;
    assign in5855_1 = {s5838[0]};
    assign in5855_2 = {s5839[0]};
    Full_Adder KS_5855(s5855, c5855, in5855_1, in5855_2, s5837[0]);
    wire[3:0] s5856, in5856_1, in5856_2;
    wire c5856;
    assign in5856_1 = {s4549[1],s4541[2],c2939,s4587[0]};
    assign in5856_2 = {s4550[1],s4542[2],s2941[2],s4588[0]};
    CLA_4 KS_5856(s5856, c5856, in5856_1, in5856_2);
    wire[3:0] s5857, in5857_1, in5857_2;
    wire c5857;
    assign in5857_1 = {s4551[1],s4543[2],c2943,s4589[0]};
    assign in5857_2 = {s4552[1],s4544[2],s4540[3],s4590[0]};
    CLA_4 KS_5857(s5857, c5857, in5857_1, in5857_2);
    wire[3:0] s5858, in5858_1, in5858_2;
    wire c5858;
    assign in5858_1 = {s4553[1],s4545[2],s4541[3],s4591[0]};
    assign in5858_2 = {s4554[1],s4546[2],s4542[3],s4592[0]};
    CLA_4 KS_5858(s5858, c5858, in5858_1, in5858_2);
    wire[3:0] s5859, in5859_1, in5859_2;
    wire c5859;
    assign in5859_1 = {s4555[1],s4547[2],s4543[3],s4593[0]};
    assign in5859_2 = {s4556[1],s4548[2],s4544[3],s4594[0]};
    CLA_4 KS_5859(s5859, c5859, in5859_1, in5859_2);
    wire[3:0] s5860, in5860_1, in5860_2;
    wire c5860;
    assign in5860_1 = {s4557[1],s4549[2],s4545[3],s4595[0]};
    assign in5860_2 = {s4558[1],s4550[2],s4546[3],s4596[0]};
    CLA_4 KS_5860(s5860, c5860, in5860_1, in5860_2);
    wire[3:0] s5861, in5861_1, in5861_2;
    wire c5861;
    assign in5861_1 = {c4559,s4551[2],s4547[3],s4597[0]};
    assign in5861_2 = {s4560[1],s4552[2],s4548[3],s4598[0]};
    CLA_4 KS_5861(s5861, c5861, in5861_1, in5861_2);
    wire[3:0] s5862, in5862_1, in5862_2;
    wire c5862;
    assign in5862_1 = {c4561,s4553[2],s4549[3],s4599[0]};
    assign in5862_2 = {s4562[1],s4554[2],s4550[3],s4600[0]};
    CLA_4 KS_5862(s5862, c5862, in5862_1, in5862_2);
    wire[3:0] s5863, in5863_1, in5863_2;
    wire c5863;
    assign in5863_1 = {c4563,s4555[2],s4551[3],s4601[0]};
    assign in5863_2 = {s4564[1],s4556[2],s4552[3],s4602[0]};
    CLA_4 KS_5863(s5863, c5863, in5863_1, in5863_2);
    wire[3:0] s5864, in5864_1, in5864_2;
    wire c5864;
    assign in5864_1 = {c4565,s4557[2],s4553[3],s4603[0]};
    assign in5864_2 = {s4566[1],s4558[2],s4554[3],s4604[0]};
    CLA_4 KS_5864(s5864, c5864, in5864_1, in5864_2);
    wire[3:0] s5865, in5865_1, in5865_2;
    wire c5865;
    assign in5865_1 = {c4567,c4560,s4555[3],s4605[0]};
    assign in5865_2 = {s4568[1],s4562[2],s4556[3],s4606[0]};
    CLA_4 KS_5865(s5865, c5865, in5865_1, in5865_2);
    wire[3:0] s5866, in5866_1, in5866_2;
    wire c5866;
    assign in5866_1 = {c4569,c4564,s4557[3],s4607[0]};
    assign in5866_2 = {s4570[1],s4566[2],s4558[3],s4608[0]};
    CLA_4 KS_5866(s5866, c5866, in5866_1, in5866_2);
    wire[0:0] s5867, in5867_1, in5867_2;
    wire c5867;
    assign in5867_1 = {c4571};
    assign in5867_2 = {s4572[1]};
    Half_Adder KS_5867(s5867, c5867, in5867_1, in5867_2);
    wire[1:0] s5868, in5868_1, in5868_2;
    wire c5868;
    assign in5868_1 = {c4573,c4568};
    assign in5868_2 = {s4574[1],s4570[2]};
    CLA_2 KS_5868(s5868, c5868, in5868_1, in5868_2);
    wire[0:0] s5869, in5869_1, in5869_2;
    wire c5869;
    assign in5869_1 = {c4575};
    assign in5869_2 = {c5833};
    Half_Adder KS_5869(s5869, c5869, in5869_1, in5869_2);
    wire[3:0] s5870, in5870_1, in5870_2;
    wire c5870;
    assign in5870_1 = {c5834,c4572,c4562,s4609[0]};
    assign in5870_2 = {c5835,s4574[2],s4566[3],s4610[0]};
    CLA_4 KS_5870(s5870, c5870, in5870_1, in5870_2);
    wire[0:0] s5871, in5871_1, in5871_2;
    wire c5871;
    assign in5871_1 = {c5836};
    assign in5871_2 = {c5837};
    Half_Adder KS_5871(s5871, c5871, in5871_1, in5871_2);
    wire[1:0] s5872, in5872_1, in5872_2;
    wire c5872;
    assign in5872_1 = {c5838,s5856[1]};
    assign in5872_2 = {c5839,s5857[1]};
    CLA_2 KS_5872(s5872, c5872, in5872_1, in5872_2);
    wire[0:0] s5873, in5873_1, in5873_2;
    wire c5873;
    assign in5873_1 = {c5840};
    assign in5873_2 = {c5841};
    Half_Adder KS_5873(s5873, c5873, in5873_1, in5873_2);
    wire[2:0] s5874, in5874_1, in5874_2;
    wire c5874;
    assign in5874_1 = {c5842,s5858[1],c4570};
    assign in5874_2 = {c5843,s5859[1],s4574[3]};
    CLA_3 KS_5874(s5874, c5874, in5874_1, in5874_2);
    wire[0:0] s5875, in5875_1, in5875_2;
    wire c5875;
    assign in5875_1 = {c5844};
    assign in5875_2 = {c5852};
    Half_Adder KS_5875(s5875, c5875, in5875_1, in5875_2);
    wire[1:0] s5876, in5876_1, in5876_2;
    wire c5876;
    assign in5876_1 = {s5856[0],s5860[1]};
    assign in5876_2 = {s5857[0],s5861[1]};
    CLA_2 KS_5876(s5876, c5876, in5876_1, in5876_2);
    wire[0:0] s5877, in5877_1, in5877_2;
    wire c5877;
    assign in5877_1 = {s5858[0]};
    assign in5877_2 = {s5859[0]};
    Half_Adder KS_5877(s5877, c5877, in5877_1, in5877_2);
    wire[3:0] s5878, in5878_1, in5878_2;
    wire c5878;
    assign in5878_1 = {s5861[0],s5862[1],s5856[2],s4611[0]};
    assign in5878_2 = {s5862[0],s5863[1],s5857[2],s4612[0]};
    CLA_4_c KS_5878(s5878, c5878, in5878_1, in5878_2, s5860[0]);
    wire[3:0] s5879, in5879_1, in5879_2;
    wire c5879;
    assign in5879_1 = {s4587[1],s4578[2],c3002,s4623[0]};
    assign in5879_2 = {s4588[1],s4579[2],s3004[2],s4624[0]};
    CLA_4 KS_5879(s5879, c5879, in5879_1, in5879_2);
    wire[3:0] s5880, in5880_1, in5880_2;
    wire c5880;
    assign in5880_1 = {s4589[1],s4580[2],c3006,s4625[0]};
    assign in5880_2 = {s4590[1],s4581[2],s3008[2],s4626[0]};
    CLA_4 KS_5880(s5880, c5880, in5880_1, in5880_2);
    wire[3:0] s5881, in5881_1, in5881_2;
    wire c5881;
    assign in5881_1 = {s4591[1],s4582[2],s4576[3],s4627[0]};
    assign in5881_2 = {s4592[1],s4583[2],s4577[3],s4628[0]};
    CLA_4 KS_5881(s5881, c5881, in5881_1, in5881_2);
    wire[3:0] s5882, in5882_1, in5882_2;
    wire c5882;
    assign in5882_1 = {s4593[1],s4584[2],s4578[3],s4629[0]};
    assign in5882_2 = {s4594[1],s4585[2],s4579[3],s4630[0]};
    CLA_4 KS_5882(s5882, c5882, in5882_1, in5882_2);
    wire[3:0] s5883, in5883_1, in5883_2;
    wire c5883;
    assign in5883_1 = {c4595,s4586[2],s4580[3],s4631[0]};
    assign in5883_2 = {s4596[1],s4587[2],s4581[3],s4632[0]};
    CLA_4 KS_5883(s5883, c5883, in5883_1, in5883_2);
    wire[3:0] s5884, in5884_1, in5884_2;
    wire c5884;
    assign in5884_1 = {c4597,s4588[2],s4582[3],s4633[0]};
    assign in5884_2 = {s4598[1],s4589[2],s4583[3],s4634[0]};
    CLA_4 KS_5884(s5884, c5884, in5884_1, in5884_2);
    wire[3:0] s5885, in5885_1, in5885_2;
    wire c5885;
    assign in5885_1 = {c4599,s4590[2],s4584[3],s4635[0]};
    assign in5885_2 = {s4600[1],s4591[2],s4585[3],s4636[0]};
    CLA_4 KS_5885(s5885, c5885, in5885_1, in5885_2);
    wire[3:0] s5886, in5886_1, in5886_2;
    wire c5886;
    assign in5886_1 = {c4601,s4592[2],s4586[3],s4637[0]};
    assign in5886_2 = {s4602[1],s4593[2],s4587[3],s4638[0]};
    CLA_4 KS_5886(s5886, c5886, in5886_1, in5886_2);
    wire[3:0] s5887, in5887_1, in5887_2;
    wire c5887;
    assign in5887_1 = {c4603,c4594,s4588[3],s4639[0]};
    assign in5887_2 = {s4604[1],s4596[2],s4589[3],s4640[0]};
    CLA_4 KS_5887(s5887, c5887, in5887_1, in5887_2);
    wire[3:0] s5888, in5888_1, in5888_2;
    wire c5888;
    assign in5888_1 = {c4605,c4598,s4590[3],s4641[0]};
    assign in5888_2 = {s4606[1],s4600[2],s4591[3],s4642[0]};
    CLA_4 KS_5888(s5888, c5888, in5888_1, in5888_2);
    wire[3:0] s5889, in5889_1, in5889_2;
    wire c5889;
    assign in5889_1 = {c4607,c4602,s4592[3],s4643[0]};
    assign in5889_2 = {s4608[1],s4604[2],s4593[3],s4644[0]};
    CLA_4 KS_5889(s5889, c5889, in5889_1, in5889_2);
    wire[0:0] s5890, in5890_1, in5890_2;
    wire c5890;
    assign in5890_1 = {c4609};
    assign in5890_2 = {s4610[1]};
    Half_Adder KS_5890(s5890, c5890, in5890_1, in5890_2);
    wire[3:0] s5891, in5891_1, in5891_2;
    wire c5891;
    assign in5891_1 = {c4611,c4606,c4596,s4645[0]};
    assign in5891_2 = {s4612[1],s4608[2],s4600[3],s4646[0]};
    CLA_4 KS_5891(s5891, c5891, in5891_1, in5891_2);
    wire[0:0] s5892, in5892_1, in5892_2;
    wire c5892;
    assign in5892_1 = {c4613};
    assign in5892_2 = {c5856};
    Half_Adder KS_5892(s5892, c5892, in5892_1, in5892_2);
    wire[1:0] s5893, in5893_1, in5893_2;
    wire c5893;
    assign in5893_1 = {c5857,c4610};
    assign in5893_2 = {c5858,s4612[2]};
    CLA_2 KS_5893(s5893, c5893, in5893_1, in5893_2);
    wire[0:0] s5894, in5894_1, in5894_2;
    wire c5894;
    assign in5894_1 = {c5859};
    assign in5894_2 = {c5860};
    Half_Adder KS_5894(s5894, c5894, in5894_1, in5894_2);
    wire[2:0] s5895, in5895_1, in5895_2;
    wire c5895;
    assign in5895_1 = {c5861,s5879[1],c4604};
    assign in5895_2 = {c5862,s5880[1],s4608[3]};
    CLA_3 KS_5895(s5895, c5895, in5895_1, in5895_2);
    wire[0:0] s5896, in5896_1, in5896_2;
    wire c5896;
    assign in5896_1 = {c5863};
    assign in5896_2 = {c5864};
    Half_Adder KS_5896(s5896, c5896, in5896_1, in5896_2);
    wire[1:0] s5897, in5897_1, in5897_2;
    wire c5897;
    assign in5897_1 = {c5865,s5881[1]};
    assign in5897_2 = {c5866,s5882[1]};
    CLA_2 KS_5897(s5897, c5897, in5897_1, in5897_2);
    wire[0:0] s5898, in5898_1, in5898_2;
    wire c5898;
    assign in5898_1 = {c5870};
    assign in5898_2 = {c5878};
    Half_Adder KS_5898(s5898, c5898, in5898_1, in5898_2);
    wire[3:0] s5899, in5899_1, in5899_2;
    wire c5899;
    assign in5899_1 = {s5879[0],s5883[1],c4612,s4647[0]};
    assign in5899_2 = {s5880[0],s5884[1],s5879[2],s4648[0]};
    CLA_4 KS_5899(s5899, c5899, in5899_1, in5899_2);
    wire[0:0] s5900, in5900_1, in5900_2;
    wire c5900;
    assign in5900_1 = {s5881[0]};
    assign in5900_2 = {s5882[0]};
    Half_Adder KS_5900(s5900, c5900, in5900_1, in5900_2);
    wire[1:0] s5901, in5901_1, in5901_2;
    wire c5901;
    assign in5901_1 = {s5884[0],s5885[1]};
    assign in5901_2 = {s5885[0],s5886[1]};
    CLA_2_c KS_5901(s5901, c5901, in5901_1, in5901_2, s5883[0]);
    wire[3:0] s5902, in5902_1, in5902_2;
    wire c5902;
    assign in5902_1 = {s4623[1],s4615[2],c3069,s4661[0]};
    assign in5902_2 = {s4624[1],s4616[2],s3071[2],s4662[0]};
    CLA_4 KS_5902(s5902, c5902, in5902_1, in5902_2);
    wire[3:0] s5903, in5903_1, in5903_2;
    wire c5903;
    assign in5903_1 = {s4625[1],s4617[2],c3073,s4663[0]};
    assign in5903_2 = {s4626[1],s4618[2],s4614[3],s4664[0]};
    CLA_4 KS_5903(s5903, c5903, in5903_1, in5903_2);
    wire[3:0] s5904, in5904_1, in5904_2;
    wire c5904;
    assign in5904_1 = {s4627[1],s4619[2],s4615[3],s4665[0]};
    assign in5904_2 = {s4628[1],s4620[2],s4616[3],s4666[0]};
    CLA_4 KS_5904(s5904, c5904, in5904_1, in5904_2);
    wire[3:0] s5905, in5905_1, in5905_2;
    wire c5905;
    assign in5905_1 = {s4629[1],s4621[2],s4617[3],s4667[0]};
    assign in5905_2 = {s4630[1],s4622[2],s4618[3],s4668[0]};
    CLA_4 KS_5905(s5905, c5905, in5905_1, in5905_2);
    wire[3:0] s5906, in5906_1, in5906_2;
    wire c5906;
    assign in5906_1 = {s4631[1],s4623[2],s4619[3],s4669[0]};
    assign in5906_2 = {s4632[1],s4624[2],s4620[3],s4670[0]};
    CLA_4 KS_5906(s5906, c5906, in5906_1, in5906_2);
    wire[3:0] s5907, in5907_1, in5907_2;
    wire c5907;
    assign in5907_1 = {c4633,s4625[2],s4621[3],s4671[0]};
    assign in5907_2 = {s4634[1],s4626[2],s4622[3],s4672[0]};
    CLA_4 KS_5907(s5907, c5907, in5907_1, in5907_2);
    wire[3:0] s5908, in5908_1, in5908_2;
    wire c5908;
    assign in5908_1 = {c4635,s4627[2],s4623[3],s4673[0]};
    assign in5908_2 = {s4636[1],s4628[2],s4624[3],s4674[0]};
    CLA_4 KS_5908(s5908, c5908, in5908_1, in5908_2);
    wire[3:0] s5909, in5909_1, in5909_2;
    wire c5909;
    assign in5909_1 = {c4637,s4629[2],s4625[3],s4675[0]};
    assign in5909_2 = {s4638[1],s4630[2],s4626[3],s4676[0]};
    CLA_4 KS_5909(s5909, c5909, in5909_1, in5909_2);
    wire[3:0] s5910, in5910_1, in5910_2;
    wire c5910;
    assign in5910_1 = {c4639,s4631[2],s4627[3],s4677[0]};
    assign in5910_2 = {s4640[1],s4632[2],s4628[3],s4678[0]};
    CLA_4 KS_5910(s5910, c5910, in5910_1, in5910_2);
    wire[3:0] s5911, in5911_1, in5911_2;
    wire c5911;
    assign in5911_1 = {c4641,c4634,s4629[3],s4679[0]};
    assign in5911_2 = {s4642[1],s4636[2],s4630[3],s4680[0]};
    CLA_4 KS_5911(s5911, c5911, in5911_1, in5911_2);
    wire[3:0] s5912, in5912_1, in5912_2;
    wire c5912;
    assign in5912_1 = {c4643,c4638,s4631[3],s4681[0]};
    assign in5912_2 = {s4644[1],s4640[2],s4632[3],s4682[0]};
    CLA_4 KS_5912(s5912, c5912, in5912_1, in5912_2);
    wire[0:0] s5913, in5913_1, in5913_2;
    wire c5913;
    assign in5913_1 = {c4645};
    assign in5913_2 = {s4646[1]};
    Half_Adder KS_5913(s5913, c5913, in5913_1, in5913_2);
    wire[1:0] s5914, in5914_1, in5914_2;
    wire c5914;
    assign in5914_1 = {c4647,c4642};
    assign in5914_2 = {s4648[1],s4644[2]};
    CLA_2 KS_5914(s5914, c5914, in5914_1, in5914_2);
    wire[0:0] s5915, in5915_1, in5915_2;
    wire c5915;
    assign in5915_1 = {c4649};
    assign in5915_2 = {c5879};
    Half_Adder KS_5915(s5915, c5915, in5915_1, in5915_2);
    wire[3:0] s5916, in5916_1, in5916_2;
    wire c5916;
    assign in5916_1 = {c5880,c4646,c4636,s4683[0]};
    assign in5916_2 = {c5881,s4648[2],s4640[3],s4684[0]};
    CLA_4 KS_5916(s5916, c5916, in5916_1, in5916_2);
    wire[0:0] s5917, in5917_1, in5917_2;
    wire c5917;
    assign in5917_1 = {c5882};
    assign in5917_2 = {c5883};
    Half_Adder KS_5917(s5917, c5917, in5917_1, in5917_2);
    wire[1:0] s5918, in5918_1, in5918_2;
    wire c5918;
    assign in5918_1 = {c5884,s5902[1]};
    assign in5918_2 = {c5885,s5903[1]};
    CLA_2 KS_5918(s5918, c5918, in5918_1, in5918_2);
    wire[0:0] s5919, in5919_1, in5919_2;
    wire c5919;
    assign in5919_1 = {c5886};
    assign in5919_2 = {c5887};
    Half_Adder KS_5919(s5919, c5919, in5919_1, in5919_2);
    wire[2:0] s5920, in5920_1, in5920_2;
    wire c5920;
    assign in5920_1 = {c5888,s5904[1],c4644};
    assign in5920_2 = {c5889,s5905[1],s4648[3]};
    CLA_3 KS_5920(s5920, c5920, in5920_1, in5920_2);
    wire[0:0] s5921, in5921_1, in5921_2;
    wire c5921;
    assign in5921_1 = {c5891};
    assign in5921_2 = {c5899};
    Half_Adder KS_5921(s5921, c5921, in5921_1, in5921_2);
    wire[1:0] s5922, in5922_1, in5922_2;
    wire c5922;
    assign in5922_1 = {s5902[0],s5906[1]};
    assign in5922_2 = {s5903[0],s5907[1]};
    CLA_2 KS_5922(s5922, c5922, in5922_1, in5922_2);
    wire[0:0] s5923, in5923_1, in5923_2;
    wire c5923;
    assign in5923_1 = {s5904[0]};
    assign in5923_2 = {s5905[0]};
    Half_Adder KS_5923(s5923, c5923, in5923_1, in5923_2);
    wire[3:0] s5924, in5924_1, in5924_2;
    wire c5924;
    assign in5924_1 = {s5907[0],s5908[1],s5902[2],s4685[0]};
    assign in5924_2 = {s5908[0],s5909[1],s5903[2],s4686[0]};
    CLA_4_c KS_5924(s5924, c5924, in5924_1, in5924_2, s5906[0]);
    wire[3:0] s5925, in5925_1, in5925_2;
    wire c5925;
    assign in5925_1 = {s4661[1],s4652[2],c3133,s4697[0]};
    assign in5925_2 = {s4662[1],s4653[2],s3135[2],s4698[0]};
    CLA_4 KS_5925(s5925, c5925, in5925_1, in5925_2);
    wire[3:0] s5926, in5926_1, in5926_2;
    wire c5926;
    assign in5926_1 = {s4663[1],s4654[2],c3137,s4699[0]};
    assign in5926_2 = {s4664[1],s4655[2],s3139[2],s4700[0]};
    CLA_4 KS_5926(s5926, c5926, in5926_1, in5926_2);
    wire[3:0] s5927, in5927_1, in5927_2;
    wire c5927;
    assign in5927_1 = {s4665[1],s4656[2],s4650[3],s4701[0]};
    assign in5927_2 = {s4666[1],s4657[2],s4651[3],s4702[0]};
    CLA_4 KS_5927(s5927, c5927, in5927_1, in5927_2);
    wire[3:0] s5928, in5928_1, in5928_2;
    wire c5928;
    assign in5928_1 = {s4667[1],s4658[2],s4652[3],s4703[0]};
    assign in5928_2 = {s4668[1],s4659[2],s4653[3],s4704[0]};
    CLA_4 KS_5928(s5928, c5928, in5928_1, in5928_2);
    wire[3:0] s5929, in5929_1, in5929_2;
    wire c5929;
    assign in5929_1 = {c4669,s4660[2],s4654[3],s4705[0]};
    assign in5929_2 = {s4670[1],s4661[2],s4655[3],s4706[0]};
    CLA_4 KS_5929(s5929, c5929, in5929_1, in5929_2);
    wire[3:0] s5930, in5930_1, in5930_2;
    wire c5930;
    assign in5930_1 = {c4671,s4662[2],s4656[3],s4707[0]};
    assign in5930_2 = {s4672[1],s4663[2],s4657[3],s4708[0]};
    CLA_4 KS_5930(s5930, c5930, in5930_1, in5930_2);
    wire[3:0] s5931, in5931_1, in5931_2;
    wire c5931;
    assign in5931_1 = {c4673,s4664[2],s4658[3],s4709[0]};
    assign in5931_2 = {s4674[1],s4665[2],s4659[3],s4710[0]};
    CLA_4 KS_5931(s5931, c5931, in5931_1, in5931_2);
    wire[3:0] s5932, in5932_1, in5932_2;
    wire c5932;
    assign in5932_1 = {c4675,s4666[2],s4660[3],s4711[0]};
    assign in5932_2 = {s4676[1],s4667[2],s4661[3],s4712[0]};
    CLA_4 KS_5932(s5932, c5932, in5932_1, in5932_2);
    wire[3:0] s5933, in5933_1, in5933_2;
    wire c5933;
    assign in5933_1 = {c4677,c4668,s4662[3],s4713[0]};
    assign in5933_2 = {s4678[1],s4670[2],s4663[3],s4714[0]};
    CLA_4 KS_5933(s5933, c5933, in5933_1, in5933_2);
    wire[3:0] s5934, in5934_1, in5934_2;
    wire c5934;
    assign in5934_1 = {c4679,c4672,s4664[3],s4715[0]};
    assign in5934_2 = {s4680[1],s4674[2],s4665[3],s4716[0]};
    CLA_4 KS_5934(s5934, c5934, in5934_1, in5934_2);
    wire[3:0] s5935, in5935_1, in5935_2;
    wire c5935;
    assign in5935_1 = {c4681,c4676,s4666[3],s4717[0]};
    assign in5935_2 = {s4682[1],s4678[2],s4667[3],s4718[0]};
    CLA_4 KS_5935(s5935, c5935, in5935_1, in5935_2);
    wire[0:0] s5936, in5936_1, in5936_2;
    wire c5936;
    assign in5936_1 = {c4683};
    assign in5936_2 = {s4684[1]};
    Half_Adder KS_5936(s5936, c5936, in5936_1, in5936_2);
    wire[3:0] s5937, in5937_1, in5937_2;
    wire c5937;
    assign in5937_1 = {c4685,c4680,c4670,s4719[0]};
    assign in5937_2 = {s4686[1],s4682[2],s4674[3],s4720[0]};
    CLA_4 KS_5937(s5937, c5937, in5937_1, in5937_2);
    wire[0:0] s5938, in5938_1, in5938_2;
    wire c5938;
    assign in5938_1 = {c4687};
    assign in5938_2 = {c5902};
    Half_Adder KS_5938(s5938, c5938, in5938_1, in5938_2);
    wire[1:0] s5939, in5939_1, in5939_2;
    wire c5939;
    assign in5939_1 = {c5903,c4684};
    assign in5939_2 = {c5904,s4686[2]};
    CLA_2 KS_5939(s5939, c5939, in5939_1, in5939_2);
    wire[0:0] s5940, in5940_1, in5940_2;
    wire c5940;
    assign in5940_1 = {c5905};
    assign in5940_2 = {c5906};
    Half_Adder KS_5940(s5940, c5940, in5940_1, in5940_2);
    wire[2:0] s5941, in5941_1, in5941_2;
    wire c5941;
    assign in5941_1 = {c5907,s5925[1],c4678};
    assign in5941_2 = {c5908,s5926[1],s4682[3]};
    CLA_3 KS_5941(s5941, c5941, in5941_1, in5941_2);
    wire[0:0] s5942, in5942_1, in5942_2;
    wire c5942;
    assign in5942_1 = {c5909};
    assign in5942_2 = {c5910};
    Half_Adder KS_5942(s5942, c5942, in5942_1, in5942_2);
    wire[1:0] s5943, in5943_1, in5943_2;
    wire c5943;
    assign in5943_1 = {c5911,s5927[1]};
    assign in5943_2 = {c5912,s5928[1]};
    CLA_2 KS_5943(s5943, c5943, in5943_1, in5943_2);
    wire[0:0] s5944, in5944_1, in5944_2;
    wire c5944;
    assign in5944_1 = {c5916};
    assign in5944_2 = {c5924};
    Half_Adder KS_5944(s5944, c5944, in5944_1, in5944_2);
    wire[3:0] s5945, in5945_1, in5945_2;
    wire c5945;
    assign in5945_1 = {s5925[0],s5929[1],c4686,s4721[0]};
    assign in5945_2 = {s5926[0],s5930[1],s5925[2],s4722[0]};
    CLA_4 KS_5945(s5945, c5945, in5945_1, in5945_2);
    wire[0:0] s5946, in5946_1, in5946_2;
    wire c5946;
    assign in5946_1 = {s5927[0]};
    assign in5946_2 = {s5928[0]};
    Half_Adder KS_5946(s5946, c5946, in5946_1, in5946_2);
    wire[1:0] s5947, in5947_1, in5947_2;
    wire c5947;
    assign in5947_1 = {s5930[0],s5931[1]};
    assign in5947_2 = {s5931[0],s5932[1]};
    CLA_2_c KS_5947(s5947, c5947, in5947_1, in5947_2, s5929[0]);
    wire[3:0] s5948, in5948_1, in5948_2;
    wire c5948;
    assign in5948_1 = {s4697[1],s4688[2],c3196,s4733[0]};
    assign in5948_2 = {s4698[1],s4689[2],s3198[2],s4734[0]};
    CLA_4 KS_5948(s5948, c5948, in5948_1, in5948_2);
    wire[3:0] s5949, in5949_1, in5949_2;
    wire c5949;
    assign in5949_1 = {s4699[1],s4690[2],c3200,s4735[0]};
    assign in5949_2 = {s4700[1],s4691[2],s3202[2],s4736[0]};
    CLA_4 KS_5949(s5949, c5949, in5949_1, in5949_2);
    wire[3:0] s5950, in5950_1, in5950_2;
    wire c5950;
    assign in5950_1 = {s4701[1],s4692[2],c3204,s4737[0]};
    assign in5950_2 = {s4702[1],s4693[2],s4688[3],s4738[0]};
    CLA_4 KS_5950(s5950, c5950, in5950_1, in5950_2);
    wire[3:0] s5951, in5951_1, in5951_2;
    wire c5951;
    assign in5951_1 = {s4703[1],s4694[2],s4689[3],s4739[0]};
    assign in5951_2 = {s4704[1],s4695[2],s4690[3],s4740[0]};
    CLA_4 KS_5951(s5951, c5951, in5951_1, in5951_2);
    wire[3:0] s5952, in5952_1, in5952_2;
    wire c5952;
    assign in5952_1 = {s4705[1],s4696[2],s4691[3],s4741[0]};
    assign in5952_2 = {s4706[1],s4697[2],s4692[3],s4742[0]};
    CLA_4 KS_5952(s5952, c5952, in5952_1, in5952_2);
    wire[3:0] s5953, in5953_1, in5953_2;
    wire c5953;
    assign in5953_1 = {c4707,s4698[2],s4693[3],s4743[0]};
    assign in5953_2 = {s4708[1],s4699[2],s4694[3],s4744[0]};
    CLA_4 KS_5953(s5953, c5953, in5953_1, in5953_2);
    wire[3:0] s5954, in5954_1, in5954_2;
    wire c5954;
    assign in5954_1 = {c4709,s4700[2],s4695[3],s4745[0]};
    assign in5954_2 = {s4710[1],s4701[2],s4696[3],s4746[0]};
    CLA_4 KS_5954(s5954, c5954, in5954_1, in5954_2);
    wire[3:0] s5955, in5955_1, in5955_2;
    wire c5955;
    assign in5955_1 = {c4711,s4702[2],s4697[3],s4747[0]};
    assign in5955_2 = {s4712[1],s4703[2],s4698[3],s4748[0]};
    CLA_4 KS_5955(s5955, c5955, in5955_1, in5955_2);
    wire[3:0] s5956, in5956_1, in5956_2;
    wire c5956;
    assign in5956_1 = {c4713,s4704[2],s4699[3],s4749[0]};
    assign in5956_2 = {s4714[1],s4705[2],s4700[3],s4750[0]};
    CLA_4 KS_5956(s5956, c5956, in5956_1, in5956_2);
    wire[3:0] s5957, in5957_1, in5957_2;
    wire c5957;
    assign in5957_1 = {c4715,c4706,s4701[3],s4751[0]};
    assign in5957_2 = {s4716[1],s4708[2],s4702[3],s4752[0]};
    CLA_4 KS_5957(s5957, c5957, in5957_1, in5957_2);
    wire[3:0] s5958, in5958_1, in5958_2;
    wire c5958;
    assign in5958_1 = {c4717,c4710,s4703[3],s4753[0]};
    assign in5958_2 = {s4718[1],s4712[2],s4704[3],s4754[0]};
    CLA_4 KS_5958(s5958, c5958, in5958_1, in5958_2);
    wire[3:0] s5959, in5959_1, in5959_2;
    wire c5959;
    assign in5959_1 = {c4719,c4714,s4705[3],s4755[0]};
    assign in5959_2 = {s4720[1],s4716[2],s4708[3],s4756[0]};
    CLA_4 KS_5959(s5959, c5959, in5959_1, in5959_2);
    wire[0:0] s5960, in5960_1, in5960_2;
    wire c5960;
    assign in5960_1 = {c4721};
    assign in5960_2 = {s4722[1]};
    Half_Adder KS_5960(s5960, c5960, in5960_1, in5960_2);
    wire[1:0] s5961, in5961_1, in5961_2;
    wire c5961;
    assign in5961_1 = {c4723,c4718};
    assign in5961_2 = {c5925,s4720[2]};
    CLA_2 KS_5961(s5961, c5961, in5961_1, in5961_2);
    wire[0:0] s5962, in5962_1, in5962_2;
    wire c5962;
    assign in5962_1 = {c5926};
    assign in5962_2 = {c5927};
    Half_Adder KS_5962(s5962, c5962, in5962_1, in5962_2);
    wire[2:0] s5963, in5963_1, in5963_2;
    wire c5963;
    assign in5963_1 = {c5928,c4722,c4712};
    assign in5963_2 = {c5929,s5948[1],s4716[3]};
    CLA_3 KS_5963(s5963, c5963, in5963_1, in5963_2);
    wire[0:0] s5964, in5964_1, in5964_2;
    wire c5964;
    assign in5964_1 = {c5930};
    assign in5964_2 = {c5931};
    Half_Adder KS_5964(s5964, c5964, in5964_1, in5964_2);
    wire[1:0] s5965, in5965_1, in5965_2;
    wire c5965;
    assign in5965_1 = {c5932,s5949[1]};
    assign in5965_2 = {c5933,s5950[1]};
    CLA_2 KS_5965(s5965, c5965, in5965_1, in5965_2);
    wire[0:0] s5966, in5966_1, in5966_2;
    wire c5966;
    assign in5966_1 = {c5934};
    assign in5966_2 = {c5935};
    Half_Adder KS_5966(s5966, c5966, in5966_1, in5966_2);
    wire[3:0] s5967, in5967_1, in5967_2;
    wire c5967;
    assign in5967_1 = {c5937,s5951[1],c4720,s4757[0]};
    assign in5967_2 = {c5945,s5952[1],s5948[2],s4758[0]};
    CLA_4 KS_5967(s5967, c5967, in5967_1, in5967_2);
    wire[0:0] s5968, in5968_1, in5968_2;
    wire c5968;
    assign in5968_1 = {s5948[0]};
    assign in5968_2 = {s5949[0]};
    Half_Adder KS_5968(s5968, c5968, in5968_1, in5968_2);
    wire[1:0] s5969, in5969_1, in5969_2;
    wire c5969;
    assign in5969_1 = {s5950[0],s5953[1]};
    assign in5969_2 = {s5951[0],s5954[1]};
    CLA_2 KS_5969(s5969, c5969, in5969_1, in5969_2);
    wire[0:0] s5970, in5970_1, in5970_2;
    wire c5970;
    assign in5970_1 = {s5953[0]};
    assign in5970_2 = {s5954[0]};
    Full_Adder KS_5970(s5970, c5970, in5970_1, in5970_2, s5952[0]);
    wire[3:0] s5971, in5971_1, in5971_2;
    wire c5971;
    assign in5971_1 = {s4733[1],s4724[2],c3254,s4770[0]};
    assign in5971_2 = {s4734[1],s4725[2],s3256[2],s4771[0]};
    CLA_4 KS_5971(s5971, c5971, in5971_1, in5971_2);
    wire[3:0] s5972, in5972_1, in5972_2;
    wire c5972;
    assign in5972_1 = {s4735[1],s4726[2],c3258,s4772[0]};
    assign in5972_2 = {s4736[1],s4727[2],s3260[2],s4773[0]};
    CLA_4 KS_5972(s5972, c5972, in5972_1, in5972_2);
    wire[3:0] s5973, in5973_1, in5973_2;
    wire c5973;
    assign in5973_1 = {s4737[1],s4728[2],c3262,s4774[0]};
    assign in5973_2 = {s4738[1],s4729[2],s4724[3],s4775[0]};
    CLA_4 KS_5973(s5973, c5973, in5973_1, in5973_2);
    wire[3:0] s5974, in5974_1, in5974_2;
    wire c5974;
    assign in5974_1 = {s4739[1],s4730[2],s4725[3],s4776[0]};
    assign in5974_2 = {s4740[1],s4731[2],s4726[3],s4777[0]};
    CLA_4 KS_5974(s5974, c5974, in5974_1, in5974_2);
    wire[3:0] s5975, in5975_1, in5975_2;
    wire c5975;
    assign in5975_1 = {s4741[1],s4732[2],s4727[3],s4778[0]};
    assign in5975_2 = {s4742[1],s4733[2],s4728[3],s4779[0]};
    CLA_4 KS_5975(s5975, c5975, in5975_1, in5975_2);
    wire[3:0] s5976, in5976_1, in5976_2;
    wire c5976;
    assign in5976_1 = {c4743,s4734[2],s4729[3],s4780[0]};
    assign in5976_2 = {s4744[1],s4735[2],s4730[3],s4781[0]};
    CLA_4 KS_5976(s5976, c5976, in5976_1, in5976_2);
    wire[3:0] s5977, in5977_1, in5977_2;
    wire c5977;
    assign in5977_1 = {c4745,s4736[2],s4731[3],s4782[0]};
    assign in5977_2 = {s4746[1],s4737[2],s4732[3],s4783[0]};
    CLA_4 KS_5977(s5977, c5977, in5977_1, in5977_2);
    wire[3:0] s5978, in5978_1, in5978_2;
    wire c5978;
    assign in5978_1 = {c4747,s4738[2],s4733[3],s4784[0]};
    assign in5978_2 = {s4748[1],s4739[2],s4734[3],s4785[0]};
    CLA_4 KS_5978(s5978, c5978, in5978_1, in5978_2);
    wire[3:0] s5979, in5979_1, in5979_2;
    wire c5979;
    assign in5979_1 = {c4749,s4740[2],s4735[3],s4786[0]};
    assign in5979_2 = {s4750[1],s4741[2],s4736[3],s4787[0]};
    CLA_4 KS_5979(s5979, c5979, in5979_1, in5979_2);
    wire[3:0] s5980, in5980_1, in5980_2;
    wire c5980;
    assign in5980_1 = {c4751,c4742,s4737[3],s4788[0]};
    assign in5980_2 = {s4752[1],s4744[2],s4738[3],s4789[0]};
    CLA_4 KS_5980(s5980, c5980, in5980_1, in5980_2);
    wire[3:0] s5981, in5981_1, in5981_2;
    wire c5981;
    assign in5981_1 = {c4753,c4746,s4739[3],s4790[0]};
    assign in5981_2 = {s4754[1],s4748[2],s4740[3],s4791[0]};
    CLA_4 KS_5981(s5981, c5981, in5981_1, in5981_2);
    wire[3:0] s5982, in5982_1, in5982_2;
    wire c5982;
    assign in5982_1 = {c4755,c4750,s4741[3],s4792[0]};
    assign in5982_2 = {s4756[1],s4752[2],s4744[3],s4793[0]};
    CLA_4 KS_5982(s5982, c5982, in5982_1, in5982_2);
    wire[0:0] s5983, in5983_1, in5983_2;
    wire c5983;
    assign in5983_1 = {c4757};
    assign in5983_2 = {s4758[1]};
    Half_Adder KS_5983(s5983, c5983, in5983_1, in5983_2);
    wire[1:0] s5984, in5984_1, in5984_2;
    wire c5984;
    assign in5984_1 = {c4759,c4754};
    assign in5984_2 = {c5948,s4756[2]};
    CLA_2 KS_5984(s5984, c5984, in5984_1, in5984_2);
    wire[0:0] s5985, in5985_1, in5985_2;
    wire c5985;
    assign in5985_1 = {c5949};
    assign in5985_2 = {c5950};
    Half_Adder KS_5985(s5985, c5985, in5985_1, in5985_2);
    wire[2:0] s5986, in5986_1, in5986_2;
    wire c5986;
    assign in5986_1 = {c5951,c4758,c4748};
    assign in5986_2 = {c5952,s5971[1],s4752[3]};
    CLA_3 KS_5986(s5986, c5986, in5986_1, in5986_2);
    wire[0:0] s5987, in5987_1, in5987_2;
    wire c5987;
    assign in5987_1 = {c5953};
    assign in5987_2 = {c5954};
    Half_Adder KS_5987(s5987, c5987, in5987_1, in5987_2);
    wire[1:0] s5988, in5988_1, in5988_2;
    wire c5988;
    assign in5988_1 = {c5955,s5972[1]};
    assign in5988_2 = {c5956,s5973[1]};
    CLA_2 KS_5988(s5988, c5988, in5988_1, in5988_2);
    wire[0:0] s5989, in5989_1, in5989_2;
    wire c5989;
    assign in5989_1 = {c5957};
    assign in5989_2 = {c5958};
    Half_Adder KS_5989(s5989, c5989, in5989_1, in5989_2);
    wire[3:0] s5990, in5990_1, in5990_2;
    wire c5990;
    assign in5990_1 = {c5959,s5974[1],c4756,s4794[0]};
    assign in5990_2 = {c5967,s5975[1],s5971[2],s4795[0]};
    CLA_4 KS_5990(s5990, c5990, in5990_1, in5990_2);
    wire[0:0] s5991, in5991_1, in5991_2;
    wire c5991;
    assign in5991_1 = {s5971[0]};
    assign in5991_2 = {s5972[0]};
    Half_Adder KS_5991(s5991, c5991, in5991_1, in5991_2);
    wire[1:0] s5992, in5992_1, in5992_2;
    wire c5992;
    assign in5992_1 = {s5973[0],s5976[1]};
    assign in5992_2 = {s5974[0],s5977[1]};
    CLA_2 KS_5992(s5992, c5992, in5992_1, in5992_2);
    wire[0:0] s5993, in5993_1, in5993_2;
    wire c5993;
    assign in5993_1 = {s5976[0]};
    assign in5993_2 = {s5977[0]};
    Full_Adder KS_5993(s5993, c5993, in5993_1, in5993_2, s5975[0]);
    wire[3:0] s5994, in5994_1, in5994_2;
    wire c5994;
    assign in5994_1 = {s4771[1],s4761[2],c3304,s4806[0]};
    assign in5994_2 = {s4772[1],s4762[2],s3306[2],s4807[0]};
    CLA_4 KS_5994(s5994, c5994, in5994_1, in5994_2);
    wire[3:0] s5995, in5995_1, in5995_2;
    wire c5995;
    assign in5995_1 = {s4773[1],s4763[2],c3308,s4808[0]};
    assign in5995_2 = {s4774[1],s4764[2],s3310[2],s4809[0]};
    CLA_4 KS_5995(s5995, c5995, in5995_1, in5995_2);
    wire[3:0] s5996, in5996_1, in5996_2;
    wire c5996;
    assign in5996_1 = {s4775[1],s4765[2],s4760[3],s4810[0]};
    assign in5996_2 = {s4776[1],s4766[2],s4761[3],s4811[0]};
    CLA_4 KS_5996(s5996, c5996, in5996_1, in5996_2);
    wire[3:0] s5997, in5997_1, in5997_2;
    wire c5997;
    assign in5997_1 = {s4777[1],s4767[2],s4762[3],s4812[0]};
    assign in5997_2 = {s4778[1],s4768[2],s4763[3],s4813[0]};
    CLA_4 KS_5997(s5997, c5997, in5997_1, in5997_2);
    wire[3:0] s5998, in5998_1, in5998_2;
    wire c5998;
    assign in5998_1 = {c4779,s4769[2],s4764[3],s4814[0]};
    assign in5998_2 = {s4780[1],s4770[2],s4765[3],s4815[0]};
    CLA_4 KS_5998(s5998, c5998, in5998_1, in5998_2);
    wire[3:0] s5999, in5999_1, in5999_2;
    wire c5999;
    assign in5999_1 = {c4781,s4771[2],s4766[3],s4816[0]};
    assign in5999_2 = {s4782[1],s4772[2],s4767[3],s4817[0]};
    CLA_4 KS_5999(s5999, c5999, in5999_1, in5999_2);
    wire[3:0] s6000, in6000_1, in6000_2;
    wire c6000;
    assign in6000_1 = {c4783,s4773[2],s4768[3],s4818[0]};
    assign in6000_2 = {s4784[1],s4774[2],s4769[3],s4819[0]};
    CLA_4 KS_6000(s6000, c6000, in6000_1, in6000_2);
    wire[3:0] s6001, in6001_1, in6001_2;
    wire c6001;
    assign in6001_1 = {c4785,s4775[2],s4770[3],s4820[0]};
    assign in6001_2 = {s4786[1],s4776[2],s4771[3],s4821[0]};
    CLA_4 KS_6001(s6001, c6001, in6001_1, in6001_2);
    wire[3:0] s6002, in6002_1, in6002_2;
    wire c6002;
    assign in6002_1 = {c4787,s4777[2],s4772[3],s4822[0]};
    assign in6002_2 = {s4788[1],s4778[2],s4773[3],s4823[0]};
    CLA_4 KS_6002(s6002, c6002, in6002_1, in6002_2);
    wire[3:0] s6003, in6003_1, in6003_2;
    wire c6003;
    assign in6003_1 = {c4789,c4780,s4774[3],s4824[0]};
    assign in6003_2 = {s4790[1],s4782[2],s4775[3],s4825[0]};
    CLA_4 KS_6003(s6003, c6003, in6003_1, in6003_2);
    wire[3:0] s6004, in6004_1, in6004_2;
    wire c6004;
    assign in6004_1 = {c4791,c4784,s4776[3],s4826[0]};
    assign in6004_2 = {s4792[1],s4786[2],s4777[3],s4827[0]};
    CLA_4 KS_6004(s6004, c6004, in6004_1, in6004_2);
    wire[3:0] s6005, in6005_1, in6005_2;
    wire c6005;
    assign in6005_1 = {c4793,c4788,c4778,s4828[0]};
    assign in6005_2 = {s4794[1],s4790[2],s4782[3],s4829[0]};
    CLA_4 KS_6005(s6005, c6005, in6005_1, in6005_2);
    wire[0:0] s6006, in6006_1, in6006_2;
    wire c6006;
    assign in6006_1 = {c4795};
    assign in6006_2 = {s4796[1]};
    Half_Adder KS_6006(s6006, c6006, in6006_1, in6006_2);
    wire[1:0] s6007, in6007_1, in6007_2;
    wire c6007;
    assign in6007_1 = {c5971,c4792};
    assign in6007_2 = {c5972,s4794[2]};
    CLA_2 KS_6007(s6007, c6007, in6007_1, in6007_2);
    wire[0:0] s6008, in6008_1, in6008_2;
    wire c6008;
    assign in6008_1 = {c5973};
    assign in6008_2 = {c5974};
    Half_Adder KS_6008(s6008, c6008, in6008_1, in6008_2);
    wire[2:0] s6009, in6009_1, in6009_2;
    wire c6009;
    assign in6009_1 = {c5975,c4796,c4786};
    assign in6009_2 = {c5976,s5994[1],s4790[3]};
    CLA_3 KS_6009(s6009, c6009, in6009_1, in6009_2);
    wire[0:0] s6010, in6010_1, in6010_2;
    wire c6010;
    assign in6010_1 = {c5977};
    assign in6010_2 = {c5978};
    Half_Adder KS_6010(s6010, c6010, in6010_1, in6010_2);
    wire[1:0] s6011, in6011_1, in6011_2;
    wire c6011;
    assign in6011_1 = {c5979,s5995[1]};
    assign in6011_2 = {c5980,s5996[1]};
    CLA_2 KS_6011(s6011, c6011, in6011_1, in6011_2);
    wire[0:0] s6012, in6012_1, in6012_2;
    wire c6012;
    assign in6012_1 = {c5981};
    assign in6012_2 = {c5982};
    Half_Adder KS_6012(s6012, c6012, in6012_1, in6012_2);
    wire[3:0] s6013, in6013_1, in6013_2;
    wire c6013;
    assign in6013_1 = {c5990,s5997[1],c4794,s4830[0]};
    assign in6013_2 = {s5994[0],s5998[1],s5994[2],s4831[0]};
    CLA_4 KS_6013(s6013, c6013, in6013_1, in6013_2);
    wire[0:0] s6014, in6014_1, in6014_2;
    wire c6014;
    assign in6014_1 = {s5995[0]};
    assign in6014_2 = {s5996[0]};
    Half_Adder KS_6014(s6014, c6014, in6014_1, in6014_2);
    wire[1:0] s6015, in6015_1, in6015_2;
    wire c6015;
    assign in6015_1 = {s5998[0],s5999[1]};
    assign in6015_2 = {s5999[0],s6000[1]};
    CLA_2_c KS_6015(s6015, c6015, in6015_1, in6015_2, s5997[0]);
    wire[3:0] s6016, in6016_1, in6016_2;
    wire c6016;
    assign in6016_1 = {s4806[1],s4798[2],c3345,s4843[0]};
    assign in6016_2 = {s4807[1],s4799[2],s3347[2],s4844[0]};
    CLA_4 KS_6016(s6016, c6016, in6016_1, in6016_2);
    wire[3:0] s6017, in6017_1, in6017_2;
    wire c6017;
    assign in6017_1 = {s4808[1],s4800[2],c3349,s4845[0]};
    assign in6017_2 = {s4809[1],s4801[2],s3351[2],s4846[0]};
    CLA_4 KS_6017(s6017, c6017, in6017_1, in6017_2);
    wire[3:0] s6018, in6018_1, in6018_2;
    wire c6018;
    assign in6018_1 = {s4810[1],s4802[2],s4797[3],s4847[0]};
    assign in6018_2 = {s4811[1],s4803[2],s4798[3],s4848[0]};
    CLA_4 KS_6018(s6018, c6018, in6018_1, in6018_2);
    wire[3:0] s6019, in6019_1, in6019_2;
    wire c6019;
    assign in6019_1 = {s4812[1],s4804[2],s4799[3],s4849[0]};
    assign in6019_2 = {s4813[1],s4805[2],s4800[3],s4850[0]};
    CLA_4 KS_6019(s6019, c6019, in6019_1, in6019_2);
    wire[3:0] s6020, in6020_1, in6020_2;
    wire c6020;
    assign in6020_1 = {s4814[1],s4806[2],s4801[3],s4851[0]};
    assign in6020_2 = {s4815[1],s4807[2],s4802[3],s4852[0]};
    CLA_4 KS_6020(s6020, c6020, in6020_1, in6020_2);
    wire[3:0] s6021, in6021_1, in6021_2;
    wire c6021;
    assign in6021_1 = {c4816,s4808[2],s4803[3],s4853[0]};
    assign in6021_2 = {s4817[1],s4809[2],s4804[3],s4854[0]};
    CLA_4 KS_6021(s6021, c6021, in6021_1, in6021_2);
    wire[3:0] s6022, in6022_1, in6022_2;
    wire c6022;
    assign in6022_1 = {c4818,s4810[2],s4805[3],s4855[0]};
    assign in6022_2 = {s4819[1],s4811[2],s4806[3],s4856[0]};
    CLA_4 KS_6022(s6022, c6022, in6022_1, in6022_2);
    wire[3:0] s6023, in6023_1, in6023_2;
    wire c6023;
    assign in6023_1 = {c4820,s4812[2],s4807[3],s4857[0]};
    assign in6023_2 = {s4821[1],s4813[2],s4808[3],s4858[0]};
    CLA_4 KS_6023(s6023, c6023, in6023_1, in6023_2);
    wire[3:0] s6024, in6024_1, in6024_2;
    wire c6024;
    assign in6024_1 = {c4822,s4814[2],s4809[3],s4859[0]};
    assign in6024_2 = {s4823[1],s4815[2],s4810[3],s4860[0]};
    CLA_4 KS_6024(s6024, c6024, in6024_1, in6024_2);
    wire[3:0] s6025, in6025_1, in6025_2;
    wire c6025;
    assign in6025_1 = {c4824,c4817,s4811[3],s4861[0]};
    assign in6025_2 = {s4825[1],s4819[2],s4812[3],s4862[0]};
    CLA_4 KS_6025(s6025, c6025, in6025_1, in6025_2);
    wire[3:0] s6026, in6026_1, in6026_2;
    wire c6026;
    assign in6026_1 = {c4826,c4821,s4813[3],s4863[0]};
    assign in6026_2 = {s4827[1],s4823[2],s4814[3],s4864[0]};
    CLA_4 KS_6026(s6026, c6026, in6026_1, in6026_2);
    wire[0:0] s6027, in6027_1, in6027_2;
    wire c6027;
    assign in6027_1 = {c4828};
    assign in6027_2 = {s4829[1]};
    Half_Adder KS_6027(s6027, c6027, in6027_1, in6027_2);
    wire[3:0] s6028, in6028_1, in6028_2;
    wire c6028;
    assign in6028_1 = {c4830,c4825,c4815,s4865[0]};
    assign in6028_2 = {s4831[1],s4827[2],s4819[3],s4866[0]};
    CLA_4 KS_6028(s6028, c6028, in6028_1, in6028_2);
    wire[0:0] s6029, in6029_1, in6029_2;
    wire c6029;
    assign in6029_1 = {c4832};
    assign in6029_2 = {c5994};
    Half_Adder KS_6029(s6029, c6029, in6029_1, in6029_2);
    wire[1:0] s6030, in6030_1, in6030_2;
    wire c6030;
    assign in6030_1 = {c5995,c4829};
    assign in6030_2 = {c5996,s4831[2]};
    CLA_2 KS_6030(s6030, c6030, in6030_1, in6030_2);
    wire[0:0] s6031, in6031_1, in6031_2;
    wire c6031;
    assign in6031_1 = {c5997};
    assign in6031_2 = {c5998};
    Half_Adder KS_6031(s6031, c6031, in6031_1, in6031_2);
    wire[2:0] s6032, in6032_1, in6032_2;
    wire c6032;
    assign in6032_1 = {c5999,s6016[1],c4823};
    assign in6032_2 = {c6000,s6017[1],s4827[3]};
    CLA_3 KS_6032(s6032, c6032, in6032_1, in6032_2);
    wire[0:0] s6033, in6033_1, in6033_2;
    wire c6033;
    assign in6033_1 = {c6001};
    assign in6033_2 = {c6002};
    Half_Adder KS_6033(s6033, c6033, in6033_1, in6033_2);
    wire[1:0] s6034, in6034_1, in6034_2;
    wire c6034;
    assign in6034_1 = {c6003,s6018[1]};
    assign in6034_2 = {c6004,s6019[1]};
    CLA_2 KS_6034(s6034, c6034, in6034_1, in6034_2);
    wire[0:0] s6035, in6035_1, in6035_2;
    wire c6035;
    assign in6035_1 = {c6005};
    assign in6035_2 = {c6013};
    Half_Adder KS_6035(s6035, c6035, in6035_1, in6035_2);
    wire[3:0] s6036, in6036_1, in6036_2;
    wire c6036;
    assign in6036_1 = {s6016[0],s6020[1],c4831,s4867[0]};
    assign in6036_2 = {s6017[0],s6021[1],s6016[2],s4868[0]};
    CLA_4 KS_6036(s6036, c6036, in6036_1, in6036_2);
    wire[0:0] s6037, in6037_1, in6037_2;
    wire c6037;
    assign in6037_1 = {s6018[0]};
    assign in6037_2 = {s6019[0]};
    Half_Adder KS_6037(s6037, c6037, in6037_1, in6037_2);
    wire[1:0] s6038, in6038_1, in6038_2;
    wire c6038;
    assign in6038_1 = {s6021[0],s6022[1]};
    assign in6038_2 = {s6022[0],s6023[1]};
    CLA_2_c KS_6038(s6038, c6038, in6038_1, in6038_2, s6020[0]);
    wire[3:0] s6039, in6039_1, in6039_2;
    wire c6039;
    assign in6039_1 = {s4844[1],s4835[2],c3378,s4879[0]};
    assign in6039_2 = {s4845[1],s4836[2],s3380[2],s4880[0]};
    CLA_4 KS_6039(s6039, c6039, in6039_1, in6039_2);
    wire[3:0] s6040, in6040_1, in6040_2;
    wire c6040;
    assign in6040_1 = {s4846[1],s4837[2],c3382,s4881[0]};
    assign in6040_2 = {s4847[1],s4838[2],s3384[2],s4882[0]};
    CLA_4 KS_6040(s6040, c6040, in6040_1, in6040_2);
    wire[3:0] s6041, in6041_1, in6041_2;
    wire c6041;
    assign in6041_1 = {s4848[1],s4839[2],s4833[3],s4883[0]};
    assign in6041_2 = {s4849[1],s4840[2],s4834[3],s4884[0]};
    CLA_4 KS_6041(s6041, c6041, in6041_1, in6041_2);
    wire[3:0] s6042, in6042_1, in6042_2;
    wire c6042;
    assign in6042_1 = {s4850[1],s4841[2],s4835[3],s4885[0]};
    assign in6042_2 = {s4851[1],s4842[2],s4836[3],s4886[0]};
    CLA_4 KS_6042(s6042, c6042, in6042_1, in6042_2);
    wire[3:0] s6043, in6043_1, in6043_2;
    wire c6043;
    assign in6043_1 = {c4852,s4843[2],s4837[3],s4887[0]};
    assign in6043_2 = {s4853[1],s4844[2],s4838[3],s4888[0]};
    CLA_4 KS_6043(s6043, c6043, in6043_1, in6043_2);
    wire[3:0] s6044, in6044_1, in6044_2;
    wire c6044;
    assign in6044_1 = {c4854,s4845[2],s4839[3],s4889[0]};
    assign in6044_2 = {s4855[1],s4846[2],s4840[3],s4890[0]};
    CLA_4 KS_6044(s6044, c6044, in6044_1, in6044_2);
    wire[3:0] s6045, in6045_1, in6045_2;
    wire c6045;
    assign in6045_1 = {c4856,s4847[2],s4841[3],s4891[0]};
    assign in6045_2 = {s4857[1],s4848[2],s4842[3],s4892[0]};
    CLA_4 KS_6045(s6045, c6045, in6045_1, in6045_2);
    wire[3:0] s6046, in6046_1, in6046_2;
    wire c6046;
    assign in6046_1 = {c4858,s4849[2],s4843[3],s4893[0]};
    assign in6046_2 = {s4859[1],s4850[2],s4844[3],s4894[0]};
    CLA_4 KS_6046(s6046, c6046, in6046_1, in6046_2);
    wire[3:0] s6047, in6047_1, in6047_2;
    wire c6047;
    assign in6047_1 = {c4860,c4851,s4845[3],s4895[0]};
    assign in6047_2 = {s4861[1],s4853[2],s4846[3],s4896[0]};
    CLA_4 KS_6047(s6047, c6047, in6047_1, in6047_2);
    wire[3:0] s6048, in6048_1, in6048_2;
    wire c6048;
    assign in6048_1 = {c4862,c4855,s4847[3],s4897[0]};
    assign in6048_2 = {s4863[1],s4857[2],s4848[3],s4898[0]};
    CLA_4 KS_6048(s6048, c6048, in6048_1, in6048_2);
    wire[3:0] s6049, in6049_1, in6049_2;
    wire c6049;
    assign in6049_1 = {c4864,c4859,s4849[3],s4899[0]};
    assign in6049_2 = {s4865[1],s4861[2],s4850[3],s4900[0]};
    CLA_4 KS_6049(s6049, c6049, in6049_1, in6049_2);
    wire[0:0] s6050, in6050_1, in6050_2;
    wire c6050;
    assign in6050_1 = {c4866};
    assign in6050_2 = {s4867[1]};
    Half_Adder KS_6050(s6050, c6050, in6050_1, in6050_2);
    wire[3:0] s6051, in6051_1, in6051_2;
    wire c6051;
    assign in6051_1 = {c4868,c4863,c4853,s4901[0]};
    assign in6051_2 = {s4869[1],s4865[2],s4857[3],s4902[0]};
    CLA_4 KS_6051(s6051, c6051, in6051_1, in6051_2);
    wire[0:0] s6052, in6052_1, in6052_2;
    wire c6052;
    assign in6052_1 = {c6016};
    assign in6052_2 = {c6017};
    Half_Adder KS_6052(s6052, c6052, in6052_1, in6052_2);
    wire[1:0] s6053, in6053_1, in6053_2;
    wire c6053;
    assign in6053_1 = {c6018,c4867};
    assign in6053_2 = {c6019,s4869[2]};
    CLA_2 KS_6053(s6053, c6053, in6053_1, in6053_2);
    wire[0:0] s6054, in6054_1, in6054_2;
    wire c6054;
    assign in6054_1 = {c6020};
    assign in6054_2 = {c6021};
    Half_Adder KS_6054(s6054, c6054, in6054_1, in6054_2);
    wire[2:0] s6055, in6055_1, in6055_2;
    wire c6055;
    assign in6055_1 = {c6022,s6039[1],c4861};
    assign in6055_2 = {c6023,s6040[1],s4865[3]};
    CLA_3 KS_6055(s6055, c6055, in6055_1, in6055_2);
    wire[0:0] s6056, in6056_1, in6056_2;
    wire c6056;
    assign in6056_1 = {c6024};
    assign in6056_2 = {c6025};
    Half_Adder KS_6056(s6056, c6056, in6056_1, in6056_2);
    wire[1:0] s6057, in6057_1, in6057_2;
    wire c6057;
    assign in6057_1 = {c6026,s6041[1]};
    assign in6057_2 = {c6028,s6042[1]};
    CLA_2 KS_6057(s6057, c6057, in6057_1, in6057_2);
    wire[0:0] s6058, in6058_1, in6058_2;
    wire c6058;
    assign in6058_1 = {c6036};
    assign in6058_2 = {s6039[0]};
    Half_Adder KS_6058(s6058, c6058, in6058_1, in6058_2);
    wire[3:0] s6059, in6059_1, in6059_2;
    wire c6059;
    assign in6059_1 = {s6040[0],s6043[1],c4869,s4903[0]};
    assign in6059_2 = {s6041[0],s6044[1],s6039[2],s4904[0]};
    CLA_4 KS_6059(s6059, c6059, in6059_1, in6059_2);
    wire[0:0] s6060, in6060_1, in6060_2;
    wire c6060;
    assign in6060_1 = {s6043[0]};
    assign in6060_2 = {s6044[0]};
    Full_Adder KS_6060(s6060, c6060, in6060_1, in6060_2, s6042[0]);
    wire[3:0] s6061, in6061_1, in6061_2;
    wire c6061;
    assign in6061_1 = {s4879[1],s4870[2],c3402,s4916[0]};
    assign in6061_2 = {s4880[1],s4871[2],s3404[2],s4917[0]};
    CLA_4 KS_6061(s6061, c6061, in6061_1, in6061_2);
    wire[3:0] s6062, in6062_1, in6062_2;
    wire c6062;
    assign in6062_1 = {s4881[1],s4872[2],c3406,s4918[0]};
    assign in6062_2 = {s4882[1],s4873[2],s3408[2],s4919[0]};
    CLA_4 KS_6062(s6062, c6062, in6062_1, in6062_2);
    wire[3:0] s6063, in6063_1, in6063_2;
    wire c6063;
    assign in6063_1 = {s4883[1],s4874[2],s4870[3],s4920[0]};
    assign in6063_2 = {s4884[1],s4875[2],s4871[3],s4921[0]};
    CLA_4 KS_6063(s6063, c6063, in6063_1, in6063_2);
    wire[3:0] s6064, in6064_1, in6064_2;
    wire c6064;
    assign in6064_1 = {s4885[1],s4876[2],s4872[3],s4922[0]};
    assign in6064_2 = {s4886[1],s4877[2],s4873[3],s4923[0]};
    CLA_4 KS_6064(s6064, c6064, in6064_1, in6064_2);
    wire[3:0] s6065, in6065_1, in6065_2;
    wire c6065;
    assign in6065_1 = {s4887[1],s4878[2],s4874[3],s4924[0]};
    assign in6065_2 = {s4888[1],s4879[2],s4875[3],s4925[0]};
    CLA_4 KS_6065(s6065, c6065, in6065_1, in6065_2);
    wire[3:0] s6066, in6066_1, in6066_2;
    wire c6066;
    assign in6066_1 = {c4889,s4880[2],s4876[3],s4926[0]};
    assign in6066_2 = {s4890[1],s4881[2],s4877[3],s4927[0]};
    CLA_4 KS_6066(s6066, c6066, in6066_1, in6066_2);
    wire[3:0] s6067, in6067_1, in6067_2;
    wire c6067;
    assign in6067_1 = {c4891,s4882[2],s4878[3],s4928[0]};
    assign in6067_2 = {s4892[1],s4883[2],s4879[3],s4929[0]};
    CLA_4 KS_6067(s6067, c6067, in6067_1, in6067_2);
    wire[3:0] s6068, in6068_1, in6068_2;
    wire c6068;
    assign in6068_1 = {c4893,s4884[2],s4880[3],s4930[0]};
    assign in6068_2 = {s4894[1],s4885[2],s4881[3],s4931[0]};
    CLA_4 KS_6068(s6068, c6068, in6068_1, in6068_2);
    wire[3:0] s6069, in6069_1, in6069_2;
    wire c6069;
    assign in6069_1 = {c4895,s4886[2],s4882[3],s4932[0]};
    assign in6069_2 = {s4896[1],s4887[2],s4883[3],s4933[0]};
    CLA_4 KS_6069(s6069, c6069, in6069_1, in6069_2);
    wire[3:0] s6070, in6070_1, in6070_2;
    wire c6070;
    assign in6070_1 = {c4897,c4888,s4884[3],s4934[0]};
    assign in6070_2 = {s4898[1],s4890[2],s4885[3],s4935[0]};
    CLA_4 KS_6070(s6070, c6070, in6070_1, in6070_2);
    wire[3:0] s6071, in6071_1, in6071_2;
    wire c6071;
    assign in6071_1 = {c4899,c4892,s4886[3],s4936[0]};
    assign in6071_2 = {s4900[1],s4894[2],s4887[3],s4937[0]};
    CLA_4 KS_6071(s6071, c6071, in6071_1, in6071_2);
    wire[1:0] s6072, in6072_1, in6072_2;
    wire c6072;
    assign in6072_1 = {c4901,c4896};
    assign in6072_2 = {s4902[1],s4898[2]};
    CLA_2 KS_6072(s6072, c6072, in6072_1, in6072_2);
    wire[0:0] s6073, in6073_1, in6073_2;
    wire c6073;
    assign in6073_1 = {c4903};
    assign in6073_2 = {s4904[1]};
    Half_Adder KS_6073(s6073, c6073, in6073_1, in6073_2);
    wire[3:0] s6074, in6074_1, in6074_2;
    wire c6074;
    assign in6074_1 = {c4905,c4900,c4890,s4938[0]};
    assign in6074_2 = {c6039,s4902[2],s4894[3],s4939[0]};
    CLA_4 KS_6074(s6074, c6074, in6074_1, in6074_2);
    wire[0:0] s6075, in6075_1, in6075_2;
    wire c6075;
    assign in6075_1 = {c6040};
    assign in6075_2 = {c6041};
    Half_Adder KS_6075(s6075, c6075, in6075_1, in6075_2);
    wire[1:0] s6076, in6076_1, in6076_2;
    wire c6076;
    assign in6076_1 = {c6042,c4904};
    assign in6076_2 = {c6043,s6061[1]};
    CLA_2 KS_6076(s6076, c6076, in6076_1, in6076_2);
    wire[0:0] s6077, in6077_1, in6077_2;
    wire c6077;
    assign in6077_1 = {c6044};
    assign in6077_2 = {c6045};
    Half_Adder KS_6077(s6077, c6077, in6077_1, in6077_2);
    wire[2:0] s6078, in6078_1, in6078_2;
    wire c6078;
    assign in6078_1 = {c6046,s6062[1],c4898};
    assign in6078_2 = {c6047,s6063[1],s4902[3]};
    CLA_3 KS_6078(s6078, c6078, in6078_1, in6078_2);
    wire[0:0] s6079, in6079_1, in6079_2;
    wire c6079;
    assign in6079_1 = {c6048};
    assign in6079_2 = {c6049};
    Half_Adder KS_6079(s6079, c6079, in6079_1, in6079_2);
    wire[1:0] s6080, in6080_1, in6080_2;
    wire c6080;
    assign in6080_1 = {c6051,s6064[1]};
    assign in6080_2 = {c6059,s6065[1]};
    CLA_2 KS_6080(s6080, c6080, in6080_1, in6080_2);
    wire[0:0] s6081, in6081_1, in6081_2;
    wire c6081;
    assign in6081_1 = {s6061[0]};
    assign in6081_2 = {s6062[0]};
    Half_Adder KS_6081(s6081, c6081, in6081_1, in6081_2);
    wire[3:0] s6082, in6082_1, in6082_2;
    wire c6082;
    assign in6082_1 = {s6063[0],s6066[1],s6061[2],s4940[0]};
    assign in6082_2 = {s6064[0],s6067[1],s6062[2],s4941[0]};
    CLA_4 KS_6082(s6082, c6082, in6082_1, in6082_2);
    wire[0:0] s6083, in6083_1, in6083_2;
    wire c6083;
    assign in6083_1 = {s6066[0]};
    assign in6083_2 = {s6067[0]};
    Full_Adder KS_6083(s6083, c6083, in6083_1, in6083_2, s6065[0]);
    wire[3:0] s6084, in6084_1, in6084_2;
    wire c6084;
    assign in6084_1 = {s4917[1],s4907[2],c3418,s4954[0]};
    assign in6084_2 = {s4918[1],s4908[2],s3420[2],s4955[0]};
    CLA_4 KS_6084(s6084, c6084, in6084_1, in6084_2);
    wire[3:0] s6085, in6085_1, in6085_2;
    wire c6085;
    assign in6085_1 = {s4919[1],s4909[2],c3422,s4956[0]};
    assign in6085_2 = {s4920[1],s4910[2],s4906[3],s4957[0]};
    CLA_4 KS_6085(s6085, c6085, in6085_1, in6085_2);
    wire[3:0] s6086, in6086_1, in6086_2;
    wire c6086;
    assign in6086_1 = {s4921[1],s4911[2],s4907[3],s4958[0]};
    assign in6086_2 = {s4922[1],s4912[2],s4908[3],s4959[0]};
    CLA_4 KS_6086(s6086, c6086, in6086_1, in6086_2);
    wire[3:0] s6087, in6087_1, in6087_2;
    wire c6087;
    assign in6087_1 = {s4923[1],s4913[2],s4909[3],s4960[0]};
    assign in6087_2 = {s4924[1],s4914[2],s4910[3],s4961[0]};
    CLA_4 KS_6087(s6087, c6087, in6087_1, in6087_2);
    wire[3:0] s6088, in6088_1, in6088_2;
    wire c6088;
    assign in6088_1 = {c4925,s4915[2],s4911[3],s4962[0]};
    assign in6088_2 = {s4926[1],s4916[2],s4912[3],s4963[0]};
    CLA_4 KS_6088(s6088, c6088, in6088_1, in6088_2);
    wire[3:0] s6089, in6089_1, in6089_2;
    wire c6089;
    assign in6089_1 = {c4927,s4917[2],s4913[3],s4964[0]};
    assign in6089_2 = {s4928[1],s4918[2],s4914[3],s4965[0]};
    CLA_4 KS_6089(s6089, c6089, in6089_1, in6089_2);
    wire[3:0] s6090, in6090_1, in6090_2;
    wire c6090;
    assign in6090_1 = {c4929,s4919[2],s4915[3],s4966[0]};
    assign in6090_2 = {s4930[1],s4920[2],s4916[3],s4967[0]};
    CLA_4 KS_6090(s6090, c6090, in6090_1, in6090_2);
    wire[3:0] s6091, in6091_1, in6091_2;
    wire c6091;
    assign in6091_1 = {c4931,s4921[2],s4917[3],s4968[0]};
    assign in6091_2 = {s4932[1],s4922[2],s4918[3],s4969[0]};
    CLA_4 KS_6091(s6091, c6091, in6091_1, in6091_2);
    wire[3:0] s6092, in6092_1, in6092_2;
    wire c6092;
    assign in6092_1 = {c4933,s4923[2],s4919[3],s4970[0]};
    assign in6092_2 = {s4934[1],s4924[2],s4920[3],s4971[0]};
    CLA_4 KS_6092(s6092, c6092, in6092_1, in6092_2);
    wire[3:0] s6093, in6093_1, in6093_2;
    wire c6093;
    assign in6093_1 = {c4935,c4926,s4921[3],s4972[0]};
    assign in6093_2 = {s4936[1],s4928[2],s4922[3],s4973[0]};
    CLA_4 KS_6093(s6093, c6093, in6093_1, in6093_2);
    wire[3:0] s6094, in6094_1, in6094_2;
    wire c6094;
    assign in6094_1 = {c4937,c4930,s4923[3],s4974[0]};
    assign in6094_2 = {s4938[1],s4932[2],s4924[3],s4975[0]};
    CLA_4 KS_6094(s6094, c6094, in6094_1, in6094_2);
    wire[1:0] s6095, in6095_1, in6095_2;
    wire c6095;
    assign in6095_1 = {c4939,c4934};
    assign in6095_2 = {s4940[1],s4936[2]};
    CLA_2 KS_6095(s6095, c6095, in6095_1, in6095_2);
    wire[0:0] s6096, in6096_1, in6096_2;
    wire c6096;
    assign in6096_1 = {c4941};
    assign in6096_2 = {s4942[1]};
    Half_Adder KS_6096(s6096, c6096, in6096_1, in6096_2);
    wire[3:0] s6097, in6097_1, in6097_2;
    wire c6097;
    assign in6097_1 = {c6061,c4938,c4928,s4976[0]};
    assign in6097_2 = {c6062,s4940[2],s4932[3],s4977[0]};
    CLA_4 KS_6097(s6097, c6097, in6097_1, in6097_2);
    wire[0:0] s6098, in6098_1, in6098_2;
    wire c6098;
    assign in6098_1 = {c6063};
    assign in6098_2 = {c6064};
    Half_Adder KS_6098(s6098, c6098, in6098_1, in6098_2);
    wire[1:0] s6099, in6099_1, in6099_2;
    wire c6099;
    assign in6099_1 = {c6065,c4942};
    assign in6099_2 = {c6066,s6084[1]};
    CLA_2 KS_6099(s6099, c6099, in6099_1, in6099_2);
    wire[0:0] s6100, in6100_1, in6100_2;
    wire c6100;
    assign in6100_1 = {c6067};
    assign in6100_2 = {c6068};
    Half_Adder KS_6100(s6100, c6100, in6100_1, in6100_2);
    wire[2:0] s6101, in6101_1, in6101_2;
    wire c6101;
    assign in6101_1 = {c6069,s6085[1],c4936};
    assign in6101_2 = {c6070,s6086[1],s4940[3]};
    CLA_3 KS_6101(s6101, c6101, in6101_1, in6101_2);
    wire[0:0] s6102, in6102_1, in6102_2;
    wire c6102;
    assign in6102_1 = {c6071};
    assign in6102_2 = {c6074};
    Half_Adder KS_6102(s6102, c6102, in6102_1, in6102_2);
    wire[1:0] s6103, in6103_1, in6103_2;
    wire c6103;
    assign in6103_1 = {c6082,s6087[1]};
    assign in6103_2 = {s6084[0],s6088[1]};
    CLA_2 KS_6103(s6103, c6103, in6103_1, in6103_2);
    wire[0:0] s6104, in6104_1, in6104_2;
    wire c6104;
    assign in6104_1 = {s6085[0]};
    assign in6104_2 = {s6086[0]};
    Half_Adder KS_6104(s6104, c6104, in6104_1, in6104_2);
    wire[3:0] s6105, in6105_1, in6105_2;
    wire c6105;
    assign in6105_1 = {s6088[0],s6089[1],s6084[2],s4978[0]};
    assign in6105_2 = {s6089[0],s6090[1],s6085[2],s4979[0]};
    CLA_4_c KS_6105(s6105, c6105, in6105_1, in6105_2, s6087[0]);
    wire[3:0] s6106, in6106_1, in6106_2;
    wire c6106;
    assign in6106_1 = {s4954[1],s4945[2],c3425,s4991[0]};
    assign in6106_2 = {s4955[1],s4946[2],s3427[2],s4992[0]};
    CLA_4 KS_6106(s6106, c6106, in6106_1, in6106_2);
    wire[3:0] s6107, in6107_1, in6107_2;
    wire c6107;
    assign in6107_1 = {s4956[1],s4947[2],c3429,s4993[0]};
    assign in6107_2 = {s4957[1],s4948[2],s4943[3],s4994[0]};
    CLA_4 KS_6107(s6107, c6107, in6107_1, in6107_2);
    wire[3:0] s6108, in6108_1, in6108_2;
    wire c6108;
    assign in6108_1 = {s4958[1],s4949[2],s4944[3],s4995[0]};
    assign in6108_2 = {s4959[1],s4950[2],s4945[3],s4996[0]};
    CLA_4 KS_6108(s6108, c6108, in6108_1, in6108_2);
    wire[3:0] s6109, in6109_1, in6109_2;
    wire c6109;
    assign in6109_1 = {s4960[1],s4951[2],s4946[3],s4997[0]};
    assign in6109_2 = {s4961[1],s4952[2],s4947[3],s4998[0]};
    CLA_4 KS_6109(s6109, c6109, in6109_1, in6109_2);
    wire[3:0] s6110, in6110_1, in6110_2;
    wire c6110;
    assign in6110_1 = {c4962,s4953[2],s4948[3],s4999[0]};
    assign in6110_2 = {s4963[1],s4954[2],s4949[3],s5000[0]};
    CLA_4 KS_6110(s6110, c6110, in6110_1, in6110_2);
    wire[3:0] s6111, in6111_1, in6111_2;
    wire c6111;
    assign in6111_1 = {c4964,s4955[2],s4950[3],s5001[0]};
    assign in6111_2 = {s4965[1],s4956[2],s4951[3],s5002[0]};
    CLA_4 KS_6111(s6111, c6111, in6111_1, in6111_2);
    wire[3:0] s6112, in6112_1, in6112_2;
    wire c6112;
    assign in6112_1 = {c4966,s4957[2],s4952[3],s5003[0]};
    assign in6112_2 = {s4967[1],s4958[2],s4953[3],s5004[0]};
    CLA_4 KS_6112(s6112, c6112, in6112_1, in6112_2);
    wire[3:0] s6113, in6113_1, in6113_2;
    wire c6113;
    assign in6113_1 = {c4968,s4959[2],s4954[3],s5005[0]};
    assign in6113_2 = {s4969[1],s4960[2],s4955[3],s5006[0]};
    CLA_4 KS_6113(s6113, c6113, in6113_1, in6113_2);
    wire[3:0] s6114, in6114_1, in6114_2;
    wire c6114;
    assign in6114_1 = {c4970,c4961,s4956[3],s5007[0]};
    assign in6114_2 = {s4971[1],s4963[2],s4957[3],s5008[0]};
    CLA_4 KS_6114(s6114, c6114, in6114_1, in6114_2);
    wire[3:0] s6115, in6115_1, in6115_2;
    wire c6115;
    assign in6115_1 = {c4972,c4965,s4958[3],s5009[0]};
    assign in6115_2 = {s4973[1],s4967[2],s4959[3],s5010[0]};
    CLA_4 KS_6115(s6115, c6115, in6115_1, in6115_2);
    wire[3:0] s6116, in6116_1, in6116_2;
    wire c6116;
    assign in6116_1 = {c4974,c4969,s4960[3],s5011[0]};
    assign in6116_2 = {s4975[1],s4971[2],s4963[3],s5012[0]};
    CLA_4 KS_6116(s6116, c6116, in6116_1, in6116_2);
    wire[0:0] s6117, in6117_1, in6117_2;
    wire c6117;
    assign in6117_1 = {c4976};
    assign in6117_2 = {s4977[1]};
    Half_Adder KS_6117(s6117, c6117, in6117_1, in6117_2);
    wire[1:0] s6118, in6118_1, in6118_2;
    wire c6118;
    assign in6118_1 = {c4978,c4973};
    assign in6118_2 = {s4979[1],s4975[2]};
    CLA_2 KS_6118(s6118, c6118, in6118_1, in6118_2);
    wire[0:0] s6119, in6119_1, in6119_2;
    wire c6119;
    assign in6119_1 = {c4980};
    assign in6119_2 = {c6084};
    Half_Adder KS_6119(s6119, c6119, in6119_1, in6119_2);
    wire[3:0] s6120, in6120_1, in6120_2;
    wire c6120;
    assign in6120_1 = {c6085,c4977,c4967,s5013[0]};
    assign in6120_2 = {c6086,s4979[2],s4971[3],s5014[0]};
    CLA_4 KS_6120(s6120, c6120, in6120_1, in6120_2);
    wire[0:0] s6121, in6121_1, in6121_2;
    wire c6121;
    assign in6121_1 = {c6087};
    assign in6121_2 = {c6088};
    Half_Adder KS_6121(s6121, c6121, in6121_1, in6121_2);
    wire[1:0] s6122, in6122_1, in6122_2;
    wire c6122;
    assign in6122_1 = {c6089,s6106[1]};
    assign in6122_2 = {c6090,s6107[1]};
    CLA_2 KS_6122(s6122, c6122, in6122_1, in6122_2);
    wire[0:0] s6123, in6123_1, in6123_2;
    wire c6123;
    assign in6123_1 = {c6091};
    assign in6123_2 = {c6092};
    Half_Adder KS_6123(s6123, c6123, in6123_1, in6123_2);
    wire[2:0] s6124, in6124_1, in6124_2;
    wire c6124;
    assign in6124_1 = {c6093,s6108[1],c4975};
    assign in6124_2 = {c6094,s6109[1],s4979[3]};
    CLA_3 KS_6124(s6124, c6124, in6124_1, in6124_2);
    wire[0:0] s6125, in6125_1, in6125_2;
    wire c6125;
    assign in6125_1 = {c6097};
    assign in6125_2 = {c6105};
    Half_Adder KS_6125(s6125, c6125, in6125_1, in6125_2);
    wire[1:0] s6126, in6126_1, in6126_2;
    wire c6126;
    assign in6126_1 = {s6106[0],s6110[1]};
    assign in6126_2 = {s6107[0],s6111[1]};
    CLA_2 KS_6126(s6126, c6126, in6126_1, in6126_2);
    wire[0:0] s6127, in6127_1, in6127_2;
    wire c6127;
    assign in6127_1 = {s6108[0]};
    assign in6127_2 = {s6109[0]};
    Half_Adder KS_6127(s6127, c6127, in6127_1, in6127_2);
    wire[3:0] s6128, in6128_1, in6128_2;
    wire c6128;
    assign in6128_1 = {s6111[0],s6112[1],s6106[2],s5015[0]};
    assign in6128_2 = {s6112[0],s6113[1],s6107[2],s5016[0]};
    CLA_4_c KS_6128(s6128, c6128, in6128_1, in6128_2, s6110[0]);
    wire[3:0] s6129, in6129_1, in6129_2;
    wire c6129;
    assign in6129_1 = {s4991[1],s4981[2],pp123[91],s5021[0]};
    assign in6129_2 = {s4992[1],s4982[2],pp124[90],s5022[0]};
    CLA_4 KS_6129(s6129, c6129, in6129_1, in6129_2);
    wire[3:0] s6130, in6130_1, in6130_2;
    wire c6130;
    assign in6130_1 = {s4993[1],s4983[2],pp125[89],s5023[0]};
    assign in6130_2 = {s4994[1],s4984[2],pp126[88],s5024[0]};
    CLA_4 KS_6130(s6130, c6130, in6130_1, in6130_2);
    wire[3:0] s6131, in6131_1, in6131_2;
    wire c6131;
    assign in6131_1 = {s4995[1],s4985[2],pp127[87],s5025[0]};
    assign in6131_2 = {s4996[1],s4986[2],s4981[3],s5026[0]};
    CLA_4 KS_6131(s6131, c6131, in6131_1, in6131_2);
    wire[3:0] s6132, in6132_1, in6132_2;
    wire c6132;
    assign in6132_1 = {s4997[1],s4987[2],s4982[3],s5027[0]};
    assign in6132_2 = {s4998[1],s4988[2],s4983[3],s5028[0]};
    CLA_4 KS_6132(s6132, c6132, in6132_1, in6132_2);
    wire[3:0] s6133, in6133_1, in6133_2;
    wire c6133;
    assign in6133_1 = {c4999,s4989[2],s4984[3],s5029[0]};
    assign in6133_2 = {s5000[1],s4990[2],s4985[3],s5030[0]};
    CLA_4 KS_6133(s6133, c6133, in6133_1, in6133_2);
    wire[3:0] s6134, in6134_1, in6134_2;
    wire c6134;
    assign in6134_1 = {c5001,s4991[2],s4986[3],s5031[0]};
    assign in6134_2 = {s5002[1],s4992[2],s4987[3],s5032[0]};
    CLA_4 KS_6134(s6134, c6134, in6134_1, in6134_2);
    wire[3:0] s6135, in6135_1, in6135_2;
    wire c6135;
    assign in6135_1 = {c5003,s4993[2],s4988[3],s5033[0]};
    assign in6135_2 = {s5004[1],s4994[2],s4989[3],s5034[0]};
    CLA_4 KS_6135(s6135, c6135, in6135_1, in6135_2);
    wire[3:0] s6136, in6136_1, in6136_2;
    wire c6136;
    assign in6136_1 = {c5005,s4995[2],s4990[3],s5035[0]};
    assign in6136_2 = {s5006[1],s4996[2],s4991[3],s5036[0]};
    CLA_4 KS_6136(s6136, c6136, in6136_1, in6136_2);
    wire[3:0] s6137, in6137_1, in6137_2;
    wire c6137;
    assign in6137_1 = {c5007,c4997,s4992[3],s5037[0]};
    assign in6137_2 = {s5008[1],s4998[2],s4993[3],s5038[0]};
    CLA_4 KS_6137(s6137, c6137, in6137_1, in6137_2);
    wire[3:0] s6138, in6138_1, in6138_2;
    wire c6138;
    assign in6138_1 = {c5009,c5000,s4994[3],s5039[0]};
    assign in6138_2 = {s5010[1],s5002[2],s4995[3],s5040[0]};
    CLA_4 KS_6138(s6138, c6138, in6138_1, in6138_2);
    wire[3:0] s6139, in6139_1, in6139_2;
    wire c6139;
    assign in6139_1 = {c5011,c5004,c4996,s5041[0]};
    assign in6139_2 = {s5012[1],s5006[2],s4998[3],s5042[0]};
    CLA_4 KS_6139(s6139, c6139, in6139_1, in6139_2);
    wire[1:0] s6140, in6140_1, in6140_2;
    wire c6140;
    assign in6140_1 = {c5013,c5008};
    assign in6140_2 = {s5014[1],s5010[2]};
    CLA_2 KS_6140(s6140, c6140, in6140_1, in6140_2);
    wire[0:0] s6141, in6141_1, in6141_2;
    wire c6141;
    assign in6141_1 = {c5015};
    assign in6141_2 = {s5016[1]};
    Half_Adder KS_6141(s6141, c6141, in6141_1, in6141_2);
    wire[3:0] s6142, in6142_1, in6142_2;
    wire c6142;
    assign in6142_1 = {c5017,c5012,c5002,s5043[0]};
    assign in6142_2 = {c6106,s5014[2],s5006[3],s5044[0]};
    CLA_4 KS_6142(s6142, c6142, in6142_1, in6142_2);
    wire[0:0] s6143, in6143_1, in6143_2;
    wire c6143;
    assign in6143_1 = {c6107};
    assign in6143_2 = {c6108};
    Half_Adder KS_6143(s6143, c6143, in6143_1, in6143_2);
    wire[1:0] s6144, in6144_1, in6144_2;
    wire c6144;
    assign in6144_1 = {c6109,c5016};
    assign in6144_2 = {c6110,s6129[1]};
    CLA_2 KS_6144(s6144, c6144, in6144_1, in6144_2);
    wire[0:0] s6145, in6145_1, in6145_2;
    wire c6145;
    assign in6145_1 = {c6111};
    assign in6145_2 = {c6112};
    Half_Adder KS_6145(s6145, c6145, in6145_1, in6145_2);
    wire[2:0] s6146, in6146_1, in6146_2;
    wire c6146;
    assign in6146_1 = {c6113,s6130[1],c5010};
    assign in6146_2 = {c6114,s6131[1],s5014[3]};
    CLA_3 KS_6146(s6146, c6146, in6146_1, in6146_2);
    wire[0:0] s6147, in6147_1, in6147_2;
    wire c6147;
    assign in6147_1 = {c6115};
    assign in6147_2 = {c6116};
    Half_Adder KS_6147(s6147, c6147, in6147_1, in6147_2);
    wire[1:0] s6148, in6148_1, in6148_2;
    wire c6148;
    assign in6148_1 = {c6120,s6132[1]};
    assign in6148_2 = {c6128,s6133[1]};
    CLA_2 KS_6148(s6148, c6148, in6148_1, in6148_2);
    wire[0:0] s6149, in6149_1, in6149_2;
    wire c6149;
    assign in6149_1 = {s6129[0]};
    assign in6149_2 = {s6130[0]};
    Half_Adder KS_6149(s6149, c6149, in6149_1, in6149_2);
    wire[3:0] s6150, in6150_1, in6150_2;
    wire c6150;
    assign in6150_1 = {s6131[0],s6134[1],s6129[2],s5045[0]};
    assign in6150_2 = {s6132[0],s6135[1],s6130[2],s5046[0]};
    CLA_4 KS_6150(s6150, c6150, in6150_1, in6150_2);
    wire[0:0] s6151, in6151_1, in6151_2;
    wire c6151;
    assign in6151_1 = {s6134[0]};
    assign in6151_2 = {s6135[0]};
    Full_Adder KS_6151(s6151, c6151, in6151_1, in6151_2, s6133[0]);
    wire[3:0] s6152, in6152_1, in6152_2;
    wire c6152;
    assign in6152_1 = {s5021[1],pp122[95],pp117[101],c5025};
    assign in6152_2 = {s5022[1],pp123[94],pp118[100],c5026};
    CLA_4 KS_6152(s6152, c6152, in6152_1, in6152_2);
    wire[3:0] s6153, in6153_1, in6153_2;
    wire c6153;
    assign in6153_1 = {s5023[1],pp124[93],pp119[99],c5027};
    assign in6153_2 = {s5024[1],pp125[92],pp120[98],c5028};
    CLA_4 KS_6153(s6153, c6153, in6153_1, in6153_2);
    wire[3:0] s6154, in6154_1, in6154_2;
    wire c6154;
    assign in6154_1 = {s5025[1],pp126[91],pp121[97],c5032};
    assign in6154_2 = {s5026[1],pp127[90],pp122[96],c5040};
    CLA_4 KS_6154(s6154, c6154, in6154_1, in6154_2);
    wire[3:0] s6155, in6155_1, in6155_2;
    wire c6155;
    assign in6155_1 = {s5027[1],s5018[2],pp123[95],s5048[0]};
    assign in6155_2 = {s5028[1],s5019[2],pp124[94],s5049[0]};
    CLA_4 KS_6155(s6155, c6155, in6155_1, in6155_2);
    wire[3:0] s6156, in6156_1, in6156_2;
    wire c6156;
    assign in6156_1 = {s5029[1],s5020[2],pp125[93],s5050[0]};
    assign in6156_2 = {s5030[1],s5021[2],pp126[92],s5051[0]};
    CLA_4 KS_6156(s6156, c6156, in6156_1, in6156_2);
    wire[3:0] s6157, in6157_1, in6157_2;
    wire c6157;
    assign in6157_1 = {c5031,s5022[2],pp127[91],s5052[0]};
    assign in6157_2 = {s5032[1],s5023[2],s5018[3],s5053[0]};
    CLA_4 KS_6157(s6157, c6157, in6157_1, in6157_2);
    wire[3:0] s6158, in6158_1, in6158_2;
    wire c6158;
    assign in6158_1 = {c5033,s5024[2],s5019[3],s5054[0]};
    assign in6158_2 = {s5034[1],s5025[2],s5020[3],s5055[0]};
    CLA_4 KS_6158(s6158, c6158, in6158_1, in6158_2);
    wire[3:0] s6159, in6159_1, in6159_2;
    wire c6159;
    assign in6159_1 = {c5035,s5026[2],s5021[3],s5056[0]};
    assign in6159_2 = {s5036[1],s5027[2],s5022[3],s5057[0]};
    CLA_4 KS_6159(s6159, c6159, in6159_1, in6159_2);
    wire[3:0] s6160, in6160_1, in6160_2;
    wire c6160;
    assign in6160_1 = {c5037,s5028[2],s5023[3],s5058[0]};
    assign in6160_2 = {s5038[1],s5029[2],s5024[3],s5059[0]};
    CLA_4 KS_6160(s6160, c6160, in6160_1, in6160_2);
    wire[3:0] s6161, in6161_1, in6161_2;
    wire c6161;
    assign in6161_1 = {c5039,c5030,s5025[3],s5060[0]};
    assign in6161_2 = {s5040[1],s5032[2],s5026[3],s5061[0]};
    CLA_4 KS_6161(s6161, c6161, in6161_1, in6161_2);
    wire[3:0] s6162, in6162_1, in6162_2;
    wire c6162;
    assign in6162_1 = {c5041,c5034,s5027[3],s5062[0]};
    assign in6162_2 = {s5042[1],s5036[2],s5028[3],s5063[0]};
    CLA_4 KS_6162(s6162, c6162, in6162_1, in6162_2);
    wire[3:0] s6163, in6163_1, in6163_2;
    wire c6163;
    assign in6163_1 = {c5043,c5038,c5029,s5064[0]};
    assign in6163_2 = {s5044[1],s5040[2],s5032[3],s5065[0]};
    CLA_4 KS_6163(s6163, c6163, in6163_1, in6163_2);
    wire[0:0] s6164, in6164_1, in6164_2;
    wire c6164;
    assign in6164_1 = {c5045};
    assign in6164_2 = {s5046[1]};
    Half_Adder KS_6164(s6164, c6164, in6164_1, in6164_2);
    wire[1:0] s6165, in6165_1, in6165_2;
    wire c6165;
    assign in6165_1 = {c5047,c5042};
    assign in6165_2 = {c6129,s5044[2]};
    CLA_2 KS_6165(s6165, c6165, in6165_1, in6165_2);
    wire[0:0] s6166, in6166_1, in6166_2;
    wire c6166;
    assign in6166_1 = {c6130};
    assign in6166_2 = {c6131};
    Half_Adder KS_6166(s6166, c6166, in6166_1, in6166_2);
    wire[2:0] s6167, in6167_1, in6167_2;
    wire c6167;
    assign in6167_1 = {c6132,c5046,c5036};
    assign in6167_2 = {c6133,s6152[1],s5040[3]};
    CLA_3 KS_6167(s6167, c6167, in6167_1, in6167_2);
    wire[0:0] s6168, in6168_1, in6168_2;
    wire c6168;
    assign in6168_1 = {c6134};
    assign in6168_2 = {c6135};
    Half_Adder KS_6168(s6168, c6168, in6168_1, in6168_2);
    wire[1:0] s6169, in6169_1, in6169_2;
    wire c6169;
    assign in6169_1 = {c6136,s6153[1]};
    assign in6169_2 = {c6137,s6154[1]};
    CLA_2 KS_6169(s6169, c6169, in6169_1, in6169_2);
    wire[0:0] s6170, in6170_1, in6170_2;
    wire c6170;
    assign in6170_1 = {c6138};
    assign in6170_2 = {c6139};
    Half_Adder KS_6170(s6170, c6170, in6170_1, in6170_2);
    wire[3:0] s6171, in6171_1, in6171_2;
    wire c6171;
    assign in6171_1 = {c6142,s6155[1],c5044,s5066[0]};
    assign in6171_2 = {c6150,s6156[1],s6152[2],s5067[0]};
    CLA_4 KS_6171(s6171, c6171, in6171_1, in6171_2);
    wire[0:0] s6172, in6172_1, in6172_2;
    wire c6172;
    assign in6172_1 = {s6152[0]};
    assign in6172_2 = {s6153[0]};
    Half_Adder KS_6172(s6172, c6172, in6172_1, in6172_2);
    wire[1:0] s6173, in6173_1, in6173_2;
    wire c6173;
    assign in6173_1 = {s6154[0],s6157[1]};
    assign in6173_2 = {s6155[0],s6158[1]};
    CLA_2 KS_6173(s6173, c6173, in6173_1, in6173_2);
    wire[0:0] s6174, in6174_1, in6174_2;
    wire c6174;
    assign in6174_1 = {s6157[0]};
    assign in6174_2 = {s6158[0]};
    Full_Adder KS_6174(s6174, c6174, in6174_1, in6174_2, s6156[0]);
    wire[3:0] s6175, in6175_1, in6175_2;
    wire c6175;
    assign in6175_1 = {pp123[97],pp116[105],pp113[109],pp123[100]};
    assign in6175_2 = {pp124[96],pp117[104],pp114[108],pp124[99]};
    CLA_4 KS_6175(s6175, c6175, in6175_1, in6175_2);
    wire[3:0] s6176, in6176_1, in6176_2;
    wire c6176;
    assign in6176_1 = {pp125[95],pp118[103],pp115[107],pp125[98]};
    assign in6176_2 = {pp126[94],pp119[102],pp116[106],pp126[97]};
    CLA_4 KS_6176(s6176, c6176, in6176_1, in6176_2);
    wire[3:0] s6177, in6177_1, in6177_2;
    wire c6177;
    assign in6177_1 = {pp127[93],pp120[101],pp117[105],pp127[96]};
    assign in6177_2 = {s5048[1],pp121[100],pp118[104],c5048};
    CLA_4 KS_6177(s6177, c6177, in6177_1, in6177_2);
    wire[3:0] s6178, in6178_1, in6178_2;
    wire c6178;
    assign in6178_1 = {s5049[1],pp122[99],pp119[103],c5049};
    assign in6178_2 = {s5050[1],pp123[98],pp120[102],c5050};
    CLA_4 KS_6178(s6178, c6178, in6178_1, in6178_2);
    wire[3:0] s6179, in6179_1, in6179_2;
    wire c6179;
    assign in6179_1 = {s5051[1],pp124[97],pp121[101],c5051};
    assign in6179_2 = {s5052[1],pp125[96],pp122[100],c5052};
    CLA_4 KS_6179(s6179, c6179, in6179_1, in6179_2);
    wire[3:0] s6180, in6180_1, in6180_2;
    wire c6180;
    assign in6180_1 = {s5053[1],pp126[95],pp123[99],c5053};
    assign in6180_2 = {s5054[1],pp127[94],pp124[98],c5054};
    CLA_4 KS_6180(s6180, c6180, in6180_1, in6180_2);
    wire[3:0] s6181, in6181_1, in6181_2;
    wire c6181;
    assign in6181_1 = {s5055[1],s5048[2],pp125[97],c5058};
    assign in6181_2 = {s5056[1],s5049[2],pp126[96],c5066};
    CLA_4 KS_6181(s6181, c6181, in6181_1, in6181_2);
    wire[3:0] s6182, in6182_1, in6182_2;
    wire c6182;
    assign in6182_1 = {c5057,s5050[2],pp127[95],s5069[0]};
    assign in6182_2 = {s5058[1],s5051[2],s5048[3],s5070[0]};
    CLA_4 KS_6182(s6182, c6182, in6182_1, in6182_2);
    wire[3:0] s6183, in6183_1, in6183_2;
    wire c6183;
    assign in6183_1 = {c5059,s5052[2],s5049[3],s5071[0]};
    assign in6183_2 = {s5060[1],s5053[2],s5050[3],s5072[0]};
    CLA_4 KS_6183(s6183, c6183, in6183_1, in6183_2);
    wire[3:0] s6184, in6184_1, in6184_2;
    wire c6184;
    assign in6184_1 = {c5061,s5054[2],s5051[3],s5073[0]};
    assign in6184_2 = {s5062[1],s5055[2],s5052[3],s5074[0]};
    CLA_4 KS_6184(s6184, c6184, in6184_1, in6184_2);
    wire[3:0] s6185, in6185_1, in6185_2;
    wire c6185;
    assign in6185_1 = {c5063,c5056,s5053[3],s5075[0]};
    assign in6185_2 = {s5064[1],s5058[2],s5054[3],s5076[0]};
    CLA_4 KS_6185(s6185, c6185, in6185_1, in6185_2);
    wire[1:0] s6186, in6186_1, in6186_2;
    wire c6186;
    assign in6186_1 = {c5065,c5060};
    assign in6186_2 = {s5066[1],s5062[2]};
    CLA_2 KS_6186(s6186, c6186, in6186_1, in6186_2);
    wire[0:0] s6187, in6187_1, in6187_2;
    wire c6187;
    assign in6187_1 = {c5067};
    assign in6187_2 = {s5068[1]};
    Half_Adder KS_6187(s6187, c6187, in6187_1, in6187_2);
    wire[3:0] s6188, in6188_1, in6188_2;
    wire c6188;
    assign in6188_1 = {c6152,c5064,c5055,s5077[0]};
    assign in6188_2 = {c6153,s5066[2],s5058[3],s5078[0]};
    CLA_4 KS_6188(s6188, c6188, in6188_1, in6188_2);
    wire[0:0] s6189, in6189_1, in6189_2;
    wire c6189;
    assign in6189_1 = {c6154};
    assign in6189_2 = {c6155};
    Half_Adder KS_6189(s6189, c6189, in6189_1, in6189_2);
    wire[1:0] s6190, in6190_1, in6190_2;
    wire c6190;
    assign in6190_1 = {c6156,c5068};
    assign in6190_2 = {c6157,s6175[1]};
    CLA_2 KS_6190(s6190, c6190, in6190_1, in6190_2);
    wire[0:0] s6191, in6191_1, in6191_2;
    wire c6191;
    assign in6191_1 = {c6158};
    assign in6191_2 = {c6159};
    Half_Adder KS_6191(s6191, c6191, in6191_1, in6191_2);
    wire[2:0] s6192, in6192_1, in6192_2;
    wire c6192;
    assign in6192_1 = {c6160,s6176[1],c5062};
    assign in6192_2 = {c6161,s6177[1],s5066[3]};
    CLA_3 KS_6192(s6192, c6192, in6192_1, in6192_2);
    wire[0:0] s6193, in6193_1, in6193_2;
    wire c6193;
    assign in6193_1 = {c6162};
    assign in6193_2 = {c6163};
    Half_Adder KS_6193(s6193, c6193, in6193_1, in6193_2);
    wire[1:0] s6194, in6194_1, in6194_2;
    wire c6194;
    assign in6194_1 = {c6171,s6178[1]};
    assign in6194_2 = {s6175[0],s6179[1]};
    CLA_2 KS_6194(s6194, c6194, in6194_1, in6194_2);
    wire[0:0] s6195, in6195_1, in6195_2;
    wire c6195;
    assign in6195_1 = {s6176[0]};
    assign in6195_2 = {s6177[0]};
    Half_Adder KS_6195(s6195, c6195, in6195_1, in6195_2);
    wire[3:0] s6196, in6196_1, in6196_2;
    wire c6196;
    assign in6196_1 = {s6179[0],s6180[1],s6175[2],s5079[0]};
    assign in6196_2 = {s6180[0],s6181[1],s6176[2],s5080[0]};
    CLA_4_c KS_6196(s6196, c6196, in6196_1, in6196_2, s6178[0]);
    wire[3:0] s6197, in6197_1, in6197_2;
    wire c6197;
    assign in6197_1 = {pp115[109],pp110[115],pp107[119],pp109[118]};
    assign in6197_2 = {pp116[108],pp111[114],pp108[118],pp110[117]};
    CLA_4 KS_6197(s6197, c6197, in6197_1, in6197_2);
    wire[3:0] s6198, in6198_1, in6198_2;
    wire c6198;
    assign in6198_1 = {pp117[107],pp112[113],pp109[117],pp111[116]};
    assign in6198_2 = {pp118[106],pp113[112],pp110[116],pp112[115]};
    CLA_4 KS_6198(s6198, c6198, in6198_1, in6198_2);
    wire[3:0] s6199, in6199_1, in6199_2;
    wire c6199;
    assign in6199_1 = {pp119[105],pp114[111],pp111[115],pp113[114]};
    assign in6199_2 = {pp120[104],pp115[110],pp112[114],pp114[113]};
    CLA_4 KS_6199(s6199, c6199, in6199_1, in6199_2);
    wire[3:0] s6200, in6200_1, in6200_2;
    wire c6200;
    assign in6200_1 = {pp121[103],pp116[109],pp113[113],pp115[112]};
    assign in6200_2 = {pp122[102],pp117[108],pp114[112],pp116[111]};
    CLA_4 KS_6200(s6200, c6200, in6200_1, in6200_2);
    wire[3:0] s6201, in6201_1, in6201_2;
    wire c6201;
    assign in6201_1 = {pp123[101],pp118[107],pp115[111],pp117[110]};
    assign in6201_2 = {pp124[100],pp119[106],pp116[110],pp118[109]};
    CLA_4 KS_6201(s6201, c6201, in6201_1, in6201_2);
    wire[3:0] s6202, in6202_1, in6202_2;
    wire c6202;
    assign in6202_1 = {pp125[99],pp120[105],pp117[109],pp119[108]};
    assign in6202_2 = {pp126[98],pp121[104],pp118[108],pp120[107]};
    CLA_4 KS_6202(s6202, c6202, in6202_1, in6202_2);
    wire[3:0] s6203, in6203_1, in6203_2;
    wire c6203;
    assign in6203_1 = {pp127[97],pp122[103],pp119[107],pp121[106]};
    assign in6203_2 = {s5069[1],pp123[102],pp120[106],pp122[105]};
    CLA_4 KS_6203(s6203, c6203, in6203_1, in6203_2);
    wire[3:0] s6204, in6204_1, in6204_2;
    wire c6204;
    assign in6204_1 = {s5070[1],pp124[101],pp121[105],pp123[104]};
    assign in6204_2 = {s5071[1],pp125[100],pp122[104],pp124[103]};
    CLA_4 KS_6204(s6204, c6204, in6204_1, in6204_2);
    wire[3:0] s6205, in6205_1, in6205_2;
    wire c6205;
    assign in6205_1 = {s5072[1],pp126[99],pp123[103],pp125[102]};
    assign in6205_2 = {s5073[1],pp127[98],pp124[102],pp126[101]};
    CLA_4 KS_6205(s6205, c6205, in6205_1, in6205_2);
    wire[3:0] s6206, in6206_1, in6206_2;
    wire c6206;
    assign in6206_1 = {c5074,s5069[2],pp125[101],pp127[100]};
    assign in6206_2 = {s5075[1],s5070[2],pp126[100],c5069};
    CLA_4 KS_6206(s6206, c6206, in6206_1, in6206_2);
    wire[3:0] s6207, in6207_1, in6207_2;
    wire c6207;
    assign in6207_1 = {c5076,s5071[2],pp127[99],c5070};
    assign in6207_2 = {s5077[1],s5072[2],s5069[3],c5071};
    CLA_4 KS_6207(s6207, c6207, in6207_1, in6207_2);
    wire[3:0] s6208, in6208_1, in6208_2;
    wire c6208;
    assign in6208_1 = {c5078,c5073,s5070[3],c5075};
    assign in6208_2 = {s5079[1],s5075[2],s5071[3],s5082[0]};
    CLA_4 KS_6208(s6208, c6208, in6208_1, in6208_2);
    wire[0:0] s6209, in6209_1, in6209_2;
    wire c6209;
    assign in6209_1 = {c5080};
    assign in6209_2 = {s5081[1]};
    Half_Adder KS_6209(s6209, c6209, in6209_1, in6209_2);
    wire[1:0] s6210, in6210_1, in6210_2;
    wire c6210;
    assign in6210_1 = {c6175,c5077};
    assign in6210_2 = {c6176,s5079[2]};
    CLA_2 KS_6210(s6210, c6210, in6210_1, in6210_2);
    wire[0:0] s6211, in6211_1, in6211_2;
    wire c6211;
    assign in6211_1 = {c6177};
    assign in6211_2 = {c6178};
    Half_Adder KS_6211(s6211, c6211, in6211_1, in6211_2);
    wire[2:0] s6212, in6212_1, in6212_2;
    wire c6212;
    assign in6212_1 = {c6179,c5081,c5072};
    assign in6212_2 = {c6180,s6197[1],s5075[3]};
    CLA_3 KS_6212(s6212, c6212, in6212_1, in6212_2);
    wire[0:0] s6213, in6213_1, in6213_2;
    wire c6213;
    assign in6213_1 = {c6181};
    assign in6213_2 = {c6182};
    Half_Adder KS_6213(s6213, c6213, in6213_1, in6213_2);
    wire[1:0] s6214, in6214_1, in6214_2;
    wire c6214;
    assign in6214_1 = {c6183,s6198[1]};
    assign in6214_2 = {c6184,s6199[1]};
    CLA_2 KS_6214(s6214, c6214, in6214_1, in6214_2);
    wire[0:0] s6215, in6215_1, in6215_2;
    wire c6215;
    assign in6215_1 = {c6185};
    assign in6215_2 = {c6188};
    Half_Adder KS_6215(s6215, c6215, in6215_1, in6215_2);
    wire[3:0] s6216, in6216_1, in6216_2;
    wire c6216;
    assign in6216_1 = {c6196,s6200[1],c5079,s5083[0]};
    assign in6216_2 = {s6197[0],s6201[1],s6197[2],s5084[0]};
    CLA_4 KS_6216(s6216, c6216, in6216_1, in6216_2);
    wire[0:0] s6217, in6217_1, in6217_2;
    wire c6217;
    assign in6217_1 = {s6198[0]};
    assign in6217_2 = {s6199[0]};
    Half_Adder KS_6217(s6217, c6217, in6217_1, in6217_2);
    wire[1:0] s6218, in6218_1, in6218_2;
    wire c6218;
    assign in6218_1 = {s6201[0],s6202[1]};
    assign in6218_2 = {s6202[0],s6203[1]};
    CLA_2_c KS_6218(s6218, c6218, in6218_1, in6218_2, s6200[0]);
    wire[3:0] s6219, in6219_1, in6219_2;
    wire c6219;
    assign in6219_1 = {pp105[123],pp104[125],pp103[127],pp104[127]};
    assign in6219_2 = {pp106[122],pp105[124],pp104[126],pp105[126]};
    CLA_4 KS_6219(s6219, c6219, in6219_1, in6219_2);
    wire[3:0] s6220, in6220_1, in6220_2;
    wire c6220;
    assign in6220_1 = {pp107[121],pp106[123],pp105[125],pp106[125]};
    assign in6220_2 = {pp108[120],pp107[122],pp106[124],pp107[124]};
    CLA_4 KS_6220(s6220, c6220, in6220_1, in6220_2);
    wire[3:0] s6221, in6221_1, in6221_2;
    wire c6221;
    assign in6221_1 = {pp109[119],pp108[121],pp107[123],pp108[123]};
    assign in6221_2 = {pp110[118],pp109[120],pp108[122],pp109[122]};
    CLA_4 KS_6221(s6221, c6221, in6221_1, in6221_2);
    wire[3:0] s6222, in6222_1, in6222_2;
    wire c6222;
    assign in6222_1 = {pp111[117],pp110[119],pp109[121],pp110[121]};
    assign in6222_2 = {pp112[116],pp111[118],pp110[120],pp111[120]};
    CLA_4 KS_6222(s6222, c6222, in6222_1, in6222_2);
    wire[3:0] s6223, in6223_1, in6223_2;
    wire c6223;
    assign in6223_1 = {pp113[115],pp112[117],pp111[119],pp112[119]};
    assign in6223_2 = {pp114[114],pp113[116],pp112[118],pp113[118]};
    CLA_4 KS_6223(s6223, c6223, in6223_1, in6223_2);
    wire[3:0] s6224, in6224_1, in6224_2;
    wire c6224;
    assign in6224_1 = {pp115[113],pp114[115],pp113[117],pp114[117]};
    assign in6224_2 = {pp116[112],pp115[114],pp114[116],pp115[116]};
    CLA_4 KS_6224(s6224, c6224, in6224_1, in6224_2);
    wire[3:0] s6225, in6225_1, in6225_2;
    wire c6225;
    assign in6225_1 = {pp117[111],pp116[113],pp115[115],pp116[115]};
    assign in6225_2 = {pp118[110],pp117[112],pp116[114],pp117[114]};
    CLA_4 KS_6225(s6225, c6225, in6225_1, in6225_2);
    wire[3:0] s6226, in6226_1, in6226_2;
    wire c6226;
    assign in6226_1 = {pp119[109],pp118[111],pp117[113],pp118[113]};
    assign in6226_2 = {pp120[108],pp119[110],pp118[112],pp119[112]};
    CLA_4 KS_6226(s6226, c6226, in6226_1, in6226_2);
    wire[3:0] s6227, in6227_1, in6227_2;
    wire c6227;
    assign in6227_1 = {pp121[107],pp120[109],pp119[111],pp120[111]};
    assign in6227_2 = {pp122[106],pp121[108],pp120[110],pp121[110]};
    CLA_4 KS_6227(s6227, c6227, in6227_1, in6227_2);
    wire[2:0] s6228, in6228_1, in6228_2;
    wire c6228;
    assign in6228_1 = {pp123[105],pp122[107],pp121[109]};
    assign in6228_2 = {pp124[104],pp123[106],pp122[108]};
    CLA_3 KS_6228(s6228, c6228, in6228_1, in6228_2);
    wire[3:0] s6229, in6229_1, in6229_2;
    wire c6229;
    assign in6229_1 = {pp125[103],pp124[105],pp123[107],pp122[109]};
    assign in6229_2 = {pp126[102],pp125[104],pp124[106],pp123[108]};
    CLA_4 KS_6229(s6229, c6229, in6229_1, in6229_2);
    wire[0:0] s6230, in6230_1, in6230_2;
    wire c6230;
    assign in6230_1 = {pp127[101]};
    assign in6230_2 = {s5082[1]};
    Half_Adder KS_6230(s6230, c6230, in6230_1, in6230_2);
    wire[1:0] s6231, in6231_1, in6231_2;
    wire c6231;
    assign in6231_1 = {c5083,pp126[103]};
    assign in6231_2 = {s5084[1],pp127[102]};
    CLA_2 KS_6231(s6231, c6231, in6231_1, in6231_2);
    wire[0:0] s6232, in6232_1, in6232_2;
    wire c6232;
    assign in6232_1 = {c5085};
    assign in6232_2 = {c6197};
    Half_Adder KS_6232(s6232, c6232, in6232_1, in6232_2);
    wire[2:0] s6233, in6233_1, in6233_2;
    wire c6233;
    assign in6233_1 = {c6198,c5082,pp125[105]};
    assign in6233_2 = {c6199,s5084[2],pp126[104]};
    CLA_3 KS_6233(s6233, c6233, in6233_1, in6233_2);
    wire[0:0] s6234, in6234_1, in6234_2;
    wire c6234;
    assign in6234_1 = {c6200};
    assign in6234_2 = {c6201};
    Half_Adder KS_6234(s6234, c6234, in6234_1, in6234_2);
    wire[1:0] s6235, in6235_1, in6235_2;
    wire c6235;
    assign in6235_1 = {c6202,s6219[1]};
    assign in6235_2 = {c6203,s6220[1]};
    CLA_2 KS_6235(s6235, c6235, in6235_1, in6235_2);
    wire[0:0] s6236, in6236_1, in6236_2;
    wire c6236;
    assign in6236_1 = {c6204};
    assign in6236_2 = {c6205};
    Half_Adder KS_6236(s6236, c6236, in6236_1, in6236_2);
    wire[3:0] s6237, in6237_1, in6237_2;
    wire c6237;
    assign in6237_1 = {c6206,s6221[1],pp127[103],pp124[107]};
    assign in6237_2 = {c6207,s6222[1],c5084,pp125[106]};
    CLA_4 KS_6237(s6237, c6237, in6237_1, in6237_2);
    wire[0:0] s6238, in6238_1, in6238_2;
    wire c6238;
    assign in6238_1 = {c6208};
    assign in6238_2 = {c6216};
    Half_Adder KS_6238(s6238, c6238, in6238_1, in6238_2);
    wire[1:0] s6239, in6239_1, in6239_2;
    wire c6239;
    assign in6239_1 = {s6219[0],s6223[1]};
    assign in6239_2 = {s6220[0],s6224[1]};
    CLA_2 KS_6239(s6239, c6239, in6239_1, in6239_2);
    wire[0:0] s6240, in6240_1, in6240_2;
    wire c6240;
    assign in6240_1 = {s6221[0]};
    assign in6240_2 = {s6222[0]};
    Half_Adder KS_6240(s6240, c6240, in6240_1, in6240_2);
    wire[2:0] s6241, in6241_1, in6241_2;
    wire c6241;
    assign in6241_1 = {s6224[0],s6225[1],s6219[2]};
    assign in6241_2 = {s6225[0],s6226[1],s6220[2]};
    CLA_3_c KS_6241(s6241, c6241, in6241_1, in6241_2, s6223[0]);
    wire[3:0] s6242, in6242_1, in6242_2;
    wire c6242;
    assign in6242_1 = {pp105[127],pp106[127],pp107[127],pp108[127]};
    assign in6242_2 = {pp106[126],pp107[126],pp108[126],pp109[126]};
    CLA_4 KS_6242(s6242, c6242, in6242_1, in6242_2);
    wire[3:0] s6243, in6243_1, in6243_2;
    wire c6243;
    assign in6243_1 = {pp107[125],pp108[125],pp109[125],pp110[125]};
    assign in6243_2 = {pp108[124],pp109[124],pp110[124],pp111[124]};
    CLA_4 KS_6243(s6243, c6243, in6243_1, in6243_2);
    wire[3:0] s6244, in6244_1, in6244_2;
    wire c6244;
    assign in6244_1 = {pp109[123],pp110[123],pp111[123],pp112[123]};
    assign in6244_2 = {pp110[122],pp111[122],pp112[122],pp113[122]};
    CLA_4 KS_6244(s6244, c6244, in6244_1, in6244_2);
    wire[3:0] s6245, in6245_1, in6245_2;
    wire c6245;
    assign in6245_1 = {pp111[121],pp112[121],pp113[121],pp114[121]};
    assign in6245_2 = {pp112[120],pp113[120],pp114[120],pp115[120]};
    CLA_4 KS_6245(s6245, c6245, in6245_1, in6245_2);
    wire[3:0] s6246, in6246_1, in6246_2;
    wire c6246;
    assign in6246_1 = {pp113[119],pp114[119],pp115[119],pp116[119]};
    assign in6246_2 = {pp114[118],pp115[118],pp116[118],pp117[118]};
    CLA_4 KS_6246(s6246, c6246, in6246_1, in6246_2);
    wire[2:0] s6247, in6247_1, in6247_2;
    wire c6247;
    assign in6247_1 = {pp115[117],pp116[117],pp117[117]};
    assign in6247_2 = {pp116[116],pp117[116],pp118[116]};
    CLA_3 KS_6247(s6247, c6247, in6247_1, in6247_2);
    wire[1:0] s6248, in6248_1, in6248_2;
    wire c6248;
    assign in6248_1 = {pp117[115],pp118[115]};
    assign in6248_2 = {pp118[114],pp119[114]};
    CLA_2 KS_6248(s6248, c6248, in6248_1, in6248_2);
    wire[0:0] s6249, in6249_1, in6249_2;
    wire c6249;
    assign in6249_1 = {pp119[113]};
    assign in6249_2 = {pp120[112]};
    Half_Adder KS_6249(s6249, c6249, in6249_1, in6249_2);
    wire[3:0] s6250, in6250_1, in6250_2;
    wire c6250;
    assign in6250_1 = {pp121[111],pp120[113],pp119[115],pp118[117]};
    assign in6250_2 = {pp122[110],pp121[112],pp120[114],pp119[116]};
    CLA_4 KS_6250(s6250, c6250, in6250_1, in6250_2);
    wire[0:0] s6251, in6251_1, in6251_2;
    wire c6251;
    assign in6251_1 = {pp123[109]};
    assign in6251_2 = {pp124[108]};
    Half_Adder KS_6251(s6251, c6251, in6251_1, in6251_2);
    wire[1:0] s6252, in6252_1, in6252_2;
    wire c6252;
    assign in6252_1 = {pp125[107],pp122[111]};
    assign in6252_2 = {pp126[106],pp123[110]};
    CLA_2 KS_6252(s6252, c6252, in6252_1, in6252_2);
    wire[0:0] s6253, in6253_1, in6253_2;
    wire c6253;
    assign in6253_1 = {pp127[105]};
    assign in6253_2 = {c6219};
    Half_Adder KS_6253(s6253, c6253, in6253_1, in6253_2);
    wire[2:0] s6254, in6254_1, in6254_2;
    wire c6254;
    assign in6254_1 = {c6220,pp124[109],pp121[113]};
    assign in6254_2 = {c6221,pp125[108],pp122[112]};
    CLA_3 KS_6254(s6254, c6254, in6254_1, in6254_2);
    wire[0:0] s6255, in6255_1, in6255_2;
    wire c6255;
    assign in6255_1 = {c6222};
    assign in6255_2 = {c6223};
    Half_Adder KS_6255(s6255, c6255, in6255_1, in6255_2);
    wire[1:0] s6256, in6256_1, in6256_2;
    wire c6256;
    assign in6256_1 = {c6224,pp126[107]};
    assign in6256_2 = {c6225,pp127[106]};
    CLA_2 KS_6256(s6256, c6256, in6256_1, in6256_2);
    wire[0:0] s6257, in6257_1, in6257_2;
    wire c6257;
    assign in6257_1 = {c6226};
    assign in6257_2 = {c6227};
    Half_Adder KS_6257(s6257, c6257, in6257_1, in6257_2);
    wire[3:0] s6258, in6258_1, in6258_2;
    wire c6258;
    assign in6258_1 = {c6237,s6242[1],pp123[111],pp120[115]};
    assign in6258_2 = {s6242[0],s6243[1],pp124[110],pp121[114]};
    CLA_4_c KS_6258(s6258, c6258, in6258_1, in6258_2, c6229);
    wire[3:0] s6259, in6259_1, in6259_2;
    wire c6259;
    assign in6259_1 = {pp109[127],pp110[127],pp111[127],pp112[127]};
    assign in6259_2 = {pp110[126],pp111[126],pp112[126],pp113[126]};
    CLA_4 KS_6259(s6259, c6259, in6259_1, in6259_2);
    wire[2:0] s6260, in6260_1, in6260_2;
    wire c6260;
    assign in6260_1 = {pp111[125],pp112[125],pp113[125]};
    assign in6260_2 = {pp112[124],pp113[124],pp114[124]};
    CLA_3 KS_6260(s6260, c6260, in6260_1, in6260_2);
    wire[1:0] s6261, in6261_1, in6261_2;
    wire c6261;
    assign in6261_1 = {pp113[123],pp114[123]};
    assign in6261_2 = {pp114[122],pp115[122]};
    CLA_2 KS_6261(s6261, c6261, in6261_1, in6261_2);
    wire[0:0] s6262, in6262_1, in6262_2;
    wire c6262;
    assign in6262_1 = {pp115[121]};
    assign in6262_2 = {pp116[120]};
    Half_Adder KS_6262(s6262, c6262, in6262_1, in6262_2);
    wire[3:0] s6263, in6263_1, in6263_2;
    wire c6263;
    assign in6263_1 = {pp117[119],pp116[121],pp115[123],pp114[125]};
    assign in6263_2 = {pp118[118],pp117[120],pp116[122],pp115[124]};
    CLA_4 KS_6263(s6263, c6263, in6263_1, in6263_2);
    wire[0:0] s6264, in6264_1, in6264_2;
    wire c6264;
    assign in6264_1 = {pp119[117]};
    assign in6264_2 = {pp120[116]};
    Half_Adder KS_6264(s6264, c6264, in6264_1, in6264_2);
    wire[1:0] s6265, in6265_1, in6265_2;
    wire c6265;
    assign in6265_1 = {pp121[115],pp118[119]};
    assign in6265_2 = {pp122[114],pp119[118]};
    CLA_2 KS_6265(s6265, c6265, in6265_1, in6265_2);
    wire[0:0] s6266, in6266_1, in6266_2;
    wire c6266;
    assign in6266_1 = {pp123[113]};
    assign in6266_2 = {pp124[112]};
    Half_Adder KS_6266(s6266, c6266, in6266_1, in6266_2);
    wire[2:0] s6267, in6267_1, in6267_2;
    wire c6267;
    assign in6267_1 = {pp126[110],pp120[117],pp117[121]};
    assign in6267_2 = {pp127[109],pp121[116],pp118[120]};
    CLA_3_c KS_6267(s6267, c6267, in6267_1, in6267_2, pp125[111]);
    wire[0:0] s6268, in6268_1, in6268_2;
    wire c6268;
    assign in6268_1 = {pp113[127]};
    assign in6268_2 = {pp114[126]};
    Half_Adder KS_6268(s6268, c6268, in6268_1, in6268_2);

    /*Stage 5*/
    wire[3:0] s6269, in6269_1, in6269_2;
    wire c6269;
    assign in6269_1 = {pp0[10],pp0[11],pp0[12],pp0[13]};
    assign in6269_2 = {pp1[9],pp1[10],pp1[11],pp1[12]};
    CLA_4 KS_6269(s6269, c6269, in6269_1, in6269_2);
    wire[3:0] s6270, in6270_1, in6270_2;
    wire c6270;
    assign in6270_1 = {pp2[9],pp2[10],pp2[11],pp0[14]};
    assign in6270_2 = {pp3[8],pp3[9],pp3[10],pp1[13]};
    CLA_4 KS_6270(s6270, c6270, in6270_1, in6270_2);
    wire[3:0] s6271, in6271_1, in6271_2;
    wire c6271;
    assign in6271_1 = {pp4[8],pp4[9],pp2[12],pp0[15]};
    assign in6271_2 = {pp5[7],pp5[8],pp3[11],pp1[14]};
    CLA_4 KS_6271(s6271, c6271, in6271_1, in6271_2);
    wire[3:0] s6272, in6272_1, in6272_2;
    wire c6272;
    assign in6272_1 = {pp6[7],pp4[10],pp2[13],pp2[14]};
    assign in6272_2 = {pp7[6],pp5[9],pp3[12],pp3[13]};
    CLA_4 KS_6272(s6272, c6272, in6272_1, in6272_2);
    wire[3:0] s6273, in6273_1, in6273_2;
    wire c6273;
    assign in6273_1 = {pp6[8],pp4[11],pp4[12],pp4[13]};
    assign in6273_2 = {pp7[7],pp5[10],pp5[11],pp5[12]};
    CLA_4 KS_6273(s6273, c6273, in6273_1, in6273_2);
    wire[3:0] s6274, in6274_1, in6274_2;
    wire c6274;
    assign in6274_1 = {pp9[5],pp6[9],pp6[10],pp6[11]};
    assign in6274_2 = {pp10[4],pp7[8],pp7[9],pp7[10]};
    CLA_4_c KS_6274(s6274, c6274, in6274_1, in6274_2, pp8[6]);
    wire[3:0] s6275, in6275_1, in6275_2;
    wire c6275;
    assign in6275_1 = {pp8[7],pp8[8],pp8[9],pp6[12]};
    assign in6275_2 = {pp9[6],pp9[7],pp9[8],pp7[11]};
    CLA_4 KS_6275(s6275, c6275, in6275_1, in6275_2);
    wire[3:0] s6276, in6276_1, in6276_2;
    wire c6276;
    assign in6276_1 = {pp11[4],pp10[6],pp10[7],pp8[10]};
    assign in6276_2 = {pp12[3],pp11[5],pp11[6],pp9[9]};
    CLA_4_c KS_6276(s6276, c6276, in6276_1, in6276_2, pp10[5]);
    wire[3:0] s6277, in6277_1, in6277_2;
    wire c6277;
    assign in6277_1 = {pp13[3],pp12[5],pp10[8],pp8[11]};
    assign in6277_2 = {pp14[2],pp13[4],pp11[7],pp9[10]};
    CLA_4_c KS_6277(s6277, c6277, in6277_1, in6277_2, pp12[4]);
    wire[3:0] s6278, in6278_1, in6278_2;
    wire c6278;
    assign in6278_1 = {pp15[2],pp12[6],pp10[9],pp11[9]};
    assign in6278_2 = {pp16[1],pp13[5],pp11[8],pp12[8]};
    CLA_4_c KS_6278(s6278, c6278, in6278_1, in6278_2, pp14[3]);
    wire[3:0] s6279, in6279_1, in6279_2;
    wire c6279;
    assign in6279_1 = {pp14[4],pp12[7],pp13[7],pp13[8]};
    assign in6279_2 = {pp15[3],pp13[6],pp14[6],pp14[7]};
    CLA_4 KS_6279(s6279, c6279, in6279_1, in6279_2);
    wire[3:0] s6280, in6280_1, in6280_2;
    wire c6280;
    assign in6280_1 = {pp16[2],pp14[5],pp15[5],pp15[6]};
    assign in6280_2 = {pp17[1],pp15[4],pp16[4],pp16[5]};
    CLA_4 KS_6280(s6280, c6280, in6280_1, in6280_2);
    wire[3:0] s6281, in6281_1, in6281_2;
    wire c6281;
    assign in6281_1 = {s5086[2],pp16[3],pp17[3],pp17[4]};
    assign in6281_2 = {s5087[1],pp17[2],pp18[2],pp18[3]};
    CLA_4_c KS_6281(s6281, c6281, in6281_1, in6281_2, pp18[0]);
    wire[3:0] s6282, in6282_1, in6282_2;
    wire c6282;
    assign in6282_1 = {pp18[1],pp19[1],pp19[2],pp15[7]};
    assign in6282_2 = {pp19[0],pp20[0],pp20[1],pp16[6]};
    CLA_4 KS_6282(s6282, c6282, in6282_1, in6282_2);
    wire[3:0] s6283, in6283_1, in6283_2;
    wire c6283;
    assign in6283_1 = {s5087[2],c5086,pp21[0],pp17[5]};
    assign in6283_2 = {s5088[1],s5087[3],c5087,pp18[4]};
    CLA_4_c KS_6283(s6283, c6283, in6283_1, in6283_2, s5086[3]);
    wire[3:0] s6284, in6284_1, in6284_2;
    wire c6284;
    assign in6284_1 = {s5088[2],s5088[3],pp19[3],pp17[6]};
    assign in6284_2 = {s5089[1],s5089[2],pp20[2],pp18[5]};
    CLA_4 KS_6284(s6284, c6284, in6284_1, in6284_2);
    wire[3:0] s6285, in6285_1, in6285_2;
    wire c6285;
    assign in6285_1 = {s5090[1],pp21[1],pp19[4],pp21[3]};
    assign in6285_2 = {s5091[1],pp22[0],pp20[3],pp22[2]};
    CLA_4 KS_6285(s6285, c6285, in6285_1, in6285_2);
    wire[3:0] s6286, in6286_1, in6286_2;
    wire c6286;
    assign in6286_1 = {c5088,pp21[2],pp23[1],pp23[2]};
    assign in6286_2 = {s5089[3],pp22[1],pp24[0],pp24[1]};
    CLA_4 KS_6286(s6286, c6286, in6286_1, in6286_2);
    wire[3:0] s6287, in6287_1, in6287_2;
    wire c6287;
    assign in6287_1 = {s5090[2],pp23[0],c5090,pp25[0]};
    assign in6287_2 = {s5091[2],c5089,c5091,c5092};
    CLA_4 KS_6287(s6287, c6287, in6287_1, in6287_2);
    wire[3:0] s6288, in6288_1, in6288_2;
    wire c6288;
    assign in6288_1 = {s5092[1],s5090[3],s5092[3],c5093};
    assign in6288_2 = {s5093[1],s5091[3],s5093[3],s5094[3]};
    CLA_4 KS_6288(s6288, c6288, in6288_1, in6288_2);
    wire[3:0] s6289, in6289_1, in6289_2;
    wire c6289;
    assign in6289_1 = {s5095[0],s5092[2],s5094[2],s5095[3]};
    assign in6289_2 = {c6279,s5093[2],s5095[2],s5096[2]};
    CLA_4_c KS_6289(s6289, c6289, in6289_1, in6289_2, s5094[0]);
    wire[3:0] s6290, in6290_1, in6290_2;
    wire c6290;
    assign in6290_1 = {s5095[1],s5096[1],s5097[2],pp25[1]};
    assign in6290_2 = {s5096[0],s5097[1],s5098[1],pp26[0]};
    CLA_4_c KS_6290(s6290, c6290, in6290_1, in6290_2, s5094[1]);
    wire[3:0] s6291, in6291_1, in6291_2;
    wire c6291;
    assign in6291_1 = {s5098[0],s5099[1],c5094,pp27[0]};
    assign in6291_2 = {s5099[0],s5100[1],c5095,s3430[0]};
    CLA_4 KS_6291(s6291, c6291, in6291_1, in6291_2);
    wire[3:0] s6292, in6292_1, in6292_2;
    wire c6292;
    assign in6292_1 = {s5101[1],s5096[3],c5096,c5100};
    assign in6292_2 = {s5102[0],s5097[3],c5097,c5101};
    CLA_4 KS_6292(s6292, c6292, in6292_1, in6292_2);
    wire[3:0] s6293, in6293_1, in6293_2;
    wire c6293;
    assign in6293_1 = {s5098[2],s5098[3],s5102[3],c5102};
    assign in6293_2 = {s5099[2],s5099[3],s5103[3],c5103};
    CLA_4 KS_6293(s6293, c6293, in6293_1, in6293_2);
    wire[3:0] s6294, in6294_1, in6294_2;
    wire c6294;
    assign in6294_1 = {s5100[2],s5100[3],s5104[3],c5104};
    assign in6294_2 = {s5101[2],s5101[3],s5105[2],s5105[3]};
    CLA_4 KS_6294(s6294, c6294, in6294_1, in6294_2);
    wire[3:0] s6295, in6295_1, in6295_2;
    wire c6295;
    assign in6295_1 = {s5102[1],s5102[2],s5106[2],s5106[3]};
    assign in6295_2 = {s5103[1],s5103[2],s5107[2],s5107[3]};
    CLA_4 KS_6295(s6295, c6295, in6295_1, in6295_2);
    wire[3:0] s6296, in6296_1, in6296_2;
    wire c6296;
    assign in6296_1 = {s5104[1],s5104[2],s5108[1],s5108[2]};
    assign in6296_2 = {s5105[0],s5105[1],s5109[1],s5109[2]};
    CLA_4 KS_6296(s6296, c6296, in6296_1, in6296_2);
    wire[3:0] s6297, in6297_1, in6297_2;
    wire c6297;
    assign in6297_1 = {s5106[0],s5106[1],s5110[0],s5110[1]};
    assign in6297_2 = {s5107[0],s5107[1],s5111[0],s5111[1]};
    CLA_4 KS_6297(s6297, c6297, in6297_1, in6297_2);
    wire[3:0] s6298, in6298_1, in6298_2;
    wire c6298;
    assign in6298_1 = {c6287,s5108[0],s5112[0],s5112[1]};
    assign in6298_2 = {c6288,s5109[0],s5113[0],s5113[1]};
    CLA_4_c KS_6298(s6298, c6298, in6298_1, in6298_2, c6286);
    wire[3:0] s6299, in6299_1, in6299_2;
    wire c6299;
    assign in6299_1 = {s5114[1],c5105,s3434[0],s5116[3]};
    assign in6299_2 = {s5115[1],c5106,s3435[0],s5117[3]};
    CLA_4 KS_6299(s6299, c6299, in6299_1, in6299_2);
    wire[3:0] s6300, in6300_1, in6300_2;
    wire c6300;
    assign in6300_1 = {c5107,c5108,s5118[2],c5117};
    assign in6300_2 = {s5108[3],c5109,s5119[2],s5118[3]};
    CLA_4 KS_6300(s6300, c6300, in6300_1, in6300_2);
    wire[3:0] s6301, in6301_1, in6301_2;
    wire c6301;
    assign in6301_1 = {s5109[3],s5110[3],s5120[2],s5119[3]};
    assign in6301_2 = {s5110[2],s5111[3],s5121[1],s5120[3]};
    CLA_4 KS_6301(s6301, c6301, in6301_1, in6301_2);
    wire[3:0] s6302, in6302_1, in6302_2;
    wire c6302;
    assign in6302_1 = {s5111[2],s5112[3],s5122[0],s5121[2]};
    assign in6302_2 = {s5112[2],s5113[3],s5123[0],s5122[1]};
    CLA_4 KS_6302(s6302, c6302, in6302_1, in6302_2);
    wire[3:0] s6303, in6303_1, in6303_2;
    wire c6303;
    assign in6303_1 = {s5113[2],s5114[3],s5124[0],s5123[1]};
    assign in6303_2 = {s5114[2],s5115[3],s5125[0],s5124[1]};
    CLA_4 KS_6303(s6303, c6303, in6303_1, in6303_2);
    wire[3:0] s6304, in6304_1, in6304_2;
    wire c6304;
    assign in6304_1 = {s5115[2],s5116[2],s5126[0],s5125[1]};
    assign in6304_2 = {s5116[1],s5117[2],s5127[0],s5126[1]};
    CLA_4 KS_6304(s6304, c6304, in6304_1, in6304_2);
    wire[3:0] s6305, in6305_1, in6305_2;
    wire c6305;
    assign in6305_1 = {s5117[1],s5118[1],s5128[0],s5127[1]};
    assign in6305_2 = {s5118[0],s5119[1],s5129[0],s5128[1]};
    CLA_4 KS_6305(s6305, c6305, in6305_1, in6305_2);
    wire[0:0] s6306, in6306_1, in6306_2;
    wire c6306;
    assign in6306_1 = {s5119[0]};
    assign in6306_2 = {s5120[0]};
    Half_Adder KS_6306(s6306, c6306, in6306_1, in6306_2);
    wire[1:0] s6307, in6307_1, in6307_2;
    wire c6307;
    assign in6307_1 = {c6293,s5120[1]};
    assign in6307_2 = {c6294,s5121[0]};
    CLA_2 KS_6307(s6307, c6307, in6307_1, in6307_2);
    wire[0:0] s6308, in6308_1, in6308_2;
    wire c6308;
    assign in6308_1 = {c6295};
    assign in6308_2 = {c6296};
    Half_Adder KS_6308(s6308, c6308, in6308_1, in6308_2);
    wire[3:0] s6309, in6309_1, in6309_2;
    wire c6309;
    assign in6309_1 = {c6298,s6299[2],s5130[0],s5129[1]};
    assign in6309_2 = {s6299[1],s6300[1],s5131[0],s5130[1]};
    CLA_4_c KS_6309(s6309, c6309, in6309_1, in6309_2, c6297);
    wire[3:0] s6310, in6310_1, in6310_2;
    wire c6310;
    assign in6310_1 = {c5118,s3443[0],s5136[0],s5137[1]};
    assign in6310_2 = {c5119,s3444[0],s5137[0],s5138[1]};
    CLA_4 KS_6310(s6310, c6310, in6310_1, in6310_2);
    wire[3:0] s6311, in6311_1, in6311_2;
    wire c6311;
    assign in6311_1 = {c5120,s3445[0],s5138[0],s5139[1]};
    assign in6311_2 = {s5121[3],c5121,s5139[0],s5140[1]};
    CLA_4 KS_6311(s6311, c6311, in6311_1, in6311_2);
    wire[3:0] s6312, in6312_1, in6312_2;
    wire c6312;
    assign in6312_1 = {s5122[2],s5122[3],s5140[0],s5141[1]};
    assign in6312_2 = {s5123[2],s5123[3],s5141[0],s5142[1]};
    CLA_4 KS_6312(s6312, c6312, in6312_1, in6312_2);
    wire[3:0] s6313, in6313_1, in6313_2;
    wire c6313;
    assign in6313_1 = {s5124[2],s5124[3],s5142[0],s5143[1]};
    assign in6313_2 = {s5125[2],s5125[3],s5143[0],c5144};
    CLA_4 KS_6313(s6313, c6313, in6313_1, in6313_2);
    wire[3:0] s6314, in6314_1, in6314_2;
    wire c6314;
    assign in6314_1 = {s5126[2],s5126[3],s5144[0],s5145[1]};
    assign in6314_2 = {s5127[2],s5127[3],s5145[0],c5146};
    CLA_4 KS_6314(s6314, c6314, in6314_1, in6314_2);
    wire[3:0] s6315, in6315_1, in6315_2;
    wire c6315;
    assign in6315_1 = {s5128[2],s5128[3],s5146[0],s5147[1]};
    assign in6315_2 = {s5129[2],s5129[3],s5147[0],c5148};
    CLA_4 KS_6315(s6315, c6315, in6315_1, in6315_2);
    wire[2:0] s6316, in6316_1, in6316_2;
    wire c6316;
    assign in6316_1 = {s5130[2],s5130[3],s5148[0]};
    assign in6316_2 = {s5131[2],s5131[3],s5149[0]};
    CLA_3 KS_6316(s6316, c6316, in6316_1, in6316_2);
    wire[0:0] s6317, in6317_1, in6317_2;
    wire c6317;
    assign in6317_1 = {s5132[0]};
    assign in6317_2 = {s5133[0]};
    Half_Adder KS_6317(s6317, c6317, in6317_1, in6317_2);
    wire[1:0] s6318, in6318_1, in6318_2;
    wire c6318;
    assign in6318_1 = {c6300,s5132[1]};
    assign in6318_2 = {c6301,s5133[1]};
    CLA_2 KS_6318(s6318, c6318, in6318_1, in6318_2);
    wire[0:0] s6319, in6319_1, in6319_2;
    wire c6319;
    assign in6319_1 = {c6302};
    assign in6319_2 = {c6303};
    Half_Adder KS_6319(s6319, c6319, in6319_1, in6319_2);
    wire[3:0] s6320, in6320_1, in6320_2;
    wire c6320;
    assign in6320_1 = {c6304,s6310[1],s5150[0],s5149[1]};
    assign in6320_2 = {c6305,s6311[1],s5151[0],c5150};
    CLA_4 KS_6320(s6320, c6320, in6320_1, in6320_2);
    wire[0:0] s6321, in6321_1, in6321_2;
    wire c6321;
    assign in6321_1 = {s6310[0]};
    assign in6321_2 = {s6311[0]};
    Full_Adder KS_6321(s6321, c6321, in6321_1, in6321_2, c6309);
    wire[3:0] s6322, in6322_1, in6322_2;
    wire c6322;
    assign in6322_1 = {c5133,s3461[0],s5159[0],s5159[1]};
    assign in6322_2 = {s5134[2],s5134[3],s5160[0],s5160[1]};
    CLA_4 KS_6322(s6322, c6322, in6322_1, in6322_2);
    wire[3:0] s6323, in6323_1, in6323_2;
    wire c6323;
    assign in6323_1 = {s5135[2],s5135[3],s5161[0],s5161[1]};
    assign in6323_2 = {s5136[2],s5136[3],s5162[0],s5162[1]};
    CLA_4 KS_6323(s6323, c6323, in6323_1, in6323_2);
    wire[3:0] s6324, in6324_1, in6324_2;
    wire c6324;
    assign in6324_1 = {s5137[2],s5137[3],s5163[0],s5163[1]};
    assign in6324_2 = {s5138[2],s5138[3],s5164[0],c5164};
    CLA_4 KS_6324(s6324, c6324, in6324_1, in6324_2);
    wire[3:0] s6325, in6325_1, in6325_2;
    wire c6325;
    assign in6325_1 = {s5139[2],s5139[3],s5165[0],s5165[1]};
    assign in6325_2 = {s5140[2],s5140[3],s5166[0],c5166};
    CLA_4 KS_6325(s6325, c6325, in6325_1, in6325_2);
    wire[3:0] s6326, in6326_1, in6326_2;
    wire c6326;
    assign in6326_1 = {s5141[2],s5141[3],s5167[0],s5167[1]};
    assign in6326_2 = {s5142[2],s5142[3],s5168[0],c5168};
    CLA_4 KS_6326(s6326, c6326, in6326_1, in6326_2);
    wire[3:0] s6327, in6327_1, in6327_2;
    wire c6327;
    assign in6327_1 = {s5143[2],s5143[3],s5169[0],s5169[1]};
    assign in6327_2 = {s5145[2],s5145[3],s5170[0],c5170};
    CLA_4 KS_6327(s6327, c6327, in6327_1, in6327_2);
    wire[0:0] s6328, in6328_1, in6328_2;
    wire c6328;
    assign in6328_1 = {s5147[2]};
    assign in6328_2 = {s5149[2]};
    Half_Adder KS_6328(s6328, c6328, in6328_1, in6328_2);
    wire[3:0] s6329, in6329_1, in6329_2;
    wire c6329;
    assign in6329_1 = {s5151[2],s5147[3],s5171[0],s5171[1]};
    assign in6329_2 = {c6310,c5149,s5172[0],c5172};
    CLA_4 KS_6329(s6329, c6329, in6329_1, in6329_2);
    wire[0:0] s6330, in6330_1, in6330_2;
    wire c6330;
    assign in6330_1 = {c6311};
    assign in6330_2 = {c6312};
    Half_Adder KS_6330(s6330, c6330, in6330_1, in6330_2);
    wire[1:0] s6331, in6331_1, in6331_2;
    wire c6331;
    assign in6331_1 = {c6313,s5151[3]};
    assign in6331_2 = {c6314,s6322[1]};
    CLA_2 KS_6331(s6331, c6331, in6331_1, in6331_2);
    wire[0:0] s6332, in6332_1, in6332_2;
    wire c6332;
    assign in6332_1 = {c6320};
    assign in6332_2 = {s6322[0]};
    Full_Adder KS_6332(s6332, c6332, in6332_1, in6332_2, c6315);
    wire[3:0] s6333, in6333_1, in6333_2;
    wire c6333;
    assign in6333_1 = {s5153[2],s3484[0],s5182[0],s5182[1]};
    assign in6333_2 = {s5154[2],s5152[3],s5183[0],s5183[1]};
    CLA_4 KS_6333(s6333, c6333, in6333_1, in6333_2);
    wire[3:0] s6334, in6334_1, in6334_2;
    wire c6334;
    assign in6334_1 = {s5155[2],s5153[3],s5184[0],s5184[1]};
    assign in6334_2 = {s5156[2],s5154[3],s5185[0],s5185[1]};
    CLA_4 KS_6334(s6334, c6334, in6334_1, in6334_2);
    wire[3:0] s6335, in6335_1, in6335_2;
    wire c6335;
    assign in6335_1 = {s5157[2],s5155[3],s5186[0],s5186[1]};
    assign in6335_2 = {s5158[2],s5156[3],s5187[0],c5187};
    CLA_4 KS_6335(s6335, c6335, in6335_1, in6335_2);
    wire[3:0] s6336, in6336_1, in6336_2;
    wire c6336;
    assign in6336_1 = {s5159[2],s5157[3],s5188[0],s5188[1]};
    assign in6336_2 = {s5160[2],s5158[3],s5189[0],c5189};
    CLA_4 KS_6336(s6336, c6336, in6336_1, in6336_2);
    wire[3:0] s6337, in6337_1, in6337_2;
    wire c6337;
    assign in6337_1 = {s5161[2],s5159[3],s5190[0],s5190[1]};
    assign in6337_2 = {s5162[2],s5160[3],s5191[0],c5191};
    CLA_4 KS_6337(s6337, c6337, in6337_1, in6337_2);
    wire[3:0] s6338, in6338_1, in6338_2;
    wire c6338;
    assign in6338_1 = {s5163[2],s5161[3],s5192[0],s5192[1]};
    assign in6338_2 = {c5165,s5162[3],s5193[0],c5193};
    CLA_4 KS_6338(s6338, c6338, in6338_1, in6338_2);
    wire[0:0] s6339, in6339_1, in6339_2;
    wire c6339;
    assign in6339_1 = {s5167[2]};
    assign in6339_2 = {c5169};
    Half_Adder KS_6339(s6339, c6339, in6339_1, in6339_2);
    wire[3:0] s6340, in6340_1, in6340_2;
    wire c6340;
    assign in6340_1 = {s5171[2],s5163[3],s5194[0],s5194[1]};
    assign in6340_2 = {c5173,c5167,s5195[0],c5195};
    CLA_4 KS_6340(s6340, c6340, in6340_1, in6340_2);
    wire[0:0] s6341, in6341_1, in6341_2;
    wire c6341;
    assign in6341_1 = {c6322};
    assign in6341_2 = {c6323};
    Half_Adder KS_6341(s6341, c6341, in6341_1, in6341_2);
    wire[1:0] s6342, in6342_1, in6342_2;
    wire c6342;
    assign in6342_1 = {c6324,s5171[3]};
    assign in6342_2 = {c6325,s6333[1]};
    CLA_2 KS_6342(s6342, c6342, in6342_1, in6342_2);
    wire[0:0] s6343, in6343_1, in6343_2;
    wire c6343;
    assign in6343_1 = {c6326};
    assign in6343_2 = {c6327};
    Half_Adder KS_6343(s6343, c6343, in6343_1, in6343_2);
    wire[2:0] s6344, in6344_1, in6344_2;
    wire c6344;
    assign in6344_1 = {s6333[0],s6334[1],s5196[0]};
    assign in6344_2 = {s6334[0],s6335[1],s5197[0]};
    CLA_3_c KS_6344(s6344, c6344, in6344_1, in6344_2, c6329);
    wire[3:0] s6345, in6345_1, in6345_2;
    wire c6345;
    assign in6345_1 = {s5176[2],s3513[0],s5204[0],s5205[1]};
    assign in6345_2 = {s5177[2],s5175[3],s5205[0],s5206[1]};
    CLA_4 KS_6345(s6345, c6345, in6345_1, in6345_2);
    wire[3:0] s6346, in6346_1, in6346_2;
    wire c6346;
    assign in6346_1 = {s5178[2],s5176[3],s5206[0],s5207[1]};
    assign in6346_2 = {s5179[2],s5177[3],s5207[0],s5208[1]};
    CLA_4 KS_6346(s6346, c6346, in6346_1, in6346_2);
    wire[3:0] s6347, in6347_1, in6347_2;
    wire c6347;
    assign in6347_1 = {s5180[2],s5178[3],s5208[0],s5209[1]};
    assign in6347_2 = {s5181[2],s5179[3],s5209[0],c5210};
    CLA_4 KS_6347(s6347, c6347, in6347_1, in6347_2);
    wire[3:0] s6348, in6348_1, in6348_2;
    wire c6348;
    assign in6348_1 = {s5182[2],s5180[3],s5210[0],s5211[1]};
    assign in6348_2 = {s5183[2],s5181[3],s5211[0],c5212};
    CLA_4 KS_6348(s6348, c6348, in6348_1, in6348_2);
    wire[3:0] s6349, in6349_1, in6349_2;
    wire c6349;
    assign in6349_1 = {s5184[2],s5182[3],s5212[0],s5213[1]};
    assign in6349_2 = {s5185[2],s5183[3],s5213[0],c5214};
    CLA_4 KS_6349(s6349, c6349, in6349_1, in6349_2);
    wire[3:0] s6350, in6350_1, in6350_2;
    wire c6350;
    assign in6350_1 = {s5186[2],s5184[3],s5214[0],s5215[1]};
    assign in6350_2 = {c5188,s5185[3],s5215[0],c5216};
    CLA_4 KS_6350(s6350, c6350, in6350_1, in6350_2);
    wire[0:0] s6351, in6351_1, in6351_2;
    wire c6351;
    assign in6351_1 = {s5190[2]};
    assign in6351_2 = {c5192};
    Half_Adder KS_6351(s6351, c6351, in6351_1, in6351_2);
    wire[2:0] s6352, in6352_1, in6352_2;
    wire c6352;
    assign in6352_1 = {s5194[2],s5186[3],s5216[0]};
    assign in6352_2 = {c5196,c5190,s5217[0]};
    CLA_3 KS_6352(s6352, c6352, in6352_1, in6352_2);
    wire[0:0] s6353, in6353_1, in6353_2;
    wire c6353;
    assign in6353_1 = {c6333};
    assign in6353_2 = {c6334};
    Half_Adder KS_6353(s6353, c6353, in6353_1, in6353_2);
    wire[1:0] s6354, in6354_1, in6354_2;
    wire c6354;
    assign in6354_1 = {c6335,s5194[3]};
    assign in6354_2 = {c6336,s6345[1]};
    CLA_2 KS_6354(s6354, c6354, in6354_1, in6354_2);
    wire[0:0] s6355, in6355_1, in6355_2;
    wire c6355;
    assign in6355_1 = {c6337};
    assign in6355_2 = {c6338};
    Half_Adder KS_6355(s6355, c6355, in6355_1, in6355_2);
    wire[3:0] s6356, in6356_1, in6356_2;
    wire c6356;
    assign in6356_1 = {s6345[0],s6346[1],s5218[0],s5217[1]};
    assign in6356_2 = {s6346[0],s6347[1],s5219[0],c5218};
    CLA_4_c KS_6356(s6356, c6356, in6356_1, in6356_2, c6340);
    wire[3:0] s6357, in6357_1, in6357_2;
    wire c6357;
    assign in6357_1 = {s5199[2],s3546[0],s5226[0],s5227[1]};
    assign in6357_2 = {s5200[2],s5198[3],s5227[0],s5228[1]};
    CLA_4 KS_6357(s6357, c6357, in6357_1, in6357_2);
    wire[3:0] s6358, in6358_1, in6358_2;
    wire c6358;
    assign in6358_1 = {s5201[2],s5199[3],s5228[0],s5229[1]};
    assign in6358_2 = {s5202[2],s5200[3],s5229[0],s5230[1]};
    CLA_4 KS_6358(s6358, c6358, in6358_1, in6358_2);
    wire[3:0] s6359, in6359_1, in6359_2;
    wire c6359;
    assign in6359_1 = {s5203[2],s5201[3],s5230[0],s5231[1]};
    assign in6359_2 = {s5204[2],s5202[3],s5231[0],c5232};
    CLA_4 KS_6359(s6359, c6359, in6359_1, in6359_2);
    wire[3:0] s6360, in6360_1, in6360_2;
    wire c6360;
    assign in6360_1 = {s5205[2],s5203[3],s5232[0],s5233[1]};
    assign in6360_2 = {s5206[2],s5204[3],s5233[0],c5234};
    CLA_4 KS_6360(s6360, c6360, in6360_1, in6360_2);
    wire[3:0] s6361, in6361_1, in6361_2;
    wire c6361;
    assign in6361_1 = {s5207[2],s5205[3],s5234[0],s5235[1]};
    assign in6361_2 = {s5208[2],s5206[3],s5235[0],c5236};
    CLA_4 KS_6361(s6361, c6361, in6361_1, in6361_2);
    wire[3:0] s6362, in6362_1, in6362_2;
    wire c6362;
    assign in6362_1 = {s5209[2],s5207[3],s5236[0],s5237[1]};
    assign in6362_2 = {c5211,s5208[3],s5237[0],c5238};
    CLA_4 KS_6362(s6362, c6362, in6362_1, in6362_2);
    wire[0:0] s6363, in6363_1, in6363_2;
    wire c6363;
    assign in6363_1 = {s5213[2]};
    assign in6363_2 = {c5215};
    Half_Adder KS_6363(s6363, c6363, in6363_1, in6363_2);
    wire[2:0] s6364, in6364_1, in6364_2;
    wire c6364;
    assign in6364_1 = {s5217[2],s5209[3],s5238[0]};
    assign in6364_2 = {c5219,c5213,s5239[0]};
    CLA_3 KS_6364(s6364, c6364, in6364_1, in6364_2);
    wire[0:0] s6365, in6365_1, in6365_2;
    wire c6365;
    assign in6365_1 = {c6345};
    assign in6365_2 = {c6346};
    Half_Adder KS_6365(s6365, c6365, in6365_1, in6365_2);
    wire[1:0] s6366, in6366_1, in6366_2;
    wire c6366;
    assign in6366_1 = {c6347,s5217[3]};
    assign in6366_2 = {c6348,s6357[1]};
    CLA_2 KS_6366(s6366, c6366, in6366_1, in6366_2);
    wire[0:0] s6367, in6367_1, in6367_2;
    wire c6367;
    assign in6367_1 = {c6349};
    assign in6367_2 = {c6350};
    Half_Adder KS_6367(s6367, c6367, in6367_1, in6367_2);
    wire[3:0] s6368, in6368_1, in6368_2;
    wire c6368;
    assign in6368_1 = {s6357[0],s6358[1],s5240[0],s5239[1]};
    assign in6368_2 = {s6358[0],s6359[1],s5241[0],c5240};
    CLA_4_c KS_6368(s6368, c6368, in6368_1, in6368_2, c6356);
    wire[3:0] s6369, in6369_1, in6369_2;
    wire c6369;
    assign in6369_1 = {s5221[2],s3581[0],s5248[0],s5248[1]};
    assign in6369_2 = {s5222[2],s5220[3],s5249[0],s5249[1]};
    CLA_4 KS_6369(s6369, c6369, in6369_1, in6369_2);
    wire[3:0] s6370, in6370_1, in6370_2;
    wire c6370;
    assign in6370_1 = {s5223[2],s5221[3],s5250[0],s5250[1]};
    assign in6370_2 = {s5224[2],s5222[3],s5251[0],s5251[1]};
    CLA_4 KS_6370(s6370, c6370, in6370_1, in6370_2);
    wire[3:0] s6371, in6371_1, in6371_2;
    wire c6371;
    assign in6371_1 = {s5225[2],s5223[3],s5252[0],s5252[1]};
    assign in6371_2 = {s5226[2],s5224[3],s5253[0],c5253};
    CLA_4 KS_6371(s6371, c6371, in6371_1, in6371_2);
    wire[3:0] s6372, in6372_1, in6372_2;
    wire c6372;
    assign in6372_1 = {s5227[2],s5225[3],s5254[0],s5254[1]};
    assign in6372_2 = {s5228[2],s5226[3],s5255[0],c5255};
    CLA_4 KS_6372(s6372, c6372, in6372_1, in6372_2);
    wire[3:0] s6373, in6373_1, in6373_2;
    wire c6373;
    assign in6373_1 = {s5229[2],s5227[3],s5256[0],s5256[1]};
    assign in6373_2 = {s5230[2],s5228[3],s5257[0],c5257};
    CLA_4 KS_6373(s6373, c6373, in6373_1, in6373_2);
    wire[3:0] s6374, in6374_1, in6374_2;
    wire c6374;
    assign in6374_1 = {s5231[2],s5229[3],s5258[0],s5258[1]};
    assign in6374_2 = {c5233,s5230[3],s5259[0],c5259};
    CLA_4 KS_6374(s6374, c6374, in6374_1, in6374_2);
    wire[0:0] s6375, in6375_1, in6375_2;
    wire c6375;
    assign in6375_1 = {s5235[2]};
    assign in6375_2 = {c5237};
    Half_Adder KS_6375(s6375, c6375, in6375_1, in6375_2);
    wire[3:0] s6376, in6376_1, in6376_2;
    wire c6376;
    assign in6376_1 = {s5239[2],s5231[3],s5260[0],s5260[1]};
    assign in6376_2 = {c5241,c5235,s5261[0],c5261};
    CLA_4 KS_6376(s6376, c6376, in6376_1, in6376_2);
    wire[0:0] s6377, in6377_1, in6377_2;
    wire c6377;
    assign in6377_1 = {c6357};
    assign in6377_2 = {c6358};
    Half_Adder KS_6377(s6377, c6377, in6377_1, in6377_2);
    wire[1:0] s6378, in6378_1, in6378_2;
    wire c6378;
    assign in6378_1 = {c6359,s5239[3]};
    assign in6378_2 = {c6360,s6369[1]};
    CLA_2 KS_6378(s6378, c6378, in6378_1, in6378_2);
    wire[0:0] s6379, in6379_1, in6379_2;
    wire c6379;
    assign in6379_1 = {c6361};
    assign in6379_2 = {c6362};
    Half_Adder KS_6379(s6379, c6379, in6379_1, in6379_2);
    wire[2:0] s6380, in6380_1, in6380_2;
    wire c6380;
    assign in6380_1 = {s6369[0],s6370[1],s5262[0]};
    assign in6380_2 = {s6370[0],s6371[1],s5263[0]};
    CLA_3_c KS_6380(s6380, c6380, in6380_1, in6380_2, c6368);
    wire[3:0] s6381, in6381_1, in6381_2;
    wire c6381;
    assign in6381_1 = {s5243[2],s3618[0],s5270[0],s5271[1]};
    assign in6381_2 = {s5244[2],s5242[3],s5271[0],s5272[1]};
    CLA_4 KS_6381(s6381, c6381, in6381_1, in6381_2);
    wire[3:0] s6382, in6382_1, in6382_2;
    wire c6382;
    assign in6382_1 = {s5245[2],s5243[3],s5272[0],s5273[1]};
    assign in6382_2 = {s5246[2],s5244[3],s5273[0],s5274[1]};
    CLA_4 KS_6382(s6382, c6382, in6382_1, in6382_2);
    wire[3:0] s6383, in6383_1, in6383_2;
    wire c6383;
    assign in6383_1 = {s5247[2],s5245[3],s5274[0],s5275[1]};
    assign in6383_2 = {s5248[2],s5246[3],s5275[0],c5276};
    CLA_4 KS_6383(s6383, c6383, in6383_1, in6383_2);
    wire[3:0] s6384, in6384_1, in6384_2;
    wire c6384;
    assign in6384_1 = {s5249[2],s5247[3],s5276[0],s5277[1]};
    assign in6384_2 = {s5250[2],s5248[3],s5277[0],c5278};
    CLA_4 KS_6384(s6384, c6384, in6384_1, in6384_2);
    wire[3:0] s6385, in6385_1, in6385_2;
    wire c6385;
    assign in6385_1 = {s5251[2],s5249[3],s5278[0],s5279[1]};
    assign in6385_2 = {s5252[2],s5250[3],s5279[0],c5280};
    CLA_4 KS_6385(s6385, c6385, in6385_1, in6385_2);
    wire[3:0] s6386, in6386_1, in6386_2;
    wire c6386;
    assign in6386_1 = {s5254[2],s5251[3],s5280[0],s5281[1]};
    assign in6386_2 = {c5256,s5252[3],s5281[0],c5282};
    CLA_4 KS_6386(s6386, c6386, in6386_1, in6386_2);
    wire[0:0] s6387, in6387_1, in6387_2;
    wire c6387;
    assign in6387_1 = {s5258[2]};
    assign in6387_2 = {c5260};
    Half_Adder KS_6387(s6387, c6387, in6387_1, in6387_2);
    wire[2:0] s6388, in6388_1, in6388_2;
    wire c6388;
    assign in6388_1 = {s5262[2],s5254[3],s5282[0]};
    assign in6388_2 = {c6369,c5258,s5283[0]};
    CLA_3 KS_6388(s6388, c6388, in6388_1, in6388_2);
    wire[0:0] s6389, in6389_1, in6389_2;
    wire c6389;
    assign in6389_1 = {c6370};
    assign in6389_2 = {c6371};
    Half_Adder KS_6389(s6389, c6389, in6389_1, in6389_2);
    wire[1:0] s6390, in6390_1, in6390_2;
    wire c6390;
    assign in6390_1 = {c6372,s5262[3]};
    assign in6390_2 = {c6373,s6381[1]};
    CLA_2 KS_6390(s6390, c6390, in6390_1, in6390_2);
    wire[0:0] s6391, in6391_1, in6391_2;
    wire c6391;
    assign in6391_1 = {c6376};
    assign in6391_2 = {s6381[0]};
    Full_Adder KS_6391(s6391, c6391, in6391_1, in6391_2, c6374);
    wire[3:0] s6392, in6392_1, in6392_2;
    wire c6392;
    assign in6392_1 = {s5266[2],s3656[0],s5293[0],s5293[1]};
    assign in6392_2 = {s5267[2],s5264[3],s5294[0],s5294[1]};
    CLA_4 KS_6392(s6392, c6392, in6392_1, in6392_2);
    wire[3:0] s6393, in6393_1, in6393_2;
    wire c6393;
    assign in6393_1 = {s5268[2],s5265[3],s5295[0],s5295[1]};
    assign in6393_2 = {s5269[2],s5266[3],s5296[0],s5296[1]};
    CLA_4 KS_6393(s6393, c6393, in6393_1, in6393_2);
    wire[3:0] s6394, in6394_1, in6394_2;
    wire c6394;
    assign in6394_1 = {s5270[2],s5267[3],s5297[0],s5297[1]};
    assign in6394_2 = {s5271[2],s5268[3],s5298[0],c5298};
    CLA_4 KS_6394(s6394, c6394, in6394_1, in6394_2);
    wire[3:0] s6395, in6395_1, in6395_2;
    wire c6395;
    assign in6395_1 = {s5272[2],s5269[3],s5299[0],s5299[1]};
    assign in6395_2 = {s5273[2],s5270[3],s5300[0],c5300};
    CLA_4 KS_6395(s6395, c6395, in6395_1, in6395_2);
    wire[3:0] s6396, in6396_1, in6396_2;
    wire c6396;
    assign in6396_1 = {s5274[2],s5271[3],s5301[0],s5301[1]};
    assign in6396_2 = {c5275,s5272[3],s5302[0],c5302};
    CLA_4 KS_6396(s6396, c6396, in6396_1, in6396_2);
    wire[3:0] s6397, in6397_1, in6397_2;
    wire c6397;
    assign in6397_1 = {s5277[2],s5273[3],s5303[0],s5303[1]};
    assign in6397_2 = {c5279,s5274[3],s5304[0],c5304};
    CLA_4 KS_6397(s6397, c6397, in6397_1, in6397_2);
    wire[0:0] s6398, in6398_1, in6398_2;
    wire c6398;
    assign in6398_1 = {s5281[2]};
    assign in6398_2 = {c5283};
    Half_Adder KS_6398(s6398, c6398, in6398_1, in6398_2);
    wire[3:0] s6399, in6399_1, in6399_2;
    wire c6399;
    assign in6399_1 = {s5285[2],s5277[3],s5305[0],s5305[1]};
    assign in6399_2 = {c6381,c5281,s5306[0],c5306};
    CLA_4 KS_6399(s6399, c6399, in6399_1, in6399_2);
    wire[0:0] s6400, in6400_1, in6400_2;
    wire c6400;
    assign in6400_1 = {c6382};
    assign in6400_2 = {c6383};
    Half_Adder KS_6400(s6400, c6400, in6400_1, in6400_2);
    wire[1:0] s6401, in6401_1, in6401_2;
    wire c6401;
    assign in6401_1 = {c6385,s5285[3]};
    assign in6401_2 = {c6386,s6392[1]};
    CLA_2_c KS_6401(s6401, c6401, in6401_1, in6401_2, c6384);
    wire[3:0] s6402, in6402_1, in6402_2;
    wire c6402;
    assign in6402_1 = {s5288[2],s3694[0],s5316[0],s5316[1]};
    assign in6402_2 = {s5289[2],s5286[3],s5317[0],s5317[1]};
    CLA_4 KS_6402(s6402, c6402, in6402_1, in6402_2);
    wire[3:0] s6403, in6403_1, in6403_2;
    wire c6403;
    assign in6403_1 = {s5290[2],s5287[3],s5318[0],s5318[1]};
    assign in6403_2 = {s5291[2],s5288[3],s5319[0],s5319[1]};
    CLA_4 KS_6403(s6403, c6403, in6403_1, in6403_2);
    wire[3:0] s6404, in6404_1, in6404_2;
    wire c6404;
    assign in6404_1 = {s5292[2],s5289[3],s5320[0],s5320[1]};
    assign in6404_2 = {s5293[2],s5290[3],s5321[0],c5321};
    CLA_4 KS_6404(s6404, c6404, in6404_1, in6404_2);
    wire[3:0] s6405, in6405_1, in6405_2;
    wire c6405;
    assign in6405_1 = {s5294[2],s5291[3],s5322[0],s5322[1]};
    assign in6405_2 = {s5295[2],s5292[3],s5323[0],c5323};
    CLA_4 KS_6405(s6405, c6405, in6405_1, in6405_2);
    wire[3:0] s6406, in6406_1, in6406_2;
    wire c6406;
    assign in6406_1 = {s5296[2],s5293[3],s5324[0],s5324[1]};
    assign in6406_2 = {c5297,s5294[3],s5325[0],c5325};
    CLA_4 KS_6406(s6406, c6406, in6406_1, in6406_2);
    wire[3:0] s6407, in6407_1, in6407_2;
    wire c6407;
    assign in6407_1 = {s5299[2],s5295[3],s5326[0],s5326[1]};
    assign in6407_2 = {c5301,s5296[3],s5327[0],c5327};
    CLA_4 KS_6407(s6407, c6407, in6407_1, in6407_2);
    wire[0:0] s6408, in6408_1, in6408_2;
    wire c6408;
    assign in6408_1 = {s5303[2]};
    assign in6408_2 = {c5305};
    Half_Adder KS_6408(s6408, c6408, in6408_1, in6408_2);
    wire[3:0] s6409, in6409_1, in6409_2;
    wire c6409;
    assign in6409_1 = {s5307[2],s5299[3],s5328[0],s5328[1]};
    assign in6409_2 = {c6392,c5303,s5329[0],c5329};
    CLA_4 KS_6409(s6409, c6409, in6409_1, in6409_2);
    wire[0:0] s6410, in6410_1, in6410_2;
    wire c6410;
    assign in6410_1 = {c6393};
    assign in6410_2 = {c6394};
    Half_Adder KS_6410(s6410, c6410, in6410_1, in6410_2);
    wire[1:0] s6411, in6411_1, in6411_2;
    wire c6411;
    assign in6411_1 = {c6395,s5307[3]};
    assign in6411_2 = {c6396,s6402[1]};
    CLA_2 KS_6411(s6411, c6411, in6411_1, in6411_2);
    wire[0:0] s6412, in6412_1, in6412_2;
    wire c6412;
    assign in6412_1 = {c6399};
    assign in6412_2 = {s6402[0]};
    Full_Adder KS_6412(s6412, c6412, in6412_1, in6412_2, c6397);
    wire[3:0] s6413, in6413_1, in6413_2;
    wire c6413;
    assign in6413_1 = {s5310[2],s3731[0],s5338[0],s5339[1]};
    assign in6413_2 = {s5311[2],s5309[3],s5339[0],s5340[1]};
    CLA_4 KS_6413(s6413, c6413, in6413_1, in6413_2);
    wire[3:0] s6414, in6414_1, in6414_2;
    wire c6414;
    assign in6414_1 = {s5312[2],s5310[3],s5340[0],s5341[1]};
    assign in6414_2 = {s5313[2],s5311[3],s5341[0],s5342[1]};
    CLA_4 KS_6414(s6414, c6414, in6414_1, in6414_2);
    wire[3:0] s6415, in6415_1, in6415_2;
    wire c6415;
    assign in6415_1 = {s5314[2],s5312[3],s5342[0],s5343[1]};
    assign in6415_2 = {s5315[2],s5313[3],s5343[0],c5344};
    CLA_4 KS_6415(s6415, c6415, in6415_1, in6415_2);
    wire[3:0] s6416, in6416_1, in6416_2;
    wire c6416;
    assign in6416_1 = {s5316[2],s5314[3],s5344[0],s5345[1]};
    assign in6416_2 = {s5317[2],s5315[3],s5345[0],c5346};
    CLA_4 KS_6416(s6416, c6416, in6416_1, in6416_2);
    wire[3:0] s6417, in6417_1, in6417_2;
    wire c6417;
    assign in6417_1 = {s5318[2],s5316[3],s5346[0],s5347[1]};
    assign in6417_2 = {s5319[2],s5317[3],s5347[0],c5348};
    CLA_4 KS_6417(s6417, c6417, in6417_1, in6417_2);
    wire[3:0] s6418, in6418_1, in6418_2;
    wire c6418;
    assign in6418_1 = {s5320[2],s5318[3],s5348[0],s5349[1]};
    assign in6418_2 = {c5322,s5319[3],s5349[0],c5350};
    CLA_4 KS_6418(s6418, c6418, in6418_1, in6418_2);
    wire[0:0] s6419, in6419_1, in6419_2;
    wire c6419;
    assign in6419_1 = {s5324[2]};
    assign in6419_2 = {c5326};
    Half_Adder KS_6419(s6419, c6419, in6419_1, in6419_2);
    wire[2:0] s6420, in6420_1, in6420_2;
    wire c6420;
    assign in6420_1 = {s5328[2],s5320[3],s5350[0]};
    assign in6420_2 = {c5330,c5324,s5351[0]};
    CLA_3 KS_6420(s6420, c6420, in6420_1, in6420_2);
    wire[0:0] s6421, in6421_1, in6421_2;
    wire c6421;
    assign in6421_1 = {c6402};
    assign in6421_2 = {c6403};
    Half_Adder KS_6421(s6421, c6421, in6421_1, in6421_2);
    wire[1:0] s6422, in6422_1, in6422_2;
    wire c6422;
    assign in6422_1 = {c6404,s5328[3]};
    assign in6422_2 = {c6405,s6413[1]};
    CLA_2 KS_6422(s6422, c6422, in6422_1, in6422_2);
    wire[0:0] s6423, in6423_1, in6423_2;
    wire c6423;
    assign in6423_1 = {c6406};
    assign in6423_2 = {c6407};
    Half_Adder KS_6423(s6423, c6423, in6423_1, in6423_2);
    wire[3:0] s6424, in6424_1, in6424_2;
    wire c6424;
    assign in6424_1 = {s6413[0],s6414[1],s5352[0],s5351[1]};
    assign in6424_2 = {s6414[0],s6415[1],s5353[0],c5352};
    CLA_4_c KS_6424(s6424, c6424, in6424_1, in6424_2, c6409);
    wire[3:0] s6425, in6425_1, in6425_2;
    wire c6425;
    assign in6425_1 = {s5333[2],s3768[0],s5360[0],s5361[1]};
    assign in6425_2 = {s5334[2],s5332[3],s5361[0],s5362[1]};
    CLA_4 KS_6425(s6425, c6425, in6425_1, in6425_2);
    wire[3:0] s6426, in6426_1, in6426_2;
    wire c6426;
    assign in6426_1 = {s5335[2],s5333[3],s5362[0],s5363[1]};
    assign in6426_2 = {s5336[2],s5334[3],s5363[0],s5364[1]};
    CLA_4 KS_6426(s6426, c6426, in6426_1, in6426_2);
    wire[3:0] s6427, in6427_1, in6427_2;
    wire c6427;
    assign in6427_1 = {s5337[2],s5335[3],s5364[0],s5365[1]};
    assign in6427_2 = {s5338[2],s5336[3],s5365[0],c5366};
    CLA_4 KS_6427(s6427, c6427, in6427_1, in6427_2);
    wire[3:0] s6428, in6428_1, in6428_2;
    wire c6428;
    assign in6428_1 = {s5339[2],s5337[3],s5366[0],s5367[1]};
    assign in6428_2 = {s5340[2],s5338[3],s5367[0],c5368};
    CLA_4 KS_6428(s6428, c6428, in6428_1, in6428_2);
    wire[3:0] s6429, in6429_1, in6429_2;
    wire c6429;
    assign in6429_1 = {s5341[2],s5339[3],s5368[0],s5369[1]};
    assign in6429_2 = {s5342[2],s5340[3],s5369[0],c5370};
    CLA_4 KS_6429(s6429, c6429, in6429_1, in6429_2);
    wire[3:0] s6430, in6430_1, in6430_2;
    wire c6430;
    assign in6430_1 = {s5343[2],s5341[3],s5370[0],s5371[1]};
    assign in6430_2 = {c5345,s5342[3],s5371[0],c5372};
    CLA_4 KS_6430(s6430, c6430, in6430_1, in6430_2);
    wire[0:0] s6431, in6431_1, in6431_2;
    wire c6431;
    assign in6431_1 = {s5347[2]};
    assign in6431_2 = {c5349};
    Half_Adder KS_6431(s6431, c6431, in6431_1, in6431_2);
    wire[2:0] s6432, in6432_1, in6432_2;
    wire c6432;
    assign in6432_1 = {s5351[2],s5343[3],s5372[0]};
    assign in6432_2 = {c5353,c5347,s5373[0]};
    CLA_3 KS_6432(s6432, c6432, in6432_1, in6432_2);
    wire[0:0] s6433, in6433_1, in6433_2;
    wire c6433;
    assign in6433_1 = {c6413};
    assign in6433_2 = {c6414};
    Half_Adder KS_6433(s6433, c6433, in6433_1, in6433_2);
    wire[1:0] s6434, in6434_1, in6434_2;
    wire c6434;
    assign in6434_1 = {c6415,s5351[3]};
    assign in6434_2 = {c6416,s6425[1]};
    CLA_2 KS_6434(s6434, c6434, in6434_1, in6434_2);
    wire[0:0] s6435, in6435_1, in6435_2;
    wire c6435;
    assign in6435_1 = {c6417};
    assign in6435_2 = {c6418};
    Half_Adder KS_6435(s6435, c6435, in6435_1, in6435_2);
    wire[3:0] s6436, in6436_1, in6436_2;
    wire c6436;
    assign in6436_1 = {s6425[0],s6426[1],s5374[0],s5373[1]};
    assign in6436_2 = {s6426[0],s6427[1],s5375[0],c5374};
    CLA_4_c KS_6436(s6436, c6436, in6436_1, in6436_2, c6424);
    wire[3:0] s6437, in6437_1, in6437_2;
    wire c6437;
    assign in6437_1 = {s5355[2],s3805[0],s5382[0],s5383[1]};
    assign in6437_2 = {s5356[2],s5354[3],s5383[0],s5384[1]};
    CLA_4 KS_6437(s6437, c6437, in6437_1, in6437_2);
    wire[3:0] s6438, in6438_1, in6438_2;
    wire c6438;
    assign in6438_1 = {s5357[2],s5355[3],s5384[0],s5385[1]};
    assign in6438_2 = {s5358[2],s5356[3],s5385[0],s5386[1]};
    CLA_4 KS_6438(s6438, c6438, in6438_1, in6438_2);
    wire[3:0] s6439, in6439_1, in6439_2;
    wire c6439;
    assign in6439_1 = {s5359[2],s5357[3],s5386[0],s5387[1]};
    assign in6439_2 = {s5360[2],s5358[3],s5387[0],c5388};
    CLA_4 KS_6439(s6439, c6439, in6439_1, in6439_2);
    wire[3:0] s6440, in6440_1, in6440_2;
    wire c6440;
    assign in6440_1 = {s5361[2],s5359[3],s5388[0],s5389[1]};
    assign in6440_2 = {s5362[2],s5360[3],s5389[0],c5390};
    CLA_4 KS_6440(s6440, c6440, in6440_1, in6440_2);
    wire[3:0] s6441, in6441_1, in6441_2;
    wire c6441;
    assign in6441_1 = {s5363[2],s5361[3],s5390[0],s5391[1]};
    assign in6441_2 = {s5364[2],s5362[3],s5391[0],c5392};
    CLA_4 KS_6441(s6441, c6441, in6441_1, in6441_2);
    wire[3:0] s6442, in6442_1, in6442_2;
    wire c6442;
    assign in6442_1 = {s5365[2],s5363[3],s5392[0],s5393[1]};
    assign in6442_2 = {c5367,s5364[3],s5393[0],c5394};
    CLA_4 KS_6442(s6442, c6442, in6442_1, in6442_2);
    wire[0:0] s6443, in6443_1, in6443_2;
    wire c6443;
    assign in6443_1 = {s5369[2]};
    assign in6443_2 = {c5371};
    Half_Adder KS_6443(s6443, c6443, in6443_1, in6443_2);
    wire[2:0] s6444, in6444_1, in6444_2;
    wire c6444;
    assign in6444_1 = {s5373[2],s5365[3],s5394[0]};
    assign in6444_2 = {c5375,c5369,s5395[0]};
    CLA_3 KS_6444(s6444, c6444, in6444_1, in6444_2);
    wire[0:0] s6445, in6445_1, in6445_2;
    wire c6445;
    assign in6445_1 = {c6425};
    assign in6445_2 = {c6426};
    Half_Adder KS_6445(s6445, c6445, in6445_1, in6445_2);
    wire[1:0] s6446, in6446_1, in6446_2;
    wire c6446;
    assign in6446_1 = {c6427,s5373[3]};
    assign in6446_2 = {c6428,s6437[1]};
    CLA_2 KS_6446(s6446, c6446, in6446_1, in6446_2);
    wire[0:0] s6447, in6447_1, in6447_2;
    wire c6447;
    assign in6447_1 = {c6429};
    assign in6447_2 = {c6430};
    Half_Adder KS_6447(s6447, c6447, in6447_1, in6447_2);
    wire[3:0] s6448, in6448_1, in6448_2;
    wire c6448;
    assign in6448_1 = {s6437[0],s6438[1],s5396[0],s5395[1]};
    assign in6448_2 = {s6438[0],s6439[1],s5397[0],c5396};
    CLA_4_c KS_6448(s6448, c6448, in6448_1, in6448_2, c6436);
    wire[3:0] s6449, in6449_1, in6449_2;
    wire c6449;
    assign in6449_1 = {s5377[2],s3842[0],s5404[0],s5405[1]};
    assign in6449_2 = {s5378[2],s5376[3],s5405[0],s5406[1]};
    CLA_4 KS_6449(s6449, c6449, in6449_1, in6449_2);
    wire[3:0] s6450, in6450_1, in6450_2;
    wire c6450;
    assign in6450_1 = {s5379[2],s5377[3],s5406[0],s5407[1]};
    assign in6450_2 = {s5380[2],s5378[3],s5407[0],s5408[1]};
    CLA_4 KS_6450(s6450, c6450, in6450_1, in6450_2);
    wire[3:0] s6451, in6451_1, in6451_2;
    wire c6451;
    assign in6451_1 = {s5381[2],s5379[3],s5408[0],s5409[1]};
    assign in6451_2 = {s5382[2],s5380[3],s5409[0],c5410};
    CLA_4 KS_6451(s6451, c6451, in6451_1, in6451_2);
    wire[3:0] s6452, in6452_1, in6452_2;
    wire c6452;
    assign in6452_1 = {s5383[2],s5381[3],s5410[0],s5411[1]};
    assign in6452_2 = {s5384[2],s5382[3],s5411[0],c5412};
    CLA_4 KS_6452(s6452, c6452, in6452_1, in6452_2);
    wire[3:0] s6453, in6453_1, in6453_2;
    wire c6453;
    assign in6453_1 = {s5385[2],s5383[3],s5412[0],s5413[1]};
    assign in6453_2 = {s5386[2],s5384[3],s5413[0],c5414};
    CLA_4 KS_6453(s6453, c6453, in6453_1, in6453_2);
    wire[3:0] s6454, in6454_1, in6454_2;
    wire c6454;
    assign in6454_1 = {s5387[2],s5385[3],s5414[0],s5415[1]};
    assign in6454_2 = {c5389,s5386[3],s5415[0],c5416};
    CLA_4 KS_6454(s6454, c6454, in6454_1, in6454_2);
    wire[0:0] s6455, in6455_1, in6455_2;
    wire c6455;
    assign in6455_1 = {s5391[2]};
    assign in6455_2 = {c5393};
    Half_Adder KS_6455(s6455, c6455, in6455_1, in6455_2);
    wire[2:0] s6456, in6456_1, in6456_2;
    wire c6456;
    assign in6456_1 = {s5395[2],s5387[3],s5416[0]};
    assign in6456_2 = {c5397,c5391,s5417[0]};
    CLA_3 KS_6456(s6456, c6456, in6456_1, in6456_2);
    wire[0:0] s6457, in6457_1, in6457_2;
    wire c6457;
    assign in6457_1 = {c6437};
    assign in6457_2 = {c6438};
    Half_Adder KS_6457(s6457, c6457, in6457_1, in6457_2);
    wire[1:0] s6458, in6458_1, in6458_2;
    wire c6458;
    assign in6458_1 = {c6439,s5395[3]};
    assign in6458_2 = {c6440,s6449[1]};
    CLA_2 KS_6458(s6458, c6458, in6458_1, in6458_2);
    wire[0:0] s6459, in6459_1, in6459_2;
    wire c6459;
    assign in6459_1 = {c6441};
    assign in6459_2 = {c6442};
    Half_Adder KS_6459(s6459, c6459, in6459_1, in6459_2);
    wire[3:0] s6460, in6460_1, in6460_2;
    wire c6460;
    assign in6460_1 = {s6449[0],s6450[1],s5418[0],s5417[1]};
    assign in6460_2 = {s6450[0],s6451[1],s5419[0],c5418};
    CLA_4_c KS_6460(s6460, c6460, in6460_1, in6460_2, c6448);
    wire[3:0] s6461, in6461_1, in6461_2;
    wire c6461;
    assign in6461_1 = {s5399[2],s3878[0],s5427[0],s5428[1]};
    assign in6461_2 = {s5400[2],s5398[3],s5428[0],s5429[1]};
    CLA_4 KS_6461(s6461, c6461, in6461_1, in6461_2);
    wire[3:0] s6462, in6462_1, in6462_2;
    wire c6462;
    assign in6462_1 = {s5401[2],s5399[3],s5429[0],s5430[1]};
    assign in6462_2 = {s5402[2],s5400[3],s5430[0],c5431};
    CLA_4 KS_6462(s6462, c6462, in6462_1, in6462_2);
    wire[3:0] s6463, in6463_1, in6463_2;
    wire c6463;
    assign in6463_1 = {s5403[2],s5401[3],s5431[0],s5432[1]};
    assign in6463_2 = {s5404[2],s5402[3],s5432[0],c5433};
    CLA_4 KS_6463(s6463, c6463, in6463_1, in6463_2);
    wire[3:0] s6464, in6464_1, in6464_2;
    wire c6464;
    assign in6464_1 = {s5405[2],s5403[3],s5433[0],s5434[1]};
    assign in6464_2 = {s5406[2],s5404[3],s5434[0],c5435};
    CLA_4 KS_6464(s6464, c6464, in6464_1, in6464_2);
    wire[3:0] s6465, in6465_1, in6465_2;
    wire c6465;
    assign in6465_1 = {s5407[2],s5405[3],s5435[0],s5436[1]};
    assign in6465_2 = {s5408[2],s5406[3],s5436[0],c5437};
    CLA_4 KS_6465(s6465, c6465, in6465_1, in6465_2);
    wire[3:0] s6466, in6466_1, in6466_2;
    wire c6466;
    assign in6466_1 = {s5409[2],s5407[3],s5437[0],s5438[1]};
    assign in6466_2 = {c5411,s5408[3],s5438[0],c5439};
    CLA_4 KS_6466(s6466, c6466, in6466_1, in6466_2);
    wire[0:0] s6467, in6467_1, in6467_2;
    wire c6467;
    assign in6467_1 = {s5413[2]};
    assign in6467_2 = {c5415};
    Half_Adder KS_6467(s6467, c6467, in6467_1, in6467_2);
    wire[2:0] s6468, in6468_1, in6468_2;
    wire c6468;
    assign in6468_1 = {s5417[2],s5409[3],s5439[0]};
    assign in6468_2 = {c5419,c5413,s5440[0]};
    CLA_3 KS_6468(s6468, c6468, in6468_1, in6468_2);
    wire[0:0] s6469, in6469_1, in6469_2;
    wire c6469;
    assign in6469_1 = {c6449};
    assign in6469_2 = {c6450};
    Half_Adder KS_6469(s6469, c6469, in6469_1, in6469_2);
    wire[1:0] s6470, in6470_1, in6470_2;
    wire c6470;
    assign in6470_1 = {c6451,s5417[3]};
    assign in6470_2 = {c6452,s6461[1]};
    CLA_2 KS_6470(s6470, c6470, in6470_1, in6470_2);
    wire[0:0] s6471, in6471_1, in6471_2;
    wire c6471;
    assign in6471_1 = {c6453};
    assign in6471_2 = {c6454};
    Half_Adder KS_6471(s6471, c6471, in6471_1, in6471_2);
    wire[3:0] s6472, in6472_1, in6472_2;
    wire c6472;
    assign in6472_1 = {s6461[0],s6462[1],s5441[0],s5440[1]};
    assign in6472_2 = {s6462[0],s6463[1],s5442[0],c5441};
    CLA_4_c KS_6472(s6472, c6472, in6472_1, in6472_2, c6460);
    wire[3:0] s6473, in6473_1, in6473_2;
    wire c6473;
    assign in6473_1 = {s5421[2],s3914[0],s5450[0],s5451[1]};
    assign in6473_2 = {s5422[2],s5420[3],s5451[0],s5452[1]};
    CLA_4 KS_6473(s6473, c6473, in6473_1, in6473_2);
    wire[3:0] s6474, in6474_1, in6474_2;
    wire c6474;
    assign in6474_1 = {s5423[2],s5421[3],s5452[0],s5453[1]};
    assign in6474_2 = {s5424[2],s5422[3],s5453[0],c5454};
    CLA_4 KS_6474(s6474, c6474, in6474_1, in6474_2);
    wire[3:0] s6475, in6475_1, in6475_2;
    wire c6475;
    assign in6475_1 = {s5425[2],s5423[3],s5454[0],s5455[1]};
    assign in6475_2 = {s5426[2],s5424[3],s5455[0],c5456};
    CLA_4 KS_6475(s6475, c6475, in6475_1, in6475_2);
    wire[3:0] s6476, in6476_1, in6476_2;
    wire c6476;
    assign in6476_1 = {s5427[2],s5425[3],s5456[0],s5457[1]};
    assign in6476_2 = {s5428[2],s5426[3],s5457[0],c5458};
    CLA_4 KS_6476(s6476, c6476, in6476_1, in6476_2);
    wire[3:0] s6477, in6477_1, in6477_2;
    wire c6477;
    assign in6477_1 = {s5429[2],s5427[3],s5458[0],s5459[1]};
    assign in6477_2 = {s5430[2],s5428[3],s5459[0],c5460};
    CLA_4 KS_6477(s6477, c6477, in6477_1, in6477_2);
    wire[3:0] s6478, in6478_1, in6478_2;
    wire c6478;
    assign in6478_1 = {s5432[2],s5429[3],s5460[0],s5461[1]};
    assign in6478_2 = {c5434,s5430[3],s5461[0],c5462};
    CLA_4 KS_6478(s6478, c6478, in6478_1, in6478_2);
    wire[0:0] s6479, in6479_1, in6479_2;
    wire c6479;
    assign in6479_1 = {s5436[2]};
    assign in6479_2 = {c5438};
    Half_Adder KS_6479(s6479, c6479, in6479_1, in6479_2);
    wire[2:0] s6480, in6480_1, in6480_2;
    wire c6480;
    assign in6480_1 = {s5440[2],s5432[3],s5462[0]};
    assign in6480_2 = {c5442,c5436,s5463[0]};
    CLA_3 KS_6480(s6480, c6480, in6480_1, in6480_2);
    wire[0:0] s6481, in6481_1, in6481_2;
    wire c6481;
    assign in6481_1 = {c6461};
    assign in6481_2 = {c6462};
    Half_Adder KS_6481(s6481, c6481, in6481_1, in6481_2);
    wire[1:0] s6482, in6482_1, in6482_2;
    wire c6482;
    assign in6482_1 = {c6463,s5440[3]};
    assign in6482_2 = {c6464,s6473[1]};
    CLA_2 KS_6482(s6482, c6482, in6482_1, in6482_2);
    wire[0:0] s6483, in6483_1, in6483_2;
    wire c6483;
    assign in6483_1 = {c6465};
    assign in6483_2 = {c6466};
    Half_Adder KS_6483(s6483, c6483, in6483_1, in6483_2);
    wire[3:0] s6484, in6484_1, in6484_2;
    wire c6484;
    assign in6484_1 = {s6473[0],s6474[1],s5464[0],s5463[1]};
    assign in6484_2 = {s6474[0],s6475[1],s5465[0],c5464};
    CLA_4_c KS_6484(s6484, c6484, in6484_1, in6484_2, c6472);
    wire[3:0] s6485, in6485_1, in6485_2;
    wire c6485;
    assign in6485_1 = {s5445[2],s3952[0],s5473[0],s5474[1]};
    assign in6485_2 = {s5446[2],s5443[3],s5474[0],s5475[1]};
    CLA_4 KS_6485(s6485, c6485, in6485_1, in6485_2);
    wire[3:0] s6486, in6486_1, in6486_2;
    wire c6486;
    assign in6486_1 = {s5447[2],s5444[3],s5475[0],s5476[1]};
    assign in6486_2 = {s5448[2],s5445[3],s5476[0],c5477};
    CLA_4 KS_6486(s6486, c6486, in6486_1, in6486_2);
    wire[3:0] s6487, in6487_1, in6487_2;
    wire c6487;
    assign in6487_1 = {s5449[2],s5446[3],s5477[0],s5478[1]};
    assign in6487_2 = {s5450[2],s5447[3],s5478[0],c5479};
    CLA_4 KS_6487(s6487, c6487, in6487_1, in6487_2);
    wire[3:0] s6488, in6488_1, in6488_2;
    wire c6488;
    assign in6488_1 = {s5451[2],s5448[3],s5479[0],s5480[1]};
    assign in6488_2 = {s5452[2],s5449[3],s5480[0],c5481};
    CLA_4 KS_6488(s6488, c6488, in6488_1, in6488_2);
    wire[3:0] s6489, in6489_1, in6489_2;
    wire c6489;
    assign in6489_1 = {s5453[2],s5450[3],s5481[0],s5482[1]};
    assign in6489_2 = {c5455,s5451[3],s5482[0],c5483};
    CLA_4 KS_6489(s6489, c6489, in6489_1, in6489_2);
    wire[3:0] s6490, in6490_1, in6490_2;
    wire c6490;
    assign in6490_1 = {s5457[2],s5452[3],s5483[0],s5484[1]};
    assign in6490_2 = {c5459,s5453[3],s5484[0],c5485};
    CLA_4 KS_6490(s6490, c6490, in6490_1, in6490_2);
    wire[0:0] s6491, in6491_1, in6491_2;
    wire c6491;
    assign in6491_1 = {s5461[2]};
    assign in6491_2 = {c5463};
    Half_Adder KS_6491(s6491, c6491, in6491_1, in6491_2);
    wire[2:0] s6492, in6492_1, in6492_2;
    wire c6492;
    assign in6492_1 = {s5465[2],s5457[3],s5485[0]};
    assign in6492_2 = {c6473,c5461,s5486[0]};
    CLA_3 KS_6492(s6492, c6492, in6492_1, in6492_2);
    wire[0:0] s6493, in6493_1, in6493_2;
    wire c6493;
    assign in6493_1 = {c6474};
    assign in6493_2 = {c6475};
    Half_Adder KS_6493(s6493, c6493, in6493_1, in6493_2);
    wire[1:0] s6494, in6494_1, in6494_2;
    wire c6494;
    assign in6494_1 = {c6476,s5465[3]};
    assign in6494_2 = {c6477,s6485[1]};
    CLA_2 KS_6494(s6494, c6494, in6494_1, in6494_2);
    wire[0:0] s6495, in6495_1, in6495_2;
    wire c6495;
    assign in6495_1 = {c6484};
    assign in6495_2 = {s6485[0]};
    Full_Adder KS_6495(s6495, c6495, in6495_1, in6495_2, c6478);
    wire[3:0] s6496, in6496_1, in6496_2;
    wire c6496;
    assign in6496_1 = {s5467[2],s3988[0],s5496[0],s5497[1]};
    assign in6496_2 = {s5468[2],s5466[3],s5497[0],s5498[1]};
    CLA_4 KS_6496(s6496, c6496, in6496_1, in6496_2);
    wire[3:0] s6497, in6497_1, in6497_2;
    wire c6497;
    assign in6497_1 = {s5469[2],s5467[3],s5498[0],s5499[1]};
    assign in6497_2 = {s5470[2],s5468[3],s5499[0],c5500};
    CLA_4 KS_6497(s6497, c6497, in6497_1, in6497_2);
    wire[3:0] s6498, in6498_1, in6498_2;
    wire c6498;
    assign in6498_1 = {s5471[2],s5469[3],s5500[0],s5501[1]};
    assign in6498_2 = {s5472[2],s5470[3],s5501[0],c5502};
    CLA_4 KS_6498(s6498, c6498, in6498_1, in6498_2);
    wire[3:0] s6499, in6499_1, in6499_2;
    wire c6499;
    assign in6499_1 = {s5473[2],s5471[3],s5502[0],s5503[1]};
    assign in6499_2 = {s5474[2],s5472[3],s5503[0],c5504};
    CLA_4 KS_6499(s6499, c6499, in6499_1, in6499_2);
    wire[3:0] s6500, in6500_1, in6500_2;
    wire c6500;
    assign in6500_1 = {s5475[2],s5473[3],s5504[0],s5505[1]};
    assign in6500_2 = {s5476[2],s5474[3],s5505[0],c5506};
    CLA_4 KS_6500(s6500, c6500, in6500_1, in6500_2);
    wire[3:0] s6501, in6501_1, in6501_2;
    wire c6501;
    assign in6501_1 = {s5478[2],s5475[3],s5506[0],s5507[1]};
    assign in6501_2 = {c5480,s5476[3],s5507[0],c5508};
    CLA_4 KS_6501(s6501, c6501, in6501_1, in6501_2);
    wire[0:0] s6502, in6502_1, in6502_2;
    wire c6502;
    assign in6502_1 = {s5482[2]};
    assign in6502_2 = {c5484};
    Half_Adder KS_6502(s6502, c6502, in6502_1, in6502_2);
    wire[2:0] s6503, in6503_1, in6503_2;
    wire c6503;
    assign in6503_1 = {s5486[2],s5478[3],s5508[0]};
    assign in6503_2 = {c5488,c5482,s5509[0]};
    CLA_3 KS_6503(s6503, c6503, in6503_1, in6503_2);
    wire[0:0] s6504, in6504_1, in6504_2;
    wire c6504;
    assign in6504_1 = {c6485};
    assign in6504_2 = {c6486};
    Half_Adder KS_6504(s6504, c6504, in6504_1, in6504_2);
    wire[1:0] s6505, in6505_1, in6505_2;
    wire c6505;
    assign in6505_1 = {c6487,s5486[3]};
    assign in6505_2 = {c6488,s6496[1]};
    CLA_2 KS_6505(s6505, c6505, in6505_1, in6505_2);
    wire[0:0] s6506, in6506_1, in6506_2;
    wire c6506;
    assign in6506_1 = {c6490};
    assign in6506_2 = {s6496[0]};
    Full_Adder KS_6506(s6506, c6506, in6506_1, in6506_2, c6489);
    wire[3:0] s6507, in6507_1, in6507_2;
    wire c6507;
    assign in6507_1 = {s5490[2],s4024[0],s5519[0],s5520[1]};
    assign in6507_2 = {s5491[2],s5489[3],s5520[0],s5521[1]};
    CLA_4 KS_6507(s6507, c6507, in6507_1, in6507_2);
    wire[3:0] s6508, in6508_1, in6508_2;
    wire c6508;
    assign in6508_1 = {s5492[2],s5490[3],s5521[0],s5522[1]};
    assign in6508_2 = {s5493[2],s5491[3],s5522[0],c5523};
    CLA_4 KS_6508(s6508, c6508, in6508_1, in6508_2);
    wire[3:0] s6509, in6509_1, in6509_2;
    wire c6509;
    assign in6509_1 = {s5494[2],s5492[3],s5523[0],s5524[1]};
    assign in6509_2 = {s5495[2],s5493[3],s5524[0],c5525};
    CLA_4 KS_6509(s6509, c6509, in6509_1, in6509_2);
    wire[3:0] s6510, in6510_1, in6510_2;
    wire c6510;
    assign in6510_1 = {s5496[2],s5494[3],s5525[0],s5526[1]};
    assign in6510_2 = {s5497[2],s5495[3],s5526[0],c5527};
    CLA_4 KS_6510(s6510, c6510, in6510_1, in6510_2);
    wire[3:0] s6511, in6511_1, in6511_2;
    wire c6511;
    assign in6511_1 = {s5498[2],s5496[3],s5527[0],s5528[1]};
    assign in6511_2 = {s5499[2],s5497[3],s5528[0],c5529};
    CLA_4 KS_6511(s6511, c6511, in6511_1, in6511_2);
    wire[3:0] s6512, in6512_1, in6512_2;
    wire c6512;
    assign in6512_1 = {s5501[2],s5498[3],s5529[0],s5530[1]};
    assign in6512_2 = {c5503,s5499[3],s5530[0],c5531};
    CLA_4 KS_6512(s6512, c6512, in6512_1, in6512_2);
    wire[0:0] s6513, in6513_1, in6513_2;
    wire c6513;
    assign in6513_1 = {s5505[2]};
    assign in6513_2 = {c5507};
    Half_Adder KS_6513(s6513, c6513, in6513_1, in6513_2);
    wire[2:0] s6514, in6514_1, in6514_2;
    wire c6514;
    assign in6514_1 = {s5509[2],s5501[3],s5531[0]};
    assign in6514_2 = {c5511,c5505,s5532[0]};
    CLA_3 KS_6514(s6514, c6514, in6514_1, in6514_2);
    wire[0:0] s6515, in6515_1, in6515_2;
    wire c6515;
    assign in6515_1 = {c6496};
    assign in6515_2 = {c6497};
    Half_Adder KS_6515(s6515, c6515, in6515_1, in6515_2);
    wire[1:0] s6516, in6516_1, in6516_2;
    wire c6516;
    assign in6516_1 = {c6498,s5509[3]};
    assign in6516_2 = {c6499,s6507[1]};
    CLA_2 KS_6516(s6516, c6516, in6516_1, in6516_2);
    wire[0:0] s6517, in6517_1, in6517_2;
    wire c6517;
    assign in6517_1 = {c6501};
    assign in6517_2 = {s6507[0]};
    Full_Adder KS_6517(s6517, c6517, in6517_1, in6517_2, c6500);
    wire[3:0] s6518, in6518_1, in6518_2;
    wire c6518;
    assign in6518_1 = {s5513[2],s4060[0],s5542[0],s5542[1]};
    assign in6518_2 = {s5514[2],s5512[3],s5543[0],s5543[1]};
    CLA_4 KS_6518(s6518, c6518, in6518_1, in6518_2);
    wire[3:0] s6519, in6519_1, in6519_2;
    wire c6519;
    assign in6519_1 = {s5515[2],s5513[3],s5544[0],s5544[1]};
    assign in6519_2 = {s5516[2],s5514[3],s5545[0],s5545[1]};
    CLA_4 KS_6519(s6519, c6519, in6519_1, in6519_2);
    wire[3:0] s6520, in6520_1, in6520_2;
    wire c6520;
    assign in6520_1 = {s5517[2],s5515[3],s5546[0],s5546[1]};
    assign in6520_2 = {s5518[2],s5516[3],s5547[0],c5547};
    CLA_4 KS_6520(s6520, c6520, in6520_1, in6520_2);
    wire[3:0] s6521, in6521_1, in6521_2;
    wire c6521;
    assign in6521_1 = {s5519[2],s5517[3],s5548[0],s5548[1]};
    assign in6521_2 = {s5520[2],s5518[3],s5549[0],c5549};
    CLA_4 KS_6521(s6521, c6521, in6521_1, in6521_2);
    wire[3:0] s6522, in6522_1, in6522_2;
    wire c6522;
    assign in6522_1 = {s5521[2],s5519[3],s5550[0],s5550[1]};
    assign in6522_2 = {s5522[2],s5520[3],s5551[0],c5551};
    CLA_4 KS_6522(s6522, c6522, in6522_1, in6522_2);
    wire[3:0] s6523, in6523_1, in6523_2;
    wire c6523;
    assign in6523_1 = {s5524[2],s5521[3],s5552[0],s5552[1]};
    assign in6523_2 = {c5526,s5522[3],s5553[0],c5553};
    CLA_4 KS_6523(s6523, c6523, in6523_1, in6523_2);
    wire[0:0] s6524, in6524_1, in6524_2;
    wire c6524;
    assign in6524_1 = {s5528[2]};
    assign in6524_2 = {c5530};
    Half_Adder KS_6524(s6524, c6524, in6524_1, in6524_2);
    wire[3:0] s6525, in6525_1, in6525_2;
    wire c6525;
    assign in6525_1 = {s5532[2],s5524[3],s5554[0],s5554[1]};
    assign in6525_2 = {c5534,c5528,s5555[0],c5555};
    CLA_4 KS_6525(s6525, c6525, in6525_1, in6525_2);
    wire[0:0] s6526, in6526_1, in6526_2;
    wire c6526;
    assign in6526_1 = {c6507};
    assign in6526_2 = {c6508};
    Half_Adder KS_6526(s6526, c6526, in6526_1, in6526_2);
    wire[1:0] s6527, in6527_1, in6527_2;
    wire c6527;
    assign in6527_1 = {c6509,s5532[3]};
    assign in6527_2 = {c6510,s6518[1]};
    CLA_2 KS_6527(s6527, c6527, in6527_1, in6527_2);
    wire[0:0] s6528, in6528_1, in6528_2;
    wire c6528;
    assign in6528_1 = {c6512};
    assign in6528_2 = {s6518[0]};
    Full_Adder KS_6528(s6528, c6528, in6528_1, in6528_2, c6511);
    wire[3:0] s6529, in6529_1, in6529_2;
    wire c6529;
    assign in6529_1 = {s5536[2],s4096[0],s5565[0],s5565[1]};
    assign in6529_2 = {s5537[2],s5535[3],s5566[0],s5566[1]};
    CLA_4 KS_6529(s6529, c6529, in6529_1, in6529_2);
    wire[3:0] s6530, in6530_1, in6530_2;
    wire c6530;
    assign in6530_1 = {s5538[2],s5536[3],s5567[0],s5567[1]};
    assign in6530_2 = {s5539[2],s5537[3],s5568[0],s5568[1]};
    CLA_4 KS_6530(s6530, c6530, in6530_1, in6530_2);
    wire[3:0] s6531, in6531_1, in6531_2;
    wire c6531;
    assign in6531_1 = {s5540[2],s5538[3],s5569[0],s5569[1]};
    assign in6531_2 = {s5541[2],s5539[3],s5570[0],c5570};
    CLA_4 KS_6531(s6531, c6531, in6531_1, in6531_2);
    wire[3:0] s6532, in6532_1, in6532_2;
    wire c6532;
    assign in6532_1 = {s5542[2],s5540[3],s5571[0],s5571[1]};
    assign in6532_2 = {s5543[2],s5541[3],s5572[0],c5572};
    CLA_4 KS_6532(s6532, c6532, in6532_1, in6532_2);
    wire[3:0] s6533, in6533_1, in6533_2;
    wire c6533;
    assign in6533_1 = {s5544[2],s5542[3],s5573[0],s5573[1]};
    assign in6533_2 = {s5545[2],s5543[3],s5574[0],c5574};
    CLA_4 KS_6533(s6533, c6533, in6533_1, in6533_2);
    wire[3:0] s6534, in6534_1, in6534_2;
    wire c6534;
    assign in6534_1 = {s5546[2],s5544[3],s5575[0],s5575[1]};
    assign in6534_2 = {c5548,s5545[3],s5576[0],c5576};
    CLA_4 KS_6534(s6534, c6534, in6534_1, in6534_2);
    wire[0:0] s6535, in6535_1, in6535_2;
    wire c6535;
    assign in6535_1 = {s5550[2]};
    assign in6535_2 = {c5552};
    Half_Adder KS_6535(s6535, c6535, in6535_1, in6535_2);
    wire[3:0] s6536, in6536_1, in6536_2;
    wire c6536;
    assign in6536_1 = {s5554[2],s5546[3],s5577[0],s5577[1]};
    assign in6536_2 = {c5556,c5550,s5578[0],c5578};
    CLA_4 KS_6536(s6536, c6536, in6536_1, in6536_2);
    wire[0:0] s6537, in6537_1, in6537_2;
    wire c6537;
    assign in6537_1 = {c6518};
    assign in6537_2 = {c6519};
    Half_Adder KS_6537(s6537, c6537, in6537_1, in6537_2);
    wire[1:0] s6538, in6538_1, in6538_2;
    wire c6538;
    assign in6538_1 = {c6520,s5554[3]};
    assign in6538_2 = {c6521,s6529[1]};
    CLA_2 KS_6538(s6538, c6538, in6538_1, in6538_2);
    wire[0:0] s6539, in6539_1, in6539_2;
    wire c6539;
    assign in6539_1 = {c6522};
    assign in6539_2 = {c6523};
    Half_Adder KS_6539(s6539, c6539, in6539_1, in6539_2);
    wire[2:0] s6540, in6540_1, in6540_2;
    wire c6540;
    assign in6540_1 = {s6529[0],s6530[1],s5579[0]};
    assign in6540_2 = {s6530[0],s6531[1],s5580[0]};
    CLA_3_c KS_6540(s6540, c6540, in6540_1, in6540_2, c6525);
    wire[3:0] s6541, in6541_1, in6541_2;
    wire c6541;
    assign in6541_1 = {s5560[2],s4132[0],s5588[0],s5588[1]};
    assign in6541_2 = {s5561[2],s5558[3],s5589[0],s5589[1]};
    CLA_4 KS_6541(s6541, c6541, in6541_1, in6541_2);
    wire[3:0] s6542, in6542_1, in6542_2;
    wire c6542;
    assign in6542_1 = {s5562[2],s5559[3],s5590[0],s5590[1]};
    assign in6542_2 = {s5563[2],s5560[3],s5591[0],s5591[1]};
    CLA_4 KS_6542(s6542, c6542, in6542_1, in6542_2);
    wire[3:0] s6543, in6543_1, in6543_2;
    wire c6543;
    assign in6543_1 = {s5564[2],s5561[3],s5592[0],s5592[1]};
    assign in6543_2 = {s5565[2],s5562[3],s5593[0],c5593};
    CLA_4 KS_6543(s6543, c6543, in6543_1, in6543_2);
    wire[3:0] s6544, in6544_1, in6544_2;
    wire c6544;
    assign in6544_1 = {s5566[2],s5563[3],s5594[0],s5594[1]};
    assign in6544_2 = {s5567[2],s5564[3],s5595[0],c5595};
    CLA_4 KS_6544(s6544, c6544, in6544_1, in6544_2);
    wire[3:0] s6545, in6545_1, in6545_2;
    wire c6545;
    assign in6545_1 = {s5568[2],s5565[3],s5596[0],s5596[1]};
    assign in6545_2 = {c5569,s5566[3],s5597[0],c5597};
    CLA_4 KS_6545(s6545, c6545, in6545_1, in6545_2);
    wire[3:0] s6546, in6546_1, in6546_2;
    wire c6546;
    assign in6546_1 = {s5571[2],s5567[3],s5598[0],s5598[1]};
    assign in6546_2 = {c5573,s5568[3],s5599[0],c5599};
    CLA_4 KS_6546(s6546, c6546, in6546_1, in6546_2);
    wire[0:0] s6547, in6547_1, in6547_2;
    wire c6547;
    assign in6547_1 = {s5575[2]};
    assign in6547_2 = {c5577};
    Half_Adder KS_6547(s6547, c6547, in6547_1, in6547_2);
    wire[3:0] s6548, in6548_1, in6548_2;
    wire c6548;
    assign in6548_1 = {s5579[2],s5571[3],s5600[0],s5600[1]};
    assign in6548_2 = {c6529,c5575,s5601[0],c5601};
    CLA_4 KS_6548(s6548, c6548, in6548_1, in6548_2);
    wire[0:0] s6549, in6549_1, in6549_2;
    wire c6549;
    assign in6549_1 = {c6530};
    assign in6549_2 = {c6531};
    Half_Adder KS_6549(s6549, c6549, in6549_1, in6549_2);
    wire[1:0] s6550, in6550_1, in6550_2;
    wire c6550;
    assign in6550_1 = {c6532,s5579[3]};
    assign in6550_2 = {c6533,s6541[1]};
    CLA_2 KS_6550(s6550, c6550, in6550_1, in6550_2);
    wire[0:0] s6551, in6551_1, in6551_2;
    wire c6551;
    assign in6551_1 = {c6536};
    assign in6551_2 = {s6541[0]};
    Full_Adder KS_6551(s6551, c6551, in6551_1, in6551_2, c6534);
    wire[3:0] s6552, in6552_1, in6552_2;
    wire c6552;
    assign in6552_1 = {s5583[2],s4168[0],s5611[0],s5612[1]};
    assign in6552_2 = {s5584[2],s5581[3],s5612[0],s5613[1]};
    CLA_4 KS_6552(s6552, c6552, in6552_1, in6552_2);
    wire[3:0] s6553, in6553_1, in6553_2;
    wire c6553;
    assign in6553_1 = {s5585[2],s5582[3],s5613[0],s5614[1]};
    assign in6553_2 = {s5586[2],s5583[3],s5614[0],c5615};
    CLA_4 KS_6553(s6553, c6553, in6553_1, in6553_2);
    wire[3:0] s6554, in6554_1, in6554_2;
    wire c6554;
    assign in6554_1 = {s5587[2],s5584[3],s5615[0],s5616[1]};
    assign in6554_2 = {s5588[2],s5585[3],s5616[0],c5617};
    CLA_4 KS_6554(s6554, c6554, in6554_1, in6554_2);
    wire[3:0] s6555, in6555_1, in6555_2;
    wire c6555;
    assign in6555_1 = {s5589[2],s5586[3],s5617[0],s5618[1]};
    assign in6555_2 = {s5590[2],s5587[3],s5618[0],c5619};
    CLA_4 KS_6555(s6555, c6555, in6555_1, in6555_2);
    wire[3:0] s6556, in6556_1, in6556_2;
    wire c6556;
    assign in6556_1 = {s5591[2],s5588[3],s5619[0],s5620[1]};
    assign in6556_2 = {c5592,s5589[3],s5620[0],c5621};
    CLA_4 KS_6556(s6556, c6556, in6556_1, in6556_2);
    wire[3:0] s6557, in6557_1, in6557_2;
    wire c6557;
    assign in6557_1 = {s5594[2],s5590[3],s5621[0],s5622[1]};
    assign in6557_2 = {c5596,s5591[3],s5622[0],c5623};
    CLA_4 KS_6557(s6557, c6557, in6557_1, in6557_2);
    wire[0:0] s6558, in6558_1, in6558_2;
    wire c6558;
    assign in6558_1 = {s5598[2]};
    assign in6558_2 = {c5600};
    Half_Adder KS_6558(s6558, c6558, in6558_1, in6558_2);
    wire[2:0] s6559, in6559_1, in6559_2;
    wire c6559;
    assign in6559_1 = {s5602[2],s5594[3],s5623[0]};
    assign in6559_2 = {c6541,c5598,s5624[0]};
    CLA_3 KS_6559(s6559, c6559, in6559_1, in6559_2);
    wire[0:0] s6560, in6560_1, in6560_2;
    wire c6560;
    assign in6560_1 = {c6542};
    assign in6560_2 = {c6543};
    Half_Adder KS_6560(s6560, c6560, in6560_1, in6560_2);
    wire[1:0] s6561, in6561_1, in6561_2;
    wire c6561;
    assign in6561_1 = {c6544,s5602[3]};
    assign in6561_2 = {c6545,s6552[1]};
    CLA_2 KS_6561(s6561, c6561, in6561_1, in6561_2);
    wire[0:0] s6562, in6562_1, in6562_2;
    wire c6562;
    assign in6562_1 = {c6548};
    assign in6562_2 = {s6552[0]};
    Full_Adder KS_6562(s6562, c6562, in6562_1, in6562_2, c6546);
    wire[3:0] s6563, in6563_1, in6563_2;
    wire c6563;
    assign in6563_1 = {s5606[2],s4206[0],s5634[0],s5635[1]};
    assign in6563_2 = {s5607[2],s5604[3],s5635[0],s5636[1]};
    CLA_4 KS_6563(s6563, c6563, in6563_1, in6563_2);
    wire[3:0] s6564, in6564_1, in6564_2;
    wire c6564;
    assign in6564_1 = {s5608[2],s5605[3],s5636[0],s5637[1]};
    assign in6564_2 = {s5609[2],s5606[3],s5637[0],c5638};
    CLA_4 KS_6564(s6564, c6564, in6564_1, in6564_2);
    wire[3:0] s6565, in6565_1, in6565_2;
    wire c6565;
    assign in6565_1 = {s5610[2],s5607[3],s5638[0],s5639[1]};
    assign in6565_2 = {s5611[2],s5608[3],s5639[0],c5640};
    CLA_4 KS_6565(s6565, c6565, in6565_1, in6565_2);
    wire[3:0] s6566, in6566_1, in6566_2;
    wire c6566;
    assign in6566_1 = {s5612[2],s5609[3],s5640[0],s5641[1]};
    assign in6566_2 = {s5613[2],s5610[3],s5641[0],c5642};
    CLA_4 KS_6566(s6566, c6566, in6566_1, in6566_2);
    wire[3:0] s6567, in6567_1, in6567_2;
    wire c6567;
    assign in6567_1 = {s5614[2],s5611[3],s5642[0],s5643[1]};
    assign in6567_2 = {c5616,s5612[3],s5643[0],c5644};
    CLA_4 KS_6567(s6567, c6567, in6567_1, in6567_2);
    wire[3:0] s6568, in6568_1, in6568_2;
    wire c6568;
    assign in6568_1 = {s5618[2],s5613[3],s5644[0],s5645[1]};
    assign in6568_2 = {c5620,s5614[3],s5645[0],c5646};
    CLA_4 KS_6568(s6568, c6568, in6568_1, in6568_2);
    wire[0:0] s6569, in6569_1, in6569_2;
    wire c6569;
    assign in6569_1 = {s5622[2]};
    assign in6569_2 = {c5624};
    Half_Adder KS_6569(s6569, c6569, in6569_1, in6569_2);
    wire[2:0] s6570, in6570_1, in6570_2;
    wire c6570;
    assign in6570_1 = {s5626[2],s5618[3],s5646[0]};
    assign in6570_2 = {c6552,c5622,s5647[0]};
    CLA_3 KS_6570(s6570, c6570, in6570_1, in6570_2);
    wire[0:0] s6571, in6571_1, in6571_2;
    wire c6571;
    assign in6571_1 = {c6553};
    assign in6571_2 = {c6554};
    Half_Adder KS_6571(s6571, c6571, in6571_1, in6571_2);
    wire[1:0] s6572, in6572_1, in6572_2;
    wire c6572;
    assign in6572_1 = {c6556,s5626[3]};
    assign in6572_2 = {c6557,s6563[1]};
    CLA_2_c KS_6572(s6572, c6572, in6572_1, in6572_2, c6555);
    wire[3:0] s6573, in6573_1, in6573_2;
    wire c6573;
    assign in6573_1 = {s5629[2],s4244[0],s5657[0],s5658[1]};
    assign in6573_2 = {s5630[2],s5627[3],s5658[0],s5659[1]};
    CLA_4 KS_6573(s6573, c6573, in6573_1, in6573_2);
    wire[3:0] s6574, in6574_1, in6574_2;
    wire c6574;
    assign in6574_1 = {s5631[2],s5628[3],s5659[0],s5660[1]};
    assign in6574_2 = {s5632[2],s5629[3],s5660[0],c5661};
    CLA_4 KS_6574(s6574, c6574, in6574_1, in6574_2);
    wire[3:0] s6575, in6575_1, in6575_2;
    wire c6575;
    assign in6575_1 = {s5633[2],s5630[3],s5661[0],s5662[1]};
    assign in6575_2 = {s5634[2],s5631[3],s5662[0],c5663};
    CLA_4 KS_6575(s6575, c6575, in6575_1, in6575_2);
    wire[3:0] s6576, in6576_1, in6576_2;
    wire c6576;
    assign in6576_1 = {s5635[2],s5632[3],s5663[0],s5664[1]};
    assign in6576_2 = {s5636[2],s5633[3],s5664[0],c5665};
    CLA_4 KS_6576(s6576, c6576, in6576_1, in6576_2);
    wire[3:0] s6577, in6577_1, in6577_2;
    wire c6577;
    assign in6577_1 = {s5637[2],s5634[3],s5665[0],s5666[1]};
    assign in6577_2 = {c5639,s5635[3],s5666[0],c5667};
    CLA_4 KS_6577(s6577, c6577, in6577_1, in6577_2);
    wire[3:0] s6578, in6578_1, in6578_2;
    wire c6578;
    assign in6578_1 = {s5641[2],s5636[3],s5667[0],s5668[1]};
    assign in6578_2 = {c5643,s5637[3],s5668[0],c5669};
    CLA_4 KS_6578(s6578, c6578, in6578_1, in6578_2);
    wire[0:0] s6579, in6579_1, in6579_2;
    wire c6579;
    assign in6579_1 = {s5645[2]};
    assign in6579_2 = {c5647};
    Half_Adder KS_6579(s6579, c6579, in6579_1, in6579_2);
    wire[2:0] s6580, in6580_1, in6580_2;
    wire c6580;
    assign in6580_1 = {s5649[2],s5641[3],s5669[0]};
    assign in6580_2 = {c6563,c5645,s5670[0]};
    CLA_3 KS_6580(s6580, c6580, in6580_1, in6580_2);
    wire[0:0] s6581, in6581_1, in6581_2;
    wire c6581;
    assign in6581_1 = {c6564};
    assign in6581_2 = {c6565};
    Half_Adder KS_6581(s6581, c6581, in6581_1, in6581_2);
    wire[1:0] s6582, in6582_1, in6582_2;
    wire c6582;
    assign in6582_1 = {c6567,s5649[3]};
    assign in6582_2 = {c6568,s6573[1]};
    CLA_2_c KS_6582(s6582, c6582, in6582_1, in6582_2, c6566);
    wire[3:0] s6583, in6583_1, in6583_2;
    wire c6583;
    assign in6583_1 = {s5651[2],s4280[0],s5680[0],s5681[1]};
    assign in6583_2 = {s5652[2],s5650[3],s5681[0],s5682[1]};
    CLA_4 KS_6583(s6583, c6583, in6583_1, in6583_2);
    wire[3:0] s6584, in6584_1, in6584_2;
    wire c6584;
    assign in6584_1 = {s5653[2],s5651[3],s5682[0],s5683[1]};
    assign in6584_2 = {s5654[2],s5652[3],s5683[0],c5684};
    CLA_4 KS_6584(s6584, c6584, in6584_1, in6584_2);
    wire[3:0] s6585, in6585_1, in6585_2;
    wire c6585;
    assign in6585_1 = {s5655[2],s5653[3],s5684[0],s5685[1]};
    assign in6585_2 = {s5656[2],s5654[3],s5685[0],c5686};
    CLA_4 KS_6585(s6585, c6585, in6585_1, in6585_2);
    wire[3:0] s6586, in6586_1, in6586_2;
    wire c6586;
    assign in6586_1 = {s5657[2],s5655[3],s5686[0],s5687[1]};
    assign in6586_2 = {s5658[2],s5656[3],s5687[0],c5688};
    CLA_4 KS_6586(s6586, c6586, in6586_1, in6586_2);
    wire[3:0] s6587, in6587_1, in6587_2;
    wire c6587;
    assign in6587_1 = {s5659[2],s5657[3],s5688[0],s5689[1]};
    assign in6587_2 = {s5660[2],s5658[3],s5689[0],c5690};
    CLA_4 KS_6587(s6587, c6587, in6587_1, in6587_2);
    wire[3:0] s6588, in6588_1, in6588_2;
    wire c6588;
    assign in6588_1 = {s5662[2],s5659[3],s5690[0],s5691[1]};
    assign in6588_2 = {c5664,s5660[3],s5691[0],c5692};
    CLA_4 KS_6588(s6588, c6588, in6588_1, in6588_2);
    wire[0:0] s6589, in6589_1, in6589_2;
    wire c6589;
    assign in6589_1 = {s5666[2]};
    assign in6589_2 = {c5668};
    Half_Adder KS_6589(s6589, c6589, in6589_1, in6589_2);
    wire[2:0] s6590, in6590_1, in6590_2;
    wire c6590;
    assign in6590_1 = {s5670[2],s5662[3],s5692[0]};
    assign in6590_2 = {c5672,c5666,s5693[0]};
    CLA_3 KS_6590(s6590, c6590, in6590_1, in6590_2);
    wire[0:0] s6591, in6591_1, in6591_2;
    wire c6591;
    assign in6591_1 = {c6573};
    assign in6591_2 = {c6574};
    Half_Adder KS_6591(s6591, c6591, in6591_1, in6591_2);
    wire[1:0] s6592, in6592_1, in6592_2;
    wire c6592;
    assign in6592_1 = {c6575,s5670[3]};
    assign in6592_2 = {c6576,s6583[1]};
    CLA_2 KS_6592(s6592, c6592, in6592_1, in6592_2);
    wire[0:0] s6593, in6593_1, in6593_2;
    wire c6593;
    assign in6593_1 = {c6578};
    assign in6593_2 = {s6583[0]};
    Full_Adder KS_6593(s6593, c6593, in6593_1, in6593_2, c6577);
    wire[3:0] s6594, in6594_1, in6594_2;
    wire c6594;
    assign in6594_1 = {s5674[2],s4316[0],s5703[0],s5704[1]};
    assign in6594_2 = {s5675[2],s5673[3],s5704[0],s5705[1]};
    CLA_4 KS_6594(s6594, c6594, in6594_1, in6594_2);
    wire[3:0] s6595, in6595_1, in6595_2;
    wire c6595;
    assign in6595_1 = {s5676[2],s5674[3],s5705[0],s5706[1]};
    assign in6595_2 = {s5677[2],s5675[3],s5706[0],c5707};
    CLA_4 KS_6595(s6595, c6595, in6595_1, in6595_2);
    wire[3:0] s6596, in6596_1, in6596_2;
    wire c6596;
    assign in6596_1 = {s5678[2],s5676[3],s5707[0],s5708[1]};
    assign in6596_2 = {s5679[2],s5677[3],s5708[0],c5709};
    CLA_4 KS_6596(s6596, c6596, in6596_1, in6596_2);
    wire[3:0] s6597, in6597_1, in6597_2;
    wire c6597;
    assign in6597_1 = {s5680[2],s5678[3],s5709[0],s5710[1]};
    assign in6597_2 = {s5681[2],s5679[3],s5710[0],c5711};
    CLA_4 KS_6597(s6597, c6597, in6597_1, in6597_2);
    wire[3:0] s6598, in6598_1, in6598_2;
    wire c6598;
    assign in6598_1 = {s5682[2],s5680[3],s5711[0],s5712[1]};
    assign in6598_2 = {s5683[2],s5681[3],s5712[0],c5713};
    CLA_4 KS_6598(s6598, c6598, in6598_1, in6598_2);
    wire[3:0] s6599, in6599_1, in6599_2;
    wire c6599;
    assign in6599_1 = {s5685[2],s5682[3],s5713[0],s5714[1]};
    assign in6599_2 = {c5687,s5683[3],s5714[0],c5715};
    CLA_4 KS_6599(s6599, c6599, in6599_1, in6599_2);
    wire[0:0] s6600, in6600_1, in6600_2;
    wire c6600;
    assign in6600_1 = {s5689[2]};
    assign in6600_2 = {c5691};
    Half_Adder KS_6600(s6600, c6600, in6600_1, in6600_2);
    wire[2:0] s6601, in6601_1, in6601_2;
    wire c6601;
    assign in6601_1 = {s5693[2],s5685[3],s5715[0]};
    assign in6601_2 = {c5695,c5689,s5716[0]};
    CLA_3 KS_6601(s6601, c6601, in6601_1, in6601_2);
    wire[0:0] s6602, in6602_1, in6602_2;
    wire c6602;
    assign in6602_1 = {c6583};
    assign in6602_2 = {c6584};
    Half_Adder KS_6602(s6602, c6602, in6602_1, in6602_2);
    wire[1:0] s6603, in6603_1, in6603_2;
    wire c6603;
    assign in6603_1 = {c6585,s5693[3]};
    assign in6603_2 = {c6586,s6594[1]};
    CLA_2 KS_6603(s6603, c6603, in6603_1, in6603_2);
    wire[0:0] s6604, in6604_1, in6604_2;
    wire c6604;
    assign in6604_1 = {c6588};
    assign in6604_2 = {s6594[0]};
    Full_Adder KS_6604(s6604, c6604, in6604_1, in6604_2, c6587);
    wire[3:0] s6605, in6605_1, in6605_2;
    wire c6605;
    assign in6605_1 = {s5698[2],s4354[0],s5726[0],s5727[1]};
    assign in6605_2 = {s5699[2],s5696[3],s5727[0],s5728[1]};
    CLA_4 KS_6605(s6605, c6605, in6605_1, in6605_2);
    wire[3:0] s6606, in6606_1, in6606_2;
    wire c6606;
    assign in6606_1 = {s5700[2],s5697[3],s5728[0],s5729[1]};
    assign in6606_2 = {s5701[2],s5698[3],s5729[0],c5730};
    CLA_4 KS_6606(s6606, c6606, in6606_1, in6606_2);
    wire[3:0] s6607, in6607_1, in6607_2;
    wire c6607;
    assign in6607_1 = {s5702[2],s5699[3],s5730[0],s5731[1]};
    assign in6607_2 = {s5703[2],s5700[3],s5731[0],c5732};
    CLA_4 KS_6607(s6607, c6607, in6607_1, in6607_2);
    wire[3:0] s6608, in6608_1, in6608_2;
    wire c6608;
    assign in6608_1 = {s5704[2],s5701[3],s5732[0],s5733[1]};
    assign in6608_2 = {s5705[2],s5702[3],s5733[0],c5734};
    CLA_4 KS_6608(s6608, c6608, in6608_1, in6608_2);
    wire[3:0] s6609, in6609_1, in6609_2;
    wire c6609;
    assign in6609_1 = {s5706[2],s5703[3],s5734[0],s5735[1]};
    assign in6609_2 = {c5708,s5704[3],s5735[0],c5736};
    CLA_4 KS_6609(s6609, c6609, in6609_1, in6609_2);
    wire[3:0] s6610, in6610_1, in6610_2;
    wire c6610;
    assign in6610_1 = {s5710[2],s5705[3],s5736[0],s5737[1]};
    assign in6610_2 = {c5712,s5706[3],s5737[0],c5738};
    CLA_4 KS_6610(s6610, c6610, in6610_1, in6610_2);
    wire[0:0] s6611, in6611_1, in6611_2;
    wire c6611;
    assign in6611_1 = {s5714[2]};
    assign in6611_2 = {c5716};
    Half_Adder KS_6611(s6611, c6611, in6611_1, in6611_2);
    wire[2:0] s6612, in6612_1, in6612_2;
    wire c6612;
    assign in6612_1 = {s5718[2],s5710[3],s5738[0]};
    assign in6612_2 = {c6594,c5714,s5739[0]};
    CLA_3 KS_6612(s6612, c6612, in6612_1, in6612_2);
    wire[0:0] s6613, in6613_1, in6613_2;
    wire c6613;
    assign in6613_1 = {c6595};
    assign in6613_2 = {c6596};
    Half_Adder KS_6613(s6613, c6613, in6613_1, in6613_2);
    wire[1:0] s6614, in6614_1, in6614_2;
    wire c6614;
    assign in6614_1 = {c6598,s5718[3]};
    assign in6614_2 = {c6599,s6605[1]};
    CLA_2_c KS_6614(s6614, c6614, in6614_1, in6614_2, c6597);
    wire[3:0] s6615, in6615_1, in6615_2;
    wire c6615;
    assign in6615_1 = {s5720[2],s4390[0],s5749[0],s5750[1]};
    assign in6615_2 = {s5721[2],s5719[3],s5750[0],s5751[1]};
    CLA_4 KS_6615(s6615, c6615, in6615_1, in6615_2);
    wire[3:0] s6616, in6616_1, in6616_2;
    wire c6616;
    assign in6616_1 = {s5722[2],s5720[3],s5751[0],s5752[1]};
    assign in6616_2 = {s5723[2],s5721[3],s5752[0],c5753};
    CLA_4 KS_6616(s6616, c6616, in6616_1, in6616_2);
    wire[3:0] s6617, in6617_1, in6617_2;
    wire c6617;
    assign in6617_1 = {s5724[2],s5722[3],s5753[0],s5754[1]};
    assign in6617_2 = {s5725[2],s5723[3],s5754[0],c5755};
    CLA_4 KS_6617(s6617, c6617, in6617_1, in6617_2);
    wire[3:0] s6618, in6618_1, in6618_2;
    wire c6618;
    assign in6618_1 = {s5726[2],s5724[3],s5755[0],s5756[1]};
    assign in6618_2 = {s5727[2],s5725[3],s5756[0],c5757};
    CLA_4 KS_6618(s6618, c6618, in6618_1, in6618_2);
    wire[3:0] s6619, in6619_1, in6619_2;
    wire c6619;
    assign in6619_1 = {s5728[2],s5726[3],s5757[0],s5758[1]};
    assign in6619_2 = {s5729[2],s5727[3],s5758[0],c5759};
    CLA_4 KS_6619(s6619, c6619, in6619_1, in6619_2);
    wire[3:0] s6620, in6620_1, in6620_2;
    wire c6620;
    assign in6620_1 = {s5731[2],s5728[3],s5759[0],s5760[1]};
    assign in6620_2 = {c5733,s5729[3],s5760[0],c5761};
    CLA_4 KS_6620(s6620, c6620, in6620_1, in6620_2);
    wire[0:0] s6621, in6621_1, in6621_2;
    wire c6621;
    assign in6621_1 = {s5735[2]};
    assign in6621_2 = {c5737};
    Half_Adder KS_6621(s6621, c6621, in6621_1, in6621_2);
    wire[2:0] s6622, in6622_1, in6622_2;
    wire c6622;
    assign in6622_1 = {s5739[2],s5731[3],s5761[0]};
    assign in6622_2 = {c5741,c5735,s5762[0]};
    CLA_3 KS_6622(s6622, c6622, in6622_1, in6622_2);
    wire[0:0] s6623, in6623_1, in6623_2;
    wire c6623;
    assign in6623_1 = {c6605};
    assign in6623_2 = {c6606};
    Half_Adder KS_6623(s6623, c6623, in6623_1, in6623_2);
    wire[1:0] s6624, in6624_1, in6624_2;
    wire c6624;
    assign in6624_1 = {c6607,s5739[3]};
    assign in6624_2 = {c6608,s6615[1]};
    CLA_2 KS_6624(s6624, c6624, in6624_1, in6624_2);
    wire[0:0] s6625, in6625_1, in6625_2;
    wire c6625;
    assign in6625_1 = {c6610};
    assign in6625_2 = {s6615[0]};
    Full_Adder KS_6625(s6625, c6625, in6625_1, in6625_2, c6609);
    wire[3:0] s6626, in6626_1, in6626_2;
    wire c6626;
    assign in6626_1 = {s5744[2],s4428[0],s5772[0],s5773[1]};
    assign in6626_2 = {s5745[2],s5742[3],s5773[0],s5774[1]};
    CLA_4 KS_6626(s6626, c6626, in6626_1, in6626_2);
    wire[3:0] s6627, in6627_1, in6627_2;
    wire c6627;
    assign in6627_1 = {s5746[2],s5743[3],s5774[0],s5775[1]};
    assign in6627_2 = {s5747[2],s5744[3],s5775[0],c5776};
    CLA_4 KS_6627(s6627, c6627, in6627_1, in6627_2);
    wire[3:0] s6628, in6628_1, in6628_2;
    wire c6628;
    assign in6628_1 = {s5748[2],s5745[3],s5776[0],s5777[1]};
    assign in6628_2 = {s5749[2],s5746[3],s5777[0],c5778};
    CLA_4 KS_6628(s6628, c6628, in6628_1, in6628_2);
    wire[3:0] s6629, in6629_1, in6629_2;
    wire c6629;
    assign in6629_1 = {s5750[2],s5747[3],s5778[0],s5779[1]};
    assign in6629_2 = {s5751[2],s5748[3],s5779[0],c5780};
    CLA_4 KS_6629(s6629, c6629, in6629_1, in6629_2);
    wire[3:0] s6630, in6630_1, in6630_2;
    wire c6630;
    assign in6630_1 = {s5752[2],s5749[3],s5780[0],s5781[1]};
    assign in6630_2 = {c5754,s5750[3],s5781[0],c5782};
    CLA_4 KS_6630(s6630, c6630, in6630_1, in6630_2);
    wire[3:0] s6631, in6631_1, in6631_2;
    wire c6631;
    assign in6631_1 = {s5756[2],s5751[3],s5782[0],s5783[1]};
    assign in6631_2 = {c5758,s5752[3],s5783[0],c5784};
    CLA_4 KS_6631(s6631, c6631, in6631_1, in6631_2);
    wire[0:0] s6632, in6632_1, in6632_2;
    wire c6632;
    assign in6632_1 = {s5760[2]};
    assign in6632_2 = {c5762};
    Half_Adder KS_6632(s6632, c6632, in6632_1, in6632_2);
    wire[2:0] s6633, in6633_1, in6633_2;
    wire c6633;
    assign in6633_1 = {s5764[2],s5756[3],s5784[0]};
    assign in6633_2 = {c6615,c5760,s5785[0]};
    CLA_3 KS_6633(s6633, c6633, in6633_1, in6633_2);
    wire[0:0] s6634, in6634_1, in6634_2;
    wire c6634;
    assign in6634_1 = {c6616};
    assign in6634_2 = {c6617};
    Half_Adder KS_6634(s6634, c6634, in6634_1, in6634_2);
    wire[1:0] s6635, in6635_1, in6635_2;
    wire c6635;
    assign in6635_1 = {c6619,s5764[3]};
    assign in6635_2 = {c6620,s6626[1]};
    CLA_2_c KS_6635(s6635, c6635, in6635_1, in6635_2, c6618);
    wire[3:0] s6636, in6636_1, in6636_2;
    wire c6636;
    assign in6636_1 = {s5766[2],s4464[0],s5795[0],s5795[1]};
    assign in6636_2 = {s5767[2],s5765[3],s5796[0],s5796[1]};
    CLA_4 KS_6636(s6636, c6636, in6636_1, in6636_2);
    wire[3:0] s6637, in6637_1, in6637_2;
    wire c6637;
    assign in6637_1 = {s5768[2],s5766[3],s5797[0],s5797[1]};
    assign in6637_2 = {s5769[2],s5767[3],s5798[0],s5798[1]};
    CLA_4 KS_6637(s6637, c6637, in6637_1, in6637_2);
    wire[3:0] s6638, in6638_1, in6638_2;
    wire c6638;
    assign in6638_1 = {s5770[2],s5768[3],s5799[0],s5799[1]};
    assign in6638_2 = {s5771[2],s5769[3],s5800[0],c5800};
    CLA_4 KS_6638(s6638, c6638, in6638_1, in6638_2);
    wire[3:0] s6639, in6639_1, in6639_2;
    wire c6639;
    assign in6639_1 = {s5772[2],s5770[3],s5801[0],s5801[1]};
    assign in6639_2 = {s5773[2],s5771[3],s5802[0],c5802};
    CLA_4 KS_6639(s6639, c6639, in6639_1, in6639_2);
    wire[3:0] s6640, in6640_1, in6640_2;
    wire c6640;
    assign in6640_1 = {s5774[2],s5772[3],s5803[0],s5803[1]};
    assign in6640_2 = {s5775[2],s5773[3],s5804[0],c5804};
    CLA_4 KS_6640(s6640, c6640, in6640_1, in6640_2);
    wire[3:0] s6641, in6641_1, in6641_2;
    wire c6641;
    assign in6641_1 = {s5777[2],s5774[3],s5805[0],s5805[1]};
    assign in6641_2 = {c5779,s5775[3],s5806[0],c5806};
    CLA_4 KS_6641(s6641, c6641, in6641_1, in6641_2);
    wire[0:0] s6642, in6642_1, in6642_2;
    wire c6642;
    assign in6642_1 = {s5781[2]};
    assign in6642_2 = {c5783};
    Half_Adder KS_6642(s6642, c6642, in6642_1, in6642_2);
    wire[3:0] s6643, in6643_1, in6643_2;
    wire c6643;
    assign in6643_1 = {s5785[2],s5777[3],s5807[0],s5807[1]};
    assign in6643_2 = {c5787,c5781,s5808[0],c5808};
    CLA_4 KS_6643(s6643, c6643, in6643_1, in6643_2);
    wire[0:0] s6644, in6644_1, in6644_2;
    wire c6644;
    assign in6644_1 = {c6626};
    assign in6644_2 = {c6627};
    Half_Adder KS_6644(s6644, c6644, in6644_1, in6644_2);
    wire[1:0] s6645, in6645_1, in6645_2;
    wire c6645;
    assign in6645_1 = {c6628,s5785[3]};
    assign in6645_2 = {c6629,s6636[1]};
    CLA_2 KS_6645(s6645, c6645, in6645_1, in6645_2);
    wire[0:0] s6646, in6646_1, in6646_2;
    wire c6646;
    assign in6646_1 = {c6631};
    assign in6646_2 = {s6636[0]};
    Full_Adder KS_6646(s6646, c6646, in6646_1, in6646_2, c6630);
    wire[3:0] s6647, in6647_1, in6647_2;
    wire c6647;
    assign in6647_1 = {s5789[2],s4501[0],s5817[0],s5818[1]};
    assign in6647_2 = {s5790[2],s5788[3],s5818[0],s5819[1]};
    CLA_4 KS_6647(s6647, c6647, in6647_1, in6647_2);
    wire[3:0] s6648, in6648_1, in6648_2;
    wire c6648;
    assign in6648_1 = {s5791[2],s5789[3],s5819[0],s5820[1]};
    assign in6648_2 = {s5792[2],s5790[3],s5820[0],s5821[1]};
    CLA_4 KS_6648(s6648, c6648, in6648_1, in6648_2);
    wire[3:0] s6649, in6649_1, in6649_2;
    wire c6649;
    assign in6649_1 = {s5793[2],s5791[3],s5821[0],s5822[1]};
    assign in6649_2 = {s5794[2],s5792[3],s5822[0],c5823};
    CLA_4 KS_6649(s6649, c6649, in6649_1, in6649_2);
    wire[3:0] s6650, in6650_1, in6650_2;
    wire c6650;
    assign in6650_1 = {s5795[2],s5793[3],s5823[0],s5824[1]};
    assign in6650_2 = {s5796[2],s5794[3],s5824[0],c5825};
    CLA_4 KS_6650(s6650, c6650, in6650_1, in6650_2);
    wire[3:0] s6651, in6651_1, in6651_2;
    wire c6651;
    assign in6651_1 = {s5797[2],s5795[3],s5825[0],s5826[1]};
    assign in6651_2 = {s5798[2],s5796[3],s5826[0],c5827};
    CLA_4 KS_6651(s6651, c6651, in6651_1, in6651_2);
    wire[3:0] s6652, in6652_1, in6652_2;
    wire c6652;
    assign in6652_1 = {s5799[2],s5797[3],s5827[0],s5828[1]};
    assign in6652_2 = {c5801,s5798[3],s5828[0],c5829};
    CLA_4 KS_6652(s6652, c6652, in6652_1, in6652_2);
    wire[0:0] s6653, in6653_1, in6653_2;
    wire c6653;
    assign in6653_1 = {s5803[2]};
    assign in6653_2 = {c5805};
    Half_Adder KS_6653(s6653, c6653, in6653_1, in6653_2);
    wire[2:0] s6654, in6654_1, in6654_2;
    wire c6654;
    assign in6654_1 = {s5807[2],s5799[3],s5829[0]};
    assign in6654_2 = {c5809,c5803,s5830[0]};
    CLA_3 KS_6654(s6654, c6654, in6654_1, in6654_2);
    wire[0:0] s6655, in6655_1, in6655_2;
    wire c6655;
    assign in6655_1 = {c6636};
    assign in6655_2 = {c6637};
    Half_Adder KS_6655(s6655, c6655, in6655_1, in6655_2);
    wire[1:0] s6656, in6656_1, in6656_2;
    wire c6656;
    assign in6656_1 = {c6638,s5807[3]};
    assign in6656_2 = {c6639,s6647[1]};
    CLA_2 KS_6656(s6656, c6656, in6656_1, in6656_2);
    wire[0:0] s6657, in6657_1, in6657_2;
    wire c6657;
    assign in6657_1 = {c6640};
    assign in6657_2 = {c6641};
    Half_Adder KS_6657(s6657, c6657, in6657_1, in6657_2);
    wire[3:0] s6658, in6658_1, in6658_2;
    wire c6658;
    assign in6658_1 = {s6647[0],s6648[1],s5831[0],s5830[1]};
    assign in6658_2 = {s6648[0],s6649[1],s5832[0],c5831};
    CLA_4_c KS_6658(s6658, c6658, in6658_1, in6658_2, c6643);
    wire[3:0] s6659, in6659_1, in6659_2;
    wire c6659;
    assign in6659_1 = {s5813[2],s4539[0],s5840[0],s5840[1]};
    assign in6659_2 = {s5814[2],s5811[3],s5841[0],s5841[1]};
    CLA_4 KS_6659(s6659, c6659, in6659_1, in6659_2);
    wire[3:0] s6660, in6660_1, in6660_2;
    wire c6660;
    assign in6660_1 = {s5815[2],s5812[3],s5842[0],s5842[1]};
    assign in6660_2 = {s5816[2],s5813[3],s5843[0],s5843[1]};
    CLA_4 KS_6660(s6660, c6660, in6660_1, in6660_2);
    wire[3:0] s6661, in6661_1, in6661_2;
    wire c6661;
    assign in6661_1 = {s5817[2],s5814[3],s5844[0],s5844[1]};
    assign in6661_2 = {s5818[2],s5815[3],s5845[0],c5845};
    CLA_4 KS_6661(s6661, c6661, in6661_1, in6661_2);
    wire[3:0] s6662, in6662_1, in6662_2;
    wire c6662;
    assign in6662_1 = {s5819[2],s5816[3],s5846[0],s5846[1]};
    assign in6662_2 = {s5820[2],s5817[3],s5847[0],c5847};
    CLA_4 KS_6662(s6662, c6662, in6662_1, in6662_2);
    wire[3:0] s6663, in6663_1, in6663_2;
    wire c6663;
    assign in6663_1 = {s5821[2],s5818[3],s5848[0],s5848[1]};
    assign in6663_2 = {c5822,s5819[3],s5849[0],c5849};
    CLA_4 KS_6663(s6663, c6663, in6663_1, in6663_2);
    wire[3:0] s6664, in6664_1, in6664_2;
    wire c6664;
    assign in6664_1 = {s5824[2],s5820[3],s5850[0],s5850[1]};
    assign in6664_2 = {c5826,s5821[3],s5851[0],c5851};
    CLA_4 KS_6664(s6664, c6664, in6664_1, in6664_2);
    wire[0:0] s6665, in6665_1, in6665_2;
    wire c6665;
    assign in6665_1 = {s5828[2]};
    assign in6665_2 = {c5830};
    Half_Adder KS_6665(s6665, c6665, in6665_1, in6665_2);
    wire[3:0] s6666, in6666_1, in6666_2;
    wire c6666;
    assign in6666_1 = {s5832[2],s5824[3],s5852[0],s5852[1]};
    assign in6666_2 = {c6647,c5828,s5853[0],c5853};
    CLA_4 KS_6666(s6666, c6666, in6666_1, in6666_2);
    wire[0:0] s6667, in6667_1, in6667_2;
    wire c6667;
    assign in6667_1 = {c6648};
    assign in6667_2 = {c6649};
    Half_Adder KS_6667(s6667, c6667, in6667_1, in6667_2);
    wire[1:0] s6668, in6668_1, in6668_2;
    wire c6668;
    assign in6668_1 = {c6650,s5832[3]};
    assign in6668_2 = {c6651,s6659[1]};
    CLA_2 KS_6668(s6668, c6668, in6668_1, in6668_2);
    wire[0:0] s6669, in6669_1, in6669_2;
    wire c6669;
    assign in6669_1 = {c6658};
    assign in6669_2 = {s6659[0]};
    Full_Adder KS_6669(s6669, c6669, in6669_1, in6669_2, c6652);
    wire[3:0] s6670, in6670_1, in6670_2;
    wire c6670;
    assign in6670_1 = {s5834[2],s4575[0],s5863[0],s5864[1]};
    assign in6670_2 = {s5835[2],s5833[3],s5864[0],s5865[1]};
    CLA_4 KS_6670(s6670, c6670, in6670_1, in6670_2);
    wire[3:0] s6671, in6671_1, in6671_2;
    wire c6671;
    assign in6671_1 = {s5836[2],s5834[3],s5865[0],s5866[1]};
    assign in6671_2 = {s5837[2],s5835[3],s5866[0],c5867};
    CLA_4 KS_6671(s6671, c6671, in6671_1, in6671_2);
    wire[3:0] s6672, in6672_1, in6672_2;
    wire c6672;
    assign in6672_1 = {s5838[2],s5836[3],s5867[0],s5868[1]};
    assign in6672_2 = {s5839[2],s5837[3],s5868[0],c5869};
    CLA_4 KS_6672(s6672, c6672, in6672_1, in6672_2);
    wire[3:0] s6673, in6673_1, in6673_2;
    wire c6673;
    assign in6673_1 = {s5840[2],s5838[3],s5869[0],s5870[1]};
    assign in6673_2 = {s5841[2],s5839[3],s5870[0],c5871};
    CLA_4 KS_6673(s6673, c6673, in6673_1, in6673_2);
    wire[3:0] s6674, in6674_1, in6674_2;
    wire c6674;
    assign in6674_1 = {s5842[2],s5840[3],s5871[0],s5872[1]};
    assign in6674_2 = {s5843[2],s5841[3],s5872[0],c5873};
    CLA_4 KS_6674(s6674, c6674, in6674_1, in6674_2);
    wire[3:0] s6675, in6675_1, in6675_2;
    wire c6675;
    assign in6675_1 = {s5844[2],s5842[3],s5873[0],s5874[1]};
    assign in6675_2 = {c5846,s5843[3],s5874[0],c5875};
    CLA_4 KS_6675(s6675, c6675, in6675_1, in6675_2);
    wire[0:0] s6676, in6676_1, in6676_2;
    wire c6676;
    assign in6676_1 = {s5848[2]};
    assign in6676_2 = {c5850};
    Half_Adder KS_6676(s6676, c6676, in6676_1, in6676_2);
    wire[2:0] s6677, in6677_1, in6677_2;
    wire c6677;
    assign in6677_1 = {s5852[2],s5844[3],s5875[0]};
    assign in6677_2 = {c5854,c5848,s5876[0]};
    CLA_3 KS_6677(s6677, c6677, in6677_1, in6677_2);
    wire[0:0] s6678, in6678_1, in6678_2;
    wire c6678;
    assign in6678_1 = {c6659};
    assign in6678_2 = {c6660};
    Half_Adder KS_6678(s6678, c6678, in6678_1, in6678_2);
    wire[1:0] s6679, in6679_1, in6679_2;
    wire c6679;
    assign in6679_1 = {c6661,s5852[3]};
    assign in6679_2 = {c6662,s6670[1]};
    CLA_2 KS_6679(s6679, c6679, in6679_1, in6679_2);
    wire[0:0] s6680, in6680_1, in6680_2;
    wire c6680;
    assign in6680_1 = {c6663};
    assign in6680_2 = {c6664};
    Half_Adder KS_6680(s6680, c6680, in6680_1, in6680_2);
    wire[3:0] s6681, in6681_1, in6681_2;
    wire c6681;
    assign in6681_1 = {s6670[0],s6671[1],s5877[0],s5876[1]};
    assign in6681_2 = {s6671[0],s6672[1],s5878[0],c5877};
    CLA_4_c KS_6681(s6681, c6681, in6681_1, in6681_2, c6666);
    wire[3:0] s6682, in6682_1, in6682_2;
    wire c6682;
    assign in6682_1 = {s5858[2],s4613[0],s5886[0],s5887[1]};
    assign in6682_2 = {s5859[2],s5856[3],s5887[0],s5888[1]};
    CLA_4 KS_6682(s6682, c6682, in6682_1, in6682_2);
    wire[3:0] s6683, in6683_1, in6683_2;
    wire c6683;
    assign in6683_1 = {s5860[2],s5857[3],s5888[0],s5889[1]};
    assign in6683_2 = {s5861[2],s5858[3],s5889[0],c5890};
    CLA_4 KS_6683(s6683, c6683, in6683_1, in6683_2);
    wire[3:0] s6684, in6684_1, in6684_2;
    wire c6684;
    assign in6684_1 = {s5862[2],s5859[3],s5890[0],s5891[1]};
    assign in6684_2 = {s5863[2],s5860[3],s5891[0],c5892};
    CLA_4 KS_6684(s6684, c6684, in6684_1, in6684_2);
    wire[3:0] s6685, in6685_1, in6685_2;
    wire c6685;
    assign in6685_1 = {s5864[2],s5861[3],s5892[0],s5893[1]};
    assign in6685_2 = {s5865[2],s5862[3],s5893[0],c5894};
    CLA_4 KS_6685(s6685, c6685, in6685_1, in6685_2);
    wire[3:0] s6686, in6686_1, in6686_2;
    wire c6686;
    assign in6686_1 = {s5866[2],s5863[3],s5894[0],s5895[1]};
    assign in6686_2 = {c5868,s5864[3],s5895[0],c5896};
    CLA_4 KS_6686(s6686, c6686, in6686_1, in6686_2);
    wire[3:0] s6687, in6687_1, in6687_2;
    wire c6687;
    assign in6687_1 = {s5870[2],s5865[3],s5896[0],s5897[1]};
    assign in6687_2 = {c5872,s5866[3],s5897[0],c5898};
    CLA_4 KS_6687(s6687, c6687, in6687_1, in6687_2);
    wire[0:0] s6688, in6688_1, in6688_2;
    wire c6688;
    assign in6688_1 = {s5874[2]};
    assign in6688_2 = {c5876};
    Half_Adder KS_6688(s6688, c6688, in6688_1, in6688_2);
    wire[2:0] s6689, in6689_1, in6689_2;
    wire c6689;
    assign in6689_1 = {s5878[2],s5870[3],s5898[0]};
    assign in6689_2 = {c6670,c5874,s5899[0]};
    CLA_3 KS_6689(s6689, c6689, in6689_1, in6689_2);
    wire[0:0] s6690, in6690_1, in6690_2;
    wire c6690;
    assign in6690_1 = {c6671};
    assign in6690_2 = {c6672};
    Half_Adder KS_6690(s6690, c6690, in6690_1, in6690_2);
    wire[1:0] s6691, in6691_1, in6691_2;
    wire c6691;
    assign in6691_1 = {c6673,s5878[3]};
    assign in6691_2 = {c6674,s6682[1]};
    CLA_2 KS_6691(s6691, c6691, in6691_1, in6691_2);
    wire[0:0] s6692, in6692_1, in6692_2;
    wire c6692;
    assign in6692_1 = {c6681};
    assign in6692_2 = {s6682[0]};
    Full_Adder KS_6692(s6692, c6692, in6692_1, in6692_2, c6675);
    wire[3:0] s6693, in6693_1, in6693_2;
    wire c6693;
    assign in6693_1 = {s5880[2],s4649[0],s5909[0],s5910[1]};
    assign in6693_2 = {s5881[2],s5879[3],s5910[0],s5911[1]};
    CLA_4 KS_6693(s6693, c6693, in6693_1, in6693_2);
    wire[3:0] s6694, in6694_1, in6694_2;
    wire c6694;
    assign in6694_1 = {s5882[2],s5880[3],s5911[0],s5912[1]};
    assign in6694_2 = {s5883[2],s5881[3],s5912[0],c5913};
    CLA_4 KS_6694(s6694, c6694, in6694_1, in6694_2);
    wire[3:0] s6695, in6695_1, in6695_2;
    wire c6695;
    assign in6695_1 = {s5884[2],s5882[3],s5913[0],s5914[1]};
    assign in6695_2 = {s5885[2],s5883[3],s5914[0],c5915};
    CLA_4 KS_6695(s6695, c6695, in6695_1, in6695_2);
    wire[3:0] s6696, in6696_1, in6696_2;
    wire c6696;
    assign in6696_1 = {s5886[2],s5884[3],s5915[0],s5916[1]};
    assign in6696_2 = {s5887[2],s5885[3],s5916[0],c5917};
    CLA_4 KS_6696(s6696, c6696, in6696_1, in6696_2);
    wire[3:0] s6697, in6697_1, in6697_2;
    wire c6697;
    assign in6697_1 = {s5888[2],s5886[3],s5917[0],s5918[1]};
    assign in6697_2 = {s5889[2],s5887[3],s5918[0],c5919};
    CLA_4 KS_6697(s6697, c6697, in6697_1, in6697_2);
    wire[3:0] s6698, in6698_1, in6698_2;
    wire c6698;
    assign in6698_1 = {s5891[2],s5888[3],s5919[0],s5920[1]};
    assign in6698_2 = {c5893,s5889[3],s5920[0],c5921};
    CLA_4 KS_6698(s6698, c6698, in6698_1, in6698_2);
    wire[0:0] s6699, in6699_1, in6699_2;
    wire c6699;
    assign in6699_1 = {s5895[2]};
    assign in6699_2 = {c5897};
    Half_Adder KS_6699(s6699, c6699, in6699_1, in6699_2);
    wire[2:0] s6700, in6700_1, in6700_2;
    wire c6700;
    assign in6700_1 = {s5899[2],s5891[3],s5921[0]};
    assign in6700_2 = {c5901,c5895,s5922[0]};
    CLA_3 KS_6700(s6700, c6700, in6700_1, in6700_2);
    wire[0:0] s6701, in6701_1, in6701_2;
    wire c6701;
    assign in6701_1 = {c6682};
    assign in6701_2 = {c6683};
    Half_Adder KS_6701(s6701, c6701, in6701_1, in6701_2);
    wire[1:0] s6702, in6702_1, in6702_2;
    wire c6702;
    assign in6702_1 = {c6684,s5899[3]};
    assign in6702_2 = {c6685,s6693[1]};
    CLA_2 KS_6702(s6702, c6702, in6702_1, in6702_2);
    wire[0:0] s6703, in6703_1, in6703_2;
    wire c6703;
    assign in6703_1 = {c6687};
    assign in6703_2 = {s6693[0]};
    Full_Adder KS_6703(s6703, c6703, in6703_1, in6703_2, c6686);
    wire[3:0] s6704, in6704_1, in6704_2;
    wire c6704;
    assign in6704_1 = {s5904[2],s4687[0],s5932[0],s5933[1]};
    assign in6704_2 = {s5905[2],s5902[3],s5933[0],s5934[1]};
    CLA_4 KS_6704(s6704, c6704, in6704_1, in6704_2);
    wire[3:0] s6705, in6705_1, in6705_2;
    wire c6705;
    assign in6705_1 = {s5906[2],s5903[3],s5934[0],s5935[1]};
    assign in6705_2 = {s5907[2],s5904[3],s5935[0],c5936};
    CLA_4 KS_6705(s6705, c6705, in6705_1, in6705_2);
    wire[3:0] s6706, in6706_1, in6706_2;
    wire c6706;
    assign in6706_1 = {s5908[2],s5905[3],s5936[0],s5937[1]};
    assign in6706_2 = {s5909[2],s5906[3],s5937[0],c5938};
    CLA_4 KS_6706(s6706, c6706, in6706_1, in6706_2);
    wire[3:0] s6707, in6707_1, in6707_2;
    wire c6707;
    assign in6707_1 = {s5910[2],s5907[3],s5938[0],s5939[1]};
    assign in6707_2 = {s5911[2],s5908[3],s5939[0],c5940};
    CLA_4 KS_6707(s6707, c6707, in6707_1, in6707_2);
    wire[3:0] s6708, in6708_1, in6708_2;
    wire c6708;
    assign in6708_1 = {s5912[2],s5909[3],s5940[0],s5941[1]};
    assign in6708_2 = {c5914,s5910[3],s5941[0],c5942};
    CLA_4 KS_6708(s6708, c6708, in6708_1, in6708_2);
    wire[3:0] s6709, in6709_1, in6709_2;
    wire c6709;
    assign in6709_1 = {s5916[2],s5911[3],s5942[0],s5943[1]};
    assign in6709_2 = {c5918,s5912[3],s5943[0],c5944};
    CLA_4 KS_6709(s6709, c6709, in6709_1, in6709_2);
    wire[0:0] s6710, in6710_1, in6710_2;
    wire c6710;
    assign in6710_1 = {s5920[2]};
    assign in6710_2 = {c5922};
    Half_Adder KS_6710(s6710, c6710, in6710_1, in6710_2);
    wire[2:0] s6711, in6711_1, in6711_2;
    wire c6711;
    assign in6711_1 = {s5924[2],s5916[3],s5944[0]};
    assign in6711_2 = {c6693,c5920,s5945[0]};
    CLA_3 KS_6711(s6711, c6711, in6711_1, in6711_2);
    wire[0:0] s6712, in6712_1, in6712_2;
    wire c6712;
    assign in6712_1 = {c6694};
    assign in6712_2 = {c6695};
    Half_Adder KS_6712(s6712, c6712, in6712_1, in6712_2);
    wire[1:0] s6713, in6713_1, in6713_2;
    wire c6713;
    assign in6713_1 = {c6697,s5924[3]};
    assign in6713_2 = {c6698,s6704[1]};
    CLA_2_c KS_6713(s6713, c6713, in6713_1, in6713_2, c6696);
    wire[3:0] s6714, in6714_1, in6714_2;
    wire c6714;
    assign in6714_1 = {s5926[2],s4723[0],s5955[0],s5955[1]};
    assign in6714_2 = {s5927[2],s5925[3],s5956[0],s5956[1]};
    CLA_4 KS_6714(s6714, c6714, in6714_1, in6714_2);
    wire[3:0] s6715, in6715_1, in6715_2;
    wire c6715;
    assign in6715_1 = {s5928[2],s5926[3],s5957[0],s5957[1]};
    assign in6715_2 = {s5929[2],s5927[3],s5958[0],s5958[1]};
    CLA_4 KS_6715(s6715, c6715, in6715_1, in6715_2);
    wire[3:0] s6716, in6716_1, in6716_2;
    wire c6716;
    assign in6716_1 = {s5930[2],s5928[3],s5959[0],s5959[1]};
    assign in6716_2 = {s5931[2],s5929[3],s5960[0],c5960};
    CLA_4 KS_6716(s6716, c6716, in6716_1, in6716_2);
    wire[3:0] s6717, in6717_1, in6717_2;
    wire c6717;
    assign in6717_1 = {s5932[2],s5930[3],s5961[0],s5961[1]};
    assign in6717_2 = {s5933[2],s5931[3],s5962[0],c5962};
    CLA_4 KS_6717(s6717, c6717, in6717_1, in6717_2);
    wire[3:0] s6718, in6718_1, in6718_2;
    wire c6718;
    assign in6718_1 = {s5934[2],s5932[3],s5963[0],s5963[1]};
    assign in6718_2 = {s5935[2],s5933[3],s5964[0],c5964};
    CLA_4 KS_6718(s6718, c6718, in6718_1, in6718_2);
    wire[3:0] s6719, in6719_1, in6719_2;
    wire c6719;
    assign in6719_1 = {s5937[2],s5934[3],s5965[0],s5965[1]};
    assign in6719_2 = {c5939,s5935[3],s5966[0],c5966};
    CLA_4 KS_6719(s6719, c6719, in6719_1, in6719_2);
    wire[0:0] s6720, in6720_1, in6720_2;
    wire c6720;
    assign in6720_1 = {s5941[2]};
    assign in6720_2 = {c5943};
    Half_Adder KS_6720(s6720, c6720, in6720_1, in6720_2);
    wire[3:0] s6721, in6721_1, in6721_2;
    wire c6721;
    assign in6721_1 = {s5945[2],s5937[3],s5967[0],s5967[1]};
    assign in6721_2 = {c5947,c5941,s5968[0],c5968};
    CLA_4 KS_6721(s6721, c6721, in6721_1, in6721_2);
    wire[0:0] s6722, in6722_1, in6722_2;
    wire c6722;
    assign in6722_1 = {c6704};
    assign in6722_2 = {c6705};
    Half_Adder KS_6722(s6722, c6722, in6722_1, in6722_2);
    wire[1:0] s6723, in6723_1, in6723_2;
    wire c6723;
    assign in6723_1 = {c6706,s5945[3]};
    assign in6723_2 = {c6707,s6714[1]};
    CLA_2 KS_6723(s6723, c6723, in6723_1, in6723_2);
    wire[0:0] s6724, in6724_1, in6724_2;
    wire c6724;
    assign in6724_1 = {c6709};
    assign in6724_2 = {s6714[0]};
    Full_Adder KS_6724(s6724, c6724, in6724_1, in6724_2, c6708);
    wire[3:0] s6725, in6725_1, in6725_2;
    wire c6725;
    assign in6725_1 = {s5949[2],s4759[0],s5978[0],s5978[1]};
    assign in6725_2 = {s5950[2],s5948[3],s5979[0],s5979[1]};
    CLA_4 KS_6725(s6725, c6725, in6725_1, in6725_2);
    wire[3:0] s6726, in6726_1, in6726_2;
    wire c6726;
    assign in6726_1 = {s5951[2],s5949[3],s5980[0],s5980[1]};
    assign in6726_2 = {s5952[2],s5950[3],s5981[0],s5981[1]};
    CLA_4 KS_6726(s6726, c6726, in6726_1, in6726_2);
    wire[3:0] s6727, in6727_1, in6727_2;
    wire c6727;
    assign in6727_1 = {s5953[2],s5951[3],s5982[0],s5982[1]};
    assign in6727_2 = {s5954[2],s5952[3],s5983[0],c5983};
    CLA_4 KS_6727(s6727, c6727, in6727_1, in6727_2);
    wire[3:0] s6728, in6728_1, in6728_2;
    wire c6728;
    assign in6728_1 = {s5955[2],s5953[3],s5984[0],s5984[1]};
    assign in6728_2 = {s5956[2],s5954[3],s5985[0],c5985};
    CLA_4 KS_6728(s6728, c6728, in6728_1, in6728_2);
    wire[3:0] s6729, in6729_1, in6729_2;
    wire c6729;
    assign in6729_1 = {s5957[2],s5955[3],s5986[0],s5986[1]};
    assign in6729_2 = {s5958[2],s5956[3],s5987[0],c5987};
    CLA_4 KS_6729(s6729, c6729, in6729_1, in6729_2);
    wire[3:0] s6730, in6730_1, in6730_2;
    wire c6730;
    assign in6730_1 = {s5959[2],s5957[3],s5988[0],s5988[1]};
    assign in6730_2 = {c5961,s5958[3],s5989[0],c5989};
    CLA_4 KS_6730(s6730, c6730, in6730_1, in6730_2);
    wire[0:0] s6731, in6731_1, in6731_2;
    wire c6731;
    assign in6731_1 = {s5963[2]};
    assign in6731_2 = {c5965};
    Half_Adder KS_6731(s6731, c6731, in6731_1, in6731_2);
    wire[3:0] s6732, in6732_1, in6732_2;
    wire c6732;
    assign in6732_1 = {s5967[2],s5959[3],s5990[0],s5990[1]};
    assign in6732_2 = {c5969,c5963,s5991[0],c5991};
    CLA_4 KS_6732(s6732, c6732, in6732_1, in6732_2);
    wire[0:0] s6733, in6733_1, in6733_2;
    wire c6733;
    assign in6733_1 = {c6714};
    assign in6733_2 = {c6715};
    Half_Adder KS_6733(s6733, c6733, in6733_1, in6733_2);
    wire[1:0] s6734, in6734_1, in6734_2;
    wire c6734;
    assign in6734_1 = {c6716,s5967[3]};
    assign in6734_2 = {c6717,s6725[1]};
    CLA_2 KS_6734(s6734, c6734, in6734_1, in6734_2);
    wire[0:0] s6735, in6735_1, in6735_2;
    wire c6735;
    assign in6735_1 = {c6718};
    assign in6735_2 = {c6719};
    Half_Adder KS_6735(s6735, c6735, in6735_1, in6735_2);
    wire[2:0] s6736, in6736_1, in6736_2;
    wire c6736;
    assign in6736_1 = {s6725[0],s6726[1],s5992[0]};
    assign in6736_2 = {s6726[0],s6727[1],s5993[0]};
    CLA_3_c KS_6736(s6736, c6736, in6736_1, in6736_2, c6721);
    wire[3:0] s6737, in6737_1, in6737_2;
    wire c6737;
    assign in6737_1 = {s5972[2],s4796[0],s6000[0],s6001[1]};
    assign in6737_2 = {s5973[2],s5971[3],s6001[0],s6002[1]};
    CLA_4 KS_6737(s6737, c6737, in6737_1, in6737_2);
    wire[3:0] s6738, in6738_1, in6738_2;
    wire c6738;
    assign in6738_1 = {s5974[2],s5972[3],s6002[0],s6003[1]};
    assign in6738_2 = {s5975[2],s5973[3],s6003[0],s6004[1]};
    CLA_4 KS_6738(s6738, c6738, in6738_1, in6738_2);
    wire[3:0] s6739, in6739_1, in6739_2;
    wire c6739;
    assign in6739_1 = {s5976[2],s5974[3],s6004[0],s6005[1]};
    assign in6739_2 = {s5977[2],s5975[3],s6005[0],c6006};
    CLA_4 KS_6739(s6739, c6739, in6739_1, in6739_2);
    wire[3:0] s6740, in6740_1, in6740_2;
    wire c6740;
    assign in6740_1 = {s5978[2],s5976[3],s6006[0],s6007[1]};
    assign in6740_2 = {s5979[2],s5977[3],s6007[0],c6008};
    CLA_4 KS_6740(s6740, c6740, in6740_1, in6740_2);
    wire[3:0] s6741, in6741_1, in6741_2;
    wire c6741;
    assign in6741_1 = {s5980[2],s5978[3],s6008[0],s6009[1]};
    assign in6741_2 = {s5981[2],s5979[3],s6009[0],c6010};
    CLA_4 KS_6741(s6741, c6741, in6741_1, in6741_2);
    wire[3:0] s6742, in6742_1, in6742_2;
    wire c6742;
    assign in6742_1 = {s5982[2],s5980[3],s6010[0],s6011[1]};
    assign in6742_2 = {c5984,s5981[3],s6011[0],c6012};
    CLA_4 KS_6742(s6742, c6742, in6742_1, in6742_2);
    wire[0:0] s6743, in6743_1, in6743_2;
    wire c6743;
    assign in6743_1 = {s5986[2]};
    assign in6743_2 = {c5988};
    Half_Adder KS_6743(s6743, c6743, in6743_1, in6743_2);
    wire[2:0] s6744, in6744_1, in6744_2;
    wire c6744;
    assign in6744_1 = {s5990[2],s5982[3],s6012[0]};
    assign in6744_2 = {c5992,c5986,s6013[0]};
    CLA_3 KS_6744(s6744, c6744, in6744_1, in6744_2);
    wire[0:0] s6745, in6745_1, in6745_2;
    wire c6745;
    assign in6745_1 = {c6725};
    assign in6745_2 = {c6726};
    Half_Adder KS_6745(s6745, c6745, in6745_1, in6745_2);
    wire[1:0] s6746, in6746_1, in6746_2;
    wire c6746;
    assign in6746_1 = {c6727,s5990[3]};
    assign in6746_2 = {c6728,s6737[1]};
    CLA_2 KS_6746(s6746, c6746, in6746_1, in6746_2);
    wire[0:0] s6747, in6747_1, in6747_2;
    wire c6747;
    assign in6747_1 = {c6729};
    assign in6747_2 = {c6730};
    Half_Adder KS_6747(s6747, c6747, in6747_1, in6747_2);
    wire[3:0] s6748, in6748_1, in6748_2;
    wire c6748;
    assign in6748_1 = {s6737[0],s6738[1],s6014[0],s6013[1]};
    assign in6748_2 = {s6738[0],s6739[1],s6015[0],c6014};
    CLA_4_c KS_6748(s6748, c6748, in6748_1, in6748_2, c6732);
    wire[3:0] s6749, in6749_1, in6749_2;
    wire c6749;
    assign in6749_1 = {s5995[2],s4832[0],s6023[0],s6024[1]};
    assign in6749_2 = {s5996[2],s5994[3],s6024[0],s6025[1]};
    CLA_4 KS_6749(s6749, c6749, in6749_1, in6749_2);
    wire[3:0] s6750, in6750_1, in6750_2;
    wire c6750;
    assign in6750_1 = {s5997[2],s5995[3],s6025[0],s6026[1]};
    assign in6750_2 = {s5998[2],s5996[3],s6026[0],c6027};
    CLA_4 KS_6750(s6750, c6750, in6750_1, in6750_2);
    wire[3:0] s6751, in6751_1, in6751_2;
    wire c6751;
    assign in6751_1 = {s5999[2],s5997[3],s6027[0],s6028[1]};
    assign in6751_2 = {s6000[2],s5998[3],s6028[0],c6029};
    CLA_4 KS_6751(s6751, c6751, in6751_1, in6751_2);
    wire[3:0] s6752, in6752_1, in6752_2;
    wire c6752;
    assign in6752_1 = {s6001[2],s5999[3],s6029[0],s6030[1]};
    assign in6752_2 = {s6002[2],s6000[3],s6030[0],c6031};
    CLA_4 KS_6752(s6752, c6752, in6752_1, in6752_2);
    wire[3:0] s6753, in6753_1, in6753_2;
    wire c6753;
    assign in6753_1 = {s6003[2],s6001[3],s6031[0],s6032[1]};
    assign in6753_2 = {s6004[2],s6002[3],s6032[0],c6033};
    CLA_4 KS_6753(s6753, c6753, in6753_1, in6753_2);
    wire[3:0] s6754, in6754_1, in6754_2;
    wire c6754;
    assign in6754_1 = {s6005[2],s6003[3],s6033[0],s6034[1]};
    assign in6754_2 = {c6007,s6004[3],s6034[0],c6035};
    CLA_4 KS_6754(s6754, c6754, in6754_1, in6754_2);
    wire[0:0] s6755, in6755_1, in6755_2;
    wire c6755;
    assign in6755_1 = {s6009[2]};
    assign in6755_2 = {c6011};
    Half_Adder KS_6755(s6755, c6755, in6755_1, in6755_2);
    wire[2:0] s6756, in6756_1, in6756_2;
    wire c6756;
    assign in6756_1 = {s6013[2],s6005[3],s6035[0]};
    assign in6756_2 = {c6015,c6009,s6036[0]};
    CLA_3 KS_6756(s6756, c6756, in6756_1, in6756_2);
    wire[0:0] s6757, in6757_1, in6757_2;
    wire c6757;
    assign in6757_1 = {c6737};
    assign in6757_2 = {c6738};
    Half_Adder KS_6757(s6757, c6757, in6757_1, in6757_2);
    wire[1:0] s6758, in6758_1, in6758_2;
    wire c6758;
    assign in6758_1 = {c6739,s6013[3]};
    assign in6758_2 = {c6740,s6749[1]};
    CLA_2 KS_6758(s6758, c6758, in6758_1, in6758_2);
    wire[0:0] s6759, in6759_1, in6759_2;
    wire c6759;
    assign in6759_1 = {c6741};
    assign in6759_2 = {c6742};
    Half_Adder KS_6759(s6759, c6759, in6759_1, in6759_2);
    wire[3:0] s6760, in6760_1, in6760_2;
    wire c6760;
    assign in6760_1 = {s6749[0],s6750[1],s6037[0],s6036[1]};
    assign in6760_2 = {s6750[0],s6751[1],s6038[0],c6037};
    CLA_4_c KS_6760(s6760, c6760, in6760_1, in6760_2, c6748);
    wire[3:0] s6761, in6761_1, in6761_2;
    wire c6761;
    assign in6761_1 = {s6017[2],s4869[0],s6045[0],s6045[1]};
    assign in6761_2 = {s6018[2],s6016[3],s6046[0],s6046[1]};
    CLA_4 KS_6761(s6761, c6761, in6761_1, in6761_2);
    wire[3:0] s6762, in6762_1, in6762_2;
    wire c6762;
    assign in6762_1 = {s6019[2],s6017[3],s6047[0],s6047[1]};
    assign in6762_2 = {s6020[2],s6018[3],s6048[0],s6048[1]};
    CLA_4 KS_6762(s6762, c6762, in6762_1, in6762_2);
    wire[3:0] s6763, in6763_1, in6763_2;
    wire c6763;
    assign in6763_1 = {s6021[2],s6019[3],s6049[0],s6049[1]};
    assign in6763_2 = {s6022[2],s6020[3],s6050[0],c6050};
    CLA_4 KS_6763(s6763, c6763, in6763_1, in6763_2);
    wire[3:0] s6764, in6764_1, in6764_2;
    wire c6764;
    assign in6764_1 = {s6023[2],s6021[3],s6051[0],s6051[1]};
    assign in6764_2 = {s6024[2],s6022[3],s6052[0],c6052};
    CLA_4 KS_6764(s6764, c6764, in6764_1, in6764_2);
    wire[3:0] s6765, in6765_1, in6765_2;
    wire c6765;
    assign in6765_1 = {s6025[2],s6023[3],s6053[0],s6053[1]};
    assign in6765_2 = {s6026[2],s6024[3],s6054[0],c6054};
    CLA_4 KS_6765(s6765, c6765, in6765_1, in6765_2);
    wire[3:0] s6766, in6766_1, in6766_2;
    wire c6766;
    assign in6766_1 = {s6028[2],s6025[3],s6055[0],s6055[1]};
    assign in6766_2 = {c6030,s6026[3],s6056[0],c6056};
    CLA_4 KS_6766(s6766, c6766, in6766_1, in6766_2);
    wire[0:0] s6767, in6767_1, in6767_2;
    wire c6767;
    assign in6767_1 = {s6032[2]};
    assign in6767_2 = {c6034};
    Half_Adder KS_6767(s6767, c6767, in6767_1, in6767_2);
    wire[3:0] s6768, in6768_1, in6768_2;
    wire c6768;
    assign in6768_1 = {s6036[2],s6028[3],s6057[0],s6057[1]};
    assign in6768_2 = {c6038,c6032,s6058[0],c6058};
    CLA_4 KS_6768(s6768, c6768, in6768_1, in6768_2);
    wire[0:0] s6769, in6769_1, in6769_2;
    wire c6769;
    assign in6769_1 = {c6749};
    assign in6769_2 = {c6750};
    Half_Adder KS_6769(s6769, c6769, in6769_1, in6769_2);
    wire[1:0] s6770, in6770_1, in6770_2;
    wire c6770;
    assign in6770_1 = {c6751,s6036[3]};
    assign in6770_2 = {c6752,s6761[1]};
    CLA_2 KS_6770(s6770, c6770, in6770_1, in6770_2);
    wire[0:0] s6771, in6771_1, in6771_2;
    wire c6771;
    assign in6771_1 = {c6753};
    assign in6771_2 = {c6754};
    Half_Adder KS_6771(s6771, c6771, in6771_1, in6771_2);
    wire[2:0] s6772, in6772_1, in6772_2;
    wire c6772;
    assign in6772_1 = {s6761[0],s6762[1],s6059[0]};
    assign in6772_2 = {s6762[0],s6763[1],s6060[0]};
    CLA_3_c KS_6772(s6772, c6772, in6772_1, in6772_2, c6760);
    wire[3:0] s6773, in6773_1, in6773_2;
    wire c6773;
    assign in6773_1 = {s6040[2],s4905[0],s6068[0],s6068[1]};
    assign in6773_2 = {s6041[2],s6039[3],s6069[0],s6069[1]};
    CLA_4 KS_6773(s6773, c6773, in6773_1, in6773_2);
    wire[3:0] s6774, in6774_1, in6774_2;
    wire c6774;
    assign in6774_1 = {s6042[2],s6040[3],s6070[0],s6070[1]};
    assign in6774_2 = {s6043[2],s6041[3],s6071[0],s6071[1]};
    CLA_4 KS_6774(s6774, c6774, in6774_1, in6774_2);
    wire[3:0] s6775, in6775_1, in6775_2;
    wire c6775;
    assign in6775_1 = {s6044[2],s6042[3],s6072[0],s6072[1]};
    assign in6775_2 = {s6045[2],s6043[3],s6073[0],c6073};
    CLA_4 KS_6775(s6775, c6775, in6775_1, in6775_2);
    wire[3:0] s6776, in6776_1, in6776_2;
    wire c6776;
    assign in6776_1 = {s6046[2],s6044[3],s6074[0],s6074[1]};
    assign in6776_2 = {s6047[2],s6045[3],s6075[0],c6075};
    CLA_4 KS_6776(s6776, c6776, in6776_1, in6776_2);
    wire[3:0] s6777, in6777_1, in6777_2;
    wire c6777;
    assign in6777_1 = {s6048[2],s6046[3],s6076[0],s6076[1]};
    assign in6777_2 = {s6049[2],s6047[3],s6077[0],c6077};
    CLA_4 KS_6777(s6777, c6777, in6777_1, in6777_2);
    wire[3:0] s6778, in6778_1, in6778_2;
    wire c6778;
    assign in6778_1 = {s6051[2],s6048[3],s6078[0],s6078[1]};
    assign in6778_2 = {c6053,s6049[3],s6079[0],c6079};
    CLA_4 KS_6778(s6778, c6778, in6778_1, in6778_2);
    wire[0:0] s6779, in6779_1, in6779_2;
    wire c6779;
    assign in6779_1 = {s6055[2]};
    assign in6779_2 = {c6057};
    Half_Adder KS_6779(s6779, c6779, in6779_1, in6779_2);
    wire[3:0] s6780, in6780_1, in6780_2;
    wire c6780;
    assign in6780_1 = {s6059[2],s6051[3],s6080[0],s6080[1]};
    assign in6780_2 = {c6761,c6055,s6081[0],c6081};
    CLA_4 KS_6780(s6780, c6780, in6780_1, in6780_2);
    wire[0:0] s6781, in6781_1, in6781_2;
    wire c6781;
    assign in6781_1 = {c6762};
    assign in6781_2 = {c6763};
    Half_Adder KS_6781(s6781, c6781, in6781_1, in6781_2);
    wire[1:0] s6782, in6782_1, in6782_2;
    wire c6782;
    assign in6782_1 = {c6764,s6059[3]};
    assign in6782_2 = {c6765,s6773[1]};
    CLA_2 KS_6782(s6782, c6782, in6782_1, in6782_2);
    wire[0:0] s6783, in6783_1, in6783_2;
    wire c6783;
    assign in6783_1 = {c6768};
    assign in6783_2 = {s6773[0]};
    Full_Adder KS_6783(s6783, c6783, in6783_1, in6783_2, c6766);
    wire[3:0] s6784, in6784_1, in6784_2;
    wire c6784;
    assign in6784_1 = {s6063[2],s4942[0],s6090[0],s6091[1]};
    assign in6784_2 = {s6064[2],s6061[3],s6091[0],s6092[1]};
    CLA_4 KS_6784(s6784, c6784, in6784_1, in6784_2);
    wire[3:0] s6785, in6785_1, in6785_2;
    wire c6785;
    assign in6785_1 = {s6065[2],s6062[3],s6092[0],s6093[1]};
    assign in6785_2 = {s6066[2],s6063[3],s6093[0],s6094[1]};
    CLA_4 KS_6785(s6785, c6785, in6785_1, in6785_2);
    wire[3:0] s6786, in6786_1, in6786_2;
    wire c6786;
    assign in6786_1 = {s6067[2],s6064[3],s6094[0],s6095[1]};
    assign in6786_2 = {s6068[2],s6065[3],s6095[0],c6096};
    CLA_4 KS_6786(s6786, c6786, in6786_1, in6786_2);
    wire[3:0] s6787, in6787_1, in6787_2;
    wire c6787;
    assign in6787_1 = {s6069[2],s6066[3],s6096[0],s6097[1]};
    assign in6787_2 = {s6070[2],s6067[3],s6097[0],c6098};
    CLA_4 KS_6787(s6787, c6787, in6787_1, in6787_2);
    wire[3:0] s6788, in6788_1, in6788_2;
    wire c6788;
    assign in6788_1 = {s6071[2],s6068[3],s6098[0],s6099[1]};
    assign in6788_2 = {c6072,s6069[3],s6099[0],c6100};
    CLA_4 KS_6788(s6788, c6788, in6788_1, in6788_2);
    wire[3:0] s6789, in6789_1, in6789_2;
    wire c6789;
    assign in6789_1 = {s6074[2],s6070[3],s6100[0],s6101[1]};
    assign in6789_2 = {c6076,s6071[3],s6101[0],c6102};
    CLA_4 KS_6789(s6789, c6789, in6789_1, in6789_2);
    wire[0:0] s6790, in6790_1, in6790_2;
    wire c6790;
    assign in6790_1 = {s6078[2]};
    assign in6790_2 = {c6080};
    Half_Adder KS_6790(s6790, c6790, in6790_1, in6790_2);
    wire[2:0] s6791, in6791_1, in6791_2;
    wire c6791;
    assign in6791_1 = {s6082[2],s6074[3],s6102[0]};
    assign in6791_2 = {c6773,c6078,s6103[0]};
    CLA_3 KS_6791(s6791, c6791, in6791_1, in6791_2);
    wire[0:0] s6792, in6792_1, in6792_2;
    wire c6792;
    assign in6792_1 = {c6774};
    assign in6792_2 = {c6775};
    Half_Adder KS_6792(s6792, c6792, in6792_1, in6792_2);
    wire[1:0] s6793, in6793_1, in6793_2;
    wire c6793;
    assign in6793_1 = {c6776,s6082[3]};
    assign in6793_2 = {c6777,s6784[1]};
    CLA_2 KS_6793(s6793, c6793, in6793_1, in6793_2);
    wire[0:0] s6794, in6794_1, in6794_2;
    wire c6794;
    assign in6794_1 = {c6780};
    assign in6794_2 = {s6784[0]};
    Full_Adder KS_6794(s6794, c6794, in6794_1, in6794_2, c6778);
    wire[3:0] s6795, in6795_1, in6795_2;
    wire c6795;
    assign in6795_1 = {s6086[2],s4980[0],s6113[0],s6114[1]};
    assign in6795_2 = {s6087[2],s6084[3],s6114[0],s6115[1]};
    CLA_4 KS_6795(s6795, c6795, in6795_1, in6795_2);
    wire[3:0] s6796, in6796_1, in6796_2;
    wire c6796;
    assign in6796_1 = {s6088[2],s6085[3],s6115[0],s6116[1]};
    assign in6796_2 = {s6089[2],s6086[3],s6116[0],c6117};
    CLA_4 KS_6796(s6796, c6796, in6796_1, in6796_2);
    wire[3:0] s6797, in6797_1, in6797_2;
    wire c6797;
    assign in6797_1 = {s6090[2],s6087[3],s6117[0],s6118[1]};
    assign in6797_2 = {s6091[2],s6088[3],s6118[0],c6119};
    CLA_4 KS_6797(s6797, c6797, in6797_1, in6797_2);
    wire[3:0] s6798, in6798_1, in6798_2;
    wire c6798;
    assign in6798_1 = {s6092[2],s6089[3],s6119[0],s6120[1]};
    assign in6798_2 = {s6093[2],s6090[3],s6120[0],c6121};
    CLA_4 KS_6798(s6798, c6798, in6798_1, in6798_2);
    wire[3:0] s6799, in6799_1, in6799_2;
    wire c6799;
    assign in6799_1 = {s6094[2],s6091[3],s6121[0],s6122[1]};
    assign in6799_2 = {c6095,s6092[3],s6122[0],c6123};
    CLA_4 KS_6799(s6799, c6799, in6799_1, in6799_2);
    wire[3:0] s6800, in6800_1, in6800_2;
    wire c6800;
    assign in6800_1 = {s6097[2],s6093[3],s6123[0],s6124[1]};
    assign in6800_2 = {c6099,s6094[3],s6124[0],c6125};
    CLA_4 KS_6800(s6800, c6800, in6800_1, in6800_2);
    wire[0:0] s6801, in6801_1, in6801_2;
    wire c6801;
    assign in6801_1 = {s6101[2]};
    assign in6801_2 = {c6103};
    Half_Adder KS_6801(s6801, c6801, in6801_1, in6801_2);
    wire[2:0] s6802, in6802_1, in6802_2;
    wire c6802;
    assign in6802_1 = {s6105[2],s6097[3],s6125[0]};
    assign in6802_2 = {c6784,c6101,s6126[0]};
    CLA_3 KS_6802(s6802, c6802, in6802_1, in6802_2);
    wire[0:0] s6803, in6803_1, in6803_2;
    wire c6803;
    assign in6803_1 = {c6785};
    assign in6803_2 = {c6786};
    Half_Adder KS_6803(s6803, c6803, in6803_1, in6803_2);
    wire[1:0] s6804, in6804_1, in6804_2;
    wire c6804;
    assign in6804_1 = {c6788,s6105[3]};
    assign in6804_2 = {c6789,s6795[1]};
    CLA_2_c KS_6804(s6804, c6804, in6804_1, in6804_2, c6787);
    wire[3:0] s6805, in6805_1, in6805_2;
    wire c6805;
    assign in6805_1 = {s6108[2],s5017[0],s6136[0],s6136[1]};
    assign in6805_2 = {s6109[2],s6106[3],s6137[0],s6137[1]};
    CLA_4 KS_6805(s6805, c6805, in6805_1, in6805_2);
    wire[3:0] s6806, in6806_1, in6806_2;
    wire c6806;
    assign in6806_1 = {s6110[2],s6107[3],s6138[0],s6138[1]};
    assign in6806_2 = {s6111[2],s6108[3],s6139[0],s6139[1]};
    CLA_4 KS_6806(s6806, c6806, in6806_1, in6806_2);
    wire[3:0] s6807, in6807_1, in6807_2;
    wire c6807;
    assign in6807_1 = {s6112[2],s6109[3],s6140[0],s6140[1]};
    assign in6807_2 = {s6113[2],s6110[3],s6141[0],c6141};
    CLA_4 KS_6807(s6807, c6807, in6807_1, in6807_2);
    wire[3:0] s6808, in6808_1, in6808_2;
    wire c6808;
    assign in6808_1 = {s6114[2],s6111[3],s6142[0],s6142[1]};
    assign in6808_2 = {s6115[2],s6112[3],s6143[0],c6143};
    CLA_4 KS_6808(s6808, c6808, in6808_1, in6808_2);
    wire[3:0] s6809, in6809_1, in6809_2;
    wire c6809;
    assign in6809_1 = {s6116[2],s6113[3],s6144[0],s6144[1]};
    assign in6809_2 = {c6118,s6114[3],s6145[0],c6145};
    CLA_4 KS_6809(s6809, c6809, in6809_1, in6809_2);
    wire[3:0] s6810, in6810_1, in6810_2;
    wire c6810;
    assign in6810_1 = {s6120[2],s6115[3],s6146[0],s6146[1]};
    assign in6810_2 = {c6122,s6116[3],s6147[0],c6147};
    CLA_4 KS_6810(s6810, c6810, in6810_1, in6810_2);
    wire[0:0] s6811, in6811_1, in6811_2;
    wire c6811;
    assign in6811_1 = {s6124[2]};
    assign in6811_2 = {c6126};
    Half_Adder KS_6811(s6811, c6811, in6811_1, in6811_2);
    wire[3:0] s6812, in6812_1, in6812_2;
    wire c6812;
    assign in6812_1 = {s6128[2],s6120[3],s6148[0],s6148[1]};
    assign in6812_2 = {c6795,c6124,s6149[0],c6149};
    CLA_4 KS_6812(s6812, c6812, in6812_1, in6812_2);
    wire[0:0] s6813, in6813_1, in6813_2;
    wire c6813;
    assign in6813_1 = {c6796};
    assign in6813_2 = {c6797};
    Half_Adder KS_6813(s6813, c6813, in6813_1, in6813_2);
    wire[1:0] s6814, in6814_1, in6814_2;
    wire c6814;
    assign in6814_1 = {c6799,s6128[3]};
    assign in6814_2 = {c6800,s6805[1]};
    CLA_2_c KS_6814(s6814, c6814, in6814_1, in6814_2, c6798);
    wire[3:0] s6815, in6815_1, in6815_2;
    wire c6815;
    assign in6815_1 = {s6131[2],s5047[0],s6159[0],s6159[1]};
    assign in6815_2 = {s6132[2],s6129[3],s6160[0],s6160[1]};
    CLA_4 KS_6815(s6815, c6815, in6815_1, in6815_2);
    wire[3:0] s6816, in6816_1, in6816_2;
    wire c6816;
    assign in6816_1 = {s6133[2],s6130[3],s6161[0],s6161[1]};
    assign in6816_2 = {s6134[2],s6131[3],s6162[0],s6162[1]};
    CLA_4 KS_6816(s6816, c6816, in6816_1, in6816_2);
    wire[3:0] s6817, in6817_1, in6817_2;
    wire c6817;
    assign in6817_1 = {s6135[2],s6132[3],s6163[0],s6163[1]};
    assign in6817_2 = {s6136[2],s6133[3],s6164[0],c6164};
    CLA_4 KS_6817(s6817, c6817, in6817_1, in6817_2);
    wire[3:0] s6818, in6818_1, in6818_2;
    wire c6818;
    assign in6818_1 = {s6137[2],s6134[3],s6165[0],s6165[1]};
    assign in6818_2 = {s6138[2],s6135[3],s6166[0],c6166};
    CLA_4 KS_6818(s6818, c6818, in6818_1, in6818_2);
    wire[3:0] s6819, in6819_1, in6819_2;
    wire c6819;
    assign in6819_1 = {s6139[2],s6136[3],s6167[0],s6167[1]};
    assign in6819_2 = {c6140,s6137[3],s6168[0],c6168};
    CLA_4 KS_6819(s6819, c6819, in6819_1, in6819_2);
    wire[3:0] s6820, in6820_1, in6820_2;
    wire c6820;
    assign in6820_1 = {s6142[2],s6138[3],s6169[0],s6169[1]};
    assign in6820_2 = {c6144,s6139[3],s6170[0],c6170};
    CLA_4 KS_6820(s6820, c6820, in6820_1, in6820_2);
    wire[0:0] s6821, in6821_1, in6821_2;
    wire c6821;
    assign in6821_1 = {s6146[2]};
    assign in6821_2 = {c6148};
    Half_Adder KS_6821(s6821, c6821, in6821_1, in6821_2);
    wire[3:0] s6822, in6822_1, in6822_2;
    wire c6822;
    assign in6822_1 = {s6150[2],s6142[3],s6171[0],s6171[1]};
    assign in6822_2 = {c6805,c6146,s6172[0],c6172};
    CLA_4 KS_6822(s6822, c6822, in6822_1, in6822_2);
    wire[0:0] s6823, in6823_1, in6823_2;
    wire c6823;
    assign in6823_1 = {c6806};
    assign in6823_2 = {c6807};
    Half_Adder KS_6823(s6823, c6823, in6823_1, in6823_2);
    wire[1:0] s6824, in6824_1, in6824_2;
    wire c6824;
    assign in6824_1 = {c6808,s6150[3]};
    assign in6824_2 = {c6809,s6815[1]};
    CLA_2 KS_6824(s6824, c6824, in6824_1, in6824_2);
    wire[0:0] s6825, in6825_1, in6825_2;
    wire c6825;
    assign in6825_1 = {c6812};
    assign in6825_2 = {s6815[0]};
    Full_Adder KS_6825(s6825, c6825, in6825_1, in6825_2, c6810);
    wire[3:0] s6826, in6826_1, in6826_2;
    wire c6826;
    assign in6826_1 = {s6153[2],s5068[0],s6181[0],s6182[1]};
    assign in6826_2 = {s6154[2],s6152[3],s6182[0],s6183[1]};
    CLA_4 KS_6826(s6826, c6826, in6826_1, in6826_2);
    wire[3:0] s6827, in6827_1, in6827_2;
    wire c6827;
    assign in6827_1 = {s6155[2],s6153[3],s6183[0],s6184[1]};
    assign in6827_2 = {s6156[2],s6154[3],s6184[0],s6185[1]};
    CLA_4 KS_6827(s6827, c6827, in6827_1, in6827_2);
    wire[3:0] s6828, in6828_1, in6828_2;
    wire c6828;
    assign in6828_1 = {s6157[2],s6155[3],s6185[0],s6186[1]};
    assign in6828_2 = {s6158[2],s6156[3],s6186[0],c6187};
    CLA_4 KS_6828(s6828, c6828, in6828_1, in6828_2);
    wire[3:0] s6829, in6829_1, in6829_2;
    wire c6829;
    assign in6829_1 = {s6159[2],s6157[3],s6187[0],s6188[1]};
    assign in6829_2 = {s6160[2],s6158[3],s6188[0],c6189};
    CLA_4 KS_6829(s6829, c6829, in6829_1, in6829_2);
    wire[3:0] s6830, in6830_1, in6830_2;
    wire c6830;
    assign in6830_1 = {s6161[2],s6159[3],s6189[0],s6190[1]};
    assign in6830_2 = {s6162[2],s6160[3],s6190[0],c6191};
    CLA_4 KS_6830(s6830, c6830, in6830_1, in6830_2);
    wire[3:0] s6831, in6831_1, in6831_2;
    wire c6831;
    assign in6831_1 = {s6163[2],s6161[3],s6191[0],s6192[1]};
    assign in6831_2 = {c6165,s6162[3],s6192[0],c6193};
    CLA_4 KS_6831(s6831, c6831, in6831_1, in6831_2);
    wire[0:0] s6832, in6832_1, in6832_2;
    wire c6832;
    assign in6832_1 = {s6167[2]};
    assign in6832_2 = {c6169};
    Half_Adder KS_6832(s6832, c6832, in6832_1, in6832_2);
    wire[2:0] s6833, in6833_1, in6833_2;
    wire c6833;
    assign in6833_1 = {s6171[2],s6163[3],s6193[0]};
    assign in6833_2 = {c6173,c6167,s6194[0]};
    CLA_3 KS_6833(s6833, c6833, in6833_1, in6833_2);
    wire[0:0] s6834, in6834_1, in6834_2;
    wire c6834;
    assign in6834_1 = {c6815};
    assign in6834_2 = {c6816};
    Half_Adder KS_6834(s6834, c6834, in6834_1, in6834_2);
    wire[1:0] s6835, in6835_1, in6835_2;
    wire c6835;
    assign in6835_1 = {c6817,s6171[3]};
    assign in6835_2 = {c6818,s6826[1]};
    CLA_2 KS_6835(s6835, c6835, in6835_1, in6835_2);
    wire[0:0] s6836, in6836_1, in6836_2;
    wire c6836;
    assign in6836_1 = {c6819};
    assign in6836_2 = {c6820};
    Half_Adder KS_6836(s6836, c6836, in6836_1, in6836_2);
    wire[3:0] s6837, in6837_1, in6837_2;
    wire c6837;
    assign in6837_1 = {s6826[0],s6827[1],s6195[0],s6194[1]};
    assign in6837_2 = {s6827[0],s6828[1],s6196[0],c6195};
    CLA_4_c KS_6837(s6837, c6837, in6837_1, in6837_2, c6822);
    wire[3:0] s6838, in6838_1, in6838_2;
    wire c6838;
    assign in6838_1 = {s6177[2],s5081[0],s6203[0],s6204[1]};
    assign in6838_2 = {s6178[2],s6175[3],s6204[0],s6205[1]};
    CLA_4 KS_6838(s6838, c6838, in6838_1, in6838_2);
    wire[3:0] s6839, in6839_1, in6839_2;
    wire c6839;
    assign in6839_1 = {s6179[2],s6176[3],s6205[0],s6206[1]};
    assign in6839_2 = {s6180[2],s6177[3],s6206[0],s6207[1]};
    CLA_4 KS_6839(s6839, c6839, in6839_1, in6839_2);
    wire[3:0] s6840, in6840_1, in6840_2;
    wire c6840;
    assign in6840_1 = {s6181[2],s6178[3],s6207[0],s6208[1]};
    assign in6840_2 = {s6182[2],s6179[3],s6208[0],c6209};
    CLA_4 KS_6840(s6840, c6840, in6840_1, in6840_2);
    wire[3:0] s6841, in6841_1, in6841_2;
    wire c6841;
    assign in6841_1 = {s6183[2],s6180[3],s6209[0],s6210[1]};
    assign in6841_2 = {s6184[2],s6181[3],s6210[0],c6211};
    CLA_4 KS_6841(s6841, c6841, in6841_1, in6841_2);
    wire[3:0] s6842, in6842_1, in6842_2;
    wire c6842;
    assign in6842_1 = {s6185[2],s6182[3],s6211[0],s6212[1]};
    assign in6842_2 = {c6186,s6183[3],s6212[0],c6213};
    CLA_4 KS_6842(s6842, c6842, in6842_1, in6842_2);
    wire[3:0] s6843, in6843_1, in6843_2;
    wire c6843;
    assign in6843_1 = {s6188[2],s6184[3],s6213[0],s6214[1]};
    assign in6843_2 = {c6190,s6185[3],s6214[0],c6215};
    CLA_4 KS_6843(s6843, c6843, in6843_1, in6843_2);
    wire[0:0] s6844, in6844_1, in6844_2;
    wire c6844;
    assign in6844_1 = {s6192[2]};
    assign in6844_2 = {c6194};
    Half_Adder KS_6844(s6844, c6844, in6844_1, in6844_2);
    wire[2:0] s6845, in6845_1, in6845_2;
    wire c6845;
    assign in6845_1 = {s6196[2],s6188[3],s6215[0]};
    assign in6845_2 = {c6826,c6192,s6216[0]};
    CLA_3 KS_6845(s6845, c6845, in6845_1, in6845_2);
    wire[0:0] s6846, in6846_1, in6846_2;
    wire c6846;
    assign in6846_1 = {c6827};
    assign in6846_2 = {c6828};
    Half_Adder KS_6846(s6846, c6846, in6846_1, in6846_2);
    wire[1:0] s6847, in6847_1, in6847_2;
    wire c6847;
    assign in6847_1 = {c6829,s6196[3]};
    assign in6847_2 = {c6830,s6838[1]};
    CLA_2 KS_6847(s6847, c6847, in6847_1, in6847_2);
    wire[0:0] s6848, in6848_1, in6848_2;
    wire c6848;
    assign in6848_1 = {c6837};
    assign in6848_2 = {s6838[0]};
    Full_Adder KS_6848(s6848, c6848, in6848_1, in6848_2, c6831);
    wire[3:0] s6849, in6849_1, in6849_2;
    wire c6849;
    assign in6849_1 = {s6198[2],s5085[0],s6226[0],s6227[1]};
    assign in6849_2 = {s6199[2],s6197[3],s6227[0],s6228[1]};
    CLA_4 KS_6849(s6849, c6849, in6849_1, in6849_2);
    wire[3:0] s6850, in6850_1, in6850_2;
    wire c6850;
    assign in6850_1 = {s6200[2],s6198[3],s6228[0],s6229[1]};
    assign in6850_2 = {s6201[2],s6199[3],s6229[0],c6230};
    CLA_4 KS_6850(s6850, c6850, in6850_1, in6850_2);
    wire[3:0] s6851, in6851_1, in6851_2;
    wire c6851;
    assign in6851_1 = {s6202[2],s6200[3],s6230[0],s6231[1]};
    assign in6851_2 = {s6203[2],s6201[3],s6231[0],c6232};
    CLA_4 KS_6851(s6851, c6851, in6851_1, in6851_2);
    wire[3:0] s6852, in6852_1, in6852_2;
    wire c6852;
    assign in6852_1 = {s6204[2],s6202[3],s6232[0],s6233[1]};
    assign in6852_2 = {s6205[2],s6203[3],s6233[0],c6234};
    CLA_4 KS_6852(s6852, c6852, in6852_1, in6852_2);
    wire[3:0] s6853, in6853_1, in6853_2;
    wire c6853;
    assign in6853_1 = {s6206[2],s6204[3],s6234[0],s6235[1]};
    assign in6853_2 = {s6207[2],s6205[3],s6235[0],c6236};
    CLA_4 KS_6853(s6853, c6853, in6853_1, in6853_2);
    wire[3:0] s6854, in6854_1, in6854_2;
    wire c6854;
    assign in6854_1 = {s6208[2],s6206[3],s6236[0],s6237[1]};
    assign in6854_2 = {c6210,s6207[3],s6237[0],c6238};
    CLA_4 KS_6854(s6854, c6854, in6854_1, in6854_2);
    wire[0:0] s6855, in6855_1, in6855_2;
    wire c6855;
    assign in6855_1 = {s6212[2]};
    assign in6855_2 = {c6214};
    Half_Adder KS_6855(s6855, c6855, in6855_1, in6855_2);
    wire[2:0] s6856, in6856_1, in6856_2;
    wire c6856;
    assign in6856_1 = {s6216[2],s6208[3],s6238[0]};
    assign in6856_2 = {c6218,c6212,s6239[0]};
    CLA_3 KS_6856(s6856, c6856, in6856_1, in6856_2);
    wire[0:0] s6857, in6857_1, in6857_2;
    wire c6857;
    assign in6857_1 = {c6838};
    assign in6857_2 = {c6839};
    Half_Adder KS_6857(s6857, c6857, in6857_1, in6857_2);
    wire[1:0] s6858, in6858_1, in6858_2;
    wire c6858;
    assign in6858_1 = {c6840,s6216[3]};
    assign in6858_2 = {c6841,s6849[1]};
    CLA_2 KS_6858(s6858, c6858, in6858_1, in6858_2);
    wire[0:0] s6859, in6859_1, in6859_2;
    wire c6859;
    assign in6859_1 = {c6843};
    assign in6859_2 = {s6849[0]};
    Full_Adder KS_6859(s6859, c6859, in6859_1, in6859_2, c6842);
    wire[3:0] s6860, in6860_1, in6860_2;
    wire c6860;
    assign in6860_1 = {s6221[2],pp126[105],s6243[0],s6244[1]};
    assign in6860_2 = {s6222[2],pp127[104],s6244[0],s6245[1]};
    CLA_4 KS_6860(s6860, c6860, in6860_1, in6860_2);
    wire[3:0] s6861, in6861_1, in6861_2;
    wire c6861;
    assign in6861_1 = {s6223[2],s6219[3],s6245[0],s6246[1]};
    assign in6861_2 = {s6224[2],s6220[3],s6246[0],s6247[1]};
    CLA_4 KS_6861(s6861, c6861, in6861_1, in6861_2);
    wire[3:0] s6862, in6862_1, in6862_2;
    wire c6862;
    assign in6862_1 = {s6225[2],s6221[3],s6247[0],s6248[1]};
    assign in6862_2 = {s6226[2],s6222[3],s6248[0],c6249};
    CLA_4 KS_6862(s6862, c6862, in6862_1, in6862_2);
    wire[3:0] s6863, in6863_1, in6863_2;
    wire c6863;
    assign in6863_1 = {s6227[2],s6223[3],s6249[0],s6250[1]};
    assign in6863_2 = {s6228[2],s6224[3],s6250[0],c6251};
    CLA_4 KS_6863(s6863, c6863, in6863_1, in6863_2);
    wire[3:0] s6864, in6864_1, in6864_2;
    wire c6864;
    assign in6864_1 = {s6229[2],s6225[3],s6251[0],s6252[1]};
    assign in6864_2 = {c6231,s6226[3],s6252[0],c6253};
    CLA_4 KS_6864(s6864, c6864, in6864_1, in6864_2);
    wire[3:0] s6865, in6865_1, in6865_2;
    wire c6865;
    assign in6865_1 = {s6233[2],s6227[3],s6253[0],s6254[1]};
    assign in6865_2 = {c6235,c6228,s6254[0],c6255};
    CLA_4 KS_6865(s6865, c6865, in6865_1, in6865_2);
    wire[2:0] s6866, in6866_1, in6866_2;
    wire c6866;
    assign in6866_1 = {s6237[2],s6229[3],s6255[0]};
    assign in6866_2 = {c6239,c6233,s6256[0]};
    CLA_3 KS_6866(s6866, c6866, in6866_1, in6866_2);
    wire[0:0] s6867, in6867_1, in6867_2;
    wire c6867;
    assign in6867_1 = {s6241[2]};
    assign in6867_2 = {c6849};
    Half_Adder KS_6867(s6867, c6867, in6867_1, in6867_2);
    wire[1:0] s6868, in6868_1, in6868_2;
    wire c6868;
    assign in6868_1 = {c6850,s6237[3]};
    assign in6868_2 = {c6851,c6241};
    CLA_2 KS_6868(s6868, c6868, in6868_1, in6868_2);
    wire[0:0] s6869, in6869_1, in6869_2;
    wire c6869;
    assign in6869_1 = {c6853};
    assign in6869_2 = {c6854};
    Full_Adder KS_6869(s6869, c6869, in6869_1, in6869_2, c6852);
    wire[3:0] s6870, in6870_1, in6870_2;
    wire c6870;
    assign in6870_1 = {pp125[109],pp122[113],c6242,pp122[115]};
    assign in6870_2 = {pp126[108],pp123[112],c6243,pp123[114]};
    CLA_4 KS_6870(s6870, c6870, in6870_1, in6870_2);
    wire[3:0] s6871, in6871_1, in6871_2;
    wire c6871;
    assign in6871_1 = {pp127[107],pp124[111],c6244,pp124[113]};
    assign in6871_2 = {s6242[2],pp125[110],c6245,pp125[112]};
    CLA_4 KS_6871(s6871, c6871, in6871_1, in6871_2);
    wire[3:0] s6872, in6872_1, in6872_2;
    wire c6872;
    assign in6872_1 = {s6243[2],pp126[109],c6246,pp126[111]};
    assign in6872_2 = {s6244[2],pp127[108],c6250,pp127[110]};
    CLA_4 KS_6872(s6872, c6872, in6872_1, in6872_2);
    wire[3:0] s6873, in6873_1, in6873_2;
    wire c6873;
    assign in6873_1 = {s6245[2],s6242[3],c6258,s6259[1]};
    assign in6873_2 = {s6246[2],s6243[3],s6259[0],s6260[1]};
    CLA_4 KS_6873(s6873, c6873, in6873_1, in6873_2);
    wire[3:0] s6874, in6874_1, in6874_2;
    wire c6874;
    assign in6874_1 = {s6247[2],s6244[3],s6260[0],s6261[1]};
    assign in6874_2 = {c6248,s6245[3],s6261[0],c6262};
    CLA_4 KS_6874(s6874, c6874, in6874_1, in6874_2);
    wire[3:0] s6875, in6875_1, in6875_2;
    wire c6875;
    assign in6875_1 = {s6250[2],s6246[3],s6262[0],s6263[1]};
    assign in6875_2 = {c6252,c6247,s6263[0],c6264};
    CLA_4 KS_6875(s6875, c6875, in6875_1, in6875_2);
    wire[0:0] s6876, in6876_1, in6876_2;
    wire c6876;
    assign in6876_1 = {s6254[2]};
    assign in6876_2 = {c6256};
    Half_Adder KS_6876(s6876, c6876, in6876_1, in6876_2);
    wire[2:0] s6877, in6877_1, in6877_2;
    wire c6877;
    assign in6877_1 = {s6258[2],s6250[3],s6264[0]};
    assign in6877_2 = {c6860,c6254,s6265[0]};
    CLA_3 KS_6877(s6877, c6877, in6877_1, in6877_2);
    wire[0:0] s6878, in6878_1, in6878_2;
    wire c6878;
    assign in6878_1 = {c6861};
    assign in6878_2 = {c6862};
    Half_Adder KS_6878(s6878, c6878, in6878_1, in6878_2);
    wire[1:0] s6879, in6879_1, in6879_2;
    wire c6879;
    assign in6879_1 = {c6864,s6258[3]};
    assign in6879_2 = {c6865,s6870[1]};
    CLA_2_c KS_6879(s6879, c6879, in6879_1, in6879_2, c6863);
    wire[3:0] s6880, in6880_1, in6880_2;
    wire c6880;
    assign in6880_1 = {pp119[119],pp116[123],pp115[125],pp114[127]};
    assign in6880_2 = {pp120[118],pp117[122],pp116[124],pp115[126]};
    CLA_4 KS_6880(s6880, c6880, in6880_1, in6880_2);
    wire[3:0] s6881, in6881_1, in6881_2;
    wire c6881;
    assign in6881_1 = {pp121[117],pp118[121],pp117[123],pp116[125]};
    assign in6881_2 = {pp122[116],pp119[120],pp118[122],pp117[124]};
    CLA_4 KS_6881(s6881, c6881, in6881_1, in6881_2);
    wire[3:0] s6882, in6882_1, in6882_2;
    wire c6882;
    assign in6882_1 = {pp123[115],pp120[119],pp119[121],pp118[123]};
    assign in6882_2 = {pp124[114],pp121[118],pp120[120],pp119[122]};
    CLA_4 KS_6882(s6882, c6882, in6882_1, in6882_2);
    wire[3:0] s6883, in6883_1, in6883_2;
    wire c6883;
    assign in6883_1 = {pp125[113],pp122[117],pp121[119],pp120[121]};
    assign in6883_2 = {pp126[112],pp123[116],pp122[118],pp121[120]};
    CLA_4 KS_6883(s6883, c6883, in6883_1, in6883_2);
    wire[3:0] s6884, in6884_1, in6884_2;
    wire c6884;
    assign in6884_1 = {pp127[111],pp124[115],pp123[117],pp122[119]};
    assign in6884_2 = {s6259[2],pp125[114],pp124[116],pp123[118]};
    CLA_4 KS_6884(s6884, c6884, in6884_1, in6884_2);
    wire[3:0] s6885, in6885_1, in6885_2;
    wire c6885;
    assign in6885_1 = {s6260[2],pp126[113],pp125[115],pp124[117]};
    assign in6885_2 = {c6261,pp127[112],pp126[114],pp125[116]};
    CLA_4 KS_6885(s6885, c6885, in6885_1, in6885_2);
    wire[2:0] s6886, in6886_1, in6886_2;
    wire c6886;
    assign in6886_1 = {s6263[2],s6259[3],pp127[113]};
    assign in6886_2 = {c6265,c6260,c6259};
    CLA_3 KS_6886(s6886, c6886, in6886_1, in6886_2);
    wire[0:0] s6887, in6887_1, in6887_2;
    wire c6887;
    assign in6887_1 = {s6267[2]};
    assign in6887_2 = {c6870};
    Half_Adder KS_6887(s6887, c6887, in6887_1, in6887_2);
    wire[1:0] s6888, in6888_1, in6888_2;
    wire c6888;
    assign in6888_1 = {c6871,s6263[3]};
    assign in6888_2 = {c6872,c6267};
    CLA_2 KS_6888(s6888, c6888, in6888_1, in6888_2);
    wire[0:0] s6889, in6889_1, in6889_2;
    wire c6889;
    assign in6889_1 = {c6874};
    assign in6889_2 = {c6875};
    Full_Adder KS_6889(s6889, c6889, in6889_1, in6889_2, c6873);
    wire[3:0] s6890, in6890_1, in6890_2;
    wire c6890;
    assign in6890_1 = {pp115[127],pp116[127],pp117[127],pp118[127]};
    assign in6890_2 = {pp116[126],pp117[126],pp118[126],pp119[126]};
    CLA_4 KS_6890(s6890, c6890, in6890_1, in6890_2);
    wire[2:0] s6891, in6891_1, in6891_2;
    wire c6891;
    assign in6891_1 = {pp117[125],pp118[125],pp119[125]};
    assign in6891_2 = {pp118[124],pp119[124],pp120[124]};
    CLA_3 KS_6891(s6891, c6891, in6891_1, in6891_2);
    wire[1:0] s6892, in6892_1, in6892_2;
    wire c6892;
    assign in6892_1 = {pp119[123],pp120[123]};
    assign in6892_2 = {pp120[122],pp121[122]};
    CLA_2 KS_6892(s6892, c6892, in6892_1, in6892_2);
    wire[0:0] s6893, in6893_1, in6893_2;
    wire c6893;
    assign in6893_1 = {pp121[121]};
    assign in6893_2 = {pp122[120]};
    Half_Adder KS_6893(s6893, c6893, in6893_1, in6893_2);
    wire[3:0] s6894, in6894_1, in6894_2;
    wire c6894;
    assign in6894_1 = {pp123[119],pp122[121],pp121[123],pp120[125]};
    assign in6894_2 = {pp124[118],pp123[120],pp122[122],pp121[124]};
    CLA_4 KS_6894(s6894, c6894, in6894_1, in6894_2);
    wire[0:0] s6895, in6895_1, in6895_2;
    wire c6895;
    assign in6895_1 = {pp125[117]};
    assign in6895_2 = {pp126[116]};
    Half_Adder KS_6895(s6895, c6895, in6895_1, in6895_2);
    wire[1:0] s6896, in6896_1, in6896_2;
    wire c6896;
    assign in6896_1 = {pp127[115],pp124[119]};
    assign in6896_2 = {c6880,pp125[118]};
    CLA_2 KS_6896(s6896, c6896, in6896_1, in6896_2);
    wire[0:0] s6897, in6897_1, in6897_2;
    wire c6897;
    assign in6897_1 = {c6882};
    assign in6897_2 = {c6883};
    Full_Adder KS_6897(s6897, c6897, in6897_1, in6897_2, c6881);
    wire[0:0] s6898, in6898_1, in6898_2;
    wire c6898;
    assign in6898_1 = {pp119[127]};
    assign in6898_2 = {pp120[126]};
    Half_Adder KS_6898(s6898, c6898, in6898_1, in6898_2);

    /*Stage 6*/
    wire[3:0] s6899, in6899_1, in6899_2;
    wire c6899;
    assign in6899_1 = {pp0[6],pp0[7],pp0[8],pp0[9]};
    assign in6899_2 = {pp1[5],pp1[6],pp1[7],pp1[8]};
    CLA_4 KS_6899(s6899, c6899, in6899_1, in6899_2);
    wire[3:0] s6900, in6900_1, in6900_2;
    wire c6900;
    assign in6900_1 = {pp2[5],pp2[6],pp2[7],pp2[8]};
    assign in6900_2 = {pp3[4],pp3[5],pp3[6],pp3[7]};
    CLA_4 KS_6900(s6900, c6900, in6900_1, in6900_2);
    wire[3:0] s6901, in6901_1, in6901_2;
    wire c6901;
    assign in6901_1 = {pp4[4],pp4[5],pp4[6],pp4[7]};
    assign in6901_2 = {pp5[3],pp5[4],pp5[5],pp5[6]};
    CLA_4 KS_6901(s6901, c6901, in6901_1, in6901_2);
    wire[3:0] s6902, in6902_1, in6902_2;
    wire c6902;
    assign in6902_1 = {pp6[3],pp6[4],pp6[5],pp6[6]};
    assign in6902_2 = {pp7[2],pp7[3],pp7[4],pp7[5]};
    CLA_4 KS_6902(s6902, c6902, in6902_1, in6902_2);
    wire[3:0] s6903, in6903_1, in6903_2;
    wire c6903;
    assign in6903_1 = {pp9[1],pp8[3],pp8[4],pp8[5]};
    assign in6903_2 = {pp10[0],pp9[2],pp9[3],pp9[4]};
    CLA_4_c KS_6903(s6903, c6903, in6903_1, in6903_2, pp8[2]);
    wire[3:0] s6904, in6904_1, in6904_2;
    wire c6904;
    assign in6904_1 = {pp11[0],pp10[2],pp10[3],pp11[3]};
    assign in6904_2 = {s6269[1],pp11[1],pp11[2],pp12[2]};
    CLA_4_c KS_6904(s6904, c6904, in6904_1, in6904_2, pp10[1]);
    wire[3:0] s6905, in6905_1, in6905_2;
    wire c6905;
    assign in6905_1 = {s6269[2],pp12[1],pp13[1],pp13[2]};
    assign in6905_2 = {s6270[1],pp13[0],pp14[0],pp14[1]};
    CLA_4_c KS_6905(s6905, c6905, in6905_1, in6905_2, pp12[0]);
    wire[3:0] s6906, in6906_1, in6906_2;
    wire c6906;
    assign in6906_1 = {s6270[2],c6269,pp15[0],pp15[1]};
    assign in6906_2 = {s6271[1],s6270[3],c6270,pp16[0]};
    CLA_4_c KS_6906(s6906, c6906, in6906_1, in6906_2, s6269[3]);
    wire[3:0] s6907, in6907_1, in6907_2;
    wire c6907;
    assign in6907_1 = {s6272[1],s6271[3],s5086[0],pp17[0]};
    assign in6907_2 = {s6273[0],s6272[2],c6271,s5086[1]};
    CLA_4_c KS_6907(s6907, c6907, in6907_1, in6907_2, s6271[2]);
    wire[3:0] s6908, in6908_1, in6908_2;
    wire c6908;
    assign in6908_1 = {s6274[1],s6272[3],s5087[0],s5088[0]};
    assign in6908_2 = {s6275[0],s6273[2],c6272,c6273};
    CLA_4_c KS_6908(s6908, c6908, in6908_1, in6908_2, s6273[1]);
    wire[3:0] s6909, in6909_1, in6909_2;
    wire c6909;
    assign in6909_1 = {s6275[1],s6273[3],c6274,s5089[0]};
    assign in6909_2 = {s6276[1],s6274[3],s6275[3],c6275};
    CLA_4_c KS_6909(s6909, c6909, in6909_1, in6909_2, s6274[2]);
    wire[3:0] s6910, in6910_1, in6910_2;
    wire c6910;
    assign in6910_1 = {s6276[2],s6276[3],c6276,s5090[0]};
    assign in6910_2 = {s6277[1],s6277[2],s6277[3],s5091[0]};
    CLA_4_c KS_6910(s6910, c6910, in6910_1, in6910_2, s6275[2]);
    wire[3:0] s6911, in6911_1, in6911_2;
    wire c6911;
    assign in6911_1 = {s6279[0],s6278[2],c6277,s5092[0]};
    assign in6911_2 = {s6280[0],s6279[1],s6278[3],s5093[0]};
    CLA_4_c KS_6911(s6911, c6911, in6911_1, in6911_2, s6278[1]);
    wire[3:0] s6912, in6912_1, in6912_2;
    wire c6912;
    assign in6912_1 = {s6281[1],s6279[2],c6278,c6280};
    assign in6912_2 = {s6282[0],s6280[2],s6279[3],c6281};
    CLA_4_c KS_6912(s6912, c6912, in6912_1, in6912_2, s6280[1]);
    wire[3:0] s6913, in6913_1, in6913_2;
    wire c6913;
    assign in6913_1 = {s6282[1],s6280[3],s6282[3],s5097[0]};
    assign in6913_2 = {s6283[1],s6281[3],s6283[3],c6282};
    CLA_4_c KS_6913(s6913, c6913, in6913_1, in6913_2, s6281[2]);
    wire[3:0] s6914, in6914_1, in6914_2;
    wire c6914;
    assign in6914_1 = {s6283[2],s6284[2],c6283,s5100[0]};
    assign in6914_2 = {s6284[1],s6285[1],s6284[3],s5101[0]};
    CLA_4_c KS_6914(s6914, c6914, in6914_1, in6914_2, s6282[2]);
    wire[3:0] s6915, in6915_1, in6915_2;
    wire c6915;
    assign in6915_1 = {s6287[0],s6285[2],c6284,s5103[0]};
    assign in6915_2 = {s6288[0],s6286[1],s6285[3],s5104[0]};
    CLA_4_c KS_6915(s6915, c6915, in6915_1, in6915_2, s6286[0]);
    wire[3:0] s6916, in6916_1, in6916_2;
    wire c6916;
    assign in6916_1 = {s6288[1],s6286[2],c6285,c6289};
    assign in6916_2 = {s6289[1],s6287[2],s6286[3],s6290[3]};
    CLA_4_c KS_6916(s6916, c6916, in6916_1, in6916_2, s6287[1]);
    wire[3:0] s6917, in6917_1, in6917_2;
    wire c6917;
    assign in6917_1 = {s6289[2],s6287[3],s6291[2],c6290};
    assign in6917_2 = {s6290[1],s6288[3],s6292[1],s6291[3]};
    CLA_4_c KS_6917(s6917, c6917, in6917_1, in6917_2, s6288[2]);
    wire[3:0] s6918, in6918_1, in6918_2;
    wire c6918;
    assign in6918_1 = {s6290[2],s6293[0],s6292[2],s5114[0]};
    assign in6918_2 = {s6291[1],s6294[0],s6293[1],s5115[0]};
    CLA_4_c KS_6918(s6918, c6918, in6918_1, in6918_2, s6289[3]);
    wire[3:0] s6919, in6919_1, in6919_2;
    wire c6919;
    assign in6919_1 = {s6296[0],s6294[1],c6291,s5116[0]};
    assign in6919_2 = {s6297[0],s6295[1],s6292[3],s5117[0]};
    CLA_4_c KS_6919(s6919, c6919, in6919_1, in6919_2, s6295[0]);
    wire[3:0] s6920, in6920_1, in6920_2;
    wire c6920;
    assign in6920_1 = {s6296[1],s6293[2],c6292,s6300[0]};
    assign in6920_2 = {s6297[1],s6294[2],s6293[3],s6301[0]};
    CLA_4 KS_6920(s6920, c6920, in6920_1, in6920_2);
    wire[3:0] s6921, in6921_1, in6921_2;
    wire c6921;
    assign in6921_1 = {s6296[2],s6294[3],s6302[0],s6301[1]};
    assign in6921_2 = {s6297[2],s6295[3],s6303[0],s6302[1]};
    CLA_4_c KS_6921(s6921, c6921, in6921_1, in6921_2, s6295[2]);
    wire[3:0] s6922, in6922_1, in6922_2;
    wire c6922;
    assign in6922_1 = {s6297[3],s6304[0],s6303[1],s6299[3]};
    assign in6922_2 = {s6298[3],s6305[0],s6304[1],s6300[2]};
    CLA_4_c KS_6922(s6922, c6922, in6922_1, in6922_2, s6296[3]);
    wire[3:0] s6923, in6923_1, in6923_2;
    wire c6923;
    assign in6923_1 = {s6307[0],s6305[1],s6301[2],s5131[1]};
    assign in6923_2 = {s6308[0],c6306,s6302[2],c6299};
    CLA_4_c KS_6923(s6923, c6923, in6923_1, in6923_2, s6306[0]);
    wire[3:0] s6924, in6924_1, in6924_2;
    wire c6924;
    assign in6924_1 = {s6307[1],s6303[2],s6300[3],s6312[0]};
    assign in6924_2 = {c6308,s6304[2],s6301[3],s6313[0]};
    CLA_4 KS_6924(s6924, c6924, in6924_1, in6924_2);
    wire[3:0] s6925, in6925_1, in6925_2;
    wire c6925;
    assign in6925_1 = {s6305[2],s6302[3],s6314[0],s6312[1]};
    assign in6925_2 = {c6307,s6303[3],s6315[0],s6313[1]};
    CLA_4 KS_6925(s6925, c6925, in6925_1, in6925_2);
    wire[3:0] s6926, in6926_1, in6926_2;
    wire c6926;
    assign in6926_1 = {s6304[3],s6316[0],s6314[1],s6310[2]};
    assign in6926_2 = {s6305[3],s6317[0],s6315[1],s6311[2]};
    CLA_4 KS_6926(s6926, c6926, in6926_1, in6926_2);
    wire[3:0] s6927, in6927_1, in6927_2;
    wire c6927;
    assign in6927_1 = {s6319[0],s6316[1],s6312[2],s5151[1]};
    assign in6927_2 = {s6320[0],c6317,s6313[2],s6310[3]};
    CLA_4_c KS_6927(s6927, c6927, in6927_1, in6927_2, s6318[0]);
    wire[3:0] s6928, in6928_1, in6928_2;
    wire c6928;
    assign in6928_1 = {c6319,s6314[2],s6311[3],s6323[0]};
    assign in6928_2 = {s6320[1],s6315[2],s6312[3],s6324[0]};
    CLA_4_c KS_6928(s6928, c6928, in6928_1, in6928_2, s6318[1]);
    wire[3:0] s6929, in6929_1, in6929_2;
    wire c6929;
    assign in6929_1 = {s6316[2],s6313[3],s6325[0],s6323[1]};
    assign in6929_2 = {c6318,s6314[3],s6326[0],s6324[1]};
    CLA_4 KS_6929(s6929, c6929, in6929_1, in6929_2);
    wire[3:0] s6930, in6930_1, in6930_2;
    wire c6930;
    assign in6930_1 = {s6315[3],s6327[0],s6325[1],s5173[0]};
    assign in6930_2 = {c6316,s6328[0],s6326[1],s5174[0]};
    CLA_4 KS_6930(s6930, c6930, in6930_1, in6930_2);
    wire[3:0] s6931, in6931_1, in6931_2;
    wire c6931;
    assign in6931_1 = {s6330[0],s6327[1],s6322[2],s5173[1]};
    assign in6931_2 = {s6331[0],c6328,s6323[2],c5174};
    CLA_4_c KS_6931(s6931, c6931, in6931_1, in6931_2, s6329[0]);
    wire[3:0] s6932, in6932_1, in6932_2;
    wire c6932;
    assign in6932_1 = {c6330,s6324[2],s6322[3],s6335[0]};
    assign in6932_2 = {s6331[1],s6325[2],s6323[3],s6336[0]};
    CLA_4_c KS_6932(s6932, c6932, in6932_1, in6932_2, s6329[1]);
    wire[3:0] s6933, in6933_1, in6933_2;
    wire c6933;
    assign in6933_1 = {s6327[2],s6324[3],s6337[0],s6336[1]};
    assign in6933_2 = {s6329[2],s6325[3],s6338[0],s6337[1]};
    CLA_4_c KS_6933(s6933, c6933, in6933_1, in6933_2, s6326[2]);
    wire[3:0] s6934, in6934_1, in6934_2;
    wire c6934;
    assign in6934_1 = {s6326[3],s6339[0],s6338[1],s6333[2]};
    assign in6934_2 = {s6327[3],s6340[0],c6339,s6334[2]};
    CLA_4 KS_6934(s6934, c6934, in6934_1, in6934_2);
    wire[3:0] s6935, in6935_1, in6935_2;
    wire c6935;
    assign in6935_1 = {s6342[0],s6340[1],s6335[2],s5196[1]};
    assign in6935_2 = {s6343[0],c6341,s6336[2],c5197};
    CLA_4_c KS_6935(s6935, c6935, in6935_1, in6935_2, s6341[0]);
    wire[3:0] s6936, in6936_1, in6936_2;
    wire c6936;
    assign in6936_1 = {s6342[1],s6337[2],s6333[3],s6347[0]};
    assign in6936_2 = {c6343,s6338[2],s6334[3],s6348[0]};
    CLA_4 KS_6936(s6936, c6936, in6936_1, in6936_2);
    wire[3:0] s6937, in6937_1, in6937_2;
    wire c6937;
    assign in6937_1 = {s6340[2],s6335[3],s6349[0],s6348[1]};
    assign in6937_2 = {c6342,s6336[3],s6350[0],s6349[1]};
    CLA_4 KS_6937(s6937, c6937, in6937_1, in6937_2);
    wire[3:0] s6938, in6938_1, in6938_2;
    wire c6938;
    assign in6938_1 = {s6338[3],s6351[0],s6350[1],s6345[2]};
    assign in6938_2 = {s6340[3],s6352[0],c6351,s6346[2]};
    CLA_4_c KS_6938(s6938, c6938, in6938_1, in6938_2, s6337[3]);
    wire[3:0] s6939, in6939_1, in6939_2;
    wire c6939;
    assign in6939_1 = {s6354[0],s6352[1],s6347[2],s5219[1]};
    assign in6939_2 = {s6355[0],c6353,s6348[2],s6345[3]};
    CLA_4_c KS_6939(s6939, c6939, in6939_1, in6939_2, s6353[0]);
    wire[3:0] s6940, in6940_1, in6940_2;
    wire c6940;
    assign in6940_1 = {s6354[1],s6349[2],s6346[3],s6359[0]};
    assign in6940_2 = {c6355,s6350[2],s6347[3],s6360[0]};
    CLA_4 KS_6940(s6940, c6940, in6940_1, in6940_2);
    wire[3:0] s6941, in6941_1, in6941_2;
    wire c6941;
    assign in6941_1 = {s6352[2],s6348[3],s6361[0],s6360[1]};
    assign in6941_2 = {c6354,s6349[3],s6362[0],s6361[1]};
    CLA_4 KS_6941(s6941, c6941, in6941_1, in6941_2);
    wire[3:0] s6942, in6942_1, in6942_2;
    wire c6942;
    assign in6942_1 = {s6350[3],s6363[0],s6362[1],s6357[2]};
    assign in6942_2 = {c6352,s6364[0],c6363,s6358[2]};
    CLA_4 KS_6942(s6942, c6942, in6942_1, in6942_2);
    wire[3:0] s6943, in6943_1, in6943_2;
    wire c6943;
    assign in6943_1 = {s6366[0],s6364[1],s6359[2],s5241[1]};
    assign in6943_2 = {s6367[0],c6365,s6360[2],s6357[3]};
    CLA_4_c KS_6943(s6943, c6943, in6943_1, in6943_2, s6365[0]);
    wire[3:0] s6944, in6944_1, in6944_2;
    wire c6944;
    assign in6944_1 = {s6366[1],s6361[2],s6358[3],s6371[0]};
    assign in6944_2 = {c6367,s6362[2],s6359[3],s6372[0]};
    CLA_4 KS_6944(s6944, c6944, in6944_1, in6944_2);
    wire[3:0] s6945, in6945_1, in6945_2;
    wire c6945;
    assign in6945_1 = {s6364[2],s6360[3],s6373[0],s6372[1]};
    assign in6945_2 = {c6366,s6361[3],s6374[0],s6373[1]};
    CLA_4 KS_6945(s6945, c6945, in6945_1, in6945_2);
    wire[3:0] s6946, in6946_1, in6946_2;
    wire c6946;
    assign in6946_1 = {s6362[3],s6375[0],s6374[1],s6369[2]};
    assign in6946_2 = {c6364,s6376[0],c6375,s6370[2]};
    CLA_4 KS_6946(s6946, c6946, in6946_1, in6946_2);
    wire[3:0] s6947, in6947_1, in6947_2;
    wire c6947;
    assign in6947_1 = {s6378[0],s6376[1],s6371[2],s5262[1]};
    assign in6947_2 = {s6379[0],c6377,s6372[2],c5263};
    CLA_4_c KS_6947(s6947, c6947, in6947_1, in6947_2, s6377[0]);
    wire[3:0] s6948, in6948_1, in6948_2;
    wire c6948;
    assign in6948_1 = {s6378[1],s6373[2],s6369[3],s6382[0]};
    assign in6948_2 = {c6379,s6374[2],s6370[3],s6383[0]};
    CLA_4 KS_6948(s6948, c6948, in6948_1, in6948_2);
    wire[3:0] s6949, in6949_1, in6949_2;
    wire c6949;
    assign in6949_1 = {s6376[2],s6371[3],s6384[0],s6382[1]};
    assign in6949_2 = {c6378,s6372[3],s6385[0],s6383[1]};
    CLA_4 KS_6949(s6949, c6949, in6949_1, in6949_2);
    wire[3:0] s6950, in6950_1, in6950_2;
    wire c6950;
    assign in6950_1 = {s6374[3],s6386[0],s6384[1],s5284[0]};
    assign in6950_2 = {s6376[3],s6387[0],s6385[1],s5285[0]};
    CLA_4_c KS_6950(s6950, c6950, in6950_1, in6950_2, s6373[3]);
    wire[3:0] s6951, in6951_1, in6951_2;
    wire c6951;
    assign in6951_1 = {s6389[0],s6386[1],s6381[2],s5283[1]};
    assign in6951_2 = {s6390[0],c6387,s6382[2],c5284};
    CLA_4_c KS_6951(s6951, c6951, in6951_1, in6951_2, s6388[0]);
    wire[3:0] s6952, in6952_1, in6952_2;
    wire c6952;
    assign in6952_1 = {c6389,s6383[2],s5285[1],s6392[0]};
    assign in6952_2 = {s6390[1],s6384[2],s6381[3],s6393[0]};
    CLA_4_c KS_6952(s6952, c6952, in6952_1, in6952_2, s6388[1]);
    wire[3:0] s6953, in6953_1, in6953_2;
    wire c6953;
    assign in6953_1 = {s6386[2],s6382[3],s6394[0],s6393[1]};
    assign in6953_2 = {s6388[2],s6383[3],s6395[0],s6394[1]};
    CLA_4_c KS_6953(s6953, c6953, in6953_1, in6953_2, s6385[2]);
    wire[3:0] s6954, in6954_1, in6954_2;
    wire c6954;
    assign in6954_1 = {s6385[3],s6396[0],s6395[1],s5307[0]};
    assign in6954_2 = {s6386[3],s6397[0],s6396[1],s5308[0]};
    CLA_4_c KS_6954(s6954, c6954, in6954_1, in6954_2, s6384[3]);
    wire[3:0] s6955, in6955_1, in6955_2;
    wire c6955;
    assign in6955_1 = {s6399[0],s6397[1],s6392[2],s5307[1]};
    assign in6955_2 = {s6400[0],c6398,s6393[2],c5308};
    CLA_4_c KS_6955(s6955, c6955, in6955_1, in6955_2, s6398[0]);
    wire[3:0] s6956, in6956_1, in6956_2;
    wire c6956;
    assign in6956_1 = {s6399[1],s6394[2],s6392[3],s6403[0]};
    assign in6956_2 = {c6400,s6395[2],s6393[3],s6404[0]};
    CLA_4 KS_6956(s6956, c6956, in6956_1, in6956_2);
    wire[3:0] s6957, in6957_1, in6957_2;
    wire c6957;
    assign in6957_1 = {s6397[2],s6394[3],s6405[0],s6403[1]};
    assign in6957_2 = {s6399[2],s6395[3],s6406[0],s6404[1]};
    CLA_4_c KS_6957(s6957, c6957, in6957_1, in6957_2, s6396[2]);
    wire[3:0] s6958, in6958_1, in6958_2;
    wire c6958;
    assign in6958_1 = {s6396[3],s6407[0],s6405[1],s5330[0]};
    assign in6958_2 = {s6397[3],s6408[0],s6406[1],s5331[0]};
    CLA_4 KS_6958(s6958, c6958, in6958_1, in6958_2);
    wire[3:0] s6959, in6959_1, in6959_2;
    wire c6959;
    assign in6959_1 = {s6410[0],s6407[1],s6402[2],s5330[1]};
    assign in6959_2 = {s6411[0],c6408,s6403[2],c5331};
    CLA_4_c KS_6959(s6959, c6959, in6959_1, in6959_2, s6409[0]);
    wire[3:0] s6960, in6960_1, in6960_2;
    wire c6960;
    assign in6960_1 = {c6410,s6404[2],s6402[3],s6415[0]};
    assign in6960_2 = {s6411[1],s6405[2],s6403[3],s6416[0]};
    CLA_4_c KS_6960(s6960, c6960, in6960_1, in6960_2, s6409[1]);
    wire[3:0] s6961, in6961_1, in6961_2;
    wire c6961;
    assign in6961_1 = {s6407[2],s6404[3],s6417[0],s6416[1]};
    assign in6961_2 = {s6409[2],s6405[3],s6418[0],s6417[1]};
    CLA_4_c KS_6961(s6961, c6961, in6961_1, in6961_2, s6406[2]);
    wire[3:0] s6962, in6962_1, in6962_2;
    wire c6962;
    assign in6962_1 = {s6406[3],s6419[0],s6418[1],s6413[2]};
    assign in6962_2 = {s6407[3],s6420[0],c6419,s6414[2]};
    CLA_4 KS_6962(s6962, c6962, in6962_1, in6962_2);
    wire[3:0] s6963, in6963_1, in6963_2;
    wire c6963;
    assign in6963_1 = {s6422[0],s6420[1],s6415[2],s5353[1]};
    assign in6963_2 = {s6423[0],c6421,s6416[2],s6413[3]};
    CLA_4_c KS_6963(s6963, c6963, in6963_1, in6963_2, s6421[0]);
    wire[3:0] s6964, in6964_1, in6964_2;
    wire c6964;
    assign in6964_1 = {s6422[1],s6417[2],s6414[3],s6427[0]};
    assign in6964_2 = {c6423,s6418[2],s6415[3],s6428[0]};
    CLA_4 KS_6964(s6964, c6964, in6964_1, in6964_2);
    wire[3:0] s6965, in6965_1, in6965_2;
    wire c6965;
    assign in6965_1 = {s6420[2],s6416[3],s6429[0],s6428[1]};
    assign in6965_2 = {c6422,s6417[3],s6430[0],s6429[1]};
    CLA_4 KS_6965(s6965, c6965, in6965_1, in6965_2);
    wire[3:0] s6966, in6966_1, in6966_2;
    wire c6966;
    assign in6966_1 = {s6418[3],s6431[0],s6430[1],s6425[2]};
    assign in6966_2 = {c6420,s6432[0],c6431,s6426[2]};
    CLA_4 KS_6966(s6966, c6966, in6966_1, in6966_2);
    wire[3:0] s6967, in6967_1, in6967_2;
    wire c6967;
    assign in6967_1 = {s6434[0],s6432[1],s6427[2],s5375[1]};
    assign in6967_2 = {s6435[0],c6433,s6428[2],s6425[3]};
    CLA_4_c KS_6967(s6967, c6967, in6967_1, in6967_2, s6433[0]);
    wire[3:0] s6968, in6968_1, in6968_2;
    wire c6968;
    assign in6968_1 = {s6434[1],s6429[2],s6426[3],s6439[0]};
    assign in6968_2 = {c6435,s6430[2],s6427[3],s6440[0]};
    CLA_4 KS_6968(s6968, c6968, in6968_1, in6968_2);
    wire[3:0] s6969, in6969_1, in6969_2;
    wire c6969;
    assign in6969_1 = {s6432[2],s6428[3],s6441[0],s6440[1]};
    assign in6969_2 = {c6434,s6429[3],s6442[0],s6441[1]};
    CLA_4 KS_6969(s6969, c6969, in6969_1, in6969_2);
    wire[3:0] s6970, in6970_1, in6970_2;
    wire c6970;
    assign in6970_1 = {s6430[3],s6443[0],s6442[1],s6437[2]};
    assign in6970_2 = {c6432,s6444[0],c6443,s6438[2]};
    CLA_4 KS_6970(s6970, c6970, in6970_1, in6970_2);
    wire[3:0] s6971, in6971_1, in6971_2;
    wire c6971;
    assign in6971_1 = {s6446[0],s6444[1],s6439[2],s5397[1]};
    assign in6971_2 = {s6447[0],c6445,s6440[2],s6437[3]};
    CLA_4_c KS_6971(s6971, c6971, in6971_1, in6971_2, s6445[0]);
    wire[3:0] s6972, in6972_1, in6972_2;
    wire c6972;
    assign in6972_1 = {s6446[1],s6441[2],s6438[3],s6451[0]};
    assign in6972_2 = {c6447,s6442[2],s6439[3],s6452[0]};
    CLA_4 KS_6972(s6972, c6972, in6972_1, in6972_2);
    wire[3:0] s6973, in6973_1, in6973_2;
    wire c6973;
    assign in6973_1 = {s6444[2],s6440[3],s6453[0],s6452[1]};
    assign in6973_2 = {c6446,s6441[3],s6454[0],s6453[1]};
    CLA_4 KS_6973(s6973, c6973, in6973_1, in6973_2);
    wire[3:0] s6974, in6974_1, in6974_2;
    wire c6974;
    assign in6974_1 = {s6442[3],s6455[0],s6454[1],s6449[2]};
    assign in6974_2 = {c6444,s6456[0],c6455,s6450[2]};
    CLA_4 KS_6974(s6974, c6974, in6974_1, in6974_2);
    wire[3:0] s6975, in6975_1, in6975_2;
    wire c6975;
    assign in6975_1 = {s6458[0],s6456[1],s6451[2],s5419[1]};
    assign in6975_2 = {s6459[0],c6457,s6452[2],s6449[3]};
    CLA_4_c KS_6975(s6975, c6975, in6975_1, in6975_2, s6457[0]);
    wire[3:0] s6976, in6976_1, in6976_2;
    wire c6976;
    assign in6976_1 = {s6458[1],s6453[2],s6450[3],s6463[0]};
    assign in6976_2 = {c6459,s6454[2],s6451[3],s6464[0]};
    CLA_4 KS_6976(s6976, c6976, in6976_1, in6976_2);
    wire[3:0] s6977, in6977_1, in6977_2;
    wire c6977;
    assign in6977_1 = {s6456[2],s6452[3],s6465[0],s6464[1]};
    assign in6977_2 = {c6458,s6453[3],s6466[0],s6465[1]};
    CLA_4 KS_6977(s6977, c6977, in6977_1, in6977_2);
    wire[3:0] s6978, in6978_1, in6978_2;
    wire c6978;
    assign in6978_1 = {s6454[3],s6467[0],s6466[1],s6461[2]};
    assign in6978_2 = {c6456,s6468[0],c6467,s6462[2]};
    CLA_4 KS_6978(s6978, c6978, in6978_1, in6978_2);
    wire[3:0] s6979, in6979_1, in6979_2;
    wire c6979;
    assign in6979_1 = {s6470[0],s6468[1],s6463[2],s5442[1]};
    assign in6979_2 = {s6471[0],c6469,s6464[2],s6461[3]};
    CLA_4_c KS_6979(s6979, c6979, in6979_1, in6979_2, s6469[0]);
    wire[3:0] s6980, in6980_1, in6980_2;
    wire c6980;
    assign in6980_1 = {s6470[1],s6465[2],s6462[3],s6475[0]};
    assign in6980_2 = {c6471,s6466[2],s6463[3],s6476[0]};
    CLA_4 KS_6980(s6980, c6980, in6980_1, in6980_2);
    wire[3:0] s6981, in6981_1, in6981_2;
    wire c6981;
    assign in6981_1 = {s6468[2],s6464[3],s6477[0],s6476[1]};
    assign in6981_2 = {c6470,s6465[3],s6478[0],s6477[1]};
    CLA_4 KS_6981(s6981, c6981, in6981_1, in6981_2);
    wire[3:0] s6982, in6982_1, in6982_2;
    wire c6982;
    assign in6982_1 = {s6466[3],s6479[0],s6478[1],s6473[2]};
    assign in6982_2 = {c6468,s6480[0],c6479,s6474[2]};
    CLA_4 KS_6982(s6982, c6982, in6982_1, in6982_2);
    wire[3:0] s6983, in6983_1, in6983_2;
    wire c6983;
    assign in6983_1 = {s6482[0],s6480[1],s6475[2],s5465[1]};
    assign in6983_2 = {s6483[0],c6481,s6476[2],s6473[3]};
    CLA_4_c KS_6983(s6983, c6983, in6983_1, in6983_2, s6481[0]);
    wire[3:0] s6984, in6984_1, in6984_2;
    wire c6984;
    assign in6984_1 = {s6482[1],s6477[2],s6474[3],s6486[0]};
    assign in6984_2 = {c6483,s6478[2],s6475[3],s6487[0]};
    CLA_4 KS_6984(s6984, c6984, in6984_1, in6984_2);
    wire[3:0] s6985, in6985_1, in6985_2;
    wire c6985;
    assign in6985_1 = {s6480[2],s6476[3],s6488[0],s6486[1]};
    assign in6985_2 = {c6482,s6477[3],s6489[0],s6487[1]};
    CLA_4 KS_6985(s6985, c6985, in6985_1, in6985_2);
    wire[3:0] s6986, in6986_1, in6986_2;
    wire c6986;
    assign in6986_1 = {s6478[3],s6490[0],s6488[1],s5487[0]};
    assign in6986_2 = {c6480,s6491[0],s6489[1],s5488[0]};
    CLA_4 KS_6986(s6986, c6986, in6986_1, in6986_2);
    wire[3:0] s6987, in6987_1, in6987_2;
    wire c6987;
    assign in6987_1 = {s6493[0],s6490[1],s6485[2],s5486[1]};
    assign in6987_2 = {s6494[0],c6491,s6486[2],c5487};
    CLA_4_c KS_6987(s6987, c6987, in6987_1, in6987_2, s6492[0]);
    wire[3:0] s6988, in6988_1, in6988_2;
    wire c6988;
    assign in6988_1 = {c6493,s6487[2],s5488[1],s6497[0]};
    assign in6988_2 = {s6494[1],s6488[2],s6485[3],s6498[0]};
    CLA_4_c KS_6988(s6988, c6988, in6988_1, in6988_2, s6492[1]);
    wire[3:0] s6989, in6989_1, in6989_2;
    wire c6989;
    assign in6989_1 = {s6490[2],s6486[3],s6499[0],s6497[1]};
    assign in6989_2 = {s6492[2],s6487[3],s6500[0],s6498[1]};
    CLA_4_c KS_6989(s6989, c6989, in6989_1, in6989_2, s6489[2]);
    wire[3:0] s6990, in6990_1, in6990_2;
    wire c6990;
    assign in6990_1 = {s6489[3],s6501[0],s6499[1],s5510[0]};
    assign in6990_2 = {s6490[3],s6502[0],s6500[1],s5511[0]};
    CLA_4_c KS_6990(s6990, c6990, in6990_1, in6990_2, s6488[3]);
    wire[3:0] s6991, in6991_1, in6991_2;
    wire c6991;
    assign in6991_1 = {s6504[0],s6501[1],s6496[2],s5509[1]};
    assign in6991_2 = {s6505[0],c6502,s6497[2],c5510};
    CLA_4_c KS_6991(s6991, c6991, in6991_1, in6991_2, s6503[0]);
    wire[3:0] s6992, in6992_1, in6992_2;
    wire c6992;
    assign in6992_1 = {c6504,s6498[2],s5511[1],s6508[0]};
    assign in6992_2 = {s6505[1],s6499[2],s6496[3],s6509[0]};
    CLA_4_c KS_6992(s6992, c6992, in6992_1, in6992_2, s6503[1]);
    wire[3:0] s6993, in6993_1, in6993_2;
    wire c6993;
    assign in6993_1 = {s6501[2],s6497[3],s6510[0],s6508[1]};
    assign in6993_2 = {s6503[2],s6498[3],s6511[0],s6509[1]};
    CLA_4_c KS_6993(s6993, c6993, in6993_1, in6993_2, s6500[2]);
    wire[3:0] s6994, in6994_1, in6994_2;
    wire c6994;
    assign in6994_1 = {s6500[3],s6512[0],s6510[1],s5533[0]};
    assign in6994_2 = {s6501[3],s6513[0],s6511[1],s5534[0]};
    CLA_4_c KS_6994(s6994, c6994, in6994_1, in6994_2, s6499[3]);
    wire[3:0] s6995, in6995_1, in6995_2;
    wire c6995;
    assign in6995_1 = {s6515[0],s6512[1],s6507[2],s5532[1]};
    assign in6995_2 = {s6516[0],c6513,s6508[2],c5533};
    CLA_4_c KS_6995(s6995, c6995, in6995_1, in6995_2, s6514[0]);
    wire[3:0] s6996, in6996_1, in6996_2;
    wire c6996;
    assign in6996_1 = {c6515,s6509[2],s5534[1],s6519[0]};
    assign in6996_2 = {s6516[1],s6510[2],s6507[3],s6520[0]};
    CLA_4_c KS_6996(s6996, c6996, in6996_1, in6996_2, s6514[1]);
    wire[3:0] s6997, in6997_1, in6997_2;
    wire c6997;
    assign in6997_1 = {s6512[2],s6508[3],s6521[0],s6519[1]};
    assign in6997_2 = {s6514[2],s6509[3],s6522[0],s6520[1]};
    CLA_4_c KS_6997(s6997, c6997, in6997_1, in6997_2, s6511[2]);
    wire[3:0] s6998, in6998_1, in6998_2;
    wire c6998;
    assign in6998_1 = {s6511[3],s6523[0],s6521[1],s5556[0]};
    assign in6998_2 = {s6512[3],s6524[0],s6522[1],s5557[0]};
    CLA_4_c KS_6998(s6998, c6998, in6998_1, in6998_2, s6510[3]);
    wire[3:0] s6999, in6999_1, in6999_2;
    wire c6999;
    assign in6999_1 = {s6526[0],s6523[1],s6518[2],s5556[1]};
    assign in6999_2 = {s6527[0],c6524,s6519[2],c5557};
    CLA_4_c KS_6999(s6999, c6999, in6999_1, in6999_2, s6525[0]);
    wire[3:0] s7000, in7000_1, in7000_2;
    wire c7000;
    assign in7000_1 = {c6526,s6520[2],s6518[3],s6531[0]};
    assign in7000_2 = {s6527[1],s6521[2],s6519[3],s6532[0]};
    CLA_4_c KS_7000(s7000, c7000, in7000_1, in7000_2, s6525[1]);
    wire[3:0] s7001, in7001_1, in7001_2;
    wire c7001;
    assign in7001_1 = {s6523[2],s6520[3],s6533[0],s6532[1]};
    assign in7001_2 = {s6525[2],s6521[3],s6534[0],s6533[1]};
    CLA_4_c KS_7001(s7001, c7001, in7001_1, in7001_2, s6522[2]);
    wire[3:0] s7002, in7002_1, in7002_2;
    wire c7002;
    assign in7002_1 = {s6522[3],s6535[0],s6534[1],s6529[2]};
    assign in7002_2 = {s6523[3],s6536[0],c6535,s6530[2]};
    CLA_4 KS_7002(s7002, c7002, in7002_1, in7002_2);
    wire[3:0] s7003, in7003_1, in7003_2;
    wire c7003;
    assign in7003_1 = {s6538[0],s6536[1],s6531[2],s5579[1]};
    assign in7003_2 = {s6539[0],c6537,s6532[2],c5580};
    CLA_4_c KS_7003(s7003, c7003, in7003_1, in7003_2, s6537[0]);
    wire[3:0] s7004, in7004_1, in7004_2;
    wire c7004;
    assign in7004_1 = {s6538[1],s6533[2],s6529[3],s6542[0]};
    assign in7004_2 = {c6539,s6534[2],s6530[3],s6543[0]};
    CLA_4 KS_7004(s7004, c7004, in7004_1, in7004_2);
    wire[3:0] s7005, in7005_1, in7005_2;
    wire c7005;
    assign in7005_1 = {s6536[2],s6531[3],s6544[0],s6542[1]};
    assign in7005_2 = {c6538,s6532[3],s6545[0],s6543[1]};
    CLA_4 KS_7005(s7005, c7005, in7005_1, in7005_2);
    wire[3:0] s7006, in7006_1, in7006_2;
    wire c7006;
    assign in7006_1 = {s6534[3],s6546[0],s6544[1],s5602[0]};
    assign in7006_2 = {s6536[3],s6547[0],s6545[1],s5603[0]};
    CLA_4_c KS_7006(s7006, c7006, in7006_1, in7006_2, s6533[3]);
    wire[3:0] s7007, in7007_1, in7007_2;
    wire c7007;
    assign in7007_1 = {s6549[0],s6546[1],s6541[2],s5602[1]};
    assign in7007_2 = {s6550[0],c6547,s6542[2],c5603};
    CLA_4_c KS_7007(s7007, c7007, in7007_1, in7007_2, s6548[0]);
    wire[3:0] s7008, in7008_1, in7008_2;
    wire c7008;
    assign in7008_1 = {c6549,s6543[2],s6541[3],s6553[0]};
    assign in7008_2 = {s6550[1],s6544[2],s6542[3],s6554[0]};
    CLA_4_c KS_7008(s7008, c7008, in7008_1, in7008_2, s6548[1]);
    wire[3:0] s7009, in7009_1, in7009_2;
    wire c7009;
    assign in7009_1 = {s6546[2],s6543[3],s6555[0],s6553[1]};
    assign in7009_2 = {s6548[2],s6544[3],s6556[0],s6554[1]};
    CLA_4_c KS_7009(s7009, c7009, in7009_1, in7009_2, s6545[2]);
    wire[3:0] s7010, in7010_1, in7010_2;
    wire c7010;
    assign in7010_1 = {s6545[3],s6557[0],s6555[1],s5625[0]};
    assign in7010_2 = {s6546[3],s6558[0],s6556[1],s5626[0]};
    CLA_4 KS_7010(s7010, c7010, in7010_1, in7010_2);
    wire[3:0] s7011, in7011_1, in7011_2;
    wire c7011;
    assign in7011_1 = {s6560[0],s6557[1],s6552[2],s5624[1]};
    assign in7011_2 = {s6561[0],c6558,s6553[2],c5625};
    CLA_4_c KS_7011(s7011, c7011, in7011_1, in7011_2, s6559[0]);
    wire[3:0] s7012, in7012_1, in7012_2;
    wire c7012;
    assign in7012_1 = {c6560,s6554[2],s5626[1],s6563[0]};
    assign in7012_2 = {s6561[1],s6555[2],s6552[3],s6564[0]};
    CLA_4_c KS_7012(s7012, c7012, in7012_1, in7012_2, s6559[1]);
    wire[3:0] s7013, in7013_1, in7013_2;
    wire c7013;
    assign in7013_1 = {s6557[2],s6553[3],s6565[0],s6564[1]};
    assign in7013_2 = {s6559[2],s6554[3],s6566[0],s6565[1]};
    CLA_4_c KS_7013(s7013, c7013, in7013_1, in7013_2, s6556[2]);
    wire[3:0] s7014, in7014_1, in7014_2;
    wire c7014;
    assign in7014_1 = {s6556[3],s6567[0],s6566[1],s5648[0]};
    assign in7014_2 = {s6557[3],s6568[0],s6567[1],s5649[0]};
    CLA_4_c KS_7014(s7014, c7014, in7014_1, in7014_2, s6555[3]);
    wire[3:0] s7015, in7015_1, in7015_2;
    wire c7015;
    assign in7015_1 = {s6570[0],s6568[1],s6563[2],s5647[1]};
    assign in7015_2 = {s6571[0],c6569,s6564[2],c5648};
    CLA_4_c KS_7015(s7015, c7015, in7015_1, in7015_2, s6569[0]);
    wire[3:0] s7016, in7016_1, in7016_2;
    wire c7016;
    assign in7016_1 = {s6570[1],s6565[2],s5649[1],s6573[0]};
    assign in7016_2 = {c6571,s6566[2],s6563[3],s6574[0]};
    CLA_4 KS_7016(s7016, c7016, in7016_1, in7016_2);
    wire[3:0] s7017, in7017_1, in7017_2;
    wire c7017;
    assign in7017_1 = {s6568[2],s6564[3],s6575[0],s6574[1]};
    assign in7017_2 = {s6570[2],s6565[3],s6576[0],s6575[1]};
    CLA_4_c KS_7017(s7017, c7017, in7017_1, in7017_2, s6567[2]);
    wire[3:0] s7018, in7018_1, in7018_2;
    wire c7018;
    assign in7018_1 = {s6567[3],s6577[0],s6576[1],s5671[0]};
    assign in7018_2 = {s6568[3],s6578[0],s6577[1],s5672[0]};
    CLA_4_c KS_7018(s7018, c7018, in7018_1, in7018_2, s6566[3]);
    wire[3:0] s7019, in7019_1, in7019_2;
    wire c7019;
    assign in7019_1 = {s6580[0],s6578[1],s6573[2],s5670[1]};
    assign in7019_2 = {s6581[0],c6579,s6574[2],c5671};
    CLA_4_c KS_7019(s7019, c7019, in7019_1, in7019_2, s6579[0]);
    wire[3:0] s7020, in7020_1, in7020_2;
    wire c7020;
    assign in7020_1 = {s6580[1],s6575[2],s5672[1],s6584[0]};
    assign in7020_2 = {c6581,s6576[2],s6573[3],s6585[0]};
    CLA_4 KS_7020(s7020, c7020, in7020_1, in7020_2);
    wire[3:0] s7021, in7021_1, in7021_2;
    wire c7021;
    assign in7021_1 = {s6578[2],s6574[3],s6586[0],s6584[1]};
    assign in7021_2 = {s6580[2],s6575[3],s6587[0],s6585[1]};
    CLA_4_c KS_7021(s7021, c7021, in7021_1, in7021_2, s6577[2]);
    wire[3:0] s7022, in7022_1, in7022_2;
    wire c7022;
    assign in7022_1 = {s6577[3],s6588[0],s6586[1],s5694[0]};
    assign in7022_2 = {s6578[3],s6589[0],s6587[1],s5695[0]};
    CLA_4_c KS_7022(s7022, c7022, in7022_1, in7022_2, s6576[3]);
    wire[3:0] s7023, in7023_1, in7023_2;
    wire c7023;
    assign in7023_1 = {s6591[0],s6588[1],s6583[2],s5693[1]};
    assign in7023_2 = {s6592[0],c6589,s6584[2],c5694};
    CLA_4_c KS_7023(s7023, c7023, in7023_1, in7023_2, s6590[0]);
    wire[3:0] s7024, in7024_1, in7024_2;
    wire c7024;
    assign in7024_1 = {c6591,s6585[2],s5695[1],s6595[0]};
    assign in7024_2 = {s6592[1],s6586[2],s6583[3],s6596[0]};
    CLA_4_c KS_7024(s7024, c7024, in7024_1, in7024_2, s6590[1]);
    wire[3:0] s7025, in7025_1, in7025_2;
    wire c7025;
    assign in7025_1 = {s6588[2],s6584[3],s6597[0],s6595[1]};
    assign in7025_2 = {s6590[2],s6585[3],s6598[0],s6596[1]};
    CLA_4_c KS_7025(s7025, c7025, in7025_1, in7025_2, s6587[2]);
    wire[3:0] s7026, in7026_1, in7026_2;
    wire c7026;
    assign in7026_1 = {s6587[3],s6599[0],s6597[1],s5717[0]};
    assign in7026_2 = {s6588[3],s6600[0],s6598[1],s5718[0]};
    CLA_4_c KS_7026(s7026, c7026, in7026_1, in7026_2, s6586[3]);
    wire[3:0] s7027, in7027_1, in7027_2;
    wire c7027;
    assign in7027_1 = {s6602[0],s6599[1],s6594[2],s5716[1]};
    assign in7027_2 = {s6603[0],c6600,s6595[2],c5717};
    CLA_4_c KS_7027(s7027, c7027, in7027_1, in7027_2, s6601[0]);
    wire[3:0] s7028, in7028_1, in7028_2;
    wire c7028;
    assign in7028_1 = {c6602,s6596[2],s5718[1],s6605[0]};
    assign in7028_2 = {s6603[1],s6597[2],s6594[3],s6606[0]};
    CLA_4_c KS_7028(s7028, c7028, in7028_1, in7028_2, s6601[1]);
    wire[3:0] s7029, in7029_1, in7029_2;
    wire c7029;
    assign in7029_1 = {s6599[2],s6595[3],s6607[0],s6606[1]};
    assign in7029_2 = {s6601[2],s6596[3],s6608[0],s6607[1]};
    CLA_4_c KS_7029(s7029, c7029, in7029_1, in7029_2, s6598[2]);
    wire[3:0] s7030, in7030_1, in7030_2;
    wire c7030;
    assign in7030_1 = {s6598[3],s6609[0],s6608[1],s5740[0]};
    assign in7030_2 = {s6599[3],s6610[0],s6609[1],s5741[0]};
    CLA_4_c KS_7030(s7030, c7030, in7030_1, in7030_2, s6597[3]);
    wire[3:0] s7031, in7031_1, in7031_2;
    wire c7031;
    assign in7031_1 = {s6612[0],s6610[1],s6605[2],s5739[1]};
    assign in7031_2 = {s6613[0],c6611,s6606[2],c5740};
    CLA_4_c KS_7031(s7031, c7031, in7031_1, in7031_2, s6611[0]);
    wire[3:0] s7032, in7032_1, in7032_2;
    wire c7032;
    assign in7032_1 = {s6612[1],s6607[2],s5741[1],s6616[0]};
    assign in7032_2 = {c6613,s6608[2],s6605[3],s6617[0]};
    CLA_4 KS_7032(s7032, c7032, in7032_1, in7032_2);
    wire[3:0] s7033, in7033_1, in7033_2;
    wire c7033;
    assign in7033_1 = {s6610[2],s6606[3],s6618[0],s6616[1]};
    assign in7033_2 = {s6612[2],s6607[3],s6619[0],s6617[1]};
    CLA_4_c KS_7033(s7033, c7033, in7033_1, in7033_2, s6609[2]);
    wire[3:0] s7034, in7034_1, in7034_2;
    wire c7034;
    assign in7034_1 = {s6609[3],s6620[0],s6618[1],s5763[0]};
    assign in7034_2 = {s6610[3],s6621[0],s6619[1],s5764[0]};
    CLA_4_c KS_7034(s7034, c7034, in7034_1, in7034_2, s6608[3]);
    wire[3:0] s7035, in7035_1, in7035_2;
    wire c7035;
    assign in7035_1 = {s6623[0],s6620[1],s6615[2],s5762[1]};
    assign in7035_2 = {s6624[0],c6621,s6616[2],c5763};
    CLA_4_c KS_7035(s7035, c7035, in7035_1, in7035_2, s6622[0]);
    wire[3:0] s7036, in7036_1, in7036_2;
    wire c7036;
    assign in7036_1 = {c6623,s6617[2],s5764[1],s6626[0]};
    assign in7036_2 = {s6624[1],s6618[2],s6615[3],s6627[0]};
    CLA_4_c KS_7036(s7036, c7036, in7036_1, in7036_2, s6622[1]);
    wire[3:0] s7037, in7037_1, in7037_2;
    wire c7037;
    assign in7037_1 = {s6620[2],s6616[3],s6628[0],s6627[1]};
    assign in7037_2 = {s6622[2],s6617[3],s6629[0],s6628[1]};
    CLA_4_c KS_7037(s7037, c7037, in7037_1, in7037_2, s6619[2]);
    wire[3:0] s7038, in7038_1, in7038_2;
    wire c7038;
    assign in7038_1 = {s6619[3],s6630[0],s6629[1],s5786[0]};
    assign in7038_2 = {s6620[3],s6631[0],s6630[1],s5787[0]};
    CLA_4_c KS_7038(s7038, c7038, in7038_1, in7038_2, s6618[3]);
    wire[3:0] s7039, in7039_1, in7039_2;
    wire c7039;
    assign in7039_1 = {s6633[0],s6631[1],s6626[2],s5785[1]};
    assign in7039_2 = {s6634[0],c6632,s6627[2],c5786};
    CLA_4_c KS_7039(s7039, c7039, in7039_1, in7039_2, s6632[0]);
    wire[3:0] s7040, in7040_1, in7040_2;
    wire c7040;
    assign in7040_1 = {s6633[1],s6628[2],s5787[1],s6637[0]};
    assign in7040_2 = {c6634,s6629[2],s6626[3],s6638[0]};
    CLA_4 KS_7040(s7040, c7040, in7040_1, in7040_2);
    wire[3:0] s7041, in7041_1, in7041_2;
    wire c7041;
    assign in7041_1 = {s6631[2],s6627[3],s6639[0],s6637[1]};
    assign in7041_2 = {s6633[2],s6628[3],s6640[0],s6638[1]};
    CLA_4_c KS_7041(s7041, c7041, in7041_1, in7041_2, s6630[2]);
    wire[3:0] s7042, in7042_1, in7042_2;
    wire c7042;
    assign in7042_1 = {s6630[3],s6641[0],s6639[1],s5809[0]};
    assign in7042_2 = {s6631[3],s6642[0],s6640[1],s5810[0]};
    CLA_4_c KS_7042(s7042, c7042, in7042_1, in7042_2, s6629[3]);
    wire[3:0] s7043, in7043_1, in7043_2;
    wire c7043;
    assign in7043_1 = {s6644[0],s6641[1],s6636[2],s5809[1]};
    assign in7043_2 = {s6645[0],c6642,s6637[2],c5810};
    CLA_4_c KS_7043(s7043, c7043, in7043_1, in7043_2, s6643[0]);
    wire[3:0] s7044, in7044_1, in7044_2;
    wire c7044;
    assign in7044_1 = {c6644,s6638[2],s6636[3],s6649[0]};
    assign in7044_2 = {s6645[1],s6639[2],s6637[3],s6650[0]};
    CLA_4_c KS_7044(s7044, c7044, in7044_1, in7044_2, s6643[1]);
    wire[3:0] s7045, in7045_1, in7045_2;
    wire c7045;
    assign in7045_1 = {s6641[2],s6638[3],s6651[0],s6650[1]};
    assign in7045_2 = {s6643[2],s6639[3],s6652[0],s6651[1]};
    CLA_4_c KS_7045(s7045, c7045, in7045_1, in7045_2, s6640[2]);
    wire[3:0] s7046, in7046_1, in7046_2;
    wire c7046;
    assign in7046_1 = {s6640[3],s6653[0],s6652[1],s6647[2]};
    assign in7046_2 = {s6641[3],s6654[0],c6653,s6648[2]};
    CLA_4 KS_7046(s7046, c7046, in7046_1, in7046_2);
    wire[3:0] s7047, in7047_1, in7047_2;
    wire c7047;
    assign in7047_1 = {s6656[0],s6654[1],s6649[2],s5832[1]};
    assign in7047_2 = {s6657[0],c6655,s6650[2],s6647[3]};
    CLA_4_c KS_7047(s7047, c7047, in7047_1, in7047_2, s6655[0]);
    wire[3:0] s7048, in7048_1, in7048_2;
    wire c7048;
    assign in7048_1 = {s6656[1],s6651[2],s6648[3],s6660[0]};
    assign in7048_2 = {c6657,s6652[2],s6649[3],s6661[0]};
    CLA_4 KS_7048(s7048, c7048, in7048_1, in7048_2);
    wire[3:0] s7049, in7049_1, in7049_2;
    wire c7049;
    assign in7049_1 = {s6654[2],s6650[3],s6662[0],s6660[1]};
    assign in7049_2 = {c6656,s6651[3],s6663[0],s6661[1]};
    CLA_4 KS_7049(s7049, c7049, in7049_1, in7049_2);
    wire[3:0] s7050, in7050_1, in7050_2;
    wire c7050;
    assign in7050_1 = {s6652[3],s6664[0],s6662[1],s5854[0]};
    assign in7050_2 = {c6654,s6665[0],s6663[1],s5855[0]};
    CLA_4 KS_7050(s7050, c7050, in7050_1, in7050_2);
    wire[3:0] s7051, in7051_1, in7051_2;
    wire c7051;
    assign in7051_1 = {s6667[0],s6664[1],s6659[2],s5854[1]};
    assign in7051_2 = {s6668[0],c6665,s6660[2],c5855};
    CLA_4_c KS_7051(s7051, c7051, in7051_1, in7051_2, s6666[0]);
    wire[3:0] s7052, in7052_1, in7052_2;
    wire c7052;
    assign in7052_1 = {c6667,s6661[2],s6659[3],s6672[0]};
    assign in7052_2 = {s6668[1],s6662[2],s6660[3],s6673[0]};
    CLA_4_c KS_7052(s7052, c7052, in7052_1, in7052_2, s6666[1]);
    wire[3:0] s7053, in7053_1, in7053_2;
    wire c7053;
    assign in7053_1 = {s6664[2],s6661[3],s6674[0],s6673[1]};
    assign in7053_2 = {s6666[2],s6662[3],s6675[0],s6674[1]};
    CLA_4_c KS_7053(s7053, c7053, in7053_1, in7053_2, s6663[2]);
    wire[3:0] s7054, in7054_1, in7054_2;
    wire c7054;
    assign in7054_1 = {s6663[3],s6676[0],s6675[1],s6670[2]};
    assign in7054_2 = {s6664[3],s6677[0],c6676,s6671[2]};
    CLA_4 KS_7054(s7054, c7054, in7054_1, in7054_2);
    wire[3:0] s7055, in7055_1, in7055_2;
    wire c7055;
    assign in7055_1 = {s6679[0],s6677[1],s6672[2],s5878[1]};
    assign in7055_2 = {s6680[0],c6678,s6673[2],s6670[3]};
    CLA_4_c KS_7055(s7055, c7055, in7055_1, in7055_2, s6678[0]);
    wire[3:0] s7056, in7056_1, in7056_2;
    wire c7056;
    assign in7056_1 = {s6679[1],s6674[2],s6671[3],s6683[0]};
    assign in7056_2 = {c6680,s6675[2],s6672[3],s6684[0]};
    CLA_4 KS_7056(s7056, c7056, in7056_1, in7056_2);
    wire[3:0] s7057, in7057_1, in7057_2;
    wire c7057;
    assign in7057_1 = {s6677[2],s6673[3],s6685[0],s6683[1]};
    assign in7057_2 = {c6679,s6674[3],s6686[0],s6684[1]};
    CLA_4 KS_7057(s7057, c7057, in7057_1, in7057_2);
    wire[3:0] s7058, in7058_1, in7058_2;
    wire c7058;
    assign in7058_1 = {s6675[3],s6687[0],s6685[1],s5900[0]};
    assign in7058_2 = {c6677,s6688[0],s6686[1],s5901[0]};
    CLA_4 KS_7058(s7058, c7058, in7058_1, in7058_2);
    wire[3:0] s7059, in7059_1, in7059_2;
    wire c7059;
    assign in7059_1 = {s6690[0],s6687[1],s6682[2],s5899[1]};
    assign in7059_2 = {s6691[0],c6688,s6683[2],c5900};
    CLA_4_c KS_7059(s7059, c7059, in7059_1, in7059_2, s6689[0]);
    wire[3:0] s7060, in7060_1, in7060_2;
    wire c7060;
    assign in7060_1 = {c6690,s6684[2],s5901[1],s6694[0]};
    assign in7060_2 = {s6691[1],s6685[2],s6682[3],s6695[0]};
    CLA_4_c KS_7060(s7060, c7060, in7060_1, in7060_2, s6689[1]);
    wire[3:0] s7061, in7061_1, in7061_2;
    wire c7061;
    assign in7061_1 = {s6687[2],s6683[3],s6696[0],s6694[1]};
    assign in7061_2 = {s6689[2],s6684[3],s6697[0],s6695[1]};
    CLA_4_c KS_7061(s7061, c7061, in7061_1, in7061_2, s6686[2]);
    wire[3:0] s7062, in7062_1, in7062_2;
    wire c7062;
    assign in7062_1 = {s6686[3],s6698[0],s6696[1],s5923[0]};
    assign in7062_2 = {s6687[3],s6699[0],s6697[1],s5924[0]};
    CLA_4_c KS_7062(s7062, c7062, in7062_1, in7062_2, s6685[3]);
    wire[3:0] s7063, in7063_1, in7063_2;
    wire c7063;
    assign in7063_1 = {s6701[0],s6698[1],s6693[2],s5922[1]};
    assign in7063_2 = {s6702[0],c6699,s6694[2],c5923};
    CLA_4_c KS_7063(s7063, c7063, in7063_1, in7063_2, s6700[0]);
    wire[3:0] s7064, in7064_1, in7064_2;
    wire c7064;
    assign in7064_1 = {c6701,s6695[2],s5924[1],s6704[0]};
    assign in7064_2 = {s6702[1],s6696[2],s6693[3],s6705[0]};
    CLA_4_c KS_7064(s7064, c7064, in7064_1, in7064_2, s6700[1]);
    wire[3:0] s7065, in7065_1, in7065_2;
    wire c7065;
    assign in7065_1 = {s6698[2],s6694[3],s6706[0],s6705[1]};
    assign in7065_2 = {s6700[2],s6695[3],s6707[0],s6706[1]};
    CLA_4_c KS_7065(s7065, c7065, in7065_1, in7065_2, s6697[2]);
    wire[3:0] s7066, in7066_1, in7066_2;
    wire c7066;
    assign in7066_1 = {s6697[3],s6708[0],s6707[1],s5946[0]};
    assign in7066_2 = {s6698[3],s6709[0],s6708[1],s5947[0]};
    CLA_4_c KS_7066(s7066, c7066, in7066_1, in7066_2, s6696[3]);
    wire[3:0] s7067, in7067_1, in7067_2;
    wire c7067;
    assign in7067_1 = {s6711[0],s6709[1],s6704[2],s5945[1]};
    assign in7067_2 = {s6712[0],c6710,s6705[2],c5946};
    CLA_4_c KS_7067(s7067, c7067, in7067_1, in7067_2, s6710[0]);
    wire[3:0] s7068, in7068_1, in7068_2;
    wire c7068;
    assign in7068_1 = {s6711[1],s6706[2],s5947[1],s6715[0]};
    assign in7068_2 = {c6712,s6707[2],s6704[3],s6716[0]};
    CLA_4 KS_7068(s7068, c7068, in7068_1, in7068_2);
    wire[3:0] s7069, in7069_1, in7069_2;
    wire c7069;
    assign in7069_1 = {s6709[2],s6705[3],s6717[0],s6715[1]};
    assign in7069_2 = {s6711[2],s6706[3],s6718[0],s6716[1]};
    CLA_4_c KS_7069(s7069, c7069, in7069_1, in7069_2, s6708[2]);
    wire[3:0] s7070, in7070_1, in7070_2;
    wire c7070;
    assign in7070_1 = {s6708[3],s6719[0],s6717[1],s5969[0]};
    assign in7070_2 = {s6709[3],s6720[0],s6718[1],s5970[0]};
    CLA_4_c KS_7070(s7070, c7070, in7070_1, in7070_2, s6707[3]);
    wire[3:0] s7071, in7071_1, in7071_2;
    wire c7071;
    assign in7071_1 = {s6722[0],s6719[1],s6714[2],s5969[1]};
    assign in7071_2 = {s6723[0],c6720,s6715[2],c5970};
    CLA_4_c KS_7071(s7071, c7071, in7071_1, in7071_2, s6721[0]);
    wire[3:0] s7072, in7072_1, in7072_2;
    wire c7072;
    assign in7072_1 = {c6722,s6716[2],s6714[3],s6727[0]};
    assign in7072_2 = {s6723[1],s6717[2],s6715[3],s6728[0]};
    CLA_4_c KS_7072(s7072, c7072, in7072_1, in7072_2, s6721[1]);
    wire[3:0] s7073, in7073_1, in7073_2;
    wire c7073;
    assign in7073_1 = {s6719[2],s6716[3],s6729[0],s6728[1]};
    assign in7073_2 = {s6721[2],s6717[3],s6730[0],s6729[1]};
    CLA_4_c KS_7073(s7073, c7073, in7073_1, in7073_2, s6718[2]);
    wire[3:0] s7074, in7074_1, in7074_2;
    wire c7074;
    assign in7074_1 = {s6718[3],s6731[0],s6730[1],s6725[2]};
    assign in7074_2 = {s6719[3],s6732[0],c6731,s6726[2]};
    CLA_4 KS_7074(s7074, c7074, in7074_1, in7074_2);
    wire[3:0] s7075, in7075_1, in7075_2;
    wire c7075;
    assign in7075_1 = {s6734[0],s6732[1],s6727[2],s5992[1]};
    assign in7075_2 = {s6735[0],c6733,s6728[2],c5993};
    CLA_4_c KS_7075(s7075, c7075, in7075_1, in7075_2, s6733[0]);
    wire[3:0] s7076, in7076_1, in7076_2;
    wire c7076;
    assign in7076_1 = {s6734[1],s6729[2],s6725[3],s6739[0]};
    assign in7076_2 = {c6735,s6730[2],s6726[3],s6740[0]};
    CLA_4 KS_7076(s7076, c7076, in7076_1, in7076_2);
    wire[3:0] s7077, in7077_1, in7077_2;
    wire c7077;
    assign in7077_1 = {s6732[2],s6727[3],s6741[0],s6740[1]};
    assign in7077_2 = {c6734,s6728[3],s6742[0],s6741[1]};
    CLA_4 KS_7077(s7077, c7077, in7077_1, in7077_2);
    wire[3:0] s7078, in7078_1, in7078_2;
    wire c7078;
    assign in7078_1 = {s6730[3],s6743[0],s6742[1],s6737[2]};
    assign in7078_2 = {s6732[3],s6744[0],c6743,s6738[2]};
    CLA_4_c KS_7078(s7078, c7078, in7078_1, in7078_2, s6729[3]);
    wire[3:0] s7079, in7079_1, in7079_2;
    wire c7079;
    assign in7079_1 = {s6746[0],s6744[1],s6739[2],s6015[1]};
    assign in7079_2 = {s6747[0],c6745,s6740[2],s6737[3]};
    CLA_4_c KS_7079(s7079, c7079, in7079_1, in7079_2, s6745[0]);
    wire[3:0] s7080, in7080_1, in7080_2;
    wire c7080;
    assign in7080_1 = {s6746[1],s6741[2],s6738[3],s6751[0]};
    assign in7080_2 = {c6747,s6742[2],s6739[3],s6752[0]};
    CLA_4 KS_7080(s7080, c7080, in7080_1, in7080_2);
    wire[3:0] s7081, in7081_1, in7081_2;
    wire c7081;
    assign in7081_1 = {s6744[2],s6740[3],s6753[0],s6752[1]};
    assign in7081_2 = {c6746,s6741[3],s6754[0],s6753[1]};
    CLA_4 KS_7081(s7081, c7081, in7081_1, in7081_2);
    wire[3:0] s7082, in7082_1, in7082_2;
    wire c7082;
    assign in7082_1 = {s6742[3],s6755[0],s6754[1],s6749[2]};
    assign in7082_2 = {c6744,s6756[0],c6755,s6750[2]};
    CLA_4 KS_7082(s7082, c7082, in7082_1, in7082_2);
    wire[3:0] s7083, in7083_1, in7083_2;
    wire c7083;
    assign in7083_1 = {s6758[0],s6756[1],s6751[2],s6038[1]};
    assign in7083_2 = {s6759[0],c6757,s6752[2],s6749[3]};
    CLA_4_c KS_7083(s7083, c7083, in7083_1, in7083_2, s6757[0]);
    wire[3:0] s7084, in7084_1, in7084_2;
    wire c7084;
    assign in7084_1 = {s6758[1],s6753[2],s6750[3],s6763[0]};
    assign in7084_2 = {c6759,s6754[2],s6751[3],s6764[0]};
    CLA_4 KS_7084(s7084, c7084, in7084_1, in7084_2);
    wire[3:0] s7085, in7085_1, in7085_2;
    wire c7085;
    assign in7085_1 = {s6756[2],s6752[3],s6765[0],s6764[1]};
    assign in7085_2 = {c6758,s6753[3],s6766[0],s6765[1]};
    CLA_4 KS_7085(s7085, c7085, in7085_1, in7085_2);
    wire[3:0] s7086, in7086_1, in7086_2;
    wire c7086;
    assign in7086_1 = {s6754[3],s6767[0],s6766[1],s6761[2]};
    assign in7086_2 = {c6756,s6768[0],c6767,s6762[2]};
    CLA_4 KS_7086(s7086, c7086, in7086_1, in7086_2);
    wire[3:0] s7087, in7087_1, in7087_2;
    wire c7087;
    assign in7087_1 = {s6770[0],s6768[1],s6763[2],s6059[1]};
    assign in7087_2 = {s6771[0],c6769,s6764[2],c6060};
    CLA_4_c KS_7087(s7087, c7087, in7087_1, in7087_2, s6769[0]);
    wire[3:0] s7088, in7088_1, in7088_2;
    wire c7088;
    assign in7088_1 = {s6770[1],s6765[2],s6761[3],s6774[0]};
    assign in7088_2 = {c6771,s6766[2],s6762[3],s6775[0]};
    CLA_4 KS_7088(s7088, c7088, in7088_1, in7088_2);
    wire[3:0] s7089, in7089_1, in7089_2;
    wire c7089;
    assign in7089_1 = {s6768[2],s6763[3],s6776[0],s6774[1]};
    assign in7089_2 = {c6770,s6764[3],s6777[0],s6775[1]};
    CLA_4 KS_7089(s7089, c7089, in7089_1, in7089_2);
    wire[3:0] s7090, in7090_1, in7090_2;
    wire c7090;
    assign in7090_1 = {s6766[3],s6778[0],s6776[1],s6082[0]};
    assign in7090_2 = {s6768[3],s6779[0],s6777[1],s6083[0]};
    CLA_4_c KS_7090(s7090, c7090, in7090_1, in7090_2, s6765[3]);
    wire[3:0] s7091, in7091_1, in7091_2;
    wire c7091;
    assign in7091_1 = {s6781[0],s6778[1],s6773[2],s6082[1]};
    assign in7091_2 = {s6782[0],c6779,s6774[2],c6083};
    CLA_4_c KS_7091(s7091, c7091, in7091_1, in7091_2, s6780[0]);
    wire[3:0] s7092, in7092_1, in7092_2;
    wire c7092;
    assign in7092_1 = {c6781,s6775[2],s6773[3],s6785[0]};
    assign in7092_2 = {s6782[1],s6776[2],s6774[3],s6786[0]};
    CLA_4_c KS_7092(s7092, c7092, in7092_1, in7092_2, s6780[1]);
    wire[3:0] s7093, in7093_1, in7093_2;
    wire c7093;
    assign in7093_1 = {s6778[2],s6775[3],s6787[0],s6785[1]};
    assign in7093_2 = {s6780[2],s6776[3],s6788[0],s6786[1]};
    CLA_4_c KS_7093(s7093, c7093, in7093_1, in7093_2, s6777[2]);
    wire[3:0] s7094, in7094_1, in7094_2;
    wire c7094;
    assign in7094_1 = {s6777[3],s6789[0],s6787[1],s6104[0]};
    assign in7094_2 = {s6778[3],s6790[0],s6788[1],s6105[0]};
    CLA_4 KS_7094(s7094, c7094, in7094_1, in7094_2);
    wire[3:0] s7095, in7095_1, in7095_2;
    wire c7095;
    assign in7095_1 = {s6792[0],s6789[1],s6784[2],s6103[1]};
    assign in7095_2 = {s6793[0],c6790,s6785[2],c6104};
    CLA_4_c KS_7095(s7095, c7095, in7095_1, in7095_2, s6791[0]);
    wire[3:0] s7096, in7096_1, in7096_2;
    wire c7096;
    assign in7096_1 = {c6792,s6786[2],s6105[1],s6795[0]};
    assign in7096_2 = {s6793[1],s6787[2],s6784[3],s6796[0]};
    CLA_4_c KS_7096(s7096, c7096, in7096_1, in7096_2, s6791[1]);
    wire[3:0] s7097, in7097_1, in7097_2;
    wire c7097;
    assign in7097_1 = {s6789[2],s6785[3],s6797[0],s6796[1]};
    assign in7097_2 = {s6791[2],s6786[3],s6798[0],s6797[1]};
    CLA_4_c KS_7097(s7097, c7097, in7097_1, in7097_2, s6788[2]);
    wire[3:0] s7098, in7098_1, in7098_2;
    wire c7098;
    assign in7098_1 = {s6788[3],s6799[0],s6798[1],s6127[0]};
    assign in7098_2 = {s6789[3],s6800[0],s6799[1],s6128[0]};
    CLA_4_c KS_7098(s7098, c7098, in7098_1, in7098_2, s6787[3]);
    wire[3:0] s7099, in7099_1, in7099_2;
    wire c7099;
    assign in7099_1 = {s6802[0],s6800[1],s6795[2],s6126[1]};
    assign in7099_2 = {s6803[0],c6801,s6796[2],c6127};
    CLA_4_c KS_7099(s7099, c7099, in7099_1, in7099_2, s6801[0]);
    wire[3:0] s7100, in7100_1, in7100_2;
    wire c7100;
    assign in7100_1 = {s6802[1],s6797[2],s6128[1],s6805[0]};
    assign in7100_2 = {c6803,s6798[2],s6795[3],s6806[0]};
    CLA_4 KS_7100(s7100, c7100, in7100_1, in7100_2);
    wire[3:0] s7101, in7101_1, in7101_2;
    wire c7101;
    assign in7101_1 = {s6800[2],s6796[3],s6807[0],s6806[1]};
    assign in7101_2 = {s6802[2],s6797[3],s6808[0],s6807[1]};
    CLA_4_c KS_7101(s7101, c7101, in7101_1, in7101_2, s6799[2]);
    wire[3:0] s7102, in7102_1, in7102_2;
    wire c7102;
    assign in7102_1 = {s6799[3],s6809[0],s6808[1],s6150[0]};
    assign in7102_2 = {s6800[3],s6810[0],s6809[1],s6151[0]};
    CLA_4_c KS_7102(s7102, c7102, in7102_1, in7102_2, s6798[3]);
    wire[3:0] s7103, in7103_1, in7103_2;
    wire c7103;
    assign in7103_1 = {s6812[0],s6810[1],s6805[2],s6150[1]};
    assign in7103_2 = {s6813[0],c6811,s6806[2],c6151};
    CLA_4_c KS_7103(s7103, c7103, in7103_1, in7103_2, s6811[0]);
    wire[3:0] s7104, in7104_1, in7104_2;
    wire c7104;
    assign in7104_1 = {s6812[1],s6807[2],s6805[3],s6816[0]};
    assign in7104_2 = {c6813,s6808[2],s6806[3],s6817[0]};
    CLA_4 KS_7104(s7104, c7104, in7104_1, in7104_2);
    wire[3:0] s7105, in7105_1, in7105_2;
    wire c7105;
    assign in7105_1 = {s6810[2],s6807[3],s6818[0],s6816[1]};
    assign in7105_2 = {s6812[2],s6808[3],s6819[0],s6817[1]};
    CLA_4_c KS_7105(s7105, c7105, in7105_1, in7105_2, s6809[2]);
    wire[3:0] s7106, in7106_1, in7106_2;
    wire c7106;
    assign in7106_1 = {s6809[3],s6820[0],s6818[1],s6173[0]};
    assign in7106_2 = {s6810[3],s6821[0],s6819[1],s6174[0]};
    CLA_4 KS_7106(s7106, c7106, in7106_1, in7106_2);
    wire[3:0] s7107, in7107_1, in7107_2;
    wire c7107;
    assign in7107_1 = {s6823[0],s6820[1],s6815[2],s6173[1]};
    assign in7107_2 = {s6824[0],c6821,s6816[2],c6174};
    CLA_4_c KS_7107(s7107, c7107, in7107_1, in7107_2, s6822[0]);
    wire[3:0] s7108, in7108_1, in7108_2;
    wire c7108;
    assign in7108_1 = {c6823,s6817[2],s6815[3],s6828[0]};
    assign in7108_2 = {s6824[1],s6818[2],s6816[3],s6829[0]};
    CLA_4_c KS_7108(s7108, c7108, in7108_1, in7108_2, s6822[1]);
    wire[3:0] s7109, in7109_1, in7109_2;
    wire c7109;
    assign in7109_1 = {s6820[2],s6817[3],s6830[0],s6829[1]};
    assign in7109_2 = {s6822[2],s6818[3],s6831[0],s6830[1]};
    CLA_4_c KS_7109(s7109, c7109, in7109_1, in7109_2, s6819[2]);
    wire[3:0] s7110, in7110_1, in7110_2;
    wire c7110;
    assign in7110_1 = {s6819[3],s6832[0],s6831[1],s6826[2]};
    assign in7110_2 = {s6820[3],s6833[0],c6832,s6827[2]};
    CLA_4 KS_7110(s7110, c7110, in7110_1, in7110_2);
    wire[3:0] s7111, in7111_1, in7111_2;
    wire c7111;
    assign in7111_1 = {s6835[0],s6833[1],s6828[2],s6196[1]};
    assign in7111_2 = {s6836[0],c6834,s6829[2],s6826[3]};
    CLA_4_c KS_7111(s7111, c7111, in7111_1, in7111_2, s6834[0]);
    wire[3:0] s7112, in7112_1, in7112_2;
    wire c7112;
    assign in7112_1 = {s6835[1],s6830[2],s6827[3],s6839[0]};
    assign in7112_2 = {c6836,s6831[2],s6828[3],s6840[0]};
    CLA_4 KS_7112(s7112, c7112, in7112_1, in7112_2);
    wire[3:0] s7113, in7113_1, in7113_2;
    wire c7113;
    assign in7113_1 = {s6833[2],s6829[3],s6841[0],s6839[1]};
    assign in7113_2 = {c6835,s6830[3],s6842[0],s6840[1]};
    CLA_4 KS_7113(s7113, c7113, in7113_1, in7113_2);
    wire[3:0] s7114, in7114_1, in7114_2;
    wire c7114;
    assign in7114_1 = {s6831[3],s6843[0],s6841[1],s6217[0]};
    assign in7114_2 = {c6833,s6844[0],s6842[1],s6218[0]};
    CLA_4 KS_7114(s7114, c7114, in7114_1, in7114_2);
    wire[3:0] s7115, in7115_1, in7115_2;
    wire c7115;
    assign in7115_1 = {s6846[0],s6843[1],s6838[2],s6216[1]};
    assign in7115_2 = {s6847[0],c6844,s6839[2],c6217};
    CLA_4_c KS_7115(s7115, c7115, in7115_1, in7115_2, s6845[0]);
    wire[3:0] s7116, in7116_1, in7116_2;
    wire c7116;
    assign in7116_1 = {c6846,s6840[2],s6218[1],s6850[0]};
    assign in7116_2 = {s6847[1],s6841[2],s6838[3],s6851[0]};
    CLA_4_c KS_7116(s7116, c7116, in7116_1, in7116_2, s6845[1]);
    wire[3:0] s7117, in7117_1, in7117_2;
    wire c7117;
    assign in7117_1 = {s6843[2],s6839[3],s6852[0],s6850[1]};
    assign in7117_2 = {s6845[2],s6840[3],s6853[0],s6851[1]};
    CLA_4_c KS_7117(s7117, c7117, in7117_1, in7117_2, s6842[2]);
    wire[3:0] s7118, in7118_1, in7118_2;
    wire c7118;
    assign in7118_1 = {s6842[3],s6854[0],s6852[1],s6240[0]};
    assign in7118_2 = {s6843[3],s6855[0],s6853[1],s6241[0]};
    CLA_4_c KS_7118(s7118, c7118, in7118_1, in7118_2, s6841[3]);
    wire[3:0] s7119, in7119_1, in7119_2;
    wire c7119;
    assign in7119_1 = {s6857[0],s6854[1],s6849[2],s6239[1]};
    assign in7119_2 = {s6858[0],c6855,s6850[2],c6240};
    CLA_4_c KS_7119(s7119, c7119, in7119_1, in7119_2, s6856[0]);
    wire[3:0] s7120, in7120_1, in7120_2;
    wire c7120;
    assign in7120_1 = {c6857,s6851[2],s6241[1],s6860[0]};
    assign in7120_2 = {s6858[1],s6852[2],s6849[3],s6861[0]};
    CLA_4_c KS_7120(s7120, c7120, in7120_1, in7120_2, s6856[1]);
    wire[3:0] s7121, in7121_1, in7121_2;
    wire c7121;
    assign in7121_1 = {s6854[2],s6850[3],s6862[0],s6860[1]};
    assign in7121_2 = {s6856[2],s6851[3],s6863[0],s6861[1]};
    CLA_4_c KS_7121(s7121, c7121, in7121_1, in7121_2, s6853[2]);
    wire[3:0] s7122, in7122_1, in7122_2;
    wire c7122;
    assign in7122_1 = {s6853[3],s6864[0],s6862[1],s6257[0]};
    assign in7122_2 = {s6854[3],s6865[0],s6863[1],s6258[0]};
    CLA_4_c KS_7122(s7122, c7122, in7122_1, in7122_2, s6852[3]);
    wire[3:0] s7123, in7123_1, in7123_2;
    wire c7123;
    assign in7123_1 = {s6867[0],s6864[1],s6860[2],s6256[1]};
    assign in7123_2 = {s6868[0],s6865[1],s6861[2],c6257};
    CLA_4_c KS_7123(s7123, c7123, in7123_1, in7123_2, s6866[0]);
    wire[3:0] s7124, in7124_1, in7124_2;
    wire c7124;
    assign in7124_1 = {c6867,s6862[2],s6258[1],s6870[0]};
    assign in7124_2 = {s6868[1],s6863[2],s6860[3],s6871[0]};
    CLA_4_c KS_7124(s7124, c7124, in7124_1, in7124_2, s6866[1]);
    wire[3:0] s7125, in7125_1, in7125_2;
    wire c7125;
    assign in7125_1 = {s6865[2],s6861[3],s6872[0],s6871[1]};
    assign in7125_2 = {s6866[2],s6862[3],s6873[0],s6872[1]};
    CLA_4_c KS_7125(s7125, c7125, in7125_1, in7125_2, s6864[2]);
    wire[3:0] s7126, in7126_1, in7126_2;
    wire c7126;
    assign in7126_1 = {s6864[3],s6874[0],s6873[1],s6266[0]};
    assign in7126_2 = {s6865[3],s6875[0],s6874[1],s6267[0]};
    CLA_4_c KS_7126(s7126, c7126, in7126_1, in7126_2, s6863[3]);
    wire[3:0] s7127, in7127_1, in7127_2;
    wire c7127;
    assign in7127_1 = {s6877[0],s6875[1],s6870[2],s6265[1]};
    assign in7127_2 = {s6878[0],c6876,s6871[2],c6266};
    CLA_4_c KS_7127(s7127, c7127, in7127_1, in7127_2, s6876[0]);
    wire[3:0] s7128, in7128_1, in7128_2;
    wire c7128;
    assign in7128_1 = {s6877[1],s6872[2],s6267[1],s6880[0]};
    assign in7128_2 = {c6878,s6873[2],s6870[3],s6881[0]};
    CLA_4 KS_7128(s7128, c7128, in7128_1, in7128_2);
    wire[3:0] s7129, in7129_1, in7129_2;
    wire c7129;
    assign in7129_1 = {s6875[2],s6871[3],s6882[0],s6880[1]};
    assign in7129_2 = {s6877[2],s6872[3],s6883[0],s6881[1]};
    CLA_4_c KS_7129(s7129, c7129, in7129_1, in7129_2, s6874[2]);
    wire[3:0] s7130, in7130_1, in7130_2;
    wire c7130;
    assign in7130_1 = {s6874[3],s6884[0],s6882[1],c6263};
    assign in7130_2 = {s6875[3],s6885[0],s6883[1],s6268[0]};
    CLA_4_c KS_7130(s7130, c7130, in7130_1, in7130_2, s6873[3]);
    wire[3:0] s7131, in7131_1, in7131_2;
    wire c7131;
    assign in7131_1 = {s6887[0],s6884[1],s6880[2],pp126[115]};
    assign in7131_2 = {s6888[0],s6885[1],s6881[2],pp127[114]};
    CLA_4_c KS_7131(s7131, c7131, in7131_1, in7131_2, s6886[0]);
    wire[3:0] s7132, in7132_1, in7132_2;
    wire c7132;
    assign in7132_1 = {c6887,s6882[2],c6268,c6884};
    assign in7132_2 = {s6888[1],s6883[2],s6880[3],c6885};
    CLA_4_c KS_7132(s7132, c7132, in7132_1, in7132_2, s6886[1]);
    wire[3:0] s7133, in7133_1, in7133_2;
    wire c7133;
    assign in7133_1 = {s6885[2],s6881[3],s6890[0],pp126[117]};
    assign in7133_2 = {s6886[2],s6882[3],s6891[0],pp127[116]};
    CLA_4_c KS_7133(s7133, c7133, in7133_1, in7133_2, s6884[2]);
    wire[3:0] s7134, in7134_1, in7134_2;
    wire c7134;
    assign in7134_1 = {s6884[3],s6892[0],s6890[1],pp123[121]};
    assign in7134_2 = {s6885[3],s6893[0],s6891[1],pp124[120]};
    CLA_4_c KS_7134(s7134, c7134, in7134_1, in7134_2, s6883[3]);
    wire[3:0] s7135, in7135_1, in7135_2;
    wire c7135;
    assign in7135_1 = {s6895[0],s6892[1],pp125[119],pp122[123]};
    assign in7135_2 = {s6896[0],c6893,pp126[118],pp123[122]};
    CLA_4_c KS_7135(s7135, c7135, in7135_1, in7135_2, s6894[0]);
    wire[3:0] s7136, in7136_1, in7136_2;
    wire c7136;
    assign in7136_1 = {c6895,pp127[117],pp124[121],pp121[125]};
    assign in7136_2 = {s6896[1],s6890[2],pp125[120],pp122[124]};
    CLA_4_c KS_7136(s7136, c7136, in7136_1, in7136_2, s6894[1]);
    wire[3:0] s7137, in7137_1, in7137_2;
    wire c7137;
    assign in7137_1 = {c6892,pp126[119],pp123[123],pp120[127]};
    assign in7137_2 = {s6894[2],pp127[118],pp124[122],pp121[126]};
    CLA_4_c KS_7137(s7137, c7137, in7137_1, in7137_2, s6891[2]);
    wire[3:0] s7138, in7138_1, in7138_2;
    wire c7138;
    assign in7138_1 = {s6890[3],pp125[121],pp122[125],pp121[127]};
    assign in7138_2 = {c6891,pp126[120],pp123[124],pp122[126]};
    CLA_4 KS_7138(s7138, c7138, in7138_1, in7138_2);
    wire[3:0] s7139, in7139_1, in7139_2;
    wire c7139;
    assign in7139_1 = {c6890,pp124[123],pp123[125],pp122[127]};
    assign in7139_2 = {c6894,pp125[122],pp124[124],pp123[126]};
    CLA_4_c KS_7139(s7139, c7139, in7139_1, in7139_2, pp127[119]);
    wire[3:0] s7140, in7140_1, in7140_2;
    wire c7140;
    assign in7140_1 = {pp126[121],pp125[123],pp124[125],pp123[127]};
    assign in7140_2 = {pp127[120],pp126[122],pp125[124],pp124[126]};
    CLA_4 KS_7140(s7140, c7140, in7140_1, in7140_2);

    /*Stage 7*/
    wire[3:0] s7141, in7141_1, in7141_2;
    wire c7141;
    assign in7141_1 = {pp0[4],pp0[5],pp2[4],pp4[3]};
    assign in7141_2 = {pp1[3],pp1[4],pp3[3],pp5[2]};
    CLA_4 KS_7141(s7141, c7141, in7141_1, in7141_2);
    wire[3:0] s7142, in7142_1, in7142_2;
    wire c7142;
    assign in7142_1 = {pp2[3],pp4[2],pp6[1],pp6[2]};
    assign in7142_2 = {pp3[2],pp5[1],pp7[0],pp7[1]};
    CLA_4 KS_7142(s7142, c7142, in7142_1, in7142_2);
    wire[3:0] s7143, in7143_1, in7143_2;
    wire c7143;
    assign in7143_1 = {s6899[2],pp8[1],s6269[0],s6270[0]};
    assign in7143_2 = {s6900[1],pp9[0],c6899,c6900};
    CLA_4_c KS_7143(s7143, c7143, in7143_1, in7143_2, pp8[0]);
    wire[3:0] s7144, in7144_1, in7144_2;
    wire c7144;
    assign in7144_1 = {s6900[2],s6900[3],s6901[3],s6271[0]};
    assign in7144_2 = {s6901[1],s6901[2],s6902[2],c6901};
    CLA_4_c KS_7144(s7144, c7144, in7144_1, in7144_2, s6899[3]);
    wire[3:0] s7145, in7145_1, in7145_2;
    wire c7145;
    assign in7145_1 = {s6903[2],s6272[0],s6274[0],s6276[0]};
    assign in7145_2 = {s6904[1],c6902,c6903,c6904};
    CLA_4_c KS_7145(s7145, c7145, in7145_1, in7145_2, s6902[3]);
    wire[3:0] s7146, in7146_1, in7146_2;
    wire c7146;
    assign in7146_1 = {s6904[2],s6904[3],s6905[3],s6277[0]};
    assign in7146_2 = {s6905[1],s6905[2],s6906[2],c6905};
    CLA_4_c KS_7146(s7146, c7146, in7146_1, in7146_2, s6903[3]);
    wire[3:0] s7147, in7147_1, in7147_2;
    wire c7147;
    assign in7147_1 = {s6907[2],s6278[0],s6281[0],s6283[0]};
    assign in7147_2 = {s6908[1],c6906,c6907,c6908};
    CLA_4_c KS_7147(s7147, c7147, in7147_1, in7147_2, s6906[3]);
    wire[3:0] s7148, in7148_1, in7148_2;
    wire c7148;
    assign in7148_1 = {s6908[2],s6908[3],s6909[3],s6284[0]};
    assign in7148_2 = {s6909[1],s6909[2],s6910[2],c6909};
    CLA_4_c KS_7148(s7148, c7148, in7148_1, in7148_2, s6907[3]);
    wire[3:0] s7149, in7149_1, in7149_2;
    wire c7149;
    assign in7149_1 = {s6911[2],s6285[0],s6289[0],s6290[0]};
    assign in7149_2 = {s6912[1],c6910,c6911,c6912};
    CLA_4_c KS_7149(s7149, c7149, in7149_1, in7149_2, s6910[3]);
    wire[3:0] s7150, in7150_1, in7150_2;
    wire c7150;
    assign in7150_1 = {s6912[2],s6912[3],s6913[3],s6291[0]};
    assign in7150_2 = {s6913[1],s6913[2],s6914[2],c6913};
    CLA_4_c KS_7150(s7150, c7150, in7150_1, in7150_2, s6911[3]);
    wire[3:0] s7151, in7151_1, in7151_2;
    wire c7151;
    assign in7151_1 = {s6915[2],s6292[0],s6298[0],s6298[1]};
    assign in7151_2 = {s6916[1],c6914,c6915,c6916};
    CLA_4_c KS_7151(s7151, c7151, in7151_1, in7151_2, s6914[3]);
    wire[3:0] s7152, in7152_1, in7152_2;
    wire c7152;
    assign in7152_1 = {s6916[2],s6916[3],s6917[3],s6298[2]};
    assign in7152_2 = {s6917[1],s6917[2],s6918[2],c6917};
    CLA_4_c KS_7152(s7152, c7152, in7152_1, in7152_2, s6915[3]);
    wire[3:0] s7153, in7153_1, in7153_2;
    wire c7153;
    assign in7153_1 = {s6919[2],s6299[0],s6309[0],s6309[1]};
    assign in7153_2 = {s6920[1],c6918,c6919,c6920};
    CLA_4_c KS_7153(s7153, c7153, in7153_1, in7153_2, s6918[3]);
    wire[3:0] s7154, in7154_1, in7154_2;
    wire c7154;
    assign in7154_1 = {s6920[2],s6920[3],s6921[3],s6309[2]};
    assign in7154_2 = {s6921[1],s6921[2],s6922[2],c6921};
    CLA_4_c KS_7154(s7154, c7154, in7154_1, in7154_2, s6919[3]);
    wire[3:0] s7155, in7155_1, in7155_2;
    wire c7155;
    assign in7155_1 = {s6923[2],s6309[3],s6321[0],c6321};
    assign in7155_2 = {s6924[1],c6922,c6923,c6924};
    CLA_4_c KS_7155(s7155, c7155, in7155_1, in7155_2, s6922[3]);
    wire[3:0] s7156, in7156_1, in7156_2;
    wire c7156;
    assign in7156_1 = {s6924[2],s6924[3],s6925[3],s6320[2]};
    assign in7156_2 = {s6925[1],s6925[2],s6926[2],c6925};
    CLA_4_c KS_7156(s7156, c7156, in7156_1, in7156_2, s6923[3]);
    wire[3:0] s7157, in7157_1, in7157_2;
    wire c7157;
    assign in7157_1 = {s6927[2],s6320[3],s6332[0],c6332};
    assign in7157_2 = {s6928[1],c6926,c6927,c6928};
    CLA_4_c KS_7157(s7157, c7157, in7157_1, in7157_2, s6926[3]);
    wire[3:0] s7158, in7158_1, in7158_2;
    wire c7158;
    assign in7158_1 = {s6928[2],s6928[3],s6929[3],c6331};
    assign in7158_2 = {s6929[1],s6929[2],s6930[2],c6929};
    CLA_4_c KS_7158(s7158, c7158, in7158_1, in7158_2, s6927[3]);
    wire[3:0] s7159, in7159_1, in7159_2;
    wire c7159;
    assign in7159_1 = {s6931[2],s6329[3],s6344[0],s6344[1]};
    assign in7159_2 = {s6932[1],c6930,c6931,c6932};
    CLA_4_c KS_7159(s7159, c7159, in7159_1, in7159_2, s6930[3]);
    wire[3:0] s7160, in7160_1, in7160_2;
    wire c7160;
    assign in7160_1 = {s6932[2],s6932[3],s6933[3],s6344[2]};
    assign in7160_2 = {s6933[1],s6933[2],s6934[2],c6933};
    CLA_4_c KS_7160(s7160, c7160, in7160_1, in7160_2, s6931[3]);
    wire[3:0] s7161, in7161_1, in7161_2;
    wire c7161;
    assign in7161_1 = {s6935[2],c6344,s6356[0],s6356[1]};
    assign in7161_2 = {s6936[1],c6934,c6935,c6936};
    CLA_4_c KS_7161(s7161, c7161, in7161_1, in7161_2, s6934[3]);
    wire[3:0] s7162, in7162_1, in7162_2;
    wire c7162;
    assign in7162_1 = {s6936[2],s6936[3],s6937[3],s6356[2]};
    assign in7162_2 = {s6937[1],s6937[2],s6938[2],c6937};
    CLA_4_c KS_7162(s7162, c7162, in7162_1, in7162_2, s6935[3]);
    wire[3:0] s7163, in7163_1, in7163_2;
    wire c7163;
    assign in7163_1 = {s6939[2],s6356[3],s6368[0],s6368[1]};
    assign in7163_2 = {s6940[1],c6938,c6939,c6940};
    CLA_4_c KS_7163(s7163, c7163, in7163_1, in7163_2, s6938[3]);
    wire[3:0] s7164, in7164_1, in7164_2;
    wire c7164;
    assign in7164_1 = {s6940[2],s6940[3],s6941[3],s6368[2]};
    assign in7164_2 = {s6941[1],s6941[2],s6942[2],c6941};
    CLA_4_c KS_7164(s7164, c7164, in7164_1, in7164_2, s6939[3]);
    wire[3:0] s7165, in7165_1, in7165_2;
    wire c7165;
    assign in7165_1 = {s6943[2],s6368[3],s6380[0],s6380[1]};
    assign in7165_2 = {s6944[1],c6942,c6943,c6944};
    CLA_4_c KS_7165(s7165, c7165, in7165_1, in7165_2, s6942[3]);
    wire[3:0] s7166, in7166_1, in7166_2;
    wire c7166;
    assign in7166_1 = {s6944[2],s6944[3],s6945[3],s6380[2]};
    assign in7166_2 = {s6945[1],s6945[2],s6946[2],c6945};
    CLA_4_c KS_7166(s7166, c7166, in7166_1, in7166_2, s6943[3]);
    wire[3:0] s7167, in7167_1, in7167_2;
    wire c7167;
    assign in7167_1 = {s6947[2],c6380,s6391[0],c6391};
    assign in7167_2 = {s6948[1],c6946,c6947,c6948};
    CLA_4_c KS_7167(s7167, c7167, in7167_1, in7167_2, s6946[3]);
    wire[3:0] s7168, in7168_1, in7168_2;
    wire c7168;
    assign in7168_1 = {s6948[2],s6948[3],s6949[3],c6390};
    assign in7168_2 = {s6949[1],s6949[2],s6950[2],c6949};
    CLA_4_c KS_7168(s7168, c7168, in7168_1, in7168_2, s6947[3]);
    wire[3:0] s7169, in7169_1, in7169_2;
    wire c7169;
    assign in7169_1 = {s6951[2],c6388,s6401[0],s6401[1]};
    assign in7169_2 = {s6952[1],c6950,c6951,c6952};
    CLA_4_c KS_7169(s7169, c7169, in7169_1, in7169_2, s6950[3]);
    wire[3:0] s7170, in7170_1, in7170_2;
    wire c7170;
    assign in7170_1 = {s6952[2],s6952[3],s6953[3],c6401};
    assign in7170_2 = {s6953[1],s6953[2],s6954[2],c6953};
    CLA_4_c KS_7170(s7170, c7170, in7170_1, in7170_2, s6951[3]);
    wire[3:0] s7171, in7171_1, in7171_2;
    wire c7171;
    assign in7171_1 = {s6955[2],s6399[3],s6412[0],c6412};
    assign in7171_2 = {s6956[1],c6954,c6955,c6956};
    CLA_4_c KS_7171(s7171, c7171, in7171_1, in7171_2, s6954[3]);
    wire[3:0] s7172, in7172_1, in7172_2;
    wire c7172;
    assign in7172_1 = {s6956[2],s6956[3],s6957[3],c6411};
    assign in7172_2 = {s6957[1],s6957[2],s6958[2],c6957};
    CLA_4_c KS_7172(s7172, c7172, in7172_1, in7172_2, s6955[3]);
    wire[3:0] s7173, in7173_1, in7173_2;
    wire c7173;
    assign in7173_1 = {s6959[2],s6409[3],s6424[0],s6424[1]};
    assign in7173_2 = {s6960[1],c6958,c6959,c6960};
    CLA_4_c KS_7173(s7173, c7173, in7173_1, in7173_2, s6958[3]);
    wire[3:0] s7174, in7174_1, in7174_2;
    wire c7174;
    assign in7174_1 = {s6960[2],s6960[3],s6961[3],s6424[2]};
    assign in7174_2 = {s6961[1],s6961[2],s6962[2],c6961};
    CLA_4_c KS_7174(s7174, c7174, in7174_1, in7174_2, s6959[3]);
    wire[3:0] s7175, in7175_1, in7175_2;
    wire c7175;
    assign in7175_1 = {s6963[2],s6424[3],s6436[0],s6436[1]};
    assign in7175_2 = {s6964[1],c6962,c6963,c6964};
    CLA_4_c KS_7175(s7175, c7175, in7175_1, in7175_2, s6962[3]);
    wire[3:0] s7176, in7176_1, in7176_2;
    wire c7176;
    assign in7176_1 = {s6964[2],s6964[3],s6965[3],s6436[2]};
    assign in7176_2 = {s6965[1],s6965[2],s6966[2],c6965};
    CLA_4_c KS_7176(s7176, c7176, in7176_1, in7176_2, s6963[3]);
    wire[3:0] s7177, in7177_1, in7177_2;
    wire c7177;
    assign in7177_1 = {s6967[2],s6436[3],s6448[0],s6448[1]};
    assign in7177_2 = {s6968[1],c6966,c6967,c6968};
    CLA_4_c KS_7177(s7177, c7177, in7177_1, in7177_2, s6966[3]);
    wire[3:0] s7178, in7178_1, in7178_2;
    wire c7178;
    assign in7178_1 = {s6968[2],s6968[3],s6969[3],s6448[2]};
    assign in7178_2 = {s6969[1],s6969[2],s6970[2],c6969};
    CLA_4_c KS_7178(s7178, c7178, in7178_1, in7178_2, s6967[3]);
    wire[3:0] s7179, in7179_1, in7179_2;
    wire c7179;
    assign in7179_1 = {s6971[2],s6448[3],s6460[0],s6460[1]};
    assign in7179_2 = {s6972[1],c6970,c6971,c6972};
    CLA_4_c KS_7179(s7179, c7179, in7179_1, in7179_2, s6970[3]);
    wire[3:0] s7180, in7180_1, in7180_2;
    wire c7180;
    assign in7180_1 = {s6972[2],s6972[3],s6973[3],s6460[2]};
    assign in7180_2 = {s6973[1],s6973[2],s6974[2],c6973};
    CLA_4_c KS_7180(s7180, c7180, in7180_1, in7180_2, s6971[3]);
    wire[3:0] s7181, in7181_1, in7181_2;
    wire c7181;
    assign in7181_1 = {s6975[2],s6460[3],s6472[0],s6472[1]};
    assign in7181_2 = {s6976[1],c6974,c6975,c6976};
    CLA_4_c KS_7181(s7181, c7181, in7181_1, in7181_2, s6974[3]);
    wire[3:0] s7182, in7182_1, in7182_2;
    wire c7182;
    assign in7182_1 = {s6976[2],s6976[3],s6977[3],s6472[2]};
    assign in7182_2 = {s6977[1],s6977[2],s6978[2],c6977};
    CLA_4_c KS_7182(s7182, c7182, in7182_1, in7182_2, s6975[3]);
    wire[3:0] s7183, in7183_1, in7183_2;
    wire c7183;
    assign in7183_1 = {s6979[2],s6472[3],s6484[0],s6484[1]};
    assign in7183_2 = {s6980[1],c6978,c6979,c6980};
    CLA_4_c KS_7183(s7183, c7183, in7183_1, in7183_2, s6978[3]);
    wire[3:0] s7184, in7184_1, in7184_2;
    wire c7184;
    assign in7184_1 = {s6980[2],s6980[3],s6981[3],s6484[2]};
    assign in7184_2 = {s6981[1],s6981[2],s6982[2],c6981};
    CLA_4_c KS_7184(s7184, c7184, in7184_1, in7184_2, s6979[3]);
    wire[3:0] s7185, in7185_1, in7185_2;
    wire c7185;
    assign in7185_1 = {s6983[2],s6484[3],s6495[0],c6495};
    assign in7185_2 = {s6984[1],c6982,c6983,c6984};
    CLA_4_c KS_7185(s7185, c7185, in7185_1, in7185_2, s6982[3]);
    wire[3:0] s7186, in7186_1, in7186_2;
    wire c7186;
    assign in7186_1 = {s6984[2],s6984[3],s6985[3],c6494};
    assign in7186_2 = {s6985[1],s6985[2],s6986[2],c6985};
    CLA_4_c KS_7186(s7186, c7186, in7186_1, in7186_2, s6983[3]);
    wire[3:0] s7187, in7187_1, in7187_2;
    wire c7187;
    assign in7187_1 = {s6987[2],c6492,s6506[0],c6506};
    assign in7187_2 = {s6988[1],c6986,c6987,c6988};
    CLA_4_c KS_7187(s7187, c7187, in7187_1, in7187_2, s6986[3]);
    wire[3:0] s7188, in7188_1, in7188_2;
    wire c7188;
    assign in7188_1 = {s6988[2],s6988[3],s6989[3],c6505};
    assign in7188_2 = {s6989[1],s6989[2],s6990[2],c6989};
    CLA_4_c KS_7188(s7188, c7188, in7188_1, in7188_2, s6987[3]);
    wire[3:0] s7189, in7189_1, in7189_2;
    wire c7189;
    assign in7189_1 = {s6991[2],c6503,s6517[0],c6517};
    assign in7189_2 = {s6992[1],c6990,c6991,c6992};
    CLA_4_c KS_7189(s7189, c7189, in7189_1, in7189_2, s6990[3]);
    wire[3:0] s7190, in7190_1, in7190_2;
    wire c7190;
    assign in7190_1 = {s6992[2],s6992[3],s6993[3],c6516};
    assign in7190_2 = {s6993[1],s6993[2],s6994[2],c6993};
    CLA_4_c KS_7190(s7190, c7190, in7190_1, in7190_2, s6991[3]);
    wire[3:0] s7191, in7191_1, in7191_2;
    wire c7191;
    assign in7191_1 = {s6995[2],c6514,s6528[0],c6528};
    assign in7191_2 = {s6996[1],c6994,c6995,c6996};
    CLA_4_c KS_7191(s7191, c7191, in7191_1, in7191_2, s6994[3]);
    wire[3:0] s7192, in7192_1, in7192_2;
    wire c7192;
    assign in7192_1 = {s6996[2],s6996[3],s6997[3],c6527};
    assign in7192_2 = {s6997[1],s6997[2],s6998[2],c6997};
    CLA_4_c KS_7192(s7192, c7192, in7192_1, in7192_2, s6995[3]);
    wire[3:0] s7193, in7193_1, in7193_2;
    wire c7193;
    assign in7193_1 = {s6999[2],s6525[3],s6540[0],s6540[1]};
    assign in7193_2 = {s7000[1],c6998,c6999,c7000};
    CLA_4_c KS_7193(s7193, c7193, in7193_1, in7193_2, s6998[3]);
    wire[3:0] s7194, in7194_1, in7194_2;
    wire c7194;
    assign in7194_1 = {s7000[2],s7000[3],s7001[3],s6540[2]};
    assign in7194_2 = {s7001[1],s7001[2],s7002[2],c7001};
    CLA_4_c KS_7194(s7194, c7194, in7194_1, in7194_2, s6999[3]);
    wire[3:0] s7195, in7195_1, in7195_2;
    wire c7195;
    assign in7195_1 = {s7003[2],c6540,s6551[0],c6551};
    assign in7195_2 = {s7004[1],c7002,c7003,c7004};
    CLA_4_c KS_7195(s7195, c7195, in7195_1, in7195_2, s7002[3]);
    wire[3:0] s7196, in7196_1, in7196_2;
    wire c7196;
    assign in7196_1 = {s7004[2],s7004[3],s7005[3],c6550};
    assign in7196_2 = {s7005[1],s7005[2],s7006[2],c7005};
    CLA_4_c KS_7196(s7196, c7196, in7196_1, in7196_2, s7003[3]);
    wire[3:0] s7197, in7197_1, in7197_2;
    wire c7197;
    assign in7197_1 = {s7007[2],s6548[3],s6562[0],c6562};
    assign in7197_2 = {s7008[1],c7006,c7007,c7008};
    CLA_4_c KS_7197(s7197, c7197, in7197_1, in7197_2, s7006[3]);
    wire[3:0] s7198, in7198_1, in7198_2;
    wire c7198;
    assign in7198_1 = {s7008[2],s7008[3],s7009[3],c6561};
    assign in7198_2 = {s7009[1],s7009[2],s7010[2],c7009};
    CLA_4_c KS_7198(s7198, c7198, in7198_1, in7198_2, s7007[3]);
    wire[3:0] s7199, in7199_1, in7199_2;
    wire c7199;
    assign in7199_1 = {s7011[2],c6559,s6572[0],s6572[1]};
    assign in7199_2 = {s7012[1],c7010,c7011,c7012};
    CLA_4_c KS_7199(s7199, c7199, in7199_1, in7199_2, s7010[3]);
    wire[3:0] s7200, in7200_1, in7200_2;
    wire c7200;
    assign in7200_1 = {s7012[2],s7012[3],s7013[3],c6572};
    assign in7200_2 = {s7013[1],s7013[2],s7014[2],c7013};
    CLA_4_c KS_7200(s7200, c7200, in7200_1, in7200_2, s7011[3]);
    wire[3:0] s7201, in7201_1, in7201_2;
    wire c7201;
    assign in7201_1 = {s7015[2],c6570,s6582[0],s6582[1]};
    assign in7201_2 = {s7016[1],c7014,c7015,c7016};
    CLA_4_c KS_7201(s7201, c7201, in7201_1, in7201_2, s7014[3]);
    wire[3:0] s7202, in7202_1, in7202_2;
    wire c7202;
    assign in7202_1 = {s7016[2],s7016[3],s7017[3],c6582};
    assign in7202_2 = {s7017[1],s7017[2],s7018[2],c7017};
    CLA_4_c KS_7202(s7202, c7202, in7202_1, in7202_2, s7015[3]);
    wire[3:0] s7203, in7203_1, in7203_2;
    wire c7203;
    assign in7203_1 = {s7019[2],c6580,s6593[0],c6593};
    assign in7203_2 = {s7020[1],c7018,c7019,c7020};
    CLA_4_c KS_7203(s7203, c7203, in7203_1, in7203_2, s7018[3]);
    wire[3:0] s7204, in7204_1, in7204_2;
    wire c7204;
    assign in7204_1 = {s7020[2],s7020[3],s7021[3],c6592};
    assign in7204_2 = {s7021[1],s7021[2],s7022[2],c7021};
    CLA_4_c KS_7204(s7204, c7204, in7204_1, in7204_2, s7019[3]);
    wire[3:0] s7205, in7205_1, in7205_2;
    wire c7205;
    assign in7205_1 = {s7023[2],c6590,s6604[0],c6604};
    assign in7205_2 = {s7024[1],c7022,c7023,c7024};
    CLA_4_c KS_7205(s7205, c7205, in7205_1, in7205_2, s7022[3]);
    wire[3:0] s7206, in7206_1, in7206_2;
    wire c7206;
    assign in7206_1 = {s7024[2],s7024[3],s7025[3],c6603};
    assign in7206_2 = {s7025[1],s7025[2],s7026[2],c7025};
    CLA_4_c KS_7206(s7206, c7206, in7206_1, in7206_2, s7023[3]);
    wire[3:0] s7207, in7207_1, in7207_2;
    wire c7207;
    assign in7207_1 = {s7027[2],c6601,s6614[0],s6614[1]};
    assign in7207_2 = {s7028[1],c7026,c7027,c7028};
    CLA_4_c KS_7207(s7207, c7207, in7207_1, in7207_2, s7026[3]);
    wire[3:0] s7208, in7208_1, in7208_2;
    wire c7208;
    assign in7208_1 = {s7028[2],s7028[3],s7029[3],c6614};
    assign in7208_2 = {s7029[1],s7029[2],s7030[2],c7029};
    CLA_4_c KS_7208(s7208, c7208, in7208_1, in7208_2, s7027[3]);
    wire[3:0] s7209, in7209_1, in7209_2;
    wire c7209;
    assign in7209_1 = {s7031[2],c6612,s6625[0],c6625};
    assign in7209_2 = {s7032[1],c7030,c7031,c7032};
    CLA_4_c KS_7209(s7209, c7209, in7209_1, in7209_2, s7030[3]);
    wire[3:0] s7210, in7210_1, in7210_2;
    wire c7210;
    assign in7210_1 = {s7032[2],s7032[3],s7033[3],c6624};
    assign in7210_2 = {s7033[1],s7033[2],s7034[2],c7033};
    CLA_4_c KS_7210(s7210, c7210, in7210_1, in7210_2, s7031[3]);
    wire[3:0] s7211, in7211_1, in7211_2;
    wire c7211;
    assign in7211_1 = {s7035[2],c6622,s6635[0],s6635[1]};
    assign in7211_2 = {s7036[1],c7034,c7035,c7036};
    CLA_4_c KS_7211(s7211, c7211, in7211_1, in7211_2, s7034[3]);
    wire[3:0] s7212, in7212_1, in7212_2;
    wire c7212;
    assign in7212_1 = {s7036[2],s7036[3],s7037[3],c6635};
    assign in7212_2 = {s7037[1],s7037[2],s7038[2],c7037};
    CLA_4_c KS_7212(s7212, c7212, in7212_1, in7212_2, s7035[3]);
    wire[3:0] s7213, in7213_1, in7213_2;
    wire c7213;
    assign in7213_1 = {s7039[2],c6633,s6646[0],c6646};
    assign in7213_2 = {s7040[1],c7038,c7039,c7040};
    CLA_4_c KS_7213(s7213, c7213, in7213_1, in7213_2, s7038[3]);
    wire[3:0] s7214, in7214_1, in7214_2;
    wire c7214;
    assign in7214_1 = {s7040[2],s7040[3],s7041[3],c6645};
    assign in7214_2 = {s7041[1],s7041[2],s7042[2],c7041};
    CLA_4_c KS_7214(s7214, c7214, in7214_1, in7214_2, s7039[3]);
    wire[3:0] s7215, in7215_1, in7215_2;
    wire c7215;
    assign in7215_1 = {s7043[2],s6643[3],s6658[0],s6658[1]};
    assign in7215_2 = {s7044[1],c7042,c7043,c7044};
    CLA_4_c KS_7215(s7215, c7215, in7215_1, in7215_2, s7042[3]);
    wire[3:0] s7216, in7216_1, in7216_2;
    wire c7216;
    assign in7216_1 = {s7044[2],s7044[3],s7045[3],s6658[2]};
    assign in7216_2 = {s7045[1],s7045[2],s7046[2],c7045};
    CLA_4_c KS_7216(s7216, c7216, in7216_1, in7216_2, s7043[3]);
    wire[3:0] s7217, in7217_1, in7217_2;
    wire c7217;
    assign in7217_1 = {s7047[2],s6658[3],s6669[0],c6669};
    assign in7217_2 = {s7048[1],c7046,c7047,c7048};
    CLA_4_c KS_7217(s7217, c7217, in7217_1, in7217_2, s7046[3]);
    wire[3:0] s7218, in7218_1, in7218_2;
    wire c7218;
    assign in7218_1 = {s7048[2],s7048[3],s7049[3],c6668};
    assign in7218_2 = {s7049[1],s7049[2],s7050[2],c7049};
    CLA_4_c KS_7218(s7218, c7218, in7218_1, in7218_2, s7047[3]);
    wire[3:0] s7219, in7219_1, in7219_2;
    wire c7219;
    assign in7219_1 = {s7051[2],s6666[3],s6681[0],s6681[1]};
    assign in7219_2 = {s7052[1],c7050,c7051,c7052};
    CLA_4_c KS_7219(s7219, c7219, in7219_1, in7219_2, s7050[3]);
    wire[3:0] s7220, in7220_1, in7220_2;
    wire c7220;
    assign in7220_1 = {s7052[2],s7052[3],s7053[3],s6681[2]};
    assign in7220_2 = {s7053[1],s7053[2],s7054[2],c7053};
    CLA_4_c KS_7220(s7220, c7220, in7220_1, in7220_2, s7051[3]);
    wire[3:0] s7221, in7221_1, in7221_2;
    wire c7221;
    assign in7221_1 = {s7055[2],s6681[3],s6692[0],c6692};
    assign in7221_2 = {s7056[1],c7054,c7055,c7056};
    CLA_4_c KS_7221(s7221, c7221, in7221_1, in7221_2, s7054[3]);
    wire[3:0] s7222, in7222_1, in7222_2;
    wire c7222;
    assign in7222_1 = {s7056[2],s7056[3],s7057[3],c6691};
    assign in7222_2 = {s7057[1],s7057[2],s7058[2],c7057};
    CLA_4_c KS_7222(s7222, c7222, in7222_1, in7222_2, s7055[3]);
    wire[3:0] s7223, in7223_1, in7223_2;
    wire c7223;
    assign in7223_1 = {s7059[2],c6689,s6703[0],c6703};
    assign in7223_2 = {s7060[1],c7058,c7059,c7060};
    CLA_4_c KS_7223(s7223, c7223, in7223_1, in7223_2, s7058[3]);
    wire[3:0] s7224, in7224_1, in7224_2;
    wire c7224;
    assign in7224_1 = {s7060[2],s7060[3],s7061[3],c6702};
    assign in7224_2 = {s7061[1],s7061[2],s7062[2],c7061};
    CLA_4_c KS_7224(s7224, c7224, in7224_1, in7224_2, s7059[3]);
    wire[3:0] s7225, in7225_1, in7225_2;
    wire c7225;
    assign in7225_1 = {s7063[2],c6700,s6713[0],s6713[1]};
    assign in7225_2 = {s7064[1],c7062,c7063,c7064};
    CLA_4_c KS_7225(s7225, c7225, in7225_1, in7225_2, s7062[3]);
    wire[3:0] s7226, in7226_1, in7226_2;
    wire c7226;
    assign in7226_1 = {s7064[2],s7064[3],s7065[3],c6713};
    assign in7226_2 = {s7065[1],s7065[2],s7066[2],c7065};
    CLA_4_c KS_7226(s7226, c7226, in7226_1, in7226_2, s7063[3]);
    wire[3:0] s7227, in7227_1, in7227_2;
    wire c7227;
    assign in7227_1 = {s7067[2],c6711,s6724[0],c6724};
    assign in7227_2 = {s7068[1],c7066,c7067,c7068};
    CLA_4_c KS_7227(s7227, c7227, in7227_1, in7227_2, s7066[3]);
    wire[3:0] s7228, in7228_1, in7228_2;
    wire c7228;
    assign in7228_1 = {s7068[2],s7068[3],s7069[3],c6723};
    assign in7228_2 = {s7069[1],s7069[2],s7070[2],c7069};
    CLA_4_c KS_7228(s7228, c7228, in7228_1, in7228_2, s7067[3]);
    wire[3:0] s7229, in7229_1, in7229_2;
    wire c7229;
    assign in7229_1 = {s7071[2],s6721[3],s6736[0],s6736[1]};
    assign in7229_2 = {s7072[1],c7070,c7071,c7072};
    CLA_4_c KS_7229(s7229, c7229, in7229_1, in7229_2, s7070[3]);
    wire[3:0] s7230, in7230_1, in7230_2;
    wire c7230;
    assign in7230_1 = {s7072[2],s7072[3],s7073[3],s6736[2]};
    assign in7230_2 = {s7073[1],s7073[2],s7074[2],c7073};
    CLA_4_c KS_7230(s7230, c7230, in7230_1, in7230_2, s7071[3]);
    wire[3:0] s7231, in7231_1, in7231_2;
    wire c7231;
    assign in7231_1 = {s7075[2],c6736,s6748[0],s6748[1]};
    assign in7231_2 = {s7076[1],c7074,c7075,c7076};
    CLA_4_c KS_7231(s7231, c7231, in7231_1, in7231_2, s7074[3]);
    wire[3:0] s7232, in7232_1, in7232_2;
    wire c7232;
    assign in7232_1 = {s7076[2],s7076[3],s7077[3],s6748[2]};
    assign in7232_2 = {s7077[1],s7077[2],s7078[2],c7077};
    CLA_4_c KS_7232(s7232, c7232, in7232_1, in7232_2, s7075[3]);
    wire[3:0] s7233, in7233_1, in7233_2;
    wire c7233;
    assign in7233_1 = {s7079[2],s6748[3],s6760[0],s6760[1]};
    assign in7233_2 = {s7080[1],c7078,c7079,c7080};
    CLA_4_c KS_7233(s7233, c7233, in7233_1, in7233_2, s7078[3]);
    wire[3:0] s7234, in7234_1, in7234_2;
    wire c7234;
    assign in7234_1 = {s7080[2],s7080[3],s7081[3],s6760[2]};
    assign in7234_2 = {s7081[1],s7081[2],s7082[2],c7081};
    CLA_4_c KS_7234(s7234, c7234, in7234_1, in7234_2, s7079[3]);
    wire[3:0] s7235, in7235_1, in7235_2;
    wire c7235;
    assign in7235_1 = {s7083[2],s6760[3],s6772[0],s6772[1]};
    assign in7235_2 = {s7084[1],c7082,c7083,c7084};
    CLA_4_c KS_7235(s7235, c7235, in7235_1, in7235_2, s7082[3]);
    wire[3:0] s7236, in7236_1, in7236_2;
    wire c7236;
    assign in7236_1 = {s7084[2],s7084[3],s7085[3],s6772[2]};
    assign in7236_2 = {s7085[1],s7085[2],s7086[2],c7085};
    CLA_4_c KS_7236(s7236, c7236, in7236_1, in7236_2, s7083[3]);
    wire[3:0] s7237, in7237_1, in7237_2;
    wire c7237;
    assign in7237_1 = {s7087[2],c6772,s6783[0],c6783};
    assign in7237_2 = {s7088[1],c7086,c7087,c7088};
    CLA_4_c KS_7237(s7237, c7237, in7237_1, in7237_2, s7086[3]);
    wire[3:0] s7238, in7238_1, in7238_2;
    wire c7238;
    assign in7238_1 = {s7088[2],s7088[3],s7089[3],c6782};
    assign in7238_2 = {s7089[1],s7089[2],s7090[2],c7089};
    CLA_4_c KS_7238(s7238, c7238, in7238_1, in7238_2, s7087[3]);
    wire[3:0] s7239, in7239_1, in7239_2;
    wire c7239;
    assign in7239_1 = {s7091[2],s6780[3],s6794[0],c6794};
    assign in7239_2 = {s7092[1],c7090,c7091,c7092};
    CLA_4_c KS_7239(s7239, c7239, in7239_1, in7239_2, s7090[3]);
    wire[3:0] s7240, in7240_1, in7240_2;
    wire c7240;
    assign in7240_1 = {s7092[2],s7092[3],s7093[3],c6793};
    assign in7240_2 = {s7093[1],s7093[2],s7094[2],c7093};
    CLA_4_c KS_7240(s7240, c7240, in7240_1, in7240_2, s7091[3]);
    wire[3:0] s7241, in7241_1, in7241_2;
    wire c7241;
    assign in7241_1 = {s7095[2],c6791,s6804[0],s6804[1]};
    assign in7241_2 = {s7096[1],c7094,c7095,c7096};
    CLA_4_c KS_7241(s7241, c7241, in7241_1, in7241_2, s7094[3]);
    wire[3:0] s7242, in7242_1, in7242_2;
    wire c7242;
    assign in7242_1 = {s7096[2],s7096[3],s7097[3],c6804};
    assign in7242_2 = {s7097[1],s7097[2],s7098[2],c7097};
    CLA_4_c KS_7242(s7242, c7242, in7242_1, in7242_2, s7095[3]);
    wire[3:0] s7243, in7243_1, in7243_2;
    wire c7243;
    assign in7243_1 = {s7099[2],c6802,s6814[0],s6814[1]};
    assign in7243_2 = {s7100[1],c7098,c7099,c7100};
    CLA_4_c KS_7243(s7243, c7243, in7243_1, in7243_2, s7098[3]);
    wire[3:0] s7244, in7244_1, in7244_2;
    wire c7244;
    assign in7244_1 = {s7100[2],s7100[3],s7101[3],c6814};
    assign in7244_2 = {s7101[1],s7101[2],s7102[2],c7101};
    CLA_4_c KS_7244(s7244, c7244, in7244_1, in7244_2, s7099[3]);
    wire[3:0] s7245, in7245_1, in7245_2;
    wire c7245;
    assign in7245_1 = {s7103[2],s6812[3],s6825[0],c6825};
    assign in7245_2 = {s7104[1],c7102,c7103,c7104};
    CLA_4_c KS_7245(s7245, c7245, in7245_1, in7245_2, s7102[3]);
    wire[3:0] s7246, in7246_1, in7246_2;
    wire c7246;
    assign in7246_1 = {s7104[2],s7104[3],s7105[3],c6824};
    assign in7246_2 = {s7105[1],s7105[2],s7106[2],c7105};
    CLA_4_c KS_7246(s7246, c7246, in7246_1, in7246_2, s7103[3]);
    wire[3:0] s7247, in7247_1, in7247_2;
    wire c7247;
    assign in7247_1 = {s7107[2],s6822[3],s6837[0],s6837[1]};
    assign in7247_2 = {s7108[1],c7106,c7107,c7108};
    CLA_4_c KS_7247(s7247, c7247, in7247_1, in7247_2, s7106[3]);
    wire[3:0] s7248, in7248_1, in7248_2;
    wire c7248;
    assign in7248_1 = {s7108[2],s7108[3],s7109[3],s6837[2]};
    assign in7248_2 = {s7109[1],s7109[2],s7110[2],c7109};
    CLA_4_c KS_7248(s7248, c7248, in7248_1, in7248_2, s7107[3]);
    wire[3:0] s7249, in7249_1, in7249_2;
    wire c7249;
    assign in7249_1 = {s7111[2],s6837[3],s6848[0],c6848};
    assign in7249_2 = {s7112[1],c7110,c7111,c7112};
    CLA_4_c KS_7249(s7249, c7249, in7249_1, in7249_2, s7110[3]);
    wire[3:0] s7250, in7250_1, in7250_2;
    wire c7250;
    assign in7250_1 = {s7112[2],s7112[3],s7113[3],c6847};
    assign in7250_2 = {s7113[1],s7113[2],s7114[2],c7113};
    CLA_4_c KS_7250(s7250, c7250, in7250_1, in7250_2, s7111[3]);
    wire[3:0] s7251, in7251_1, in7251_2;
    wire c7251;
    assign in7251_1 = {s7115[2],c6845,s6859[0],c6859};
    assign in7251_2 = {s7116[1],c7114,c7115,c7116};
    CLA_4_c KS_7251(s7251, c7251, in7251_1, in7251_2, s7114[3]);
    wire[3:0] s7252, in7252_1, in7252_2;
    wire c7252;
    assign in7252_1 = {s7116[2],s7116[3],s7117[3],c6858};
    assign in7252_2 = {s7117[1],s7117[2],s7118[2],c7117};
    CLA_4_c KS_7252(s7252, c7252, in7252_1, in7252_2, s7115[3]);
    wire[3:0] s7253, in7253_1, in7253_2;
    wire c7253;
    assign in7253_1 = {s7119[2],c6856,s6869[0],c6869};
    assign in7253_2 = {s7120[1],c7118,c7119,c7120};
    CLA_4_c KS_7253(s7253, c7253, in7253_1, in7253_2, s7118[3]);
    wire[3:0] s7254, in7254_1, in7254_2;
    wire c7254;
    assign in7254_1 = {s7120[2],s7120[3],s7121[3],c6868};
    assign in7254_2 = {s7121[1],s7121[2],s7122[2],c7121};
    CLA_4_c KS_7254(s7254, c7254, in7254_1, in7254_2, s7119[3]);
    wire[3:0] s7255, in7255_1, in7255_2;
    wire c7255;
    assign in7255_1 = {s7123[2],c6866,s6879[0],s6879[1]};
    assign in7255_2 = {s7124[1],c7122,c7123,c7124};
    CLA_4_c KS_7255(s7255, c7255, in7255_1, in7255_2, s7122[3]);
    wire[3:0] s7256, in7256_1, in7256_2;
    wire c7256;
    assign in7256_1 = {s7124[2],s7124[3],s7125[3],c6879};
    assign in7256_2 = {s7125[1],s7125[2],s7126[2],c7125};
    CLA_4_c KS_7256(s7256, c7256, in7256_1, in7256_2, s7123[3]);
    wire[3:0] s7257, in7257_1, in7257_2;
    wire c7257;
    assign in7257_1 = {s7127[2],c6877,s6889[0],c6889};
    assign in7257_2 = {s7128[1],c7126,c7127,c7128};
    CLA_4_c KS_7257(s7257, c7257, in7257_1, in7257_2, s7126[3]);
    wire[3:0] s7258, in7258_1, in7258_2;
    wire c7258;
    assign in7258_1 = {s7128[2],s7128[3],s7129[3],c6888};
    assign in7258_2 = {s7129[1],s7129[2],s7130[2],c7129};
    CLA_4_c KS_7258(s7258, c7258, in7258_1, in7258_2, s7127[3]);
    wire[3:0] s7259, in7259_1, in7259_2;
    wire c7259;
    assign in7259_1 = {s7131[2],c6886,s6897[0],c6897};
    assign in7259_2 = {s7132[1],c7130,c7131,c7132};
    CLA_4_c KS_7259(s7259, c7259, in7259_1, in7259_2, s7130[3]);
    wire[3:0] s7260, in7260_1, in7260_2;
    wire c7260;
    assign in7260_1 = {s7132[2],s7132[3],s7133[3],c6896};
    assign in7260_2 = {s7133[1],s7133[2],s7134[2],c7133};
    CLA_4_c KS_7260(s7260, c7260, in7260_1, in7260_2, s7131[3]);
    wire[3:0] s7261, in7261_1, in7261_2;
    wire c7261;
    assign in7261_1 = {s7135[2],s6894[3],s6898[0],c6898};
    assign in7261_2 = {s7136[1],c7134,c7135,c7136};
    CLA_4_c KS_7261(s7261, c7261, in7261_1, in7261_2, s7134[3]);
    wire[3:0] s7262, in7262_1, in7262_2;
    wire c7262;
    assign in7262_1 = {s7136[2],s7136[3],s7137[3],pp127[121]};
    assign in7262_2 = {s7137[1],s7137[2],s7138[2],c7137};
    CLA_4_c KS_7262(s7262, c7262, in7262_1, in7262_2, s7135[3]);
    wire[3:0] s7263, in7263_1, in7263_2;
    wire c7263;
    assign in7263_1 = {s7138[3],pp126[123],pp125[125],pp124[127]};
    assign in7263_2 = {s7139[2],pp127[122],pp126[124],pp125[126]};
    CLA_4 KS_7263(s7263, c7263, in7263_1, in7263_2);
    wire[3:0] s7264, in7264_1, in7264_2;
    wire c7264;
    assign in7264_1 = {c7138,pp127[123],pp126[125],pp125[127]};
    assign in7264_2 = {s7139[3],c7139,pp127[124],pp126[126]};
    CLA_4 KS_7264(s7264, c7264, in7264_1, in7264_2);

    /*Stage 8*/
    wire[3:0] s7265, in7265_1, in7265_2;
    wire c7265;
    assign in7265_1 = {pp0[3],pp2[2],pp4[1],pp6[0]};
    assign in7265_2 = {pp1[2],pp3[1],pp5[0],s6899[0]};
    CLA_4 KS_7265(s7265, c7265, in7265_1, in7265_2);
    wire[3:0] s7266, in7266_1, in7266_2;
    wire c7266;
    assign in7266_1 = {s6900[0],s6901[0],s6902[0],s6902[1]};
    assign in7266_2 = {s7141[3],c7141,c7142,s6903[0]};
    CLA_4_c KS_7266(s7266, c7266, in7266_1, in7266_2, s6899[1]);
    wire[3:0] s7267, in7267_1, in7267_2;
    wire c7267;
    assign in7267_1 = {s6904[0],s6905[0],s6906[0],s6906[1]};
    assign in7267_2 = {s7143[3],c7143,c7144,s6907[0]};
    CLA_4_c KS_7267(s7267, c7267, in7267_1, in7267_2, s6903[1]);
    wire[3:0] s7268, in7268_1, in7268_2;
    wire c7268;
    assign in7268_1 = {s6908[0],s6909[0],s6910[0],s6910[1]};
    assign in7268_2 = {s7145[3],c7145,c7146,s6911[0]};
    CLA_4_c KS_7268(s7268, c7268, in7268_1, in7268_2, s6907[1]);
    wire[3:0] s7269, in7269_1, in7269_2;
    wire c7269;
    assign in7269_1 = {s6912[0],s6913[0],s6914[0],s6914[1]};
    assign in7269_2 = {s7147[3],c7147,c7148,s6915[0]};
    CLA_4_c KS_7269(s7269, c7269, in7269_1, in7269_2, s6911[1]);
    wire[3:0] s7270, in7270_1, in7270_2;
    wire c7270;
    assign in7270_1 = {s6916[0],s6917[0],s6918[0],s6918[1]};
    assign in7270_2 = {s7149[3],c7149,c7150,s6919[0]};
    CLA_4_c KS_7270(s7270, c7270, in7270_1, in7270_2, s6915[1]);
    wire[3:0] s7271, in7271_1, in7271_2;
    wire c7271;
    assign in7271_1 = {s6920[0],s6921[0],s6922[0],s6922[1]};
    assign in7271_2 = {s7151[3],c7151,c7152,s6923[0]};
    CLA_4_c KS_7271(s7271, c7271, in7271_1, in7271_2, s6919[1]);
    wire[3:0] s7272, in7272_1, in7272_2;
    wire c7272;
    assign in7272_1 = {s6924[0],s6925[0],s6926[0],s6926[1]};
    assign in7272_2 = {s7153[3],c7153,c7154,s6927[0]};
    CLA_4_c KS_7272(s7272, c7272, in7272_1, in7272_2, s6923[1]);
    wire[3:0] s7273, in7273_1, in7273_2;
    wire c7273;
    assign in7273_1 = {s6928[0],s6929[0],s6930[0],s6930[1]};
    assign in7273_2 = {s7155[3],c7155,c7156,s6931[0]};
    CLA_4_c KS_7273(s7273, c7273, in7273_1, in7273_2, s6927[1]);
    wire[3:0] s7274, in7274_1, in7274_2;
    wire c7274;
    assign in7274_1 = {s6932[0],s6933[0],s6934[0],s6934[1]};
    assign in7274_2 = {s7157[3],c7157,c7158,s6935[0]};
    CLA_4_c KS_7274(s7274, c7274, in7274_1, in7274_2, s6931[1]);
    wire[3:0] s7275, in7275_1, in7275_2;
    wire c7275;
    assign in7275_1 = {s6936[0],s6937[0],s6938[0],s6938[1]};
    assign in7275_2 = {s7159[3],c7159,c7160,s6939[0]};
    CLA_4_c KS_7275(s7275, c7275, in7275_1, in7275_2, s6935[1]);
    wire[3:0] s7276, in7276_1, in7276_2;
    wire c7276;
    assign in7276_1 = {s6940[0],s6941[0],s6942[0],s6942[1]};
    assign in7276_2 = {s7161[3],c7161,c7162,s6943[0]};
    CLA_4_c KS_7276(s7276, c7276, in7276_1, in7276_2, s6939[1]);
    wire[3:0] s7277, in7277_1, in7277_2;
    wire c7277;
    assign in7277_1 = {s6944[0],s6945[0],s6946[0],s6946[1]};
    assign in7277_2 = {s7163[3],c7163,c7164,s6947[0]};
    CLA_4_c KS_7277(s7277, c7277, in7277_1, in7277_2, s6943[1]);
    wire[3:0] s7278, in7278_1, in7278_2;
    wire c7278;
    assign in7278_1 = {s6948[0],s6949[0],s6950[0],s6950[1]};
    assign in7278_2 = {s7165[3],c7165,c7166,s6951[0]};
    CLA_4_c KS_7278(s7278, c7278, in7278_1, in7278_2, s6947[1]);
    wire[3:0] s7279, in7279_1, in7279_2;
    wire c7279;
    assign in7279_1 = {s6952[0],s6953[0],s6954[0],s6954[1]};
    assign in7279_2 = {s7167[3],c7167,c7168,s6955[0]};
    CLA_4_c KS_7279(s7279, c7279, in7279_1, in7279_2, s6951[1]);
    wire[3:0] s7280, in7280_1, in7280_2;
    wire c7280;
    assign in7280_1 = {s6956[0],s6957[0],s6958[0],s6958[1]};
    assign in7280_2 = {s7169[3],c7169,c7170,s6959[0]};
    CLA_4_c KS_7280(s7280, c7280, in7280_1, in7280_2, s6955[1]);
    wire[3:0] s7281, in7281_1, in7281_2;
    wire c7281;
    assign in7281_1 = {s6960[0],s6961[0],s6962[0],s6962[1]};
    assign in7281_2 = {s7171[3],c7171,c7172,s6963[0]};
    CLA_4_c KS_7281(s7281, c7281, in7281_1, in7281_2, s6959[1]);
    wire[3:0] s7282, in7282_1, in7282_2;
    wire c7282;
    assign in7282_1 = {s6964[0],s6965[0],s6966[0],s6966[1]};
    assign in7282_2 = {s7173[3],c7173,c7174,s6967[0]};
    CLA_4_c KS_7282(s7282, c7282, in7282_1, in7282_2, s6963[1]);
    wire[3:0] s7283, in7283_1, in7283_2;
    wire c7283;
    assign in7283_1 = {s6968[0],s6969[0],s6970[0],s6970[1]};
    assign in7283_2 = {s7175[3],c7175,c7176,s6971[0]};
    CLA_4_c KS_7283(s7283, c7283, in7283_1, in7283_2, s6967[1]);
    wire[3:0] s7284, in7284_1, in7284_2;
    wire c7284;
    assign in7284_1 = {s6972[0],s6973[0],s6974[0],s6974[1]};
    assign in7284_2 = {s7177[3],c7177,c7178,s6975[0]};
    CLA_4_c KS_7284(s7284, c7284, in7284_1, in7284_2, s6971[1]);
    wire[3:0] s7285, in7285_1, in7285_2;
    wire c7285;
    assign in7285_1 = {s6976[0],s6977[0],s6978[0],s6978[1]};
    assign in7285_2 = {s7179[3],c7179,c7180,s6979[0]};
    CLA_4_c KS_7285(s7285, c7285, in7285_1, in7285_2, s6975[1]);
    wire[3:0] s7286, in7286_1, in7286_2;
    wire c7286;
    assign in7286_1 = {s6980[0],s6981[0],s6982[0],s6982[1]};
    assign in7286_2 = {s7181[3],c7181,c7182,s6983[0]};
    CLA_4_c KS_7286(s7286, c7286, in7286_1, in7286_2, s6979[1]);
    wire[3:0] s7287, in7287_1, in7287_2;
    wire c7287;
    assign in7287_1 = {s6984[0],s6985[0],s6986[0],s6986[1]};
    assign in7287_2 = {s7183[3],c7183,c7184,s6987[0]};
    CLA_4_c KS_7287(s7287, c7287, in7287_1, in7287_2, s6983[1]);
    wire[3:0] s7288, in7288_1, in7288_2;
    wire c7288;
    assign in7288_1 = {s6988[0],s6989[0],s6990[0],s6990[1]};
    assign in7288_2 = {s7185[3],c7185,c7186,s6991[0]};
    CLA_4_c KS_7288(s7288, c7288, in7288_1, in7288_2, s6987[1]);
    wire[3:0] s7289, in7289_1, in7289_2;
    wire c7289;
    assign in7289_1 = {s6992[0],s6993[0],s6994[0],s6994[1]};
    assign in7289_2 = {s7187[3],c7187,c7188,s6995[0]};
    CLA_4_c KS_7289(s7289, c7289, in7289_1, in7289_2, s6991[1]);
    wire[3:0] s7290, in7290_1, in7290_2;
    wire c7290;
    assign in7290_1 = {s6996[0],s6997[0],s6998[0],s6998[1]};
    assign in7290_2 = {s7189[3],c7189,c7190,s6999[0]};
    CLA_4_c KS_7290(s7290, c7290, in7290_1, in7290_2, s6995[1]);
    wire[3:0] s7291, in7291_1, in7291_2;
    wire c7291;
    assign in7291_1 = {s7000[0],s7001[0],s7002[0],s7002[1]};
    assign in7291_2 = {s7191[3],c7191,c7192,s7003[0]};
    CLA_4_c KS_7291(s7291, c7291, in7291_1, in7291_2, s6999[1]);
    wire[3:0] s7292, in7292_1, in7292_2;
    wire c7292;
    assign in7292_1 = {s7004[0],s7005[0],s7006[0],s7006[1]};
    assign in7292_2 = {s7193[3],c7193,c7194,s7007[0]};
    CLA_4_c KS_7292(s7292, c7292, in7292_1, in7292_2, s7003[1]);
    wire[3:0] s7293, in7293_1, in7293_2;
    wire c7293;
    assign in7293_1 = {s7008[0],s7009[0],s7010[0],s7010[1]};
    assign in7293_2 = {s7195[3],c7195,c7196,s7011[0]};
    CLA_4_c KS_7293(s7293, c7293, in7293_1, in7293_2, s7007[1]);
    wire[3:0] s7294, in7294_1, in7294_2;
    wire c7294;
    assign in7294_1 = {s7012[0],s7013[0],s7014[0],s7014[1]};
    assign in7294_2 = {s7197[3],c7197,c7198,s7015[0]};
    CLA_4_c KS_7294(s7294, c7294, in7294_1, in7294_2, s7011[1]);
    wire[3:0] s7295, in7295_1, in7295_2;
    wire c7295;
    assign in7295_1 = {s7016[0],s7017[0],s7018[0],s7018[1]};
    assign in7295_2 = {s7199[3],c7199,c7200,s7019[0]};
    CLA_4_c KS_7295(s7295, c7295, in7295_1, in7295_2, s7015[1]);
    wire[3:0] s7296, in7296_1, in7296_2;
    wire c7296;
    assign in7296_1 = {s7020[0],s7021[0],s7022[0],s7022[1]};
    assign in7296_2 = {s7201[3],c7201,c7202,s7023[0]};
    CLA_4_c KS_7296(s7296, c7296, in7296_1, in7296_2, s7019[1]);
    wire[3:0] s7297, in7297_1, in7297_2;
    wire c7297;
    assign in7297_1 = {s7024[0],s7025[0],s7026[0],s7026[1]};
    assign in7297_2 = {s7203[3],c7203,c7204,s7027[0]};
    CLA_4_c KS_7297(s7297, c7297, in7297_1, in7297_2, s7023[1]);
    wire[3:0] s7298, in7298_1, in7298_2;
    wire c7298;
    assign in7298_1 = {s7028[0],s7029[0],s7030[0],s7030[1]};
    assign in7298_2 = {s7205[3],c7205,c7206,s7031[0]};
    CLA_4_c KS_7298(s7298, c7298, in7298_1, in7298_2, s7027[1]);
    wire[3:0] s7299, in7299_1, in7299_2;
    wire c7299;
    assign in7299_1 = {s7032[0],s7033[0],s7034[0],s7034[1]};
    assign in7299_2 = {s7207[3],c7207,c7208,s7035[0]};
    CLA_4_c KS_7299(s7299, c7299, in7299_1, in7299_2, s7031[1]);
    wire[3:0] s7300, in7300_1, in7300_2;
    wire c7300;
    assign in7300_1 = {s7036[0],s7037[0],s7038[0],s7038[1]};
    assign in7300_2 = {s7209[3],c7209,c7210,s7039[0]};
    CLA_4_c KS_7300(s7300, c7300, in7300_1, in7300_2, s7035[1]);
    wire[3:0] s7301, in7301_1, in7301_2;
    wire c7301;
    assign in7301_1 = {s7040[0],s7041[0],s7042[0],s7042[1]};
    assign in7301_2 = {s7211[3],c7211,c7212,s7043[0]};
    CLA_4_c KS_7301(s7301, c7301, in7301_1, in7301_2, s7039[1]);
    wire[3:0] s7302, in7302_1, in7302_2;
    wire c7302;
    assign in7302_1 = {s7044[0],s7045[0],s7046[0],s7046[1]};
    assign in7302_2 = {s7213[3],c7213,c7214,s7047[0]};
    CLA_4_c KS_7302(s7302, c7302, in7302_1, in7302_2, s7043[1]);
    wire[3:0] s7303, in7303_1, in7303_2;
    wire c7303;
    assign in7303_1 = {s7048[0],s7049[0],s7050[0],s7050[1]};
    assign in7303_2 = {s7215[3],c7215,c7216,s7051[0]};
    CLA_4_c KS_7303(s7303, c7303, in7303_1, in7303_2, s7047[1]);
    wire[3:0] s7304, in7304_1, in7304_2;
    wire c7304;
    assign in7304_1 = {s7052[0],s7053[0],s7054[0],s7054[1]};
    assign in7304_2 = {s7217[3],c7217,c7218,s7055[0]};
    CLA_4_c KS_7304(s7304, c7304, in7304_1, in7304_2, s7051[1]);
    wire[3:0] s7305, in7305_1, in7305_2;
    wire c7305;
    assign in7305_1 = {s7056[0],s7057[0],s7058[0],s7058[1]};
    assign in7305_2 = {s7219[3],c7219,c7220,s7059[0]};
    CLA_4_c KS_7305(s7305, c7305, in7305_1, in7305_2, s7055[1]);
    wire[3:0] s7306, in7306_1, in7306_2;
    wire c7306;
    assign in7306_1 = {s7060[0],s7061[0],s7062[0],s7062[1]};
    assign in7306_2 = {s7221[3],c7221,c7222,s7063[0]};
    CLA_4_c KS_7306(s7306, c7306, in7306_1, in7306_2, s7059[1]);
    wire[3:0] s7307, in7307_1, in7307_2;
    wire c7307;
    assign in7307_1 = {s7064[0],s7065[0],s7066[0],s7066[1]};
    assign in7307_2 = {s7223[3],c7223,c7224,s7067[0]};
    CLA_4_c KS_7307(s7307, c7307, in7307_1, in7307_2, s7063[1]);
    wire[3:0] s7308, in7308_1, in7308_2;
    wire c7308;
    assign in7308_1 = {s7068[0],s7069[0],s7070[0],s7070[1]};
    assign in7308_2 = {s7225[3],c7225,c7226,s7071[0]};
    CLA_4_c KS_7308(s7308, c7308, in7308_1, in7308_2, s7067[1]);
    wire[3:0] s7309, in7309_1, in7309_2;
    wire c7309;
    assign in7309_1 = {s7072[0],s7073[0],s7074[0],s7074[1]};
    assign in7309_2 = {s7227[3],c7227,c7228,s7075[0]};
    CLA_4_c KS_7309(s7309, c7309, in7309_1, in7309_2, s7071[1]);
    wire[3:0] s7310, in7310_1, in7310_2;
    wire c7310;
    assign in7310_1 = {s7076[0],s7077[0],s7078[0],s7078[1]};
    assign in7310_2 = {s7229[3],c7229,c7230,s7079[0]};
    CLA_4_c KS_7310(s7310, c7310, in7310_1, in7310_2, s7075[1]);
    wire[3:0] s7311, in7311_1, in7311_2;
    wire c7311;
    assign in7311_1 = {s7080[0],s7081[0],s7082[0],s7082[1]};
    assign in7311_2 = {s7231[3],c7231,c7232,s7083[0]};
    CLA_4_c KS_7311(s7311, c7311, in7311_1, in7311_2, s7079[1]);
    wire[3:0] s7312, in7312_1, in7312_2;
    wire c7312;
    assign in7312_1 = {s7084[0],s7085[0],s7086[0],s7086[1]};
    assign in7312_2 = {s7233[3],c7233,c7234,s7087[0]};
    CLA_4_c KS_7312(s7312, c7312, in7312_1, in7312_2, s7083[1]);
    wire[3:0] s7313, in7313_1, in7313_2;
    wire c7313;
    assign in7313_1 = {s7088[0],s7089[0],s7090[0],s7090[1]};
    assign in7313_2 = {s7235[3],c7235,c7236,s7091[0]};
    CLA_4_c KS_7313(s7313, c7313, in7313_1, in7313_2, s7087[1]);
    wire[3:0] s7314, in7314_1, in7314_2;
    wire c7314;
    assign in7314_1 = {s7092[0],s7093[0],s7094[0],s7094[1]};
    assign in7314_2 = {s7237[3],c7237,c7238,s7095[0]};
    CLA_4_c KS_7314(s7314, c7314, in7314_1, in7314_2, s7091[1]);
    wire[3:0] s7315, in7315_1, in7315_2;
    wire c7315;
    assign in7315_1 = {s7096[0],s7097[0],s7098[0],s7098[1]};
    assign in7315_2 = {s7239[3],c7239,c7240,s7099[0]};
    CLA_4_c KS_7315(s7315, c7315, in7315_1, in7315_2, s7095[1]);
    wire[3:0] s7316, in7316_1, in7316_2;
    wire c7316;
    assign in7316_1 = {s7100[0],s7101[0],s7102[0],s7102[1]};
    assign in7316_2 = {s7241[3],c7241,c7242,s7103[0]};
    CLA_4_c KS_7316(s7316, c7316, in7316_1, in7316_2, s7099[1]);
    wire[3:0] s7317, in7317_1, in7317_2;
    wire c7317;
    assign in7317_1 = {s7104[0],s7105[0],s7106[0],s7106[1]};
    assign in7317_2 = {s7243[3],c7243,c7244,s7107[0]};
    CLA_4_c KS_7317(s7317, c7317, in7317_1, in7317_2, s7103[1]);
    wire[3:0] s7318, in7318_1, in7318_2;
    wire c7318;
    assign in7318_1 = {s7108[0],s7109[0],s7110[0],s7110[1]};
    assign in7318_2 = {s7245[3],c7245,c7246,s7111[0]};
    CLA_4_c KS_7318(s7318, c7318, in7318_1, in7318_2, s7107[1]);
    wire[3:0] s7319, in7319_1, in7319_2;
    wire c7319;
    assign in7319_1 = {s7112[0],s7113[0],s7114[0],s7114[1]};
    assign in7319_2 = {s7247[3],c7247,c7248,s7115[0]};
    CLA_4_c KS_7319(s7319, c7319, in7319_1, in7319_2, s7111[1]);
    wire[3:0] s7320, in7320_1, in7320_2;
    wire c7320;
    assign in7320_1 = {s7116[0],s7117[0],s7118[0],s7118[1]};
    assign in7320_2 = {s7249[3],c7249,c7250,s7119[0]};
    CLA_4_c KS_7320(s7320, c7320, in7320_1, in7320_2, s7115[1]);
    wire[3:0] s7321, in7321_1, in7321_2;
    wire c7321;
    assign in7321_1 = {s7120[0],s7121[0],s7122[0],s7122[1]};
    assign in7321_2 = {s7251[3],c7251,c7252,s7123[0]};
    CLA_4_c KS_7321(s7321, c7321, in7321_1, in7321_2, s7119[1]);
    wire[3:0] s7322, in7322_1, in7322_2;
    wire c7322;
    assign in7322_1 = {s7124[0],s7125[0],s7126[0],s7126[1]};
    assign in7322_2 = {s7253[3],c7253,c7254,s7127[0]};
    CLA_4_c KS_7322(s7322, c7322, in7322_1, in7322_2, s7123[1]);
    wire[3:0] s7323, in7323_1, in7323_2;
    wire c7323;
    assign in7323_1 = {s7128[0],s7129[0],s7130[0],s7130[1]};
    assign in7323_2 = {s7255[3],c7255,c7256,s7131[0]};
    CLA_4_c KS_7323(s7323, c7323, in7323_1, in7323_2, s7127[1]);
    wire[3:0] s7324, in7324_1, in7324_2;
    wire c7324;
    assign in7324_1 = {s7132[0],s7133[0],s7134[0],s7134[1]};
    assign in7324_2 = {s7257[3],c7257,c7258,s7135[0]};
    CLA_4_c KS_7324(s7324, c7324, in7324_1, in7324_2, s7131[1]);
    wire[3:0] s7325, in7325_1, in7325_2;
    wire c7325;
    assign in7325_1 = {s7136[0],s7137[0],s7138[0],s7138[1]};
    assign in7325_2 = {s7259[3],c7259,c7260,s7139[0]};
    CLA_4_c KS_7325(s7325, c7325, in7325_1, in7325_2, s7135[1]);
    wire[3:0] s7326, in7326_1, in7326_2;
    wire c7326;
    assign in7326_1 = {s7140[0],s7140[1],s7140[2],s7140[3]};
    assign in7326_2 = {s7261[3],c7261,c7262,s7263[2]};
    CLA_4_c KS_7326(s7326, c7326, in7326_1, in7326_2, s7139[1]);
    wire[2:0] s7327, in7327_1, in7327_2;
    wire c7327;
    assign in7327_1 = {c7140,pp127[125],pp126[127]};
    assign in7327_2 = {s7263[3],c7263,pp127[126]};
    CLA_3 KS_7327(s7327, c7327, in7327_1, in7327_2);

    /*Stage 9*/
    wire[3:0] s7328, in7328_1, in7328_2;
    wire c7328;
    assign in7328_1 = {pp0[2],pp2[1],pp4[0],s7141[1]};
    assign in7328_2 = {pp1[1],pp3[0],s7141[0],s7142[0]};
    CLA_4 KS_7328(s7328, c7328, in7328_1, in7328_2);
    wire[3:0] s7329, in7329_1, in7329_2;
    wire c7329;
    assign in7329_1 = {s7142[1],s7142[2],s7142[3],s7143[1]};
    assign in7329_2 = {s7265[3],c7265,s7143[0],s7144[0]};
    CLA_4_c KS_7329(s7329, c7329, in7329_1, in7329_2, s7141[2]);
    wire[3:0] s7330, in7330_1, in7330_2;
    wire c7330;
    assign in7330_1 = {s7144[1],s7144[2],s7144[3],s7145[1]};
    assign in7330_2 = {s7266[3],c7266,s7145[0],s7146[0]};
    CLA_4_c KS_7330(s7330, c7330, in7330_1, in7330_2, s7143[2]);
    wire[3:0] s7331, in7331_1, in7331_2;
    wire c7331;
    assign in7331_1 = {s7146[1],s7146[2],s7146[3],s7147[1]};
    assign in7331_2 = {s7267[3],c7267,s7147[0],s7148[0]};
    CLA_4_c KS_7331(s7331, c7331, in7331_1, in7331_2, s7145[2]);
    wire[3:0] s7332, in7332_1, in7332_2;
    wire c7332;
    assign in7332_1 = {s7148[1],s7148[2],s7148[3],s7149[1]};
    assign in7332_2 = {s7268[3],c7268,s7149[0],s7150[0]};
    CLA_4_c KS_7332(s7332, c7332, in7332_1, in7332_2, s7147[2]);
    wire[3:0] s7333, in7333_1, in7333_2;
    wire c7333;
    assign in7333_1 = {s7150[1],s7150[2],s7150[3],s7151[1]};
    assign in7333_2 = {s7269[3],c7269,s7151[0],s7152[0]};
    CLA_4_c KS_7333(s7333, c7333, in7333_1, in7333_2, s7149[2]);
    wire[3:0] s7334, in7334_1, in7334_2;
    wire c7334;
    assign in7334_1 = {s7152[1],s7152[2],s7152[3],s7153[1]};
    assign in7334_2 = {s7270[3],c7270,s7153[0],s7154[0]};
    CLA_4_c KS_7334(s7334, c7334, in7334_1, in7334_2, s7151[2]);
    wire[3:0] s7335, in7335_1, in7335_2;
    wire c7335;
    assign in7335_1 = {s7154[1],s7154[2],s7154[3],s7155[1]};
    assign in7335_2 = {s7271[3],c7271,s7155[0],s7156[0]};
    CLA_4_c KS_7335(s7335, c7335, in7335_1, in7335_2, s7153[2]);
    wire[3:0] s7336, in7336_1, in7336_2;
    wire c7336;
    assign in7336_1 = {s7156[1],s7156[2],s7156[3],s7157[1]};
    assign in7336_2 = {s7272[3],c7272,s7157[0],s7158[0]};
    CLA_4_c KS_7336(s7336, c7336, in7336_1, in7336_2, s7155[2]);
    wire[3:0] s7337, in7337_1, in7337_2;
    wire c7337;
    assign in7337_1 = {s7158[1],s7158[2],s7158[3],s7159[1]};
    assign in7337_2 = {s7273[3],c7273,s7159[0],s7160[0]};
    CLA_4_c KS_7337(s7337, c7337, in7337_1, in7337_2, s7157[2]);
    wire[3:0] s7338, in7338_1, in7338_2;
    wire c7338;
    assign in7338_1 = {s7160[1],s7160[2],s7160[3],s7161[1]};
    assign in7338_2 = {s7274[3],c7274,s7161[0],s7162[0]};
    CLA_4_c KS_7338(s7338, c7338, in7338_1, in7338_2, s7159[2]);
    wire[3:0] s7339, in7339_1, in7339_2;
    wire c7339;
    assign in7339_1 = {s7162[1],s7162[2],s7162[3],s7163[1]};
    assign in7339_2 = {s7275[3],c7275,s7163[0],s7164[0]};
    CLA_4_c KS_7339(s7339, c7339, in7339_1, in7339_2, s7161[2]);
    wire[3:0] s7340, in7340_1, in7340_2;
    wire c7340;
    assign in7340_1 = {s7164[1],s7164[2],s7164[3],s7165[1]};
    assign in7340_2 = {s7276[3],c7276,s7165[0],s7166[0]};
    CLA_4_c KS_7340(s7340, c7340, in7340_1, in7340_2, s7163[2]);
    wire[3:0] s7341, in7341_1, in7341_2;
    wire c7341;
    assign in7341_1 = {s7166[1],s7166[2],s7166[3],s7167[1]};
    assign in7341_2 = {s7277[3],c7277,s7167[0],s7168[0]};
    CLA_4_c KS_7341(s7341, c7341, in7341_1, in7341_2, s7165[2]);
    wire[3:0] s7342, in7342_1, in7342_2;
    wire c7342;
    assign in7342_1 = {s7168[1],s7168[2],s7168[3],s7169[1]};
    assign in7342_2 = {s7278[3],c7278,s7169[0],s7170[0]};
    CLA_4_c KS_7342(s7342, c7342, in7342_1, in7342_2, s7167[2]);
    wire[3:0] s7343, in7343_1, in7343_2;
    wire c7343;
    assign in7343_1 = {s7170[1],s7170[2],s7170[3],s7171[1]};
    assign in7343_2 = {s7279[3],c7279,s7171[0],s7172[0]};
    CLA_4_c KS_7343(s7343, c7343, in7343_1, in7343_2, s7169[2]);
    wire[3:0] s7344, in7344_1, in7344_2;
    wire c7344;
    assign in7344_1 = {s7172[1],s7172[2],s7172[3],s7173[1]};
    assign in7344_2 = {s7280[3],c7280,s7173[0],s7174[0]};
    CLA_4_c KS_7344(s7344, c7344, in7344_1, in7344_2, s7171[2]);
    wire[3:0] s7345, in7345_1, in7345_2;
    wire c7345;
    assign in7345_1 = {s7174[1],s7174[2],s7174[3],s7175[1]};
    assign in7345_2 = {s7281[3],c7281,s7175[0],s7176[0]};
    CLA_4_c KS_7345(s7345, c7345, in7345_1, in7345_2, s7173[2]);
    wire[3:0] s7346, in7346_1, in7346_2;
    wire c7346;
    assign in7346_1 = {s7176[1],s7176[2],s7176[3],s7177[1]};
    assign in7346_2 = {s7282[3],c7282,s7177[0],s7178[0]};
    CLA_4_c KS_7346(s7346, c7346, in7346_1, in7346_2, s7175[2]);
    wire[3:0] s7347, in7347_1, in7347_2;
    wire c7347;
    assign in7347_1 = {s7178[1],s7178[2],s7178[3],s7179[1]};
    assign in7347_2 = {s7283[3],c7283,s7179[0],s7180[0]};
    CLA_4_c KS_7347(s7347, c7347, in7347_1, in7347_2, s7177[2]);
    wire[3:0] s7348, in7348_1, in7348_2;
    wire c7348;
    assign in7348_1 = {s7180[1],s7180[2],s7180[3],s7181[1]};
    assign in7348_2 = {s7284[3],c7284,s7181[0],s7182[0]};
    CLA_4_c KS_7348(s7348, c7348, in7348_1, in7348_2, s7179[2]);
    wire[3:0] s7349, in7349_1, in7349_2;
    wire c7349;
    assign in7349_1 = {s7182[1],s7182[2],s7182[3],s7183[1]};
    assign in7349_2 = {s7285[3],c7285,s7183[0],s7184[0]};
    CLA_4_c KS_7349(s7349, c7349, in7349_1, in7349_2, s7181[2]);
    wire[3:0] s7350, in7350_1, in7350_2;
    wire c7350;
    assign in7350_1 = {s7184[1],s7184[2],s7184[3],s7185[1]};
    assign in7350_2 = {s7286[3],c7286,s7185[0],s7186[0]};
    CLA_4_c KS_7350(s7350, c7350, in7350_1, in7350_2, s7183[2]);
    wire[3:0] s7351, in7351_1, in7351_2;
    wire c7351;
    assign in7351_1 = {s7186[1],s7186[2],s7186[3],s7187[1]};
    assign in7351_2 = {s7287[3],c7287,s7187[0],s7188[0]};
    CLA_4_c KS_7351(s7351, c7351, in7351_1, in7351_2, s7185[2]);
    wire[3:0] s7352, in7352_1, in7352_2;
    wire c7352;
    assign in7352_1 = {s7188[1],s7188[2],s7188[3],s7189[1]};
    assign in7352_2 = {s7288[3],c7288,s7189[0],s7190[0]};
    CLA_4_c KS_7352(s7352, c7352, in7352_1, in7352_2, s7187[2]);
    wire[3:0] s7353, in7353_1, in7353_2;
    wire c7353;
    assign in7353_1 = {s7190[1],s7190[2],s7190[3],s7191[1]};
    assign in7353_2 = {s7289[3],c7289,s7191[0],s7192[0]};
    CLA_4_c KS_7353(s7353, c7353, in7353_1, in7353_2, s7189[2]);
    wire[3:0] s7354, in7354_1, in7354_2;
    wire c7354;
    assign in7354_1 = {s7192[1],s7192[2],s7192[3],s7193[1]};
    assign in7354_2 = {s7290[3],c7290,s7193[0],s7194[0]};
    CLA_4_c KS_7354(s7354, c7354, in7354_1, in7354_2, s7191[2]);
    wire[3:0] s7355, in7355_1, in7355_2;
    wire c7355;
    assign in7355_1 = {s7194[1],s7194[2],s7194[3],s7195[1]};
    assign in7355_2 = {s7291[3],c7291,s7195[0],s7196[0]};
    CLA_4_c KS_7355(s7355, c7355, in7355_1, in7355_2, s7193[2]);
    wire[3:0] s7356, in7356_1, in7356_2;
    wire c7356;
    assign in7356_1 = {s7196[1],s7196[2],s7196[3],s7197[1]};
    assign in7356_2 = {s7292[3],c7292,s7197[0],s7198[0]};
    CLA_4_c KS_7356(s7356, c7356, in7356_1, in7356_2, s7195[2]);
    wire[3:0] s7357, in7357_1, in7357_2;
    wire c7357;
    assign in7357_1 = {s7198[1],s7198[2],s7198[3],s7199[1]};
    assign in7357_2 = {s7293[3],c7293,s7199[0],s7200[0]};
    CLA_4_c KS_7357(s7357, c7357, in7357_1, in7357_2, s7197[2]);
    wire[3:0] s7358, in7358_1, in7358_2;
    wire c7358;
    assign in7358_1 = {s7200[1],s7200[2],s7200[3],s7201[1]};
    assign in7358_2 = {s7294[3],c7294,s7201[0],s7202[0]};
    CLA_4_c KS_7358(s7358, c7358, in7358_1, in7358_2, s7199[2]);
    wire[3:0] s7359, in7359_1, in7359_2;
    wire c7359;
    assign in7359_1 = {s7202[1],s7202[2],s7202[3],s7203[1]};
    assign in7359_2 = {s7295[3],c7295,s7203[0],s7204[0]};
    CLA_4_c KS_7359(s7359, c7359, in7359_1, in7359_2, s7201[2]);
    wire[3:0] s7360, in7360_1, in7360_2;
    wire c7360;
    assign in7360_1 = {s7204[1],s7204[2],s7204[3],s7205[1]};
    assign in7360_2 = {s7296[3],c7296,s7205[0],s7206[0]};
    CLA_4_c KS_7360(s7360, c7360, in7360_1, in7360_2, s7203[2]);
    wire[3:0] s7361, in7361_1, in7361_2;
    wire c7361;
    assign in7361_1 = {s7206[1],s7206[2],s7206[3],s7207[1]};
    assign in7361_2 = {s7297[3],c7297,s7207[0],s7208[0]};
    CLA_4_c KS_7361(s7361, c7361, in7361_1, in7361_2, s7205[2]);
    wire[3:0] s7362, in7362_1, in7362_2;
    wire c7362;
    assign in7362_1 = {s7208[1],s7208[2],s7208[3],s7209[1]};
    assign in7362_2 = {s7298[3],c7298,s7209[0],s7210[0]};
    CLA_4_c KS_7362(s7362, c7362, in7362_1, in7362_2, s7207[2]);
    wire[3:0] s7363, in7363_1, in7363_2;
    wire c7363;
    assign in7363_1 = {s7210[1],s7210[2],s7210[3],s7211[1]};
    assign in7363_2 = {s7299[3],c7299,s7211[0],s7212[0]};
    CLA_4_c KS_7363(s7363, c7363, in7363_1, in7363_2, s7209[2]);
    wire[3:0] s7364, in7364_1, in7364_2;
    wire c7364;
    assign in7364_1 = {s7212[1],s7212[2],s7212[3],s7213[1]};
    assign in7364_2 = {s7300[3],c7300,s7213[0],s7214[0]};
    CLA_4_c KS_7364(s7364, c7364, in7364_1, in7364_2, s7211[2]);
    wire[3:0] s7365, in7365_1, in7365_2;
    wire c7365;
    assign in7365_1 = {s7214[1],s7214[2],s7214[3],s7215[1]};
    assign in7365_2 = {s7301[3],c7301,s7215[0],s7216[0]};
    CLA_4_c KS_7365(s7365, c7365, in7365_1, in7365_2, s7213[2]);
    wire[3:0] s7366, in7366_1, in7366_2;
    wire c7366;
    assign in7366_1 = {s7216[1],s7216[2],s7216[3],s7217[1]};
    assign in7366_2 = {s7302[3],c7302,s7217[0],s7218[0]};
    CLA_4_c KS_7366(s7366, c7366, in7366_1, in7366_2, s7215[2]);
    wire[3:0] s7367, in7367_1, in7367_2;
    wire c7367;
    assign in7367_1 = {s7218[1],s7218[2],s7218[3],s7219[1]};
    assign in7367_2 = {s7303[3],c7303,s7219[0],s7220[0]};
    CLA_4_c KS_7367(s7367, c7367, in7367_1, in7367_2, s7217[2]);
    wire[3:0] s7368, in7368_1, in7368_2;
    wire c7368;
    assign in7368_1 = {s7220[1],s7220[2],s7220[3],s7221[1]};
    assign in7368_2 = {s7304[3],c7304,s7221[0],s7222[0]};
    CLA_4_c KS_7368(s7368, c7368, in7368_1, in7368_2, s7219[2]);
    wire[3:0] s7369, in7369_1, in7369_2;
    wire c7369;
    assign in7369_1 = {s7222[1],s7222[2],s7222[3],s7223[1]};
    assign in7369_2 = {s7305[3],c7305,s7223[0],s7224[0]};
    CLA_4_c KS_7369(s7369, c7369, in7369_1, in7369_2, s7221[2]);
    wire[3:0] s7370, in7370_1, in7370_2;
    wire c7370;
    assign in7370_1 = {s7224[1],s7224[2],s7224[3],s7225[1]};
    assign in7370_2 = {s7306[3],c7306,s7225[0],s7226[0]};
    CLA_4_c KS_7370(s7370, c7370, in7370_1, in7370_2, s7223[2]);
    wire[3:0] s7371, in7371_1, in7371_2;
    wire c7371;
    assign in7371_1 = {s7226[1],s7226[2],s7226[3],s7227[1]};
    assign in7371_2 = {s7307[3],c7307,s7227[0],s7228[0]};
    CLA_4_c KS_7371(s7371, c7371, in7371_1, in7371_2, s7225[2]);
    wire[3:0] s7372, in7372_1, in7372_2;
    wire c7372;
    assign in7372_1 = {s7228[1],s7228[2],s7228[3],s7229[1]};
    assign in7372_2 = {s7308[3],c7308,s7229[0],s7230[0]};
    CLA_4_c KS_7372(s7372, c7372, in7372_1, in7372_2, s7227[2]);
    wire[3:0] s7373, in7373_1, in7373_2;
    wire c7373;
    assign in7373_1 = {s7230[1],s7230[2],s7230[3],s7231[1]};
    assign in7373_2 = {s7309[3],c7309,s7231[0],s7232[0]};
    CLA_4_c KS_7373(s7373, c7373, in7373_1, in7373_2, s7229[2]);
    wire[3:0] s7374, in7374_1, in7374_2;
    wire c7374;
    assign in7374_1 = {s7232[1],s7232[2],s7232[3],s7233[1]};
    assign in7374_2 = {s7310[3],c7310,s7233[0],s7234[0]};
    CLA_4_c KS_7374(s7374, c7374, in7374_1, in7374_2, s7231[2]);
    wire[3:0] s7375, in7375_1, in7375_2;
    wire c7375;
    assign in7375_1 = {s7234[1],s7234[2],s7234[3],s7235[1]};
    assign in7375_2 = {s7311[3],c7311,s7235[0],s7236[0]};
    CLA_4_c KS_7375(s7375, c7375, in7375_1, in7375_2, s7233[2]);
    wire[3:0] s7376, in7376_1, in7376_2;
    wire c7376;
    assign in7376_1 = {s7236[1],s7236[2],s7236[3],s7237[1]};
    assign in7376_2 = {s7312[3],c7312,s7237[0],s7238[0]};
    CLA_4_c KS_7376(s7376, c7376, in7376_1, in7376_2, s7235[2]);
    wire[3:0] s7377, in7377_1, in7377_2;
    wire c7377;
    assign in7377_1 = {s7238[1],s7238[2],s7238[3],s7239[1]};
    assign in7377_2 = {s7313[3],c7313,s7239[0],s7240[0]};
    CLA_4_c KS_7377(s7377, c7377, in7377_1, in7377_2, s7237[2]);
    wire[3:0] s7378, in7378_1, in7378_2;
    wire c7378;
    assign in7378_1 = {s7240[1],s7240[2],s7240[3],s7241[1]};
    assign in7378_2 = {s7314[3],c7314,s7241[0],s7242[0]};
    CLA_4_c KS_7378(s7378, c7378, in7378_1, in7378_2, s7239[2]);
    wire[3:0] s7379, in7379_1, in7379_2;
    wire c7379;
    assign in7379_1 = {s7242[1],s7242[2],s7242[3],s7243[1]};
    assign in7379_2 = {s7315[3],c7315,s7243[0],s7244[0]};
    CLA_4_c KS_7379(s7379, c7379, in7379_1, in7379_2, s7241[2]);
    wire[3:0] s7380, in7380_1, in7380_2;
    wire c7380;
    assign in7380_1 = {s7244[1],s7244[2],s7244[3],s7245[1]};
    assign in7380_2 = {s7316[3],c7316,s7245[0],s7246[0]};
    CLA_4_c KS_7380(s7380, c7380, in7380_1, in7380_2, s7243[2]);
    wire[3:0] s7381, in7381_1, in7381_2;
    wire c7381;
    assign in7381_1 = {s7246[1],s7246[2],s7246[3],s7247[1]};
    assign in7381_2 = {s7317[3],c7317,s7247[0],s7248[0]};
    CLA_4_c KS_7381(s7381, c7381, in7381_1, in7381_2, s7245[2]);
    wire[3:0] s7382, in7382_1, in7382_2;
    wire c7382;
    assign in7382_1 = {s7248[1],s7248[2],s7248[3],s7249[1]};
    assign in7382_2 = {s7318[3],c7318,s7249[0],s7250[0]};
    CLA_4_c KS_7382(s7382, c7382, in7382_1, in7382_2, s7247[2]);
    wire[3:0] s7383, in7383_1, in7383_2;
    wire c7383;
    assign in7383_1 = {s7250[1],s7250[2],s7250[3],s7251[1]};
    assign in7383_2 = {s7319[3],c7319,s7251[0],s7252[0]};
    CLA_4_c KS_7383(s7383, c7383, in7383_1, in7383_2, s7249[2]);
    wire[3:0] s7384, in7384_1, in7384_2;
    wire c7384;
    assign in7384_1 = {s7252[1],s7252[2],s7252[3],s7253[1]};
    assign in7384_2 = {s7320[3],c7320,s7253[0],s7254[0]};
    CLA_4_c KS_7384(s7384, c7384, in7384_1, in7384_2, s7251[2]);
    wire[3:0] s7385, in7385_1, in7385_2;
    wire c7385;
    assign in7385_1 = {s7254[1],s7254[2],s7254[3],s7255[1]};
    assign in7385_2 = {s7321[3],c7321,s7255[0],s7256[0]};
    CLA_4_c KS_7385(s7385, c7385, in7385_1, in7385_2, s7253[2]);
    wire[3:0] s7386, in7386_1, in7386_2;
    wire c7386;
    assign in7386_1 = {s7256[1],s7256[2],s7256[3],s7257[1]};
    assign in7386_2 = {s7322[3],c7322,s7257[0],s7258[0]};
    CLA_4_c KS_7386(s7386, c7386, in7386_1, in7386_2, s7255[2]);
    wire[3:0] s7387, in7387_1, in7387_2;
    wire c7387;
    assign in7387_1 = {s7258[1],s7258[2],s7258[3],s7259[1]};
    assign in7387_2 = {s7323[3],c7323,s7259[0],s7260[0]};
    CLA_4_c KS_7387(s7387, c7387, in7387_1, in7387_2, s7257[2]);
    wire[3:0] s7388, in7388_1, in7388_2;
    wire c7388;
    assign in7388_1 = {s7260[1],s7260[2],s7260[3],s7261[1]};
    assign in7388_2 = {s7324[3],c7324,s7261[0],s7262[0]};
    CLA_4_c KS_7388(s7388, c7388, in7388_1, in7388_2, s7259[2]);
    wire[3:0] s7389, in7389_1, in7389_2;
    wire c7389;
    assign in7389_1 = {s7262[1],s7262[2],s7262[3],s7263[1]};
    assign in7389_2 = {s7325[3],c7325,s7263[0],s7264[0]};
    CLA_4_c KS_7389(s7389, c7389, in7389_1, in7389_2, s7261[2]);
    wire[3:0] s7390, in7390_1, in7390_2;
    wire c7390;
    assign in7390_1 = {s7264[1],s7264[2],s7264[3],c7264};
    assign in7390_2 = {s7326[3],c7326,s7327[1],s7327[2]};
    CLA_4 KS_7390(s7390, c7390, in7390_1, in7390_2);


    /*Final Stage 9*/
    wire[253:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],s7265[0],s7265[1],s7265[2],c7328,s7266[0],s7266[1],s7266[2],c7329,s7267[0],s7267[1],s7267[2],c7330,s7268[0],s7268[1],s7268[2],c7331,s7269[0],s7269[1],s7269[2],c7332,s7270[0],s7270[1],s7270[2],c7333,s7271[0],s7271[1],s7271[2],c7334,s7272[0],s7272[1],s7272[2],c7335,s7273[0],s7273[1],s7273[2],c7336,s7274[0],s7274[1],s7274[2],c7337,s7275[0],s7275[1],s7275[2],c7338,s7276[0],s7276[1],s7276[2],c7339,s7277[0],s7277[1],s7277[2],c7340,s7278[0],s7278[1],s7278[2],c7341,s7279[0],s7279[1],s7279[2],c7342,s7280[0],s7280[1],s7280[2],c7343,s7281[0],s7281[1],s7281[2],c7344,s7282[0],s7282[1],s7282[2],c7345,s7283[0],s7283[1],s7283[2],c7346,s7284[0],s7284[1],s7284[2],c7347,s7285[0],s7285[1],s7285[2],c7348,s7286[0],s7286[1],s7286[2],c7349,s7287[0],s7287[1],s7287[2],c7350,s7288[0],s7288[1],s7288[2],c7351,s7289[0],s7289[1],s7289[2],c7352,s7290[0],s7290[1],s7290[2],c7353,s7291[0],s7291[1],s7291[2],c7354,s7292[0],s7292[1],s7292[2],c7355,s7293[0],s7293[1],s7293[2],c7356,s7294[0],s7294[1],s7294[2],c7357,s7295[0],s7295[1],s7295[2],c7358,s7296[0],s7296[1],s7296[2],c7359,s7297[0],s7297[1],s7297[2],c7360,s7298[0],s7298[1],s7298[2],c7361,s7299[0],s7299[1],s7299[2],c7362,s7300[0],s7300[1],s7300[2],c7363,s7301[0],s7301[1],s7301[2],c7364,s7302[0],s7302[1],s7302[2],c7365,s7303[0],s7303[1],s7303[2],c7366,s7304[0],s7304[1],s7304[2],c7367,s7305[0],s7305[1],s7305[2],c7368,s7306[0],s7306[1],s7306[2],c7369,s7307[0],s7307[1],s7307[2],c7370,s7308[0],s7308[1],s7308[2],c7371,s7309[0],s7309[1],s7309[2],c7372,s7310[0],s7310[1],s7310[2],c7373,s7311[0],s7311[1],s7311[2],c7374,s7312[0],s7312[1],s7312[2],c7375,s7313[0],s7313[1],s7313[2],c7376,s7314[0],s7314[1],s7314[2],c7377,s7315[0],s7315[1],s7315[2],c7378,s7316[0],s7316[1],s7316[2],c7379,s7317[0],s7317[1],s7317[2],c7380,s7318[0],s7318[1],s7318[2],c7381,s7319[0],s7319[1],s7319[2],c7382,s7320[0],s7320[1],s7320[2],c7383,s7321[0],s7321[1],s7321[2],c7384,s7322[0],s7322[1],s7322[2],c7385,s7323[0],s7323[1],s7323[2],c7386,s7324[0],s7324[1],s7324[2],c7387,s7325[0],s7325[1],s7325[2],c7388,s7326[0],s7326[1],s7326[2],c7389,s7327[0],s7390[2],s7390[3],c7390};
    assign in_2 = {pp1[0],s7328[0],s7328[1],s7328[2],s7328[3],s7329[0],s7329[1],s7329[2],s7329[3],s7330[0],s7330[1],s7330[2],s7330[3],s7331[0],s7331[1],s7331[2],s7331[3],s7332[0],s7332[1],s7332[2],s7332[3],s7333[0],s7333[1],s7333[2],s7333[3],s7334[0],s7334[1],s7334[2],s7334[3],s7335[0],s7335[1],s7335[2],s7335[3],s7336[0],s7336[1],s7336[2],s7336[3],s7337[0],s7337[1],s7337[2],s7337[3],s7338[0],s7338[1],s7338[2],s7338[3],s7339[0],s7339[1],s7339[2],s7339[3],s7340[0],s7340[1],s7340[2],s7340[3],s7341[0],s7341[1],s7341[2],s7341[3],s7342[0],s7342[1],s7342[2],s7342[3],s7343[0],s7343[1],s7343[2],s7343[3],s7344[0],s7344[1],s7344[2],s7344[3],s7345[0],s7345[1],s7345[2],s7345[3],s7346[0],s7346[1],s7346[2],s7346[3],s7347[0],s7347[1],s7347[2],s7347[3],s7348[0],s7348[1],s7348[2],s7348[3],s7349[0],s7349[1],s7349[2],s7349[3],s7350[0],s7350[1],s7350[2],s7350[3],s7351[0],s7351[1],s7351[2],s7351[3],s7352[0],s7352[1],s7352[2],s7352[3],s7353[0],s7353[1],s7353[2],s7353[3],s7354[0],s7354[1],s7354[2],s7354[3],s7355[0],s7355[1],s7355[2],s7355[3],s7356[0],s7356[1],s7356[2],s7356[3],s7357[0],s7357[1],s7357[2],s7357[3],s7358[0],s7358[1],s7358[2],s7358[3],s7359[0],s7359[1],s7359[2],s7359[3],s7360[0],s7360[1],s7360[2],s7360[3],s7361[0],s7361[1],s7361[2],s7361[3],s7362[0],s7362[1],s7362[2],s7362[3],s7363[0],s7363[1],s7363[2],s7363[3],s7364[0],s7364[1],s7364[2],s7364[3],s7365[0],s7365[1],s7365[2],s7365[3],s7366[0],s7366[1],s7366[2],s7366[3],s7367[0],s7367[1],s7367[2],s7367[3],s7368[0],s7368[1],s7368[2],s7368[3],s7369[0],s7369[1],s7369[2],s7369[3],s7370[0],s7370[1],s7370[2],s7370[3],s7371[0],s7371[1],s7371[2],s7371[3],s7372[0],s7372[1],s7372[2],s7372[3],s7373[0],s7373[1],s7373[2],s7373[3],s7374[0],s7374[1],s7374[2],s7374[3],s7375[0],s7375[1],s7375[2],s7375[3],s7376[0],s7376[1],s7376[2],s7376[3],s7377[0],s7377[1],s7377[2],s7377[3],s7378[0],s7378[1],s7378[2],s7378[3],s7379[0],s7379[1],s7379[2],s7379[3],s7380[0],s7380[1],s7380[2],s7380[3],s7381[0],s7381[1],s7381[2],s7381[3],s7382[0],s7382[1],s7382[2],s7382[3],s7383[0],s7383[1],s7383[2],s7383[3],s7384[0],s7384[1],s7384[2],s7384[3],s7385[0],s7385[1],s7385[2],s7385[3],s7386[0],s7386[1],s7386[2],s7386[3],s7387[0],s7387[1],s7387[2],s7387[3],s7388[0],s7388[1],s7388[2],s7388[3],s7389[0],s7389[1],s7389[2],s7389[3],s7390[0],s7390[1],1'b0,1'b0,1'b0};
    CLA_254(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = s[126];
    assign product[128] = s[127];
    assign product[129] = s[128];
    assign product[130] = s[129];
    assign product[131] = s[130];
    assign product[132] = s[131];
    assign product[133] = s[132];
    assign product[134] = s[133];
    assign product[135] = s[134];
    assign product[136] = s[135];
    assign product[137] = s[136];
    assign product[138] = s[137];
    assign product[139] = s[138];
    assign product[140] = s[139];
    assign product[141] = s[140];
    assign product[142] = s[141];
    assign product[143] = s[142];
    assign product[144] = s[143];
    assign product[145] = s[144];
    assign product[146] = s[145];
    assign product[147] = s[146];
    assign product[148] = s[147];
    assign product[149] = s[148];
    assign product[150] = s[149];
    assign product[151] = s[150];
    assign product[152] = s[151];
    assign product[153] = s[152];
    assign product[154] = s[153];
    assign product[155] = s[154];
    assign product[156] = s[155];
    assign product[157] = s[156];
    assign product[158] = s[157];
    assign product[159] = s[158];
    assign product[160] = s[159];
    assign product[161] = s[160];
    assign product[162] = s[161];
    assign product[163] = s[162];
    assign product[164] = s[163];
    assign product[165] = s[164];
    assign product[166] = s[165];
    assign product[167] = s[166];
    assign product[168] = s[167];
    assign product[169] = s[168];
    assign product[170] = s[169];
    assign product[171] = s[170];
    assign product[172] = s[171];
    assign product[173] = s[172];
    assign product[174] = s[173];
    assign product[175] = s[174];
    assign product[176] = s[175];
    assign product[177] = s[176];
    assign product[178] = s[177];
    assign product[179] = s[178];
    assign product[180] = s[179];
    assign product[181] = s[180];
    assign product[182] = s[181];
    assign product[183] = s[182];
    assign product[184] = s[183];
    assign product[185] = s[184];
    assign product[186] = s[185];
    assign product[187] = s[186];
    assign product[188] = s[187];
    assign product[189] = s[188];
    assign product[190] = s[189];
    assign product[191] = s[190];
    assign product[192] = s[191];
    assign product[193] = s[192];
    assign product[194] = s[193];
    assign product[195] = s[194];
    assign product[196] = s[195];
    assign product[197] = s[196];
    assign product[198] = s[197];
    assign product[199] = s[198];
    assign product[200] = s[199];
    assign product[201] = s[200];
    assign product[202] = s[201];
    assign product[203] = s[202];
    assign product[204] = s[203];
    assign product[205] = s[204];
    assign product[206] = s[205];
    assign product[207] = s[206];
    assign product[208] = s[207];
    assign product[209] = s[208];
    assign product[210] = s[209];
    assign product[211] = s[210];
    assign product[212] = s[211];
    assign product[213] = s[212];
    assign product[214] = s[213];
    assign product[215] = s[214];
    assign product[216] = s[215];
    assign product[217] = s[216];
    assign product[218] = s[217];
    assign product[219] = s[218];
    assign product[220] = s[219];
    assign product[221] = s[220];
    assign product[222] = s[221];
    assign product[223] = s[222];
    assign product[224] = s[223];
    assign product[225] = s[224];
    assign product[226] = s[225];
    assign product[227] = s[226];
    assign product[228] = s[227];
    assign product[229] = s[228];
    assign product[230] = s[229];
    assign product[231] = s[230];
    assign product[232] = s[231];
    assign product[233] = s[232];
    assign product[234] = s[233];
    assign product[235] = s[234];
    assign product[236] = s[235];
    assign product[237] = s[236];
    assign product[238] = s[237];
    assign product[239] = s[238];
    assign product[240] = s[239];
    assign product[241] = s[240];
    assign product[242] = s[241];
    assign product[243] = s[242];
    assign product[244] = s[243];
    assign product[245] = s[244];
    assign product[246] = s[245];
    assign product[247] = s[246];
    assign product[248] = s[247];
    assign product[249] = s[248];
    assign product[250] = s[249];
    assign product[251] = s[250];
    assign product[252] = s[251];
    assign product[253] = s[252];
    assign product[254] = s[253];
    assign product[255] = c;
endmodule

module CLA_2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2);

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in1[1] & in2[1];
    assign P[0] = in1[1] ^ in2[1];
    assign G[1] = in1[0] & in2[0];
    assign P[1] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_2_c(output [1:0] sum,
            output cout,
            input [1:0] in1, in2,
            input cin);

    wire [1:0] G; /* Generate */
    wire [1:0] P; /* Propagate */
    wire [1:0] C; /* Carry */

    assign G[0] = in1[1] & in2[1]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[0] & in2[0];

    assign P[0] = in1[1] ^ in2[1];
    assign P[1] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule


module CLA_3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_3_c(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2, input cin);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = cin;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_4(output [3:0] sum,
            output cout,
            input [3:0] in1, in2);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = 0;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA_4_c(output [3:0] sum,
            output cout,
            input [3:0] in1, in2,
            input cin);

    wire [3:0] G; /* Generate */
    wire [3:0] P; /* Propagate */
    wire [3:0] C; /* Carry */

    assign G[0] = in1[3] & in2[3]; /*Generate    Gi = Ai * Bi */
    assign G[1] = in1[2] & in2[2];
    assign G[2] = in1[1] & in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[0] = in1[3] ^ in2[3]; /*Propagate   Pi = Ai + Bi */
    assign P[1] = in1[2] ^ in2[2];
    assign P[2] = in1[1] ^ in2[1];
    assign P[3] = in1[0] ^ in2[0];

    assign C[0] = cin;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module Half_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2);
    xor(sum, in1, in2);
    and(cout, in1, in2);
endmodule

module Full_Adder(output wire sum,
                  output wire cout,
                  input wire in1,
                  input wire in2,
                  input wire cin);
    wire temp1;
    wire temp2;
    wire temp3;
    xor(sum, in1, in2, cin);
    and(temp1,in1,in2);
    and(temp2,in1,cin);
    and(temp3,in2,cin);
    or(cout,temp1,temp2,temp3);
endmodule

