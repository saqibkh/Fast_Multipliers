module multiplier_128bits_version11(product, A, B);

    output [255:0] product;
    input [127:0] A, B;

    wire [127:0] pp0;
    wire [127:0] pp1;
    wire [127:0] pp2;
    wire [127:0] pp3;
    wire [127:0] pp4;
    wire [127:0] pp5;
    wire [127:0] pp6;
    wire [127:0] pp7;
    wire [127:0] pp8;
    wire [127:0] pp9;
    wire [127:0] pp10;
    wire [127:0] pp11;
    wire [127:0] pp12;
    wire [127:0] pp13;
    wire [127:0] pp14;
    wire [127:0] pp15;
    wire [127:0] pp16;
    wire [127:0] pp17;
    wire [127:0] pp18;
    wire [127:0] pp19;
    wire [127:0] pp20;
    wire [127:0] pp21;
    wire [127:0] pp22;
    wire [127:0] pp23;
    wire [127:0] pp24;
    wire [127:0] pp25;
    wire [127:0] pp26;
    wire [127:0] pp27;
    wire [127:0] pp28;
    wire [127:0] pp29;
    wire [127:0] pp30;
    wire [127:0] pp31;
    wire [127:0] pp32;
    wire [127:0] pp33;
    wire [127:0] pp34;
    wire [127:0] pp35;
    wire [127:0] pp36;
    wire [127:0] pp37;
    wire [127:0] pp38;
    wire [127:0] pp39;
    wire [127:0] pp40;
    wire [127:0] pp41;
    wire [127:0] pp42;
    wire [127:0] pp43;
    wire [127:0] pp44;
    wire [127:0] pp45;
    wire [127:0] pp46;
    wire [127:0] pp47;
    wire [127:0] pp48;
    wire [127:0] pp49;
    wire [127:0] pp50;
    wire [127:0] pp51;
    wire [127:0] pp52;
    wire [127:0] pp53;
    wire [127:0] pp54;
    wire [127:0] pp55;
    wire [127:0] pp56;
    wire [127:0] pp57;
    wire [127:0] pp58;
    wire [127:0] pp59;
    wire [127:0] pp60;
    wire [127:0] pp61;
    wire [127:0] pp62;
    wire [127:0] pp63;
    wire [127:0] pp64;
    wire [127:0] pp65;
    wire [127:0] pp66;
    wire [127:0] pp67;
    wire [127:0] pp68;
    wire [127:0] pp69;
    wire [127:0] pp70;
    wire [127:0] pp71;
    wire [127:0] pp72;
    wire [127:0] pp73;
    wire [127:0] pp74;
    wire [127:0] pp75;
    wire [127:0] pp76;
    wire [127:0] pp77;
    wire [127:0] pp78;
    wire [127:0] pp79;
    wire [127:0] pp80;
    wire [127:0] pp81;
    wire [127:0] pp82;
    wire [127:0] pp83;
    wire [127:0] pp84;
    wire [127:0] pp85;
    wire [127:0] pp86;
    wire [127:0] pp87;
    wire [127:0] pp88;
    wire [127:0] pp89;
    wire [127:0] pp90;
    wire [127:0] pp91;
    wire [127:0] pp92;
    wire [127:0] pp93;
    wire [127:0] pp94;
    wire [127:0] pp95;
    wire [127:0] pp96;
    wire [127:0] pp97;
    wire [127:0] pp98;
    wire [127:0] pp99;
    wire [127:0] pp100;
    wire [127:0] pp101;
    wire [127:0] pp102;
    wire [127:0] pp103;
    wire [127:0] pp104;
    wire [127:0] pp105;
    wire [127:0] pp106;
    wire [127:0] pp107;
    wire [127:0] pp108;
    wire [127:0] pp109;
    wire [127:0] pp110;
    wire [127:0] pp111;
    wire [127:0] pp112;
    wire [127:0] pp113;
    wire [127:0] pp114;
    wire [127:0] pp115;
    wire [127:0] pp116;
    wire [127:0] pp117;
    wire [127:0] pp118;
    wire [127:0] pp119;
    wire [127:0] pp120;
    wire [127:0] pp121;
    wire [127:0] pp122;
    wire [127:0] pp123;
    wire [127:0] pp124;
    wire [127:0] pp125;
    wire [127:0] pp126;
    wire [127:0] pp127;


    assign pp0 = A[0] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp64 = A[64] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp65 = A[65] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp66 = A[66] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp67 = A[67] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp68 = A[68] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp69 = A[69] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp70 = A[70] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp71 = A[71] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp72 = A[72] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp73 = A[73] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp74 = A[74] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp75 = A[75] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp76 = A[76] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp77 = A[77] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp78 = A[78] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp79 = A[79] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp80 = A[80] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp81 = A[81] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp82 = A[82] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp83 = A[83] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp84 = A[84] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp85 = A[85] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp86 = A[86] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp87 = A[87] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp88 = A[88] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp89 = A[89] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp90 = A[90] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp91 = A[91] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp92 = A[92] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp93 = A[93] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp94 = A[94] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp95 = A[95] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp96 = A[96] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp97 = A[97] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp98 = A[98] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp99 = A[99] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp100 = A[100] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp101 = A[101] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp102 = A[102] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp103 = A[103] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp104 = A[104] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp105 = A[105] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp106 = A[106] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp107 = A[107] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp108 = A[108] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp109 = A[109] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp110 = A[110] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp111 = A[111] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp112 = A[112] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp113 = A[113] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp114 = A[114] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp115 = A[115] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp116 = A[116] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp117 = A[117] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp118 = A[118] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp119 = A[119] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp120 = A[120] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp121 = A[121] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp122 = A[122] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp123 = A[123] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp124 = A[124] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp125 = A[125] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp126 = A[126] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    assign pp127 = A[127] ? B: 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[127:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp10[54],pp10[55],pp10[56],pp10[57],pp10[58],pp10[59],pp10[60],pp10[61],pp10[62],pp10[63],pp10[64],pp10[65],pp10[66],pp10[67],pp10[68],pp10[69],pp10[70],pp10[71],pp10[72],pp10[73],pp10[74],pp10[75],pp10[76],pp10[77],pp10[78],pp10[79],pp10[80],pp10[81],pp10[82],pp10[83],pp10[84],pp10[85],pp10[86],pp10[87],pp10[88],pp10[89],pp0[100],pp0[101],pp0[102],pp0[103],pp0[104],pp0[105],pp0[106],pp0[107],pp0[108],pp0[109],pp10[100],pp10[101],pp10[102],pp10[103],pp10[104],pp10[105],pp10[106],pp10[107],pp10[108],pp10[109],pp10[110],pp10[111],pp10[112],pp10[113],pp10[114],pp10[115],pp10[116],pp10[117],pp10[118],pp10[119],pp10[120],pp10[121],pp10[122],pp10[123],pp10[124],pp10[125],pp10[126],pp10[127],pp11[127],pp12[127],pp13[127],pp14[127],pp15[127],pp16[127],pp17[127],pp18[127],pp19[127],pp20[127],pp21[127],pp22[127],pp23[127],pp24[127],pp25[127],pp26[127],pp27[127],pp28[127],pp29[127],pp30[127],pp31[127],pp32[127],pp33[127],pp34[127],pp35[127],pp36[127],pp37[127],pp38[127],pp39[127],pp40[127],pp41[127],pp42[127],pp43[127],pp44[127],pp45[127],pp46[127],pp47[127],pp48[127],pp49[127],pp50[127],pp51[127],pp52[127],pp53[127],pp54[127],pp55[127],pp56[127],pp57[127],pp58[127],pp59[127],pp60[127],pp61[127],pp62[127],pp63[127],pp64[127]};
    assign in1_2 = {pp11[53],pp11[54],pp11[55],pp11[56],pp11[57],pp11[58],pp11[59],pp11[60],pp11[61],pp11[62],pp11[63],pp11[64],pp11[65],pp11[66],pp11[67],pp11[68],pp11[69],pp11[70],pp11[71],pp11[72],pp11[73],pp11[74],pp11[75],pp11[76],pp11[77],pp11[78],pp11[79],pp11[80],pp11[81],pp11[82],pp11[83],pp11[84],pp11[85],pp11[86],pp11[87],pp11[88],pp10[90],pp1[100],pp1[101],pp1[102],pp1[103],pp1[104],pp1[105],pp1[106],pp1[107],pp1[108],pp100[10],pp11[100],pp11[101],pp11[102],pp11[103],pp11[104],pp11[105],pp11[106],pp11[107],pp11[108],pp11[109],pp11[110],pp11[111],pp11[112],pp11[113],pp11[114],pp11[115],pp11[116],pp11[117],pp11[118],pp11[119],pp11[120],pp11[121],pp11[122],pp11[123],pp11[124],pp11[125],pp11[126],pp12[126],pp13[126],pp14[126],pp15[126],pp16[126],pp17[126],pp18[126],pp19[126],pp20[126],pp21[126],pp22[126],pp23[126],pp24[126],pp25[126],pp26[126],pp27[126],pp28[126],pp29[126],pp30[126],pp31[126],pp32[126],pp33[126],pp34[126],pp35[126],pp36[126],pp37[126],pp38[126],pp39[126],pp40[126],pp41[126],pp42[126],pp43[126],pp44[126],pp45[126],pp46[126],pp47[126],pp48[126],pp49[126],pp50[126],pp51[126],pp52[126],pp53[126],pp54[126],pp55[126],pp56[126],pp57[126],pp58[126],pp59[126],pp60[126],pp61[126],pp62[126],pp63[126],pp64[126],pp65[126]};
    CLA_128 KS_1(s1, c1, in1_1, in1_2);
    wire[125:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp12[53],pp12[54],pp12[55],pp12[56],pp12[57],pp12[58],pp12[59],pp12[60],pp12[61],pp12[62],pp12[63],pp12[64],pp12[65],pp12[66],pp12[67],pp12[68],pp12[69],pp12[70],pp12[71],pp12[72],pp12[73],pp12[74],pp12[75],pp12[76],pp12[77],pp12[78],pp12[79],pp12[80],pp12[81],pp12[82],pp12[83],pp12[84],pp12[85],pp12[86],pp12[87],pp11[89],pp10[91],pp2[100],pp2[101],pp2[102],pp2[103],pp2[104],pp2[105],pp2[106],pp2[107],pp0[110],pp100[11],pp12[100],pp12[101],pp12[102],pp12[103],pp12[104],pp12[105],pp12[106],pp12[107],pp12[108],pp12[109],pp12[110],pp12[111],pp12[112],pp12[113],pp12[114],pp12[115],pp12[116],pp12[117],pp12[118],pp12[119],pp12[120],pp12[121],pp12[122],pp12[123],pp12[124],pp12[125],pp13[125],pp14[125],pp15[125],pp16[125],pp17[125],pp18[125],pp19[125],pp20[125],pp21[125],pp22[125],pp23[125],pp24[125],pp25[125],pp26[125],pp27[125],pp28[125],pp29[125],pp30[125],pp31[125],pp32[125],pp33[125],pp34[125],pp35[125],pp36[125],pp37[125],pp38[125],pp39[125],pp40[125],pp41[125],pp42[125],pp43[125],pp44[125],pp45[125],pp46[125],pp47[125],pp48[125],pp49[125],pp50[125],pp51[125],pp52[125],pp53[125],pp54[125],pp55[125],pp56[125],pp57[125],pp58[125],pp59[125],pp60[125],pp61[125],pp62[125],pp63[125],pp64[125],pp65[125]};
    assign in2_2 = {pp13[52],pp13[53],pp13[54],pp13[55],pp13[56],pp13[57],pp13[58],pp13[59],pp13[60],pp13[61],pp13[62],pp13[63],pp13[64],pp13[65],pp13[66],pp13[67],pp13[68],pp13[69],pp13[70],pp13[71],pp13[72],pp13[73],pp13[74],pp13[75],pp13[76],pp13[77],pp13[78],pp13[79],pp13[80],pp13[81],pp13[82],pp13[83],pp13[84],pp13[85],pp13[86],pp12[88],pp11[90],pp10[92],pp3[100],pp3[101],pp3[102],pp3[103],pp3[104],pp3[105],pp3[106],pp1[109],pp101[10],pp100[12],pp13[100],pp13[101],pp13[102],pp13[103],pp13[104],pp13[105],pp13[106],pp13[107],pp13[108],pp13[109],pp13[110],pp13[111],pp13[112],pp13[113],pp13[114],pp13[115],pp13[116],pp13[117],pp13[118],pp13[119],pp13[120],pp13[121],pp13[122],pp13[123],pp13[124],pp14[124],pp15[124],pp16[124],pp17[124],pp18[124],pp19[124],pp20[124],pp21[124],pp22[124],pp23[124],pp24[124],pp25[124],pp26[124],pp27[124],pp28[124],pp29[124],pp30[124],pp31[124],pp32[124],pp33[124],pp34[124],pp35[124],pp36[124],pp37[124],pp38[124],pp39[124],pp40[124],pp41[124],pp42[124],pp43[124],pp44[124],pp45[124],pp46[124],pp47[124],pp48[124],pp49[124],pp50[124],pp51[124],pp52[124],pp53[124],pp54[124],pp55[124],pp56[124],pp57[124],pp58[124],pp59[124],pp60[124],pp61[124],pp62[124],pp63[124],pp64[124],pp65[124],pp66[124]};
    CLA_126 KS_2(s2, c2, in2_1, in2_2);
    wire[123:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp14[52],pp14[53],pp14[54],pp14[55],pp14[56],pp14[57],pp14[58],pp14[59],pp14[60],pp14[61],pp14[62],pp14[63],pp14[64],pp14[65],pp14[66],pp14[67],pp14[68],pp14[69],pp14[70],pp14[71],pp14[72],pp14[73],pp14[74],pp14[75],pp14[76],pp14[77],pp14[78],pp14[79],pp14[80],pp14[81],pp14[82],pp14[83],pp14[84],pp14[85],pp13[87],pp12[89],pp11[91],pp10[93],pp4[100],pp4[101],pp4[102],pp4[103],pp4[104],pp4[105],pp2[108],pp0[111],pp101[11],pp100[13],pp14[100],pp14[101],pp14[102],pp14[103],pp14[104],pp14[105],pp14[106],pp14[107],pp14[108],pp14[109],pp14[110],pp14[111],pp14[112],pp14[113],pp14[114],pp14[115],pp14[116],pp14[117],pp14[118],pp14[119],pp14[120],pp14[121],pp14[122],pp14[123],pp15[123],pp16[123],pp17[123],pp18[123],pp19[123],pp20[123],pp21[123],pp22[123],pp23[123],pp24[123],pp25[123],pp26[123],pp27[123],pp28[123],pp29[123],pp30[123],pp31[123],pp32[123],pp33[123],pp34[123],pp35[123],pp36[123],pp37[123],pp38[123],pp39[123],pp40[123],pp41[123],pp42[123],pp43[123],pp44[123],pp45[123],pp46[123],pp47[123],pp48[123],pp49[123],pp50[123],pp51[123],pp52[123],pp53[123],pp54[123],pp55[123],pp56[123],pp57[123],pp58[123],pp59[123],pp60[123],pp61[123],pp62[123],pp63[123],pp64[123],pp65[123],pp66[123]};
    assign in3_2 = {pp15[51],pp15[52],pp15[53],pp15[54],pp15[55],pp15[56],pp15[57],pp15[58],pp15[59],pp15[60],pp15[61],pp15[62],pp15[63],pp15[64],pp15[65],pp15[66],pp15[67],pp15[68],pp15[69],pp15[70],pp15[71],pp15[72],pp15[73],pp15[74],pp15[75],pp15[76],pp15[77],pp15[78],pp15[79],pp15[80],pp15[81],pp15[82],pp15[83],pp15[84],pp14[86],pp13[88],pp12[90],pp11[92],pp10[94],pp5[100],pp5[101],pp5[102],pp5[103],pp5[104],pp3[107],pp1[110],pp102[10],pp101[12],pp100[14],pp15[100],pp15[101],pp15[102],pp15[103],pp15[104],pp15[105],pp15[106],pp15[107],pp15[108],pp15[109],pp15[110],pp15[111],pp15[112],pp15[113],pp15[114],pp15[115],pp15[116],pp15[117],pp15[118],pp15[119],pp15[120],pp15[121],pp15[122],pp16[122],pp17[122],pp18[122],pp19[122],pp20[122],pp21[122],pp22[122],pp23[122],pp24[122],pp25[122],pp26[122],pp27[122],pp28[122],pp29[122],pp30[122],pp31[122],pp32[122],pp33[122],pp34[122],pp35[122],pp36[122],pp37[122],pp38[122],pp39[122],pp40[122],pp41[122],pp42[122],pp43[122],pp44[122],pp45[122],pp46[122],pp47[122],pp48[122],pp49[122],pp50[122],pp51[122],pp52[122],pp53[122],pp54[122],pp55[122],pp56[122],pp57[122],pp58[122],pp59[122],pp60[122],pp61[122],pp62[122],pp63[122],pp64[122],pp65[122],pp66[122],pp67[122]};
    CLA_124 KS_3(s3, c3, in3_1, in3_2);
    wire[121:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp16[51],pp16[52],pp16[53],pp16[54],pp16[55],pp16[56],pp16[57],pp16[58],pp16[59],pp16[60],pp16[61],pp16[62],pp16[63],pp16[64],pp16[65],pp16[66],pp16[67],pp16[68],pp16[69],pp16[70],pp16[71],pp16[72],pp16[73],pp16[74],pp16[75],pp16[76],pp16[77],pp16[78],pp16[79],pp16[80],pp16[81],pp16[82],pp16[83],pp15[85],pp14[87],pp13[89],pp12[91],pp11[93],pp10[95],pp6[100],pp6[101],pp6[102],pp6[103],pp4[106],pp2[109],pp0[112],pp102[11],pp101[13],pp100[15],pp16[100],pp16[101],pp16[102],pp16[103],pp16[104],pp16[105],pp16[106],pp16[107],pp16[108],pp16[109],pp16[110],pp16[111],pp16[112],pp16[113],pp16[114],pp16[115],pp16[116],pp16[117],pp16[118],pp16[119],pp16[120],pp16[121],pp17[121],pp18[121],pp19[121],pp20[121],pp21[121],pp22[121],pp23[121],pp24[121],pp25[121],pp26[121],pp27[121],pp28[121],pp29[121],pp30[121],pp31[121],pp32[121],pp33[121],pp34[121],pp35[121],pp36[121],pp37[121],pp38[121],pp39[121],pp40[121],pp41[121],pp42[121],pp43[121],pp44[121],pp45[121],pp46[121],pp47[121],pp48[121],pp49[121],pp50[121],pp51[121],pp52[121],pp53[121],pp54[121],pp55[121],pp56[121],pp57[121],pp58[121],pp59[121],pp60[121],pp61[121],pp62[121],pp63[121],pp64[121],pp65[121],pp66[121],pp67[121]};
    assign in4_2 = {pp17[50],pp17[51],pp17[52],pp17[53],pp17[54],pp17[55],pp17[56],pp17[57],pp17[58],pp17[59],pp17[60],pp17[61],pp17[62],pp17[63],pp17[64],pp17[65],pp17[66],pp17[67],pp17[68],pp17[69],pp17[70],pp17[71],pp17[72],pp17[73],pp17[74],pp17[75],pp17[76],pp17[77],pp17[78],pp17[79],pp17[80],pp17[81],pp17[82],pp16[84],pp15[86],pp14[88],pp13[90],pp12[92],pp11[94],pp10[96],pp7[100],pp7[101],pp7[102],pp5[105],pp3[108],pp1[111],pp103[10],pp102[12],pp101[14],pp100[16],pp17[100],pp17[101],pp17[102],pp17[103],pp17[104],pp17[105],pp17[106],pp17[107],pp17[108],pp17[109],pp17[110],pp17[111],pp17[112],pp17[113],pp17[114],pp17[115],pp17[116],pp17[117],pp17[118],pp17[119],pp17[120],pp18[120],pp19[120],pp20[120],pp21[120],pp22[120],pp23[120],pp24[120],pp25[120],pp26[120],pp27[120],pp28[120],pp29[120],pp30[120],pp31[120],pp32[120],pp33[120],pp34[120],pp35[120],pp36[120],pp37[120],pp38[120],pp39[120],pp40[120],pp41[120],pp42[120],pp43[120],pp44[120],pp45[120],pp46[120],pp47[120],pp48[120],pp49[120],pp50[120],pp51[120],pp52[120],pp53[120],pp54[120],pp55[120],pp56[120],pp57[120],pp58[120],pp59[120],pp60[120],pp61[120],pp62[120],pp63[120],pp64[120],pp65[120],pp66[120],pp67[120],pp68[120]};
    CLA_122 KS_4(s4, c4, in4_1, in4_2);
    wire[119:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp18[50],pp18[51],pp18[52],pp18[53],pp18[54],pp18[55],pp18[56],pp18[57],pp18[58],pp18[59],pp18[60],pp18[61],pp18[62],pp18[63],pp18[64],pp18[65],pp18[66],pp18[67],pp18[68],pp18[69],pp18[70],pp18[71],pp18[72],pp18[73],pp18[74],pp18[75],pp18[76],pp18[77],pp18[78],pp18[79],pp18[80],pp18[81],pp17[83],pp16[85],pp15[87],pp14[89],pp13[91],pp12[93],pp11[95],pp10[97],pp8[100],pp8[101],pp6[104],pp4[107],pp2[110],pp0[113],pp103[11],pp102[13],pp101[15],pp100[17],pp18[100],pp18[101],pp18[102],pp18[103],pp18[104],pp18[105],pp18[106],pp18[107],pp18[108],pp18[109],pp18[110],pp18[111],pp18[112],pp18[113],pp18[114],pp18[115],pp18[116],pp18[117],pp18[118],pp18[119],pp19[119],pp20[119],pp21[119],pp22[119],pp23[119],pp24[119],pp25[119],pp26[119],pp27[119],pp28[119],pp29[119],pp30[119],pp31[119],pp32[119],pp33[119],pp34[119],pp35[119],pp36[119],pp37[119],pp38[119],pp39[119],pp40[119],pp41[119],pp42[119],pp43[119],pp44[119],pp45[119],pp46[119],pp47[119],pp48[119],pp49[119],pp50[119],pp51[119],pp52[119],pp53[119],pp54[119],pp55[119],pp56[119],pp57[119],pp58[119],pp59[119],pp60[119],pp61[119],pp62[119],pp63[119],pp64[119],pp65[119],pp66[119],pp67[119],pp68[119]};
    assign in5_2 = {pp19[49],pp19[50],pp19[51],pp19[52],pp19[53],pp19[54],pp19[55],pp19[56],pp19[57],pp19[58],pp19[59],pp19[60],pp19[61],pp19[62],pp19[63],pp19[64],pp19[65],pp19[66],pp19[67],pp19[68],pp19[69],pp19[70],pp19[71],pp19[72],pp19[73],pp19[74],pp19[75],pp19[76],pp19[77],pp19[78],pp19[79],pp19[80],pp18[82],pp17[84],pp16[86],pp15[88],pp14[90],pp13[92],pp12[94],pp11[96],pp10[98],pp9[100],pp7[103],pp5[106],pp3[109],pp1[112],pp104[10],pp103[12],pp102[14],pp101[16],pp100[18],pp19[100],pp19[101],pp19[102],pp19[103],pp19[104],pp19[105],pp19[106],pp19[107],pp19[108],pp19[109],pp19[110],pp19[111],pp19[112],pp19[113],pp19[114],pp19[115],pp19[116],pp19[117],pp19[118],pp20[118],pp21[118],pp22[118],pp23[118],pp24[118],pp25[118],pp26[118],pp27[118],pp28[118],pp29[118],pp30[118],pp31[118],pp32[118],pp33[118],pp34[118],pp35[118],pp36[118],pp37[118],pp38[118],pp39[118],pp40[118],pp41[118],pp42[118],pp43[118],pp44[118],pp45[118],pp46[118],pp47[118],pp48[118],pp49[118],pp50[118],pp51[118],pp52[118],pp53[118],pp54[118],pp55[118],pp56[118],pp57[118],pp58[118],pp59[118],pp60[118],pp61[118],pp62[118],pp63[118],pp64[118],pp65[118],pp66[118],pp67[118],pp68[118],pp69[118]};
    CLA_120 KS_5(s5, c5, in5_1, in5_2);
    wire[117:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp20[49],pp20[50],pp20[51],pp20[52],pp20[53],pp20[54],pp20[55],pp20[56],pp20[57],pp20[58],pp20[59],pp20[60],pp20[61],pp20[62],pp20[63],pp20[64],pp20[65],pp20[66],pp20[67],pp20[68],pp20[69],pp20[70],pp20[71],pp20[72],pp20[73],pp20[74],pp20[75],pp20[76],pp20[77],pp20[78],pp20[79],pp19[81],pp18[83],pp17[85],pp16[87],pp15[89],pp14[91],pp13[93],pp12[95],pp11[97],pp10[99],pp8[102],pp6[105],pp4[108],pp2[111],pp0[114],pp104[11],pp103[13],pp102[15],pp101[17],pp100[19],pp20[100],pp20[101],pp20[102],pp20[103],pp20[104],pp20[105],pp20[106],pp20[107],pp20[108],pp20[109],pp20[110],pp20[111],pp20[112],pp20[113],pp20[114],pp20[115],pp20[116],pp20[117],pp21[117],pp22[117],pp23[117],pp24[117],pp25[117],pp26[117],pp27[117],pp28[117],pp29[117],pp30[117],pp31[117],pp32[117],pp33[117],pp34[117],pp35[117],pp36[117],pp37[117],pp38[117],pp39[117],pp40[117],pp41[117],pp42[117],pp43[117],pp44[117],pp45[117],pp46[117],pp47[117],pp48[117],pp49[117],pp50[117],pp51[117],pp52[117],pp53[117],pp54[117],pp55[117],pp56[117],pp57[117],pp58[117],pp59[117],pp60[117],pp61[117],pp62[117],pp63[117],pp64[117],pp65[117],pp66[117],pp67[117],pp68[117],pp69[117]};
    assign in6_2 = {pp21[48],pp21[49],pp21[50],pp21[51],pp21[52],pp21[53],pp21[54],pp21[55],pp21[56],pp21[57],pp21[58],pp21[59],pp21[60],pp21[61],pp21[62],pp21[63],pp21[64],pp21[65],pp21[66],pp21[67],pp21[68],pp21[69],pp21[70],pp21[71],pp21[72],pp21[73],pp21[74],pp21[75],pp21[76],pp21[77],pp21[78],pp20[80],pp19[82],pp18[84],pp17[86],pp16[88],pp15[90],pp14[92],pp13[94],pp12[96],pp11[98],pp9[101],pp7[104],pp5[107],pp3[110],pp1[113],pp105[10],pp104[12],pp103[14],pp102[16],pp101[18],pp100[20],pp21[100],pp21[101],pp21[102],pp21[103],pp21[104],pp21[105],pp21[106],pp21[107],pp21[108],pp21[109],pp21[110],pp21[111],pp21[112],pp21[113],pp21[114],pp21[115],pp21[116],pp22[116],pp23[116],pp24[116],pp25[116],pp26[116],pp27[116],pp28[116],pp29[116],pp30[116],pp31[116],pp32[116],pp33[116],pp34[116],pp35[116],pp36[116],pp37[116],pp38[116],pp39[116],pp40[116],pp41[116],pp42[116],pp43[116],pp44[116],pp45[116],pp46[116],pp47[116],pp48[116],pp49[116],pp50[116],pp51[116],pp52[116],pp53[116],pp54[116],pp55[116],pp56[116],pp57[116],pp58[116],pp59[116],pp60[116],pp61[116],pp62[116],pp63[116],pp64[116],pp65[116],pp66[116],pp67[116],pp68[116],pp69[116],pp70[116]};
    CLA_118 KS_6(s6, c6, in6_1, in6_2);
    wire[115:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp22[48],pp22[49],pp22[50],pp22[51],pp22[52],pp22[53],pp22[54],pp22[55],pp22[56],pp22[57],pp22[58],pp22[59],pp22[60],pp22[61],pp22[62],pp22[63],pp22[64],pp22[65],pp22[66],pp22[67],pp22[68],pp22[69],pp22[70],pp22[71],pp22[72],pp22[73],pp22[74],pp22[75],pp22[76],pp22[77],pp21[79],pp20[81],pp19[83],pp18[85],pp17[87],pp16[89],pp15[91],pp14[93],pp13[95],pp12[97],pp11[99],pp8[103],pp6[106],pp4[109],pp2[112],pp0[115],pp105[11],pp104[13],pp103[15],pp102[17],pp101[19],pp100[21],pp22[100],pp22[101],pp22[102],pp22[103],pp22[104],pp22[105],pp22[106],pp22[107],pp22[108],pp22[109],pp22[110],pp22[111],pp22[112],pp22[113],pp22[114],pp22[115],pp23[115],pp24[115],pp25[115],pp26[115],pp27[115],pp28[115],pp29[115],pp30[115],pp31[115],pp32[115],pp33[115],pp34[115],pp35[115],pp36[115],pp37[115],pp38[115],pp39[115],pp40[115],pp41[115],pp42[115],pp43[115],pp44[115],pp45[115],pp46[115],pp47[115],pp48[115],pp49[115],pp50[115],pp51[115],pp52[115],pp53[115],pp54[115],pp55[115],pp56[115],pp57[115],pp58[115],pp59[115],pp60[115],pp61[115],pp62[115],pp63[115],pp64[115],pp65[115],pp66[115],pp67[115],pp68[115],pp69[115],pp70[115]};
    assign in7_2 = {pp23[47],pp23[48],pp23[49],pp23[50],pp23[51],pp23[52],pp23[53],pp23[54],pp23[55],pp23[56],pp23[57],pp23[58],pp23[59],pp23[60],pp23[61],pp23[62],pp23[63],pp23[64],pp23[65],pp23[66],pp23[67],pp23[68],pp23[69],pp23[70],pp23[71],pp23[72],pp23[73],pp23[74],pp23[75],pp23[76],pp22[78],pp21[80],pp20[82],pp19[84],pp18[86],pp17[88],pp16[90],pp15[92],pp14[94],pp13[96],pp12[98],pp9[102],pp7[105],pp5[108],pp3[111],pp1[114],pp106[10],pp105[12],pp104[14],pp103[16],pp102[18],pp101[20],pp100[22],pp23[100],pp23[101],pp23[102],pp23[103],pp23[104],pp23[105],pp23[106],pp23[107],pp23[108],pp23[109],pp23[110],pp23[111],pp23[112],pp23[113],pp23[114],pp24[114],pp25[114],pp26[114],pp27[114],pp28[114],pp29[114],pp30[114],pp31[114],pp32[114],pp33[114],pp34[114],pp35[114],pp36[114],pp37[114],pp38[114],pp39[114],pp40[114],pp41[114],pp42[114],pp43[114],pp44[114],pp45[114],pp46[114],pp47[114],pp48[114],pp49[114],pp50[114],pp51[114],pp52[114],pp53[114],pp54[114],pp55[114],pp56[114],pp57[114],pp58[114],pp59[114],pp60[114],pp61[114],pp62[114],pp63[114],pp64[114],pp65[114],pp66[114],pp67[114],pp68[114],pp69[114],pp70[114],pp71[114]};
    CLA_116 KS_7(s7, c7, in7_1, in7_2);
    wire[113:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp24[47],pp24[48],pp24[49],pp24[50],pp24[51],pp24[52],pp24[53],pp24[54],pp24[55],pp24[56],pp24[57],pp24[58],pp24[59],pp24[60],pp24[61],pp24[62],pp24[63],pp24[64],pp24[65],pp24[66],pp24[67],pp24[68],pp24[69],pp24[70],pp24[71],pp24[72],pp24[73],pp24[74],pp24[75],pp23[77],pp22[79],pp21[81],pp20[83],pp19[85],pp18[87],pp17[89],pp16[91],pp15[93],pp14[95],pp13[97],pp12[99],pp8[104],pp6[107],pp4[110],pp2[113],pp0[116],pp106[11],pp105[13],pp104[15],pp103[17],pp102[19],pp101[21],pp100[23],pp24[100],pp24[101],pp24[102],pp24[103],pp24[104],pp24[105],pp24[106],pp24[107],pp24[108],pp24[109],pp24[110],pp24[111],pp24[112],pp24[113],pp25[113],pp26[113],pp27[113],pp28[113],pp29[113],pp30[113],pp31[113],pp32[113],pp33[113],pp34[113],pp35[113],pp36[113],pp37[113],pp38[113],pp39[113],pp40[113],pp41[113],pp42[113],pp43[113],pp44[113],pp45[113],pp46[113],pp47[113],pp48[113],pp49[113],pp50[113],pp51[113],pp52[113],pp53[113],pp54[113],pp55[113],pp56[113],pp57[113],pp58[113],pp59[113],pp60[113],pp61[113],pp62[113],pp63[113],pp64[113],pp65[113],pp66[113],pp67[113],pp68[113],pp69[113],pp70[113],pp71[113]};
    assign in8_2 = {pp25[46],pp25[47],pp25[48],pp25[49],pp25[50],pp25[51],pp25[52],pp25[53],pp25[54],pp25[55],pp25[56],pp25[57],pp25[58],pp25[59],pp25[60],pp25[61],pp25[62],pp25[63],pp25[64],pp25[65],pp25[66],pp25[67],pp25[68],pp25[69],pp25[70],pp25[71],pp25[72],pp25[73],pp25[74],pp24[76],pp23[78],pp22[80],pp21[82],pp20[84],pp19[86],pp18[88],pp17[90],pp16[92],pp15[94],pp14[96],pp13[98],pp9[103],pp7[106],pp5[109],pp3[112],pp1[115],pp107[10],pp106[12],pp105[14],pp104[16],pp103[18],pp102[20],pp101[22],pp100[24],pp25[100],pp25[101],pp25[102],pp25[103],pp25[104],pp25[105],pp25[106],pp25[107],pp25[108],pp25[109],pp25[110],pp25[111],pp25[112],pp26[112],pp27[112],pp28[112],pp29[112],pp30[112],pp31[112],pp32[112],pp33[112],pp34[112],pp35[112],pp36[112],pp37[112],pp38[112],pp39[112],pp40[112],pp41[112],pp42[112],pp43[112],pp44[112],pp45[112],pp46[112],pp47[112],pp48[112],pp49[112],pp50[112],pp51[112],pp52[112],pp53[112],pp54[112],pp55[112],pp56[112],pp57[112],pp58[112],pp59[112],pp60[112],pp61[112],pp62[112],pp63[112],pp64[112],pp65[112],pp66[112],pp67[112],pp68[112],pp69[112],pp70[112],pp71[112],pp72[112]};
    CLA_114 KS_8(s8, c8, in8_1, in8_2);
    wire[111:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp26[46],pp26[47],pp26[48],pp26[49],pp26[50],pp26[51],pp26[52],pp26[53],pp26[54],pp26[55],pp26[56],pp26[57],pp26[58],pp26[59],pp26[60],pp26[61],pp26[62],pp26[63],pp26[64],pp26[65],pp26[66],pp26[67],pp26[68],pp26[69],pp26[70],pp26[71],pp26[72],pp26[73],pp25[75],pp24[77],pp23[79],pp22[81],pp21[83],pp20[85],pp19[87],pp18[89],pp17[91],pp16[93],pp15[95],pp14[97],pp13[99],pp8[105],pp6[108],pp4[111],pp2[114],pp0[117],pp107[11],pp106[13],pp105[15],pp104[17],pp103[19],pp102[21],pp101[23],pp100[25],pp26[100],pp26[101],pp26[102],pp26[103],pp26[104],pp26[105],pp26[106],pp26[107],pp26[108],pp26[109],pp26[110],pp26[111],pp27[111],pp28[111],pp29[111],pp30[111],pp31[111],pp32[111],pp33[111],pp34[111],pp35[111],pp36[111],pp37[111],pp38[111],pp39[111],pp40[111],pp41[111],pp42[111],pp43[111],pp44[111],pp45[111],pp46[111],pp47[111],pp48[111],pp49[111],pp50[111],pp51[111],pp52[111],pp53[111],pp54[111],pp55[111],pp56[111],pp57[111],pp58[111],pp59[111],pp60[111],pp61[111],pp62[111],pp63[111],pp64[111],pp65[111],pp66[111],pp67[111],pp68[111],pp69[111],pp70[111],pp71[111],pp72[111]};
    assign in9_2 = {pp27[45],pp27[46],pp27[47],pp27[48],pp27[49],pp27[50],pp27[51],pp27[52],pp27[53],pp27[54],pp27[55],pp27[56],pp27[57],pp27[58],pp27[59],pp27[60],pp27[61],pp27[62],pp27[63],pp27[64],pp27[65],pp27[66],pp27[67],pp27[68],pp27[69],pp27[70],pp27[71],pp27[72],pp26[74],pp25[76],pp24[78],pp23[80],pp22[82],pp21[84],pp20[86],pp19[88],pp18[90],pp17[92],pp16[94],pp15[96],pp14[98],pp9[104],pp7[107],pp5[110],pp3[113],pp1[116],pp108[10],pp107[12],pp106[14],pp105[16],pp104[18],pp103[20],pp102[22],pp101[24],pp100[26],pp27[100],pp27[101],pp27[102],pp27[103],pp27[104],pp27[105],pp27[106],pp27[107],pp27[108],pp27[109],pp27[110],pp28[110],pp29[110],pp30[110],pp31[110],pp32[110],pp33[110],pp34[110],pp35[110],pp36[110],pp37[110],pp38[110],pp39[110],pp40[110],pp41[110],pp42[110],pp43[110],pp44[110],pp45[110],pp46[110],pp47[110],pp48[110],pp49[110],pp50[110],pp51[110],pp52[110],pp53[110],pp54[110],pp55[110],pp56[110],pp57[110],pp58[110],pp59[110],pp60[110],pp61[110],pp62[110],pp63[110],pp64[110],pp65[110],pp66[110],pp67[110],pp68[110],pp69[110],pp70[110],pp71[110],pp72[110],pp73[110]};
    CLA_112 KS_9(s9, c9, in9_1, in9_2);
    wire[109:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp28[45],pp28[46],pp28[47],pp28[48],pp28[49],pp28[50],pp28[51],pp28[52],pp28[53],pp28[54],pp28[55],pp28[56],pp28[57],pp28[58],pp28[59],pp28[60],pp28[61],pp28[62],pp28[63],pp28[64],pp28[65],pp28[66],pp28[67],pp28[68],pp28[69],pp28[70],pp28[71],pp27[73],pp26[75],pp25[77],pp24[79],pp23[81],pp22[83],pp21[85],pp20[87],pp19[89],pp18[91],pp17[93],pp16[95],pp15[97],pp14[99],pp8[106],pp6[109],pp4[112],pp2[115],pp0[118],pp108[11],pp107[13],pp106[15],pp105[17],pp104[19],pp103[21],pp102[23],pp101[25],pp100[27],pp28[100],pp28[101],pp28[102],pp28[103],pp28[104],pp28[105],pp28[106],pp28[107],pp28[108],pp28[109],pp29[109],pp30[109],pp31[109],pp32[109],pp33[109],pp34[109],pp35[109],pp36[109],pp37[109],pp38[109],pp39[109],pp40[109],pp41[109],pp42[109],pp43[109],pp44[109],pp45[109],pp46[109],pp47[109],pp48[109],pp49[109],pp50[109],pp51[109],pp52[109],pp53[109],pp54[109],pp55[109],pp56[109],pp57[109],pp58[109],pp59[109],pp60[109],pp61[109],pp62[109],pp63[109],pp64[109],pp65[109],pp66[109],pp67[109],pp68[109],pp69[109],pp70[109],pp71[109],pp72[109],pp73[109]};
    assign in10_2 = {pp29[44],pp29[45],pp29[46],pp29[47],pp29[48],pp29[49],pp29[50],pp29[51],pp29[52],pp29[53],pp29[54],pp29[55],pp29[56],pp29[57],pp29[58],pp29[59],pp29[60],pp29[61],pp29[62],pp29[63],pp29[64],pp29[65],pp29[66],pp29[67],pp29[68],pp29[69],pp29[70],pp28[72],pp27[74],pp26[76],pp25[78],pp24[80],pp23[82],pp22[84],pp21[86],pp20[88],pp19[90],pp18[92],pp17[94],pp16[96],pp15[98],pp9[105],pp7[108],pp5[111],pp3[114],pp1[117],pp109[10],pp108[12],pp107[14],pp106[16],pp105[18],pp104[20],pp103[22],pp102[24],pp101[26],pp100[28],pp29[100],pp29[101],pp29[102],pp29[103],pp29[104],pp29[105],pp29[106],pp29[107],pp29[108],pp30[108],pp31[108],pp32[108],pp33[108],pp34[108],pp35[108],pp36[108],pp37[108],pp38[108],pp39[108],pp40[108],pp41[108],pp42[108],pp43[108],pp44[108],pp45[108],pp46[108],pp47[108],pp48[108],pp49[108],pp50[108],pp51[108],pp52[108],pp53[108],pp54[108],pp55[108],pp56[108],pp57[108],pp58[108],pp59[108],pp60[108],pp61[108],pp62[108],pp63[108],pp64[108],pp65[108],pp66[108],pp67[108],pp68[108],pp69[108],pp70[108],pp71[108],pp72[108],pp73[108],pp74[108]};
    CLA_110 KS_10(s10, c10, in10_1, in10_2);
    wire[107:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp30[44],pp30[45],pp30[46],pp30[47],pp30[48],pp30[49],pp30[50],pp30[51],pp30[52],pp30[53],pp30[54],pp30[55],pp30[56],pp30[57],pp30[58],pp30[59],pp30[60],pp30[61],pp30[62],pp30[63],pp30[64],pp30[65],pp30[66],pp30[67],pp30[68],pp30[69],pp29[71],pp28[73],pp27[75],pp26[77],pp25[79],pp24[81],pp23[83],pp22[85],pp21[87],pp20[89],pp19[91],pp18[93],pp17[95],pp16[97],pp15[99],pp8[107],pp6[110],pp4[113],pp2[116],pp0[119],pp109[11],pp108[13],pp107[15],pp106[17],pp105[19],pp104[21],pp103[23],pp102[25],pp101[27],pp100[29],pp30[100],pp30[101],pp30[102],pp30[103],pp30[104],pp30[105],pp30[106],pp30[107],pp31[107],pp32[107],pp33[107],pp34[107],pp35[107],pp36[107],pp37[107],pp38[107],pp39[107],pp40[107],pp41[107],pp42[107],pp43[107],pp44[107],pp45[107],pp46[107],pp47[107],pp48[107],pp49[107],pp50[107],pp51[107],pp52[107],pp53[107],pp54[107],pp55[107],pp56[107],pp57[107],pp58[107],pp59[107],pp60[107],pp61[107],pp62[107],pp63[107],pp64[107],pp65[107],pp66[107],pp67[107],pp68[107],pp69[107],pp70[107],pp71[107],pp72[107],pp73[107],pp74[107]};
    assign in11_2 = {pp31[43],pp31[44],pp31[45],pp31[46],pp31[47],pp31[48],pp31[49],pp31[50],pp31[51],pp31[52],pp31[53],pp31[54],pp31[55],pp31[56],pp31[57],pp31[58],pp31[59],pp31[60],pp31[61],pp31[62],pp31[63],pp31[64],pp31[65],pp31[66],pp31[67],pp31[68],pp30[70],pp29[72],pp28[74],pp27[76],pp26[78],pp25[80],pp24[82],pp23[84],pp22[86],pp21[88],pp20[90],pp19[92],pp18[94],pp17[96],pp16[98],pp9[106],pp7[109],pp5[112],pp3[115],pp1[118],pp110[10],pp109[12],pp108[14],pp107[16],pp106[18],pp105[20],pp104[22],pp103[24],pp102[26],pp101[28],pp100[30],pp31[100],pp31[101],pp31[102],pp31[103],pp31[104],pp31[105],pp31[106],pp32[106],pp33[106],pp34[106],pp35[106],pp36[106],pp37[106],pp38[106],pp39[106],pp40[106],pp41[106],pp42[106],pp43[106],pp44[106],pp45[106],pp46[106],pp47[106],pp48[106],pp49[106],pp50[106],pp51[106],pp52[106],pp53[106],pp54[106],pp55[106],pp56[106],pp57[106],pp58[106],pp59[106],pp60[106],pp61[106],pp62[106],pp63[106],pp64[106],pp65[106],pp66[106],pp67[106],pp68[106],pp69[106],pp70[106],pp71[106],pp72[106],pp73[106],pp74[106],pp75[106]};
    CLA_108 KS_11(s11, c11, in11_1, in11_2);
    wire[105:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp32[43],pp32[44],pp32[45],pp32[46],pp32[47],pp32[48],pp32[49],pp32[50],pp32[51],pp32[52],pp32[53],pp32[54],pp32[55],pp32[56],pp32[57],pp32[58],pp32[59],pp32[60],pp32[61],pp32[62],pp32[63],pp32[64],pp32[65],pp32[66],pp32[67],pp31[69],pp30[71],pp29[73],pp28[75],pp27[77],pp26[79],pp25[81],pp24[83],pp23[85],pp22[87],pp21[89],pp20[91],pp19[93],pp18[95],pp17[97],pp16[99],pp8[108],pp6[111],pp4[114],pp2[117],pp0[120],pp110[11],pp109[13],pp108[15],pp107[17],pp106[19],pp105[21],pp104[23],pp103[25],pp102[27],pp101[29],pp100[31],pp32[100],pp32[101],pp32[102],pp32[103],pp32[104],pp32[105],pp33[105],pp34[105],pp35[105],pp36[105],pp37[105],pp38[105],pp39[105],pp40[105],pp41[105],pp42[105],pp43[105],pp44[105],pp45[105],pp46[105],pp47[105],pp48[105],pp49[105],pp50[105],pp51[105],pp52[105],pp53[105],pp54[105],pp55[105],pp56[105],pp57[105],pp58[105],pp59[105],pp60[105],pp61[105],pp62[105],pp63[105],pp64[105],pp65[105],pp66[105],pp67[105],pp68[105],pp69[105],pp70[105],pp71[105],pp72[105],pp73[105],pp74[105],pp75[105]};
    assign in12_2 = {pp33[42],pp33[43],pp33[44],pp33[45],pp33[46],pp33[47],pp33[48],pp33[49],pp33[50],pp33[51],pp33[52],pp33[53],pp33[54],pp33[55],pp33[56],pp33[57],pp33[58],pp33[59],pp33[60],pp33[61],pp33[62],pp33[63],pp33[64],pp33[65],pp33[66],pp32[68],pp31[70],pp30[72],pp29[74],pp28[76],pp27[78],pp26[80],pp25[82],pp24[84],pp23[86],pp22[88],pp21[90],pp20[92],pp19[94],pp18[96],pp17[98],pp9[107],pp7[110],pp5[113],pp3[116],pp1[119],pp111[10],pp110[12],pp109[14],pp108[16],pp107[18],pp106[20],pp105[22],pp104[24],pp103[26],pp102[28],pp101[30],pp100[32],pp33[100],pp33[101],pp33[102],pp33[103],pp33[104],pp34[104],pp35[104],pp36[104],pp37[104],pp38[104],pp39[104],pp40[104],pp41[104],pp42[104],pp43[104],pp44[104],pp45[104],pp46[104],pp47[104],pp48[104],pp49[104],pp50[104],pp51[104],pp52[104],pp53[104],pp54[104],pp55[104],pp56[104],pp57[104],pp58[104],pp59[104],pp60[104],pp61[104],pp62[104],pp63[104],pp64[104],pp65[104],pp66[104],pp67[104],pp68[104],pp69[104],pp70[104],pp71[104],pp72[104],pp73[104],pp74[104],pp75[104],pp76[104]};
    CLA_106 KS_12(s12, c12, in12_1, in12_2);
    wire[103:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp34[42],pp34[43],pp34[44],pp34[45],pp34[46],pp34[47],pp34[48],pp34[49],pp34[50],pp34[51],pp34[52],pp34[53],pp34[54],pp34[55],pp34[56],pp34[57],pp34[58],pp34[59],pp34[60],pp34[61],pp34[62],pp34[63],pp34[64],pp34[65],pp33[67],pp32[69],pp31[71],pp30[73],pp29[75],pp28[77],pp27[79],pp26[81],pp25[83],pp24[85],pp23[87],pp22[89],pp21[91],pp20[93],pp19[95],pp18[97],pp17[99],pp8[109],pp6[112],pp4[115],pp2[118],pp0[121],pp111[11],pp110[13],pp109[15],pp108[17],pp107[19],pp106[21],pp105[23],pp104[25],pp103[27],pp102[29],pp101[31],pp100[33],pp34[100],pp34[101],pp34[102],pp34[103],pp35[103],pp36[103],pp37[103],pp38[103],pp39[103],pp40[103],pp41[103],pp42[103],pp43[103],pp44[103],pp45[103],pp46[103],pp47[103],pp48[103],pp49[103],pp50[103],pp51[103],pp52[103],pp53[103],pp54[103],pp55[103],pp56[103],pp57[103],pp58[103],pp59[103],pp60[103],pp61[103],pp62[103],pp63[103],pp64[103],pp65[103],pp66[103],pp67[103],pp68[103],pp69[103],pp70[103],pp71[103],pp72[103],pp73[103],pp74[103],pp75[103],pp76[103]};
    assign in13_2 = {pp35[41],pp35[42],pp35[43],pp35[44],pp35[45],pp35[46],pp35[47],pp35[48],pp35[49],pp35[50],pp35[51],pp35[52],pp35[53],pp35[54],pp35[55],pp35[56],pp35[57],pp35[58],pp35[59],pp35[60],pp35[61],pp35[62],pp35[63],pp35[64],pp34[66],pp33[68],pp32[70],pp31[72],pp30[74],pp29[76],pp28[78],pp27[80],pp26[82],pp25[84],pp24[86],pp23[88],pp22[90],pp21[92],pp20[94],pp19[96],pp18[98],pp9[108],pp7[111],pp5[114],pp3[117],pp1[120],pp112[10],pp111[12],pp110[14],pp109[16],pp108[18],pp107[20],pp106[22],pp105[24],pp104[26],pp103[28],pp102[30],pp101[32],pp100[34],pp35[100],pp35[101],pp35[102],pp36[102],pp37[102],pp38[102],pp39[102],pp40[102],pp41[102],pp42[102],pp43[102],pp44[102],pp45[102],pp46[102],pp47[102],pp48[102],pp49[102],pp50[102],pp51[102],pp52[102],pp53[102],pp54[102],pp55[102],pp56[102],pp57[102],pp58[102],pp59[102],pp60[102],pp61[102],pp62[102],pp63[102],pp64[102],pp65[102],pp66[102],pp67[102],pp68[102],pp69[102],pp70[102],pp71[102],pp72[102],pp73[102],pp74[102],pp75[102],pp76[102],pp77[102]};
    CLA_104 KS_13(s13, c13, in13_1, in13_2);
    wire[101:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp36[41],pp36[42],pp36[43],pp36[44],pp36[45],pp36[46],pp36[47],pp36[48],pp36[49],pp36[50],pp36[51],pp36[52],pp36[53],pp36[54],pp36[55],pp36[56],pp36[57],pp36[58],pp36[59],pp36[60],pp36[61],pp36[62],pp36[63],pp35[65],pp34[67],pp33[69],pp32[71],pp31[73],pp30[75],pp29[77],pp28[79],pp27[81],pp26[83],pp25[85],pp24[87],pp23[89],pp22[91],pp21[93],pp20[95],pp19[97],pp18[99],pp8[110],pp6[113],pp4[116],pp2[119],pp0[122],pp112[11],pp111[13],pp110[15],pp109[17],pp108[19],pp107[21],pp106[23],pp105[25],pp104[27],pp103[29],pp102[31],pp101[33],pp100[35],pp36[100],pp36[101],pp37[101],pp38[101],pp39[101],pp40[101],pp41[101],pp42[101],pp43[101],pp44[101],pp45[101],pp46[101],pp47[101],pp48[101],pp49[101],pp50[101],pp51[101],pp52[101],pp53[101],pp54[101],pp55[101],pp56[101],pp57[101],pp58[101],pp59[101],pp60[101],pp61[101],pp62[101],pp63[101],pp64[101],pp65[101],pp66[101],pp67[101],pp68[101],pp69[101],pp70[101],pp71[101],pp72[101],pp73[101],pp74[101],pp75[101],pp76[101],pp77[101]};
    assign in14_2 = {pp37[40],pp37[41],pp37[42],pp37[43],pp37[44],pp37[45],pp37[46],pp37[47],pp37[48],pp37[49],pp37[50],pp37[51],pp37[52],pp37[53],pp37[54],pp37[55],pp37[56],pp37[57],pp37[58],pp37[59],pp37[60],pp37[61],pp37[62],pp36[64],pp35[66],pp34[68],pp33[70],pp32[72],pp31[74],pp30[76],pp29[78],pp28[80],pp27[82],pp26[84],pp25[86],pp24[88],pp23[90],pp22[92],pp21[94],pp20[96],pp19[98],pp9[109],pp7[112],pp5[115],pp3[118],pp1[121],pp113[10],pp112[12],pp111[14],pp110[16],pp109[18],pp108[20],pp107[22],pp106[24],pp105[26],pp104[28],pp103[30],pp102[32],pp101[34],pp100[36],pp37[100],pp38[100],pp39[100],pp40[100],pp41[100],pp42[100],pp43[100],pp44[100],pp45[100],pp46[100],pp47[100],pp48[100],pp49[100],pp50[100],pp51[100],pp52[100],pp53[100],pp54[100],pp55[100],pp56[100],pp57[100],pp58[100],pp59[100],pp60[100],pp61[100],pp62[100],pp63[100],pp64[100],pp65[100],pp66[100],pp67[100],pp68[100],pp69[100],pp70[100],pp71[100],pp72[100],pp73[100],pp74[100],pp75[100],pp76[100],pp77[100],pp78[100]};
    CLA_102 KS_14(s14, c14, in14_1, in14_2);
    wire[99:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp38[40],pp38[41],pp38[42],pp38[43],pp38[44],pp38[45],pp38[46],pp38[47],pp38[48],pp38[49],pp38[50],pp38[51],pp38[52],pp38[53],pp38[54],pp38[55],pp38[56],pp38[57],pp38[58],pp38[59],pp38[60],pp38[61],pp37[63],pp36[65],pp35[67],pp34[69],pp33[71],pp32[73],pp31[75],pp30[77],pp29[79],pp28[81],pp27[83],pp26[85],pp25[87],pp24[89],pp23[91],pp22[93],pp21[95],pp20[97],pp19[99],pp8[111],pp6[114],pp4[117],pp2[120],pp0[123],pp113[11],pp112[13],pp111[15],pp110[17],pp109[19],pp108[21],pp107[23],pp106[25],pp105[27],pp104[29],pp103[31],pp102[33],pp101[35],pp100[37],pp100[38],pp100[39],pp100[40],pp100[41],pp100[42],pp100[43],pp100[44],pp100[45],pp100[46],pp100[47],pp100[48],pp100[49],pp100[50],pp100[51],pp100[52],pp100[53],pp100[54],pp100[55],pp100[56],pp100[57],pp100[58],pp100[59],pp100[60],pp100[61],pp100[62],pp100[63],pp100[64],pp100[65],pp100[66],pp100[67],pp100[68],pp100[69],pp100[70],pp100[71],pp100[72],pp100[73],pp100[74],pp100[75],pp100[76],pp100[77]};
    assign in15_2 = {pp39[39],pp39[40],pp39[41],pp39[42],pp39[43],pp39[44],pp39[45],pp39[46],pp39[47],pp39[48],pp39[49],pp39[50],pp39[51],pp39[52],pp39[53],pp39[54],pp39[55],pp39[56],pp39[57],pp39[58],pp39[59],pp39[60],pp38[62],pp37[64],pp36[66],pp35[68],pp34[70],pp33[72],pp32[74],pp31[76],pp30[78],pp29[80],pp28[82],pp27[84],pp26[86],pp25[88],pp24[90],pp23[92],pp22[94],pp21[96],pp20[98],pp9[110],pp7[113],pp5[116],pp3[119],pp1[122],pp114[10],pp113[12],pp112[14],pp111[16],pp110[18],pp109[20],pp108[22],pp107[24],pp106[26],pp105[28],pp104[30],pp103[32],pp102[34],pp101[36],pp101[37],pp101[38],pp101[39],pp101[40],pp101[41],pp101[42],pp101[43],pp101[44],pp101[45],pp101[46],pp101[47],pp101[48],pp101[49],pp101[50],pp101[51],pp101[52],pp101[53],pp101[54],pp101[55],pp101[56],pp101[57],pp101[58],pp101[59],pp101[60],pp101[61],pp101[62],pp101[63],pp101[64],pp101[65],pp101[66],pp101[67],pp101[68],pp101[69],pp101[70],pp101[71],pp101[72],pp101[73],pp101[74],pp101[75],pp101[76]};
    CLA_100 KS_15(s15, c15, in15_1, in15_2);
    wire[97:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp40[39],pp40[40],pp40[41],pp40[42],pp40[43],pp40[44],pp40[45],pp40[46],pp40[47],pp40[48],pp40[49],pp40[50],pp40[51],pp40[52],pp40[53],pp40[54],pp40[55],pp40[56],pp40[57],pp40[58],pp40[59],pp39[61],pp38[63],pp37[65],pp36[67],pp35[69],pp34[71],pp33[73],pp32[75],pp31[77],pp30[79],pp29[81],pp28[83],pp27[85],pp26[87],pp25[89],pp24[91],pp23[93],pp22[95],pp21[97],pp20[99],pp8[112],pp6[115],pp4[118],pp2[121],pp0[124],pp114[11],pp113[13],pp112[15],pp111[17],pp110[19],pp109[21],pp108[23],pp107[25],pp106[27],pp105[29],pp104[31],pp103[33],pp102[35],pp102[36],pp102[37],pp102[38],pp102[39],pp102[40],pp102[41],pp102[42],pp102[43],pp102[44],pp102[45],pp102[46],pp102[47],pp102[48],pp102[49],pp102[50],pp102[51],pp102[52],pp102[53],pp102[54],pp102[55],pp102[56],pp102[57],pp102[58],pp102[59],pp102[60],pp102[61],pp102[62],pp102[63],pp102[64],pp102[65],pp102[66],pp102[67],pp102[68],pp102[69],pp102[70],pp102[71],pp102[72],pp102[73],pp102[74]};
    assign in16_2 = {pp41[38],pp41[39],pp41[40],pp41[41],pp41[42],pp41[43],pp41[44],pp41[45],pp41[46],pp41[47],pp41[48],pp41[49],pp41[50],pp41[51],pp41[52],pp41[53],pp41[54],pp41[55],pp41[56],pp41[57],pp41[58],pp40[60],pp39[62],pp38[64],pp37[66],pp36[68],pp35[70],pp34[72],pp33[74],pp32[76],pp31[78],pp30[80],pp29[82],pp28[84],pp27[86],pp26[88],pp25[90],pp24[92],pp23[94],pp22[96],pp21[98],pp9[111],pp7[114],pp5[117],pp3[120],pp1[123],pp115[10],pp114[12],pp113[14],pp112[16],pp111[18],pp110[20],pp109[22],pp108[24],pp107[26],pp106[28],pp105[30],pp104[32],pp103[34],pp103[35],pp103[36],pp103[37],pp103[38],pp103[39],pp103[40],pp103[41],pp103[42],pp103[43],pp103[44],pp103[45],pp103[46],pp103[47],pp103[48],pp103[49],pp103[50],pp103[51],pp103[52],pp103[53],pp103[54],pp103[55],pp103[56],pp103[57],pp103[58],pp103[59],pp103[60],pp103[61],pp103[62],pp103[63],pp103[64],pp103[65],pp103[66],pp103[67],pp103[68],pp103[69],pp103[70],pp103[71],pp103[72],pp103[73]};
    CLA_98 KS_16(s16, c16, in16_1, in16_2);
    wire[95:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp42[38],pp42[39],pp42[40],pp42[41],pp42[42],pp42[43],pp42[44],pp42[45],pp42[46],pp42[47],pp42[48],pp42[49],pp42[50],pp42[51],pp42[52],pp42[53],pp42[54],pp42[55],pp42[56],pp42[57],pp41[59],pp40[61],pp39[63],pp38[65],pp37[67],pp36[69],pp35[71],pp34[73],pp33[75],pp32[77],pp31[79],pp30[81],pp29[83],pp28[85],pp27[87],pp26[89],pp25[91],pp24[93],pp23[95],pp22[97],pp21[99],pp8[113],pp6[116],pp4[119],pp2[122],pp0[125],pp115[11],pp114[13],pp113[15],pp112[17],pp111[19],pp110[21],pp109[23],pp108[25],pp107[27],pp106[29],pp105[31],pp104[33],pp104[34],pp104[35],pp104[36],pp104[37],pp104[38],pp104[39],pp104[40],pp104[41],pp104[42],pp104[43],pp104[44],pp104[45],pp104[46],pp104[47],pp104[48],pp104[49],pp104[50],pp104[51],pp104[52],pp104[53],pp104[54],pp104[55],pp104[56],pp104[57],pp104[58],pp104[59],pp104[60],pp104[61],pp104[62],pp104[63],pp104[64],pp104[65],pp104[66],pp104[67],pp104[68],pp104[69],pp104[70],pp104[71]};
    assign in17_2 = {pp43[37],pp43[38],pp43[39],pp43[40],pp43[41],pp43[42],pp43[43],pp43[44],pp43[45],pp43[46],pp43[47],pp43[48],pp43[49],pp43[50],pp43[51],pp43[52],pp43[53],pp43[54],pp43[55],pp43[56],pp42[58],pp41[60],pp40[62],pp39[64],pp38[66],pp37[68],pp36[70],pp35[72],pp34[74],pp33[76],pp32[78],pp31[80],pp30[82],pp29[84],pp28[86],pp27[88],pp26[90],pp25[92],pp24[94],pp23[96],pp22[98],pp9[112],pp7[115],pp5[118],pp3[121],pp1[124],pp116[10],pp115[12],pp114[14],pp113[16],pp112[18],pp111[20],pp110[22],pp109[24],pp108[26],pp107[28],pp106[30],pp105[32],pp105[33],pp105[34],pp105[35],pp105[36],pp105[37],pp105[38],pp105[39],pp105[40],pp105[41],pp105[42],pp105[43],pp105[44],pp105[45],pp105[46],pp105[47],pp105[48],pp105[49],pp105[50],pp105[51],pp105[52],pp105[53],pp105[54],pp105[55],pp105[56],pp105[57],pp105[58],pp105[59],pp105[60],pp105[61],pp105[62],pp105[63],pp105[64],pp105[65],pp105[66],pp105[67],pp105[68],pp105[69],pp105[70]};
    CLA_96 KS_17(s17, c17, in17_1, in17_2);
    wire[93:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp44[37],pp44[38],pp44[39],pp44[40],pp44[41],pp44[42],pp44[43],pp44[44],pp44[45],pp44[46],pp44[47],pp44[48],pp44[49],pp44[50],pp44[51],pp44[52],pp44[53],pp44[54],pp44[55],pp43[57],pp42[59],pp41[61],pp40[63],pp39[65],pp38[67],pp37[69],pp36[71],pp35[73],pp34[75],pp33[77],pp32[79],pp31[81],pp30[83],pp29[85],pp28[87],pp27[89],pp26[91],pp25[93],pp24[95],pp23[97],pp22[99],pp8[114],pp6[117],pp4[120],pp2[123],pp0[126],pp116[11],pp115[13],pp114[15],pp113[17],pp112[19],pp111[21],pp110[23],pp109[25],pp108[27],pp107[29],pp106[31],pp106[32],pp106[33],pp106[34],pp106[35],pp106[36],pp106[37],pp106[38],pp106[39],pp106[40],pp106[41],pp106[42],pp106[43],pp106[44],pp106[45],pp106[46],pp106[47],pp106[48],pp106[49],pp106[50],pp106[51],pp106[52],pp106[53],pp106[54],pp106[55],pp106[56],pp106[57],pp106[58],pp106[59],pp106[60],pp106[61],pp106[62],pp106[63],pp106[64],pp106[65],pp106[66],pp106[67],pp106[68]};
    assign in18_2 = {pp45[36],pp45[37],pp45[38],pp45[39],pp45[40],pp45[41],pp45[42],pp45[43],pp45[44],pp45[45],pp45[46],pp45[47],pp45[48],pp45[49],pp45[50],pp45[51],pp45[52],pp45[53],pp45[54],pp44[56],pp43[58],pp42[60],pp41[62],pp40[64],pp39[66],pp38[68],pp37[70],pp36[72],pp35[74],pp34[76],pp33[78],pp32[80],pp31[82],pp30[84],pp29[86],pp28[88],pp27[90],pp26[92],pp25[94],pp24[96],pp23[98],pp9[113],pp7[116],pp5[119],pp3[122],pp1[125],pp117[10],pp116[12],pp115[14],pp114[16],pp113[18],pp112[20],pp111[22],pp110[24],pp109[26],pp108[28],pp107[30],pp107[31],pp107[32],pp107[33],pp107[34],pp107[35],pp107[36],pp107[37],pp107[38],pp107[39],pp107[40],pp107[41],pp107[42],pp107[43],pp107[44],pp107[45],pp107[46],pp107[47],pp107[48],pp107[49],pp107[50],pp107[51],pp107[52],pp107[53],pp107[54],pp107[55],pp107[56],pp107[57],pp107[58],pp107[59],pp107[60],pp107[61],pp107[62],pp107[63],pp107[64],pp107[65],pp107[66],pp107[67]};
    CLA_94 KS_18(s18, c18, in18_1, in18_2);
    wire[91:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp46[36],pp46[37],pp46[38],pp46[39],pp46[40],pp46[41],pp46[42],pp46[43],pp46[44],pp46[45],pp46[46],pp46[47],pp46[48],pp46[49],pp46[50],pp46[51],pp46[52],pp46[53],pp45[55],pp44[57],pp43[59],pp42[61],pp41[63],pp40[65],pp39[67],pp38[69],pp37[71],pp36[73],pp35[75],pp34[77],pp33[79],pp32[81],pp31[83],pp30[85],pp29[87],pp28[89],pp27[91],pp26[93],pp25[95],pp24[97],pp23[99],pp8[115],pp6[118],pp4[121],pp2[124],pp0[127],pp117[11],pp116[13],pp115[15],pp114[17],pp113[19],pp112[21],pp111[23],pp110[25],pp109[27],pp108[29],pp108[30],pp108[31],pp108[32],pp108[33],pp108[34],pp108[35],pp108[36],pp108[37],pp108[38],pp108[39],pp108[40],pp108[41],pp108[42],pp108[43],pp108[44],pp108[45],pp108[46],pp108[47],pp108[48],pp108[49],pp108[50],pp108[51],pp108[52],pp108[53],pp108[54],pp108[55],pp108[56],pp108[57],pp108[58],pp108[59],pp108[60],pp108[61],pp108[62],pp108[63],pp108[64],pp108[65]};
    assign in19_2 = {pp47[35],pp47[36],pp47[37],pp47[38],pp47[39],pp47[40],pp47[41],pp47[42],pp47[43],pp47[44],pp47[45],pp47[46],pp47[47],pp47[48],pp47[49],pp47[50],pp47[51],pp47[52],pp46[54],pp45[56],pp44[58],pp43[60],pp42[62],pp41[64],pp40[66],pp39[68],pp38[70],pp37[72],pp36[74],pp35[76],pp34[78],pp33[80],pp32[82],pp31[84],pp30[86],pp29[88],pp28[90],pp27[92],pp26[94],pp25[96],pp24[98],pp9[114],pp7[117],pp5[120],pp3[123],pp1[126],pp118[10],pp117[12],pp116[14],pp115[16],pp114[18],pp113[20],pp112[22],pp111[24],pp110[26],pp109[28],pp109[29],pp109[30],pp109[31],pp109[32],pp109[33],pp109[34],pp109[35],pp109[36],pp109[37],pp109[38],pp109[39],pp109[40],pp109[41],pp109[42],pp109[43],pp109[44],pp109[45],pp109[46],pp109[47],pp109[48],pp109[49],pp109[50],pp109[51],pp109[52],pp109[53],pp109[54],pp109[55],pp109[56],pp109[57],pp109[58],pp109[59],pp109[60],pp109[61],pp109[62],pp109[63],pp109[64]};
    CLA_92 KS_19(s19, c19, in19_1, in19_2);
    wire[89:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp48[35],pp48[36],pp48[37],pp48[38],pp48[39],pp48[40],pp48[41],pp48[42],pp48[43],pp48[44],pp48[45],pp48[46],pp48[47],pp48[48],pp48[49],pp48[50],pp48[51],pp47[53],pp46[55],pp45[57],pp44[59],pp43[61],pp42[63],pp41[65],pp40[67],pp39[69],pp38[71],pp37[73],pp36[75],pp35[77],pp34[79],pp33[81],pp32[83],pp31[85],pp30[87],pp29[89],pp28[91],pp27[93],pp26[95],pp25[97],pp24[99],pp8[116],pp6[119],pp4[122],pp2[125],pp1[127],pp118[11],pp117[13],pp116[15],pp115[17],pp114[19],pp113[21],pp112[23],pp111[25],pp110[27],pp110[28],pp110[29],pp110[30],pp110[31],pp110[32],pp110[33],pp110[34],pp110[35],pp110[36],pp110[37],pp110[38],pp110[39],pp110[40],pp110[41],pp110[42],pp110[43],pp110[44],pp110[45],pp110[46],pp110[47],pp110[48],pp110[49],pp110[50],pp110[51],pp110[52],pp110[53],pp110[54],pp110[55],pp110[56],pp110[57],pp110[58],pp110[59],pp110[60],pp110[61],pp110[62]};
    assign in20_2 = {pp49[34],pp49[35],pp49[36],pp49[37],pp49[38],pp49[39],pp49[40],pp49[41],pp49[42],pp49[43],pp49[44],pp49[45],pp49[46],pp49[47],pp49[48],pp49[49],pp49[50],pp48[52],pp47[54],pp46[56],pp45[58],pp44[60],pp43[62],pp42[64],pp41[66],pp40[68],pp39[70],pp38[72],pp37[74],pp36[76],pp35[78],pp34[80],pp33[82],pp32[84],pp31[86],pp30[88],pp29[90],pp28[92],pp27[94],pp26[96],pp25[98],pp9[115],pp7[118],pp5[121],pp3[124],pp2[126],pp119[10],pp118[12],pp117[14],pp116[16],pp115[18],pp114[20],pp113[22],pp112[24],pp111[26],pp111[27],pp111[28],pp111[29],pp111[30],pp111[31],pp111[32],pp111[33],pp111[34],pp111[35],pp111[36],pp111[37],pp111[38],pp111[39],pp111[40],pp111[41],pp111[42],pp111[43],pp111[44],pp111[45],pp111[46],pp111[47],pp111[48],pp111[49],pp111[50],pp111[51],pp111[52],pp111[53],pp111[54],pp111[55],pp111[56],pp111[57],pp111[58],pp111[59],pp111[60],pp111[61]};
    CLA_90 KS_20(s20, c20, in20_1, in20_2);
    wire[87:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp50[34],pp50[35],pp50[36],pp50[37],pp50[38],pp50[39],pp50[40],pp50[41],pp50[42],pp50[43],pp50[44],pp50[45],pp50[46],pp50[47],pp50[48],pp50[49],pp49[51],pp48[53],pp47[55],pp46[57],pp45[59],pp44[61],pp43[63],pp42[65],pp41[67],pp40[69],pp39[71],pp38[73],pp37[75],pp36[77],pp35[79],pp34[81],pp33[83],pp32[85],pp31[87],pp30[89],pp29[91],pp28[93],pp27[95],pp26[97],pp25[99],pp8[117],pp6[120],pp4[123],pp3[125],pp2[127],pp119[11],pp118[13],pp117[15],pp116[17],pp115[19],pp114[21],pp113[23],pp112[25],pp112[26],pp112[27],pp112[28],pp112[29],pp112[30],pp112[31],pp112[32],pp112[33],pp112[34],pp112[35],pp112[36],pp112[37],pp112[38],pp112[39],pp112[40],pp112[41],pp112[42],pp112[43],pp112[44],pp112[45],pp112[46],pp112[47],pp112[48],pp112[49],pp112[50],pp112[51],pp112[52],pp112[53],pp112[54],pp112[55],pp112[56],pp112[57],pp112[58],pp112[59]};
    assign in21_2 = {pp51[33],pp51[34],pp51[35],pp51[36],pp51[37],pp51[38],pp51[39],pp51[40],pp51[41],pp51[42],pp51[43],pp51[44],pp51[45],pp51[46],pp51[47],pp51[48],pp50[50],pp49[52],pp48[54],pp47[56],pp46[58],pp45[60],pp44[62],pp43[64],pp42[66],pp41[68],pp40[70],pp39[72],pp38[74],pp37[76],pp36[78],pp35[80],pp34[82],pp33[84],pp32[86],pp31[88],pp30[90],pp29[92],pp28[94],pp27[96],pp26[98],pp9[116],pp7[119],pp5[122],pp4[124],pp3[126],pp120[10],pp119[12],pp118[14],pp117[16],pp116[18],pp115[20],pp114[22],pp113[24],pp113[25],pp113[26],pp113[27],pp113[28],pp113[29],pp113[30],pp113[31],pp113[32],pp113[33],pp113[34],pp113[35],pp113[36],pp113[37],pp113[38],pp113[39],pp113[40],pp113[41],pp113[42],pp113[43],pp113[44],pp113[45],pp113[46],pp113[47],pp113[48],pp113[49],pp113[50],pp113[51],pp113[52],pp113[53],pp113[54],pp113[55],pp113[56],pp113[57],pp113[58]};
    CLA_88 KS_21(s21, c21, in21_1, in21_2);
    wire[85:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp52[33],pp52[34],pp52[35],pp52[36],pp52[37],pp52[38],pp52[39],pp52[40],pp52[41],pp52[42],pp52[43],pp52[44],pp52[45],pp52[46],pp52[47],pp51[49],pp50[51],pp49[53],pp48[55],pp47[57],pp46[59],pp45[61],pp44[63],pp43[65],pp42[67],pp41[69],pp40[71],pp39[73],pp38[75],pp37[77],pp36[79],pp35[81],pp34[83],pp33[85],pp32[87],pp31[89],pp30[91],pp29[93],pp28[95],pp27[97],pp26[99],pp8[118],pp6[121],pp5[123],pp4[125],pp3[127],pp120[11],pp119[13],pp118[15],pp117[17],pp116[19],pp115[21],pp114[23],pp114[24],pp114[25],pp114[26],pp114[27],pp114[28],pp114[29],pp114[30],pp114[31],pp114[32],pp114[33],pp114[34],pp114[35],pp114[36],pp114[37],pp114[38],pp114[39],pp114[40],pp114[41],pp114[42],pp114[43],pp114[44],pp114[45],pp114[46],pp114[47],pp114[48],pp114[49],pp114[50],pp114[51],pp114[52],pp114[53],pp114[54],pp114[55],pp114[56]};
    assign in22_2 = {pp53[32],pp53[33],pp53[34],pp53[35],pp53[36],pp53[37],pp53[38],pp53[39],pp53[40],pp53[41],pp53[42],pp53[43],pp53[44],pp53[45],pp53[46],pp52[48],pp51[50],pp50[52],pp49[54],pp48[56],pp47[58],pp46[60],pp45[62],pp44[64],pp43[66],pp42[68],pp41[70],pp40[72],pp39[74],pp38[76],pp37[78],pp36[80],pp35[82],pp34[84],pp33[86],pp32[88],pp31[90],pp30[92],pp29[94],pp28[96],pp27[98],pp9[117],pp7[120],pp6[122],pp5[124],pp4[126],pp121[10],pp120[12],pp119[14],pp118[16],pp117[18],pp116[20],pp115[22],pp115[23],pp115[24],pp115[25],pp115[26],pp115[27],pp115[28],pp115[29],pp115[30],pp115[31],pp115[32],pp115[33],pp115[34],pp115[35],pp115[36],pp115[37],pp115[38],pp115[39],pp115[40],pp115[41],pp115[42],pp115[43],pp115[44],pp115[45],pp115[46],pp115[47],pp115[48],pp115[49],pp115[50],pp115[51],pp115[52],pp115[53],pp115[54],pp115[55]};
    CLA_86 KS_22(s22, c22, in22_1, in22_2);
    wire[83:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp54[32],pp54[33],pp54[34],pp54[35],pp54[36],pp54[37],pp54[38],pp54[39],pp54[40],pp54[41],pp54[42],pp54[43],pp54[44],pp54[45],pp53[47],pp52[49],pp51[51],pp50[53],pp49[55],pp48[57],pp47[59],pp46[61],pp45[63],pp44[65],pp43[67],pp42[69],pp41[71],pp40[73],pp39[75],pp38[77],pp37[79],pp36[81],pp35[83],pp34[85],pp33[87],pp32[89],pp31[91],pp30[93],pp29[95],pp28[97],pp27[99],pp8[119],pp7[121],pp6[123],pp5[125],pp4[127],pp121[11],pp120[13],pp119[15],pp118[17],pp117[19],pp116[21],pp116[22],pp116[23],pp116[24],pp116[25],pp116[26],pp116[27],pp116[28],pp116[29],pp116[30],pp116[31],pp116[32],pp116[33],pp116[34],pp116[35],pp116[36],pp116[37],pp116[38],pp116[39],pp116[40],pp116[41],pp116[42],pp116[43],pp116[44],pp116[45],pp116[46],pp116[47],pp116[48],pp116[49],pp116[50],pp116[51],pp116[52],pp116[53]};
    assign in23_2 = {pp55[31],pp55[32],pp55[33],pp55[34],pp55[35],pp55[36],pp55[37],pp55[38],pp55[39],pp55[40],pp55[41],pp55[42],pp55[43],pp55[44],pp54[46],pp53[48],pp52[50],pp51[52],pp50[54],pp49[56],pp48[58],pp47[60],pp46[62],pp45[64],pp44[66],pp43[68],pp42[70],pp41[72],pp40[74],pp39[76],pp38[78],pp37[80],pp36[82],pp35[84],pp34[86],pp33[88],pp32[90],pp31[92],pp30[94],pp29[96],pp28[98],pp9[118],pp8[120],pp7[122],pp6[124],pp5[126],pp122[10],pp121[12],pp120[14],pp119[16],pp118[18],pp117[20],pp117[21],pp117[22],pp117[23],pp117[24],pp117[25],pp117[26],pp117[27],pp117[28],pp117[29],pp117[30],pp117[31],pp117[32],pp117[33],pp117[34],pp117[35],pp117[36],pp117[37],pp117[38],pp117[39],pp117[40],pp117[41],pp117[42],pp117[43],pp117[44],pp117[45],pp117[46],pp117[47],pp117[48],pp117[49],pp117[50],pp117[51],pp117[52]};
    CLA_84 KS_23(s23, c23, in23_1, in23_2);
    wire[81:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp56[31],pp56[32],pp56[33],pp56[34],pp56[35],pp56[36],pp56[37],pp56[38],pp56[39],pp56[40],pp56[41],pp56[42],pp56[43],pp55[45],pp54[47],pp53[49],pp52[51],pp51[53],pp50[55],pp49[57],pp48[59],pp47[61],pp46[63],pp45[65],pp44[67],pp43[69],pp42[71],pp41[73],pp40[75],pp39[77],pp38[79],pp37[81],pp36[83],pp35[85],pp34[87],pp33[89],pp32[91],pp31[93],pp30[95],pp29[97],pp28[99],pp9[119],pp8[121],pp7[123],pp6[125],pp5[127],pp122[11],pp121[13],pp120[15],pp119[17],pp118[19],pp118[20],pp118[21],pp118[22],pp118[23],pp118[24],pp118[25],pp118[26],pp118[27],pp118[28],pp118[29],pp118[30],pp118[31],pp118[32],pp118[33],pp118[34],pp118[35],pp118[36],pp118[37],pp118[38],pp118[39],pp118[40],pp118[41],pp118[42],pp118[43],pp118[44],pp118[45],pp118[46],pp118[47],pp118[48],pp118[49],pp118[50]};
    assign in24_2 = {pp57[30],pp57[31],pp57[32],pp57[33],pp57[34],pp57[35],pp57[36],pp57[37],pp57[38],pp57[39],pp57[40],pp57[41],pp57[42],pp56[44],pp55[46],pp54[48],pp53[50],pp52[52],pp51[54],pp50[56],pp49[58],pp48[60],pp47[62],pp46[64],pp45[66],pp44[68],pp43[70],pp42[72],pp41[74],pp40[76],pp39[78],pp38[80],pp37[82],pp36[84],pp35[86],pp34[88],pp33[90],pp32[92],pp31[94],pp30[96],pp29[98],pp29[99],pp9[120],pp8[122],pp7[124],pp6[126],pp123[10],pp122[12],pp121[14],pp120[16],pp119[18],pp119[19],pp119[20],pp119[21],pp119[22],pp119[23],pp119[24],pp119[25],pp119[26],pp119[27],pp119[28],pp119[29],pp119[30],pp119[31],pp119[32],pp119[33],pp119[34],pp119[35],pp119[36],pp119[37],pp119[38],pp119[39],pp119[40],pp119[41],pp119[42],pp119[43],pp119[44],pp119[45],pp119[46],pp119[47],pp119[48],pp119[49]};
    CLA_82 KS_24(s24, c24, in24_1, in24_2);
    wire[79:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp58[30],pp58[31],pp58[32],pp58[33],pp58[34],pp58[35],pp58[36],pp58[37],pp58[38],pp58[39],pp58[40],pp58[41],pp57[43],pp56[45],pp55[47],pp54[49],pp53[51],pp52[53],pp51[55],pp50[57],pp49[59],pp48[61],pp47[63],pp46[65],pp45[67],pp44[69],pp43[71],pp42[73],pp41[75],pp40[77],pp39[79],pp38[81],pp37[83],pp36[85],pp35[87],pp34[89],pp33[91],pp32[93],pp31[95],pp30[97],pp30[98],pp30[99],pp9[121],pp8[123],pp7[125],pp6[127],pp123[11],pp122[13],pp121[15],pp120[17],pp120[18],pp120[19],pp120[20],pp120[21],pp120[22],pp120[23],pp120[24],pp120[25],pp120[26],pp120[27],pp120[28],pp120[29],pp120[30],pp120[31],pp120[32],pp120[33],pp120[34],pp120[35],pp120[36],pp120[37],pp120[38],pp120[39],pp120[40],pp120[41],pp120[42],pp120[43],pp120[44],pp120[45],pp120[46],pp120[47]};
    assign in25_2 = {pp59[29],pp59[30],pp59[31],pp59[32],pp59[33],pp59[34],pp59[35],pp59[36],pp59[37],pp59[38],pp59[39],pp59[40],pp58[42],pp57[44],pp56[46],pp55[48],pp54[50],pp53[52],pp52[54],pp51[56],pp50[58],pp49[60],pp48[62],pp47[64],pp46[66],pp45[68],pp44[70],pp43[72],pp42[74],pp41[76],pp40[78],pp39[80],pp38[82],pp37[84],pp36[86],pp35[88],pp34[90],pp33[92],pp32[94],pp31[96],pp31[97],pp31[98],pp31[99],pp9[122],pp8[124],pp7[126],pp124[10],pp123[12],pp122[14],pp121[16],pp121[17],pp121[18],pp121[19],pp121[20],pp121[21],pp121[22],pp121[23],pp121[24],pp121[25],pp121[26],pp121[27],pp121[28],pp121[29],pp121[30],pp121[31],pp121[32],pp121[33],pp121[34],pp121[35],pp121[36],pp121[37],pp121[38],pp121[39],pp121[40],pp121[41],pp121[42],pp121[43],pp121[44],pp121[45],pp121[46]};
    CLA_80 KS_25(s25, c25, in25_1, in25_2);
    wire[77:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp60[29],pp60[30],pp60[31],pp60[32],pp60[33],pp60[34],pp60[35],pp60[36],pp60[37],pp60[38],pp60[39],pp59[41],pp58[43],pp57[45],pp56[47],pp55[49],pp54[51],pp53[53],pp52[55],pp51[57],pp50[59],pp49[61],pp48[63],pp47[65],pp46[67],pp45[69],pp44[71],pp43[73],pp42[75],pp41[77],pp40[79],pp39[81],pp38[83],pp37[85],pp36[87],pp35[89],pp34[91],pp33[93],pp32[95],pp32[96],pp32[97],pp32[98],pp32[99],pp9[123],pp8[125],pp7[127],pp124[11],pp123[13],pp122[15],pp122[16],pp122[17],pp122[18],pp122[19],pp122[20],pp122[21],pp122[22],pp122[23],pp122[24],pp122[25],pp122[26],pp122[27],pp122[28],pp122[29],pp122[30],pp122[31],pp122[32],pp122[33],pp122[34],pp122[35],pp122[36],pp122[37],pp122[38],pp122[39],pp122[40],pp122[41],pp122[42],pp122[43],pp122[44]};
    assign in26_2 = {pp61[28],pp61[29],pp61[30],pp61[31],pp61[32],pp61[33],pp61[34],pp61[35],pp61[36],pp61[37],pp61[38],pp60[40],pp59[42],pp58[44],pp57[46],pp56[48],pp55[50],pp54[52],pp53[54],pp52[56],pp51[58],pp50[60],pp49[62],pp48[64],pp47[66],pp46[68],pp45[70],pp44[72],pp43[74],pp42[76],pp41[78],pp40[80],pp39[82],pp38[84],pp37[86],pp36[88],pp35[90],pp34[92],pp33[94],pp33[95],pp33[96],pp33[97],pp33[98],pp33[99],pp9[124],pp8[126],pp125[10],pp124[12],pp123[14],pp123[15],pp123[16],pp123[17],pp123[18],pp123[19],pp123[20],pp123[21],pp123[22],pp123[23],pp123[24],pp123[25],pp123[26],pp123[27],pp123[28],pp123[29],pp123[30],pp123[31],pp123[32],pp123[33],pp123[34],pp123[35],pp123[36],pp123[37],pp123[38],pp123[39],pp123[40],pp123[41],pp123[42],pp123[43]};
    CLA_78 KS_26(s26, c26, in26_1, in26_2);
    wire[75:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp62[28],pp62[29],pp62[30],pp62[31],pp62[32],pp62[33],pp62[34],pp62[35],pp62[36],pp62[37],pp61[39],pp60[41],pp59[43],pp58[45],pp57[47],pp56[49],pp55[51],pp54[53],pp53[55],pp52[57],pp51[59],pp50[61],pp49[63],pp48[65],pp47[67],pp46[69],pp45[71],pp44[73],pp43[75],pp42[77],pp41[79],pp40[81],pp39[83],pp38[85],pp37[87],pp36[89],pp35[91],pp34[93],pp34[94],pp34[95],pp34[96],pp34[97],pp34[98],pp34[99],pp9[125],pp8[127],pp125[11],pp124[13],pp124[14],pp124[15],pp124[16],pp124[17],pp124[18],pp124[19],pp124[20],pp124[21],pp124[22],pp124[23],pp124[24],pp124[25],pp124[26],pp124[27],pp124[28],pp124[29],pp124[30],pp124[31],pp124[32],pp124[33],pp124[34],pp124[35],pp124[36],pp124[37],pp124[38],pp124[39],pp124[40],pp124[41]};
    assign in27_2 = {pp63[27],pp63[28],pp63[29],pp63[30],pp63[31],pp63[32],pp63[33],pp63[34],pp63[35],pp63[36],pp62[38],pp61[40],pp60[42],pp59[44],pp58[46],pp57[48],pp56[50],pp55[52],pp54[54],pp53[56],pp52[58],pp51[60],pp50[62],pp49[64],pp48[66],pp47[68],pp46[70],pp45[72],pp44[74],pp43[76],pp42[78],pp41[80],pp40[82],pp39[84],pp38[86],pp37[88],pp36[90],pp35[92],pp35[93],pp35[94],pp35[95],pp35[96],pp35[97],pp35[98],pp35[99],pp9[126],pp126[10],pp125[12],pp125[13],pp125[14],pp125[15],pp125[16],pp125[17],pp125[18],pp125[19],pp125[20],pp125[21],pp125[22],pp125[23],pp125[24],pp125[25],pp125[26],pp125[27],pp125[28],pp125[29],pp125[30],pp125[31],pp125[32],pp125[33],pp125[34],pp125[35],pp125[36],pp125[37],pp125[38],pp125[39],pp125[40]};
    CLA_76 KS_27(s27, c27, in27_1, in27_2);
    wire[73:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp64[27],pp64[28],pp64[29],pp64[30],pp64[31],pp64[32],pp64[33],pp64[34],pp64[35],pp63[37],pp62[39],pp61[41],pp60[43],pp59[45],pp58[47],pp57[49],pp56[51],pp55[53],pp54[55],pp53[57],pp52[59],pp51[61],pp50[63],pp49[65],pp48[67],pp47[69],pp46[71],pp45[73],pp44[75],pp43[77],pp42[79],pp41[81],pp40[83],pp39[85],pp38[87],pp37[89],pp36[91],pp36[92],pp36[93],pp36[94],pp36[95],pp36[96],pp36[97],pp36[98],pp36[99],pp9[127],pp126[11],pp126[12],pp126[13],pp126[14],pp126[15],pp126[16],pp126[17],pp126[18],pp126[19],pp126[20],pp126[21],pp126[22],pp126[23],pp126[24],pp126[25],pp126[26],pp126[27],pp126[28],pp126[29],pp126[30],pp126[31],pp126[32],pp126[33],pp126[34],pp126[35],pp126[36],pp126[37],pp126[38]};
    assign in28_2 = {pp65[26],pp65[27],pp65[28],pp65[29],pp65[30],pp65[31],pp65[32],pp65[33],pp65[34],pp64[36],pp63[38],pp62[40],pp61[42],pp60[44],pp59[46],pp58[48],pp57[50],pp56[52],pp55[54],pp54[56],pp53[58],pp52[60],pp51[62],pp50[64],pp49[66],pp48[68],pp47[70],pp46[72],pp45[74],pp44[76],pp43[78],pp42[80],pp41[82],pp40[84],pp39[86],pp38[88],pp37[90],pp37[91],pp37[92],pp37[93],pp37[94],pp37[95],pp37[96],pp37[97],pp37[98],pp37[99],pp127[10],pp127[11],pp127[12],pp127[13],pp127[14],pp127[15],pp127[16],pp127[17],pp127[18],pp127[19],pp127[20],pp127[21],pp127[22],pp127[23],pp127[24],pp127[25],pp127[26],pp127[27],pp127[28],pp127[29],pp127[30],pp127[31],pp127[32],pp127[33],pp127[34],pp127[35],pp127[36],pp127[37]};
    CLA_74 KS_28(s28, c28, in28_1, in28_2);
    wire[71:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp66[26],pp66[27],pp66[28],pp66[29],pp66[30],pp66[31],pp66[32],pp66[33],pp65[35],pp64[37],pp63[39],pp62[41],pp61[43],pp60[45],pp59[47],pp58[49],pp57[51],pp56[53],pp55[55],pp54[57],pp53[59],pp52[61],pp51[63],pp50[65],pp49[67],pp48[69],pp47[71],pp46[73],pp45[75],pp44[77],pp43[79],pp42[81],pp41[83],pp40[85],pp39[87],pp38[89],pp38[90],pp38[91],pp38[92],pp38[93],pp38[94],pp38[95],pp38[96],pp38[97],pp38[98],pp38[99],pp39[99],pp40[99],pp41[99],pp42[99],pp43[99],pp44[99],pp45[99],pp46[99],pp47[99],pp48[99],pp49[99],pp50[99],pp51[99],pp52[99],pp53[99],pp54[99],pp55[99],pp56[99],pp57[99],pp58[99],pp59[99],pp60[99],pp61[99],pp62[99],pp63[99],pp64[99]};
    assign in29_2 = {pp67[25],pp67[26],pp67[27],pp67[28],pp67[29],pp67[30],pp67[31],pp67[32],pp66[34],pp65[36],pp64[38],pp63[40],pp62[42],pp61[44],pp60[46],pp59[48],pp58[50],pp57[52],pp56[54],pp55[56],pp54[58],pp53[60],pp52[62],pp51[64],pp50[66],pp49[68],pp48[70],pp47[72],pp46[74],pp45[76],pp44[78],pp43[80],pp42[82],pp41[84],pp40[86],pp39[88],pp39[89],pp39[90],pp39[91],pp39[92],pp39[93],pp39[94],pp39[95],pp39[96],pp39[97],pp39[98],pp40[98],pp41[98],pp42[98],pp43[98],pp44[98],pp45[98],pp46[98],pp47[98],pp48[98],pp49[98],pp50[98],pp51[98],pp52[98],pp53[98],pp54[98],pp55[98],pp56[98],pp57[98],pp58[98],pp59[98],pp60[98],pp61[98],pp62[98],pp63[98],pp64[98],pp65[98]};
    CLA_72 KS_29(s29, c29, in29_1, in29_2);
    wire[69:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp68[25],pp68[26],pp68[27],pp68[28],pp68[29],pp68[30],pp68[31],pp67[33],pp66[35],pp65[37],pp64[39],pp63[41],pp62[43],pp61[45],pp60[47],pp59[49],pp58[51],pp57[53],pp56[55],pp55[57],pp54[59],pp53[61],pp52[63],pp51[65],pp50[67],pp49[69],pp48[71],pp47[73],pp46[75],pp45[77],pp44[79],pp43[81],pp42[83],pp41[85],pp40[87],pp40[88],pp40[89],pp40[90],pp40[91],pp40[92],pp40[93],pp40[94],pp40[95],pp40[96],pp40[97],pp41[97],pp42[97],pp43[97],pp44[97],pp45[97],pp46[97],pp47[97],pp48[97],pp49[97],pp50[97],pp51[97],pp52[97],pp53[97],pp54[97],pp55[97],pp56[97],pp57[97],pp58[97],pp59[97],pp60[97],pp61[97],pp62[97],pp63[97],pp64[97],pp65[97]};
    assign in30_2 = {pp69[24],pp69[25],pp69[26],pp69[27],pp69[28],pp69[29],pp69[30],pp68[32],pp67[34],pp66[36],pp65[38],pp64[40],pp63[42],pp62[44],pp61[46],pp60[48],pp59[50],pp58[52],pp57[54],pp56[56],pp55[58],pp54[60],pp53[62],pp52[64],pp51[66],pp50[68],pp49[70],pp48[72],pp47[74],pp46[76],pp45[78],pp44[80],pp43[82],pp42[84],pp41[86],pp41[87],pp41[88],pp41[89],pp41[90],pp41[91],pp41[92],pp41[93],pp41[94],pp41[95],pp41[96],pp42[96],pp43[96],pp44[96],pp45[96],pp46[96],pp47[96],pp48[96],pp49[96],pp50[96],pp51[96],pp52[96],pp53[96],pp54[96],pp55[96],pp56[96],pp57[96],pp58[96],pp59[96],pp60[96],pp61[96],pp62[96],pp63[96],pp64[96],pp65[96],pp66[96]};
    CLA_70 KS_30(s30, c30, in30_1, in30_2);
    wire[67:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp70[24],pp70[25],pp70[26],pp70[27],pp70[28],pp70[29],pp69[31],pp68[33],pp67[35],pp66[37],pp65[39],pp64[41],pp63[43],pp62[45],pp61[47],pp60[49],pp59[51],pp58[53],pp57[55],pp56[57],pp55[59],pp54[61],pp53[63],pp52[65],pp51[67],pp50[69],pp49[71],pp48[73],pp47[75],pp46[77],pp45[79],pp44[81],pp43[83],pp42[85],pp42[86],pp42[87],pp42[88],pp42[89],pp42[90],pp42[91],pp42[92],pp42[93],pp42[94],pp42[95],pp43[95],pp44[95],pp45[95],pp46[95],pp47[95],pp48[95],pp49[95],pp50[95],pp51[95],pp52[95],pp53[95],pp54[95],pp55[95],pp56[95],pp57[95],pp58[95],pp59[95],pp60[95],pp61[95],pp62[95],pp63[95],pp64[95],pp65[95],pp66[95]};
    assign in31_2 = {pp71[23],pp71[24],pp71[25],pp71[26],pp71[27],pp71[28],pp70[30],pp69[32],pp68[34],pp67[36],pp66[38],pp65[40],pp64[42],pp63[44],pp62[46],pp61[48],pp60[50],pp59[52],pp58[54],pp57[56],pp56[58],pp55[60],pp54[62],pp53[64],pp52[66],pp51[68],pp50[70],pp49[72],pp48[74],pp47[76],pp46[78],pp45[80],pp44[82],pp43[84],pp43[85],pp43[86],pp43[87],pp43[88],pp43[89],pp43[90],pp43[91],pp43[92],pp43[93],pp43[94],pp44[94],pp45[94],pp46[94],pp47[94],pp48[94],pp49[94],pp50[94],pp51[94],pp52[94],pp53[94],pp54[94],pp55[94],pp56[94],pp57[94],pp58[94],pp59[94],pp60[94],pp61[94],pp62[94],pp63[94],pp64[94],pp65[94],pp66[94],pp67[94]};
    CLA_68 KS_31(s31, c31, in31_1, in31_2);
    wire[65:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp72[23],pp72[24],pp72[25],pp72[26],pp72[27],pp71[29],pp70[31],pp69[33],pp68[35],pp67[37],pp66[39],pp65[41],pp64[43],pp63[45],pp62[47],pp61[49],pp60[51],pp59[53],pp58[55],pp57[57],pp56[59],pp55[61],pp54[63],pp53[65],pp52[67],pp51[69],pp50[71],pp49[73],pp48[75],pp47[77],pp46[79],pp45[81],pp44[83],pp44[84],pp44[85],pp44[86],pp44[87],pp44[88],pp44[89],pp44[90],pp44[91],pp44[92],pp44[93],pp45[93],pp46[93],pp47[93],pp48[93],pp49[93],pp50[93],pp51[93],pp52[93],pp53[93],pp54[93],pp55[93],pp56[93],pp57[93],pp58[93],pp59[93],pp60[93],pp61[93],pp62[93],pp63[93],pp64[93],pp65[93],pp66[93],pp67[93]};
    assign in32_2 = {pp73[22],pp73[23],pp73[24],pp73[25],pp73[26],pp72[28],pp71[30],pp70[32],pp69[34],pp68[36],pp67[38],pp66[40],pp65[42],pp64[44],pp63[46],pp62[48],pp61[50],pp60[52],pp59[54],pp58[56],pp57[58],pp56[60],pp55[62],pp54[64],pp53[66],pp52[68],pp51[70],pp50[72],pp49[74],pp48[76],pp47[78],pp46[80],pp45[82],pp45[83],pp45[84],pp45[85],pp45[86],pp45[87],pp45[88],pp45[89],pp45[90],pp45[91],pp45[92],pp46[92],pp47[92],pp48[92],pp49[92],pp50[92],pp51[92],pp52[92],pp53[92],pp54[92],pp55[92],pp56[92],pp57[92],pp58[92],pp59[92],pp60[92],pp61[92],pp62[92],pp63[92],pp64[92],pp65[92],pp66[92],pp67[92],pp68[92]};
    CLA_66 KS_32(s32, c32, in32_1, in32_2);
    wire[63:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp74[22],pp74[23],pp74[24],pp74[25],pp73[27],pp72[29],pp71[31],pp70[33],pp69[35],pp68[37],pp67[39],pp66[41],pp65[43],pp64[45],pp63[47],pp62[49],pp61[51],pp60[53],pp59[55],pp58[57],pp57[59],pp56[61],pp55[63],pp54[65],pp53[67],pp52[69],pp51[71],pp50[73],pp49[75],pp48[77],pp47[79],pp46[81],pp46[82],pp46[83],pp46[84],pp46[85],pp46[86],pp46[87],pp46[88],pp46[89],pp46[90],pp46[91],pp47[91],pp48[91],pp49[91],pp50[91],pp51[91],pp52[91],pp53[91],pp54[91],pp55[91],pp56[91],pp57[91],pp58[91],pp59[91],pp60[91],pp61[91],pp62[91],pp63[91],pp64[91],pp65[91],pp66[91],pp67[91],pp68[91]};
    assign in33_2 = {pp75[21],pp75[22],pp75[23],pp75[24],pp74[26],pp73[28],pp72[30],pp71[32],pp70[34],pp69[36],pp68[38],pp67[40],pp66[42],pp65[44],pp64[46],pp63[48],pp62[50],pp61[52],pp60[54],pp59[56],pp58[58],pp57[60],pp56[62],pp55[64],pp54[66],pp53[68],pp52[70],pp51[72],pp50[74],pp49[76],pp48[78],pp47[80],pp47[81],pp47[82],pp47[83],pp47[84],pp47[85],pp47[86],pp47[87],pp47[88],pp47[89],pp47[90],pp48[90],pp49[90],pp50[90],pp51[90],pp52[90],pp53[90],pp54[90],pp55[90],pp56[90],pp57[90],pp58[90],pp59[90],pp60[90],pp61[90],pp62[90],pp63[90],pp64[90],pp65[90],pp66[90],pp67[90],pp68[90],pp69[90]};
    CLA_64 KS_33(s33, c33, in33_1, in33_2);
    wire[61:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp76[21],pp76[22],pp76[23],pp75[25],pp74[27],pp73[29],pp72[31],pp71[33],pp70[35],pp69[37],pp68[39],pp67[41],pp66[43],pp65[45],pp64[47],pp63[49],pp62[51],pp61[53],pp60[55],pp59[57],pp58[59],pp57[61],pp56[63],pp55[65],pp54[67],pp53[69],pp52[71],pp51[73],pp50[75],pp49[77],pp48[79],pp48[80],pp48[81],pp48[82],pp48[83],pp48[84],pp48[85],pp48[86],pp48[87],pp48[88],pp48[89],pp49[89],pp50[89],pp51[89],pp52[89],pp53[89],pp54[89],pp55[89],pp56[89],pp57[89],pp58[89],pp59[89],pp60[89],pp61[89],pp62[89],pp63[89],pp64[89],pp65[89],pp66[89],pp67[89],pp68[89],pp69[89]};
    assign in34_2 = {pp77[20],pp77[21],pp77[22],pp76[24],pp75[26],pp74[28],pp73[30],pp72[32],pp71[34],pp70[36],pp69[38],pp68[40],pp67[42],pp66[44],pp65[46],pp64[48],pp63[50],pp62[52],pp61[54],pp60[56],pp59[58],pp58[60],pp57[62],pp56[64],pp55[66],pp54[68],pp53[70],pp52[72],pp51[74],pp50[76],pp49[78],pp49[79],pp49[80],pp49[81],pp49[82],pp49[83],pp49[84],pp49[85],pp49[86],pp49[87],pp49[88],pp50[88],pp51[88],pp52[88],pp53[88],pp54[88],pp55[88],pp56[88],pp57[88],pp58[88],pp59[88],pp60[88],pp61[88],pp62[88],pp63[88],pp64[88],pp65[88],pp66[88],pp67[88],pp68[88],pp69[88],pp70[88]};
    CLA_62 KS_34(s34, c34, in34_1, in34_2);
    wire[59:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp78[20],pp78[21],pp77[23],pp76[25],pp75[27],pp74[29],pp73[31],pp72[33],pp71[35],pp70[37],pp69[39],pp68[41],pp67[43],pp66[45],pp65[47],pp64[49],pp63[51],pp62[53],pp61[55],pp60[57],pp59[59],pp58[61],pp57[63],pp56[65],pp55[67],pp54[69],pp53[71],pp52[73],pp51[75],pp50[77],pp50[78],pp50[79],pp50[80],pp50[81],pp50[82],pp50[83],pp50[84],pp50[85],pp50[86],pp50[87],pp51[87],pp52[87],pp53[87],pp54[87],pp55[87],pp56[87],pp57[87],pp58[87],pp59[87],pp60[87],pp61[87],pp62[87],pp63[87],pp64[87],pp65[87],pp66[87],pp67[87],pp68[87],pp69[87],pp70[87]};
    assign in35_2 = {pp79[19],pp79[20],pp78[22],pp77[24],pp76[26],pp75[28],pp74[30],pp73[32],pp72[34],pp71[36],pp70[38],pp69[40],pp68[42],pp67[44],pp66[46],pp65[48],pp64[50],pp63[52],pp62[54],pp61[56],pp60[58],pp59[60],pp58[62],pp57[64],pp56[66],pp55[68],pp54[70],pp53[72],pp52[74],pp51[76],pp51[77],pp51[78],pp51[79],pp51[80],pp51[81],pp51[82],pp51[83],pp51[84],pp51[85],pp51[86],pp52[86],pp53[86],pp54[86],pp55[86],pp56[86],pp57[86],pp58[86],pp59[86],pp60[86],pp61[86],pp62[86],pp63[86],pp64[86],pp65[86],pp66[86],pp67[86],pp68[86],pp69[86],pp70[86],pp71[86]};
    CLA_60 KS_35(s35, c35, in35_1, in35_2);
    wire[57:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp80[19],pp79[21],pp78[23],pp77[25],pp76[27],pp75[29],pp74[31],pp73[33],pp72[35],pp71[37],pp70[39],pp69[41],pp68[43],pp67[45],pp66[47],pp65[49],pp64[51],pp63[53],pp62[55],pp61[57],pp60[59],pp59[61],pp58[63],pp57[65],pp56[67],pp55[69],pp54[71],pp53[73],pp52[75],pp52[76],pp52[77],pp52[78],pp52[79],pp52[80],pp52[81],pp52[82],pp52[83],pp52[84],pp52[85],pp53[85],pp54[85],pp55[85],pp56[85],pp57[85],pp58[85],pp59[85],pp60[85],pp61[85],pp62[85],pp63[85],pp64[85],pp65[85],pp66[85],pp67[85],pp68[85],pp69[85],pp70[85],pp71[85]};
    assign in36_2 = {pp81[18],pp80[20],pp79[22],pp78[24],pp77[26],pp76[28],pp75[30],pp74[32],pp73[34],pp72[36],pp71[38],pp70[40],pp69[42],pp68[44],pp67[46],pp66[48],pp65[50],pp64[52],pp63[54],pp62[56],pp61[58],pp60[60],pp59[62],pp58[64],pp57[66],pp56[68],pp55[70],pp54[72],pp53[74],pp53[75],pp53[76],pp53[77],pp53[78],pp53[79],pp53[80],pp53[81],pp53[82],pp53[83],pp53[84],pp54[84],pp55[84],pp56[84],pp57[84],pp58[84],pp59[84],pp60[84],pp61[84],pp62[84],pp63[84],pp64[84],pp65[84],pp66[84],pp67[84],pp68[84],pp69[84],pp70[84],pp71[84],pp72[84]};
    CLA_58 KS_36(s36, c36, in36_1, in36_2);
    wire[55:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp81[19],pp80[21],pp79[23],pp78[25],pp77[27],pp76[29],pp75[31],pp74[33],pp73[35],pp72[37],pp71[39],pp70[41],pp69[43],pp68[45],pp67[47],pp66[49],pp65[51],pp64[53],pp63[55],pp62[57],pp61[59],pp60[61],pp59[63],pp58[65],pp57[67],pp56[69],pp55[71],pp54[73],pp54[74],pp54[75],pp54[76],pp54[77],pp54[78],pp54[79],pp54[80],pp54[81],pp54[82],pp54[83],pp55[83],pp56[83],pp57[83],pp58[83],pp59[83],pp60[83],pp61[83],pp62[83],pp63[83],pp64[83],pp65[83],pp66[83],pp67[83],pp68[83],pp69[83],pp70[83],pp71[83],pp72[83]};
    assign in37_2 = {pp82[18],pp81[20],pp80[22],pp79[24],pp78[26],pp77[28],pp76[30],pp75[32],pp74[34],pp73[36],pp72[38],pp71[40],pp70[42],pp69[44],pp68[46],pp67[48],pp66[50],pp65[52],pp64[54],pp63[56],pp62[58],pp61[60],pp60[62],pp59[64],pp58[66],pp57[68],pp56[70],pp55[72],pp55[73],pp55[74],pp55[75],pp55[76],pp55[77],pp55[78],pp55[79],pp55[80],pp55[81],pp55[82],pp56[82],pp57[82],pp58[82],pp59[82],pp60[82],pp61[82],pp62[82],pp63[82],pp64[82],pp65[82],pp66[82],pp67[82],pp68[82],pp69[82],pp70[82],pp71[82],pp72[82],pp73[82]};
    CLA_56 KS_37(s37, c37, in37_1, in37_2);
    wire[53:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp82[19],pp81[21],pp80[23],pp79[25],pp78[27],pp77[29],pp76[31],pp75[33],pp74[35],pp73[37],pp72[39],pp71[41],pp70[43],pp69[45],pp68[47],pp67[49],pp66[51],pp65[53],pp64[55],pp63[57],pp62[59],pp61[61],pp60[63],pp59[65],pp58[67],pp57[69],pp56[71],pp56[72],pp56[73],pp56[74],pp56[75],pp56[76],pp56[77],pp56[78],pp56[79],pp56[80],pp56[81],pp57[81],pp58[81],pp59[81],pp60[81],pp61[81],pp62[81],pp63[81],pp64[81],pp65[81],pp66[81],pp67[81],pp68[81],pp69[81],pp70[81],pp71[81],pp72[81],pp73[81]};
    assign in38_2 = {pp83[18],pp82[20],pp81[22],pp80[24],pp79[26],pp78[28],pp77[30],pp76[32],pp75[34],pp74[36],pp73[38],pp72[40],pp71[42],pp70[44],pp69[46],pp68[48],pp67[50],pp66[52],pp65[54],pp64[56],pp63[58],pp62[60],pp61[62],pp60[64],pp59[66],pp58[68],pp57[70],pp57[71],pp57[72],pp57[73],pp57[74],pp57[75],pp57[76],pp57[77],pp57[78],pp57[79],pp57[80],pp58[80],pp59[80],pp60[80],pp61[80],pp62[80],pp63[80],pp64[80],pp65[80],pp66[80],pp67[80],pp68[80],pp69[80],pp70[80],pp71[80],pp72[80],pp73[80],pp74[80]};
    CLA_54 KS_38(s38, c38, in38_1, in38_2);
    wire[51:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp83[19],pp82[21],pp81[23],pp80[25],pp79[27],pp78[29],pp77[31],pp76[33],pp75[35],pp74[37],pp73[39],pp72[41],pp71[43],pp70[45],pp69[47],pp68[49],pp67[51],pp66[53],pp65[55],pp64[57],pp63[59],pp62[61],pp61[63],pp60[65],pp59[67],pp58[69],pp58[70],pp58[71],pp58[72],pp58[73],pp58[74],pp58[75],pp58[76],pp58[77],pp58[78],pp58[79],pp59[79],pp60[79],pp61[79],pp62[79],pp63[79],pp64[79],pp65[79],pp66[79],pp67[79],pp68[79],pp69[79],pp70[79],pp71[79],pp72[79],pp73[79],pp74[79]};
    assign in39_2 = {pp84[18],pp83[20],pp82[22],pp81[24],pp80[26],pp79[28],pp78[30],pp77[32],pp76[34],pp75[36],pp74[38],pp73[40],pp72[42],pp71[44],pp70[46],pp69[48],pp68[50],pp67[52],pp66[54],pp65[56],pp64[58],pp63[60],pp62[62],pp61[64],pp60[66],pp59[68],pp59[69],pp59[70],pp59[71],pp59[72],pp59[73],pp59[74],pp59[75],pp59[76],pp59[77],pp59[78],pp60[78],pp61[78],pp62[78],pp63[78],pp64[78],pp65[78],pp66[78],pp67[78],pp68[78],pp69[78],pp70[78],pp71[78],pp72[78],pp73[78],pp74[78],pp75[78]};
    CLA_52 KS_39(s39, c39, in39_1, in39_2);
    wire[49:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp84[19],pp83[21],pp82[23],pp81[25],pp80[27],pp79[29],pp78[31],pp77[33],pp76[35],pp75[37],pp74[39],pp73[41],pp72[43],pp71[45],pp70[47],pp69[49],pp68[51],pp67[53],pp66[55],pp65[57],pp64[59],pp63[61],pp62[63],pp61[65],pp60[67],pp60[68],pp60[69],pp60[70],pp60[71],pp60[72],pp60[73],pp60[74],pp60[75],pp60[76],pp60[77],pp61[77],pp62[77],pp63[77],pp64[77],pp65[77],pp66[77],pp67[77],pp68[77],pp69[77],pp70[77],pp71[77],pp72[77],pp73[77],pp74[77],pp75[77]};
    assign in40_2 = {pp85[18],pp84[20],pp83[22],pp82[24],pp81[26],pp80[28],pp79[30],pp78[32],pp77[34],pp76[36],pp75[38],pp74[40],pp73[42],pp72[44],pp71[46],pp70[48],pp69[50],pp68[52],pp67[54],pp66[56],pp65[58],pp64[60],pp63[62],pp62[64],pp61[66],pp61[67],pp61[68],pp61[69],pp61[70],pp61[71],pp61[72],pp61[73],pp61[74],pp61[75],pp61[76],pp62[76],pp63[76],pp64[76],pp65[76],pp66[76],pp67[76],pp68[76],pp69[76],pp70[76],pp71[76],pp72[76],pp73[76],pp74[76],pp75[76],pp76[76]};
    CLA_50 KS_40(s40, c40, in40_1, in40_2);
    wire[47:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp85[19],pp84[21],pp83[23],pp82[25],pp81[27],pp80[29],pp79[31],pp78[33],pp77[35],pp76[37],pp75[39],pp74[41],pp73[43],pp72[45],pp71[47],pp70[49],pp69[51],pp68[53],pp67[55],pp66[57],pp65[59],pp64[61],pp63[63],pp62[65],pp62[66],pp62[67],pp62[68],pp62[69],pp62[70],pp62[71],pp62[72],pp62[73],pp62[74],pp62[75],pp63[75],pp64[75],pp65[75],pp66[75],pp67[75],pp68[75],pp69[75],pp70[75],pp71[75],pp72[75],pp73[75],pp74[75],pp75[75],pp76[75]};
    assign in41_2 = {pp86[18],pp85[20],pp84[22],pp83[24],pp82[26],pp81[28],pp80[30],pp79[32],pp78[34],pp77[36],pp76[38],pp75[40],pp74[42],pp73[44],pp72[46],pp71[48],pp70[50],pp69[52],pp68[54],pp67[56],pp66[58],pp65[60],pp64[62],pp63[64],pp63[65],pp63[66],pp63[67],pp63[68],pp63[69],pp63[70],pp63[71],pp63[72],pp63[73],pp63[74],pp64[74],pp65[74],pp66[74],pp67[74],pp68[74],pp69[74],pp70[74],pp71[74],pp72[74],pp73[74],pp74[74],pp75[74],pp76[74],pp77[74]};
    CLA_48 KS_41(s41, c41, in41_1, in41_2);
    wire[45:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp86[19],pp85[21],pp84[23],pp83[25],pp82[27],pp81[29],pp80[31],pp79[33],pp78[35],pp77[37],pp76[39],pp75[41],pp74[43],pp73[45],pp72[47],pp71[49],pp70[51],pp69[53],pp68[55],pp67[57],pp66[59],pp65[61],pp64[63],pp64[64],pp64[65],pp64[66],pp64[67],pp64[68],pp64[69],pp64[70],pp64[71],pp64[72],pp64[73],pp65[73],pp66[73],pp67[73],pp68[73],pp69[73],pp70[73],pp71[73],pp72[73],pp73[73],pp74[73],pp75[73],pp76[73],pp77[73]};
    assign in42_2 = {pp87[18],pp86[20],pp85[22],pp84[24],pp83[26],pp82[28],pp81[30],pp80[32],pp79[34],pp78[36],pp77[38],pp76[40],pp75[42],pp74[44],pp73[46],pp72[48],pp71[50],pp70[52],pp69[54],pp68[56],pp67[58],pp66[60],pp65[62],pp65[63],pp65[64],pp65[65],pp65[66],pp65[67],pp65[68],pp65[69],pp65[70],pp65[71],pp65[72],pp66[72],pp67[72],pp68[72],pp69[72],pp70[72],pp71[72],pp72[72],pp73[72],pp74[72],pp75[72],pp76[72],pp77[72],pp78[72]};
    CLA_46 KS_42(s42, c42, in42_1, in42_2);
    wire[43:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp87[19],pp86[21],pp85[23],pp84[25],pp83[27],pp82[29],pp81[31],pp80[33],pp79[35],pp78[37],pp77[39],pp76[41],pp75[43],pp74[45],pp73[47],pp72[49],pp71[51],pp70[53],pp69[55],pp68[57],pp67[59],pp66[61],pp66[62],pp66[63],pp66[64],pp66[65],pp66[66],pp66[67],pp66[68],pp66[69],pp66[70],pp66[71],pp67[71],pp68[71],pp69[71],pp70[71],pp71[71],pp72[71],pp73[71],pp74[71],pp75[71],pp76[71],pp77[71],pp78[71]};
    assign in43_2 = {pp88[18],pp87[20],pp86[22],pp85[24],pp84[26],pp83[28],pp82[30],pp81[32],pp80[34],pp79[36],pp78[38],pp77[40],pp76[42],pp75[44],pp74[46],pp73[48],pp72[50],pp71[52],pp70[54],pp69[56],pp68[58],pp67[60],pp67[61],pp67[62],pp67[63],pp67[64],pp67[65],pp67[66],pp67[67],pp67[68],pp67[69],pp67[70],pp68[70],pp69[70],pp70[70],pp71[70],pp72[70],pp73[70],pp74[70],pp75[70],pp76[70],pp77[70],pp78[70],pp79[70]};
    CLA_44 KS_43(s43, c43, in43_1, in43_2);
    wire[41:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp88[19],pp87[21],pp86[23],pp85[25],pp84[27],pp83[29],pp82[31],pp81[33],pp80[35],pp79[37],pp78[39],pp77[41],pp76[43],pp75[45],pp74[47],pp73[49],pp72[51],pp71[53],pp70[55],pp69[57],pp68[59],pp68[60],pp68[61],pp68[62],pp68[63],pp68[64],pp68[65],pp68[66],pp68[67],pp68[68],pp68[69],pp69[69],pp70[69],pp71[69],pp72[69],pp73[69],pp74[69],pp75[69],pp76[69],pp77[69],pp78[69],pp79[69]};
    assign in44_2 = {pp89[18],pp88[20],pp87[22],pp86[24],pp85[26],pp84[28],pp83[30],pp82[32],pp81[34],pp80[36],pp79[38],pp78[40],pp77[42],pp76[44],pp75[46],pp74[48],pp73[50],pp72[52],pp71[54],pp70[56],pp69[58],pp69[59],pp69[60],pp69[61],pp69[62],pp69[63],pp69[64],pp69[65],pp69[66],pp69[67],pp69[68],pp70[68],pp71[68],pp72[68],pp73[68],pp74[68],pp75[68],pp76[68],pp77[68],pp78[68],pp79[68],pp80[68]};
    CLA_42 KS_44(s44, c44, in44_1, in44_2);
    wire[39:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp89[19],pp88[21],pp87[23],pp86[25],pp85[27],pp84[29],pp83[31],pp82[33],pp81[35],pp80[37],pp79[39],pp78[41],pp77[43],pp76[45],pp75[47],pp74[49],pp73[51],pp72[53],pp71[55],pp70[57],pp70[58],pp70[59],pp70[60],pp70[61],pp70[62],pp70[63],pp70[64],pp70[65],pp70[66],pp70[67],pp71[67],pp72[67],pp73[67],pp74[67],pp75[67],pp76[67],pp77[67],pp78[67],pp79[67],pp80[67]};
    assign in45_2 = {pp90[18],pp89[20],pp88[22],pp87[24],pp86[26],pp85[28],pp84[30],pp83[32],pp82[34],pp81[36],pp80[38],pp79[40],pp78[42],pp77[44],pp76[46],pp75[48],pp74[50],pp73[52],pp72[54],pp71[56],pp71[57],pp71[58],pp71[59],pp71[60],pp71[61],pp71[62],pp71[63],pp71[64],pp71[65],pp71[66],pp72[66],pp73[66],pp74[66],pp75[66],pp76[66],pp77[66],pp78[66],pp79[66],pp80[66],pp81[66]};
    CLA_40 KS_45(s45, c45, in45_1, in45_2);
    wire[37:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp90[19],pp89[21],pp88[23],pp87[25],pp86[27],pp85[29],pp84[31],pp83[33],pp82[35],pp81[37],pp80[39],pp79[41],pp78[43],pp77[45],pp76[47],pp75[49],pp74[51],pp73[53],pp72[55],pp72[56],pp72[57],pp72[58],pp72[59],pp72[60],pp72[61],pp72[62],pp72[63],pp72[64],pp72[65],pp73[65],pp74[65],pp75[65],pp76[65],pp77[65],pp78[65],pp79[65],pp80[65],pp81[65]};
    assign in46_2 = {pp91[18],pp90[20],pp89[22],pp88[24],pp87[26],pp86[28],pp85[30],pp84[32],pp83[34],pp82[36],pp81[38],pp80[40],pp79[42],pp78[44],pp77[46],pp76[48],pp75[50],pp74[52],pp73[54],pp73[55],pp73[56],pp73[57],pp73[58],pp73[59],pp73[60],pp73[61],pp73[62],pp73[63],pp73[64],pp74[64],pp75[64],pp76[64],pp77[64],pp78[64],pp79[64],pp80[64],pp81[64],pp82[64]};
    CLA_38 KS_46(s46, c46, in46_1, in46_2);
    wire[35:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp91[19],pp90[21],pp89[23],pp88[25],pp87[27],pp86[29],pp85[31],pp84[33],pp83[35],pp82[37],pp81[39],pp80[41],pp79[43],pp78[45],pp77[47],pp76[49],pp75[51],pp74[53],pp74[54],pp74[55],pp74[56],pp74[57],pp74[58],pp74[59],pp74[60],pp74[61],pp74[62],pp74[63],pp75[63],pp76[63],pp77[63],pp78[63],pp79[63],pp80[63],pp81[63],pp82[63]};
    assign in47_2 = {pp92[18],pp91[20],pp90[22],pp89[24],pp88[26],pp87[28],pp86[30],pp85[32],pp84[34],pp83[36],pp82[38],pp81[40],pp80[42],pp79[44],pp78[46],pp77[48],pp76[50],pp75[52],pp75[53],pp75[54],pp75[55],pp75[56],pp75[57],pp75[58],pp75[59],pp75[60],pp75[61],pp75[62],pp76[62],pp77[62],pp78[62],pp79[62],pp80[62],pp81[62],pp82[62],pp83[62]};
    CLA_36 KS_47(s47, c47, in47_1, in47_2);
    wire[33:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp92[19],pp91[21],pp90[23],pp89[25],pp88[27],pp87[29],pp86[31],pp85[33],pp84[35],pp83[37],pp82[39],pp81[41],pp80[43],pp79[45],pp78[47],pp77[49],pp76[51],pp76[52],pp76[53],pp76[54],pp76[55],pp76[56],pp76[57],pp76[58],pp76[59],pp76[60],pp76[61],pp77[61],pp78[61],pp79[61],pp80[61],pp81[61],pp82[61],pp83[61]};
    assign in48_2 = {pp93[18],pp92[20],pp91[22],pp90[24],pp89[26],pp88[28],pp87[30],pp86[32],pp85[34],pp84[36],pp83[38],pp82[40],pp81[42],pp80[44],pp79[46],pp78[48],pp77[50],pp77[51],pp77[52],pp77[53],pp77[54],pp77[55],pp77[56],pp77[57],pp77[58],pp77[59],pp77[60],pp78[60],pp79[60],pp80[60],pp81[60],pp82[60],pp83[60],pp84[60]};
    CLA_34 KS_48(s48, c48, in48_1, in48_2);
    wire[31:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp93[19],pp92[21],pp91[23],pp90[25],pp89[27],pp88[29],pp87[31],pp86[33],pp85[35],pp84[37],pp83[39],pp82[41],pp81[43],pp80[45],pp79[47],pp78[49],pp78[50],pp78[51],pp78[52],pp78[53],pp78[54],pp78[55],pp78[56],pp78[57],pp78[58],pp78[59],pp79[59],pp80[59],pp81[59],pp82[59],pp83[59],pp84[59]};
    assign in49_2 = {pp94[18],pp93[20],pp92[22],pp91[24],pp90[26],pp89[28],pp88[30],pp87[32],pp86[34],pp85[36],pp84[38],pp83[40],pp82[42],pp81[44],pp80[46],pp79[48],pp79[49],pp79[50],pp79[51],pp79[52],pp79[53],pp79[54],pp79[55],pp79[56],pp79[57],pp79[58],pp80[58],pp81[58],pp82[58],pp83[58],pp84[58],pp85[58]};
    CLA_32 KS_49(s49, c49, in49_1, in49_2);
    wire[29:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp94[19],pp93[21],pp92[23],pp91[25],pp90[27],pp89[29],pp88[31],pp87[33],pp86[35],pp85[37],pp84[39],pp83[41],pp82[43],pp81[45],pp80[47],pp80[48],pp80[49],pp80[50],pp80[51],pp80[52],pp80[53],pp80[54],pp80[55],pp80[56],pp80[57],pp81[57],pp82[57],pp83[57],pp84[57],pp85[57]};
    assign in50_2 = {pp95[18],pp94[20],pp93[22],pp92[24],pp91[26],pp90[28],pp89[30],pp88[32],pp87[34],pp86[36],pp85[38],pp84[40],pp83[42],pp82[44],pp81[46],pp81[47],pp81[48],pp81[49],pp81[50],pp81[51],pp81[52],pp81[53],pp81[54],pp81[55],pp81[56],pp82[56],pp83[56],pp84[56],pp85[56],pp86[56]};
    CLA_30 KS_50(s50, c50, in50_1, in50_2);
    wire[27:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp95[19],pp94[21],pp93[23],pp92[25],pp91[27],pp90[29],pp89[31],pp88[33],pp87[35],pp86[37],pp85[39],pp84[41],pp83[43],pp82[45],pp82[46],pp82[47],pp82[48],pp82[49],pp82[50],pp82[51],pp82[52],pp82[53],pp82[54],pp82[55],pp83[55],pp84[55],pp85[55],pp86[55]};
    assign in51_2 = {pp96[18],pp95[20],pp94[22],pp93[24],pp92[26],pp91[28],pp90[30],pp89[32],pp88[34],pp87[36],pp86[38],pp85[40],pp84[42],pp83[44],pp83[45],pp83[46],pp83[47],pp83[48],pp83[49],pp83[50],pp83[51],pp83[52],pp83[53],pp83[54],pp84[54],pp85[54],pp86[54],pp87[54]};
    CLA_28 KS_51(s51, c51, in51_1, in51_2);
    wire[25:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp96[19],pp95[21],pp94[23],pp93[25],pp92[27],pp91[29],pp90[31],pp89[33],pp88[35],pp87[37],pp86[39],pp85[41],pp84[43],pp84[44],pp84[45],pp84[46],pp84[47],pp84[48],pp84[49],pp84[50],pp84[51],pp84[52],pp84[53],pp85[53],pp86[53],pp87[53]};
    assign in52_2 = {pp97[18],pp96[20],pp95[22],pp94[24],pp93[26],pp92[28],pp91[30],pp90[32],pp89[34],pp88[36],pp87[38],pp86[40],pp85[42],pp85[43],pp85[44],pp85[45],pp85[46],pp85[47],pp85[48],pp85[49],pp85[50],pp85[51],pp85[52],pp86[52],pp87[52],pp88[52]};
    CLA_26 KS_52(s52, c52, in52_1, in52_2);
    wire[23:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp97[19],pp96[21],pp95[23],pp94[25],pp93[27],pp92[29],pp91[31],pp90[33],pp89[35],pp88[37],pp87[39],pp86[41],pp86[42],pp86[43],pp86[44],pp86[45],pp86[46],pp86[47],pp86[48],pp86[49],pp86[50],pp86[51],pp87[51],pp88[51]};
    assign in53_2 = {pp98[18],pp97[20],pp96[22],pp95[24],pp94[26],pp93[28],pp92[30],pp91[32],pp90[34],pp89[36],pp88[38],pp87[40],pp87[41],pp87[42],pp87[43],pp87[44],pp87[45],pp87[46],pp87[47],pp87[48],pp87[49],pp87[50],pp88[50],pp89[50]};
    CLA_24 KS_53(s53, c53, in53_1, in53_2);
    wire[21:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp98[19],pp97[21],pp96[23],pp95[25],pp94[27],pp93[29],pp92[31],pp91[33],pp90[35],pp89[37],pp88[39],pp88[40],pp88[41],pp88[42],pp88[43],pp88[44],pp88[45],pp88[46],pp88[47],pp88[48],pp88[49],pp89[49]};
    assign in54_2 = {pp99[18],pp98[20],pp97[22],pp96[24],pp95[26],pp94[28],pp93[30],pp92[32],pp91[34],pp90[36],pp89[38],pp89[39],pp89[40],pp89[41],pp89[42],pp89[43],pp89[44],pp89[45],pp89[46],pp89[47],pp89[48],pp90[48]};
    CLA_22 KS_54(s54, c54, in54_1, in54_2);
    wire[19:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp99[19],pp98[21],pp97[23],pp96[25],pp95[27],pp94[29],pp93[31],pp92[33],pp91[35],pp90[37],pp90[38],pp90[39],pp90[40],pp90[41],pp90[42],pp90[43],pp90[44],pp90[45],pp90[46],pp90[47]};
    assign in55_2 = {pp109[9],pp99[20],pp98[22],pp97[24],pp96[26],pp95[28],pp94[30],pp93[32],pp92[34],pp91[36],pp91[37],pp91[38],pp91[39],pp91[40],pp91[41],pp91[42],pp91[43],pp91[44],pp91[45],pp91[46]};
    CLA_20 KS_55(s55, c55, in55_1, in55_2);
    wire[17:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp110[9],pp99[21],pp98[23],pp97[25],pp96[27],pp95[29],pp94[31],pp93[33],pp92[35],pp92[36],pp92[37],pp92[38],pp92[39],pp92[40],pp92[41],pp92[42],pp92[43],pp92[44]};
    assign in56_2 = {pp111[8],pp111[9],pp99[22],pp98[24],pp97[26],pp96[28],pp95[30],pp94[32],pp93[34],pp93[35],pp93[36],pp93[37],pp93[38],pp93[39],pp93[40],pp93[41],pp93[42],pp93[43]};
    CLA_18 KS_56(s56, c56, in56_1, in56_2);
    wire[15:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp112[8],pp112[9],pp99[23],pp98[25],pp97[27],pp96[29],pp95[31],pp94[33],pp94[34],pp94[35],pp94[36],pp94[37],pp94[38],pp94[39],pp94[40],pp94[41]};
    assign in57_2 = {pp113[7],pp113[8],pp113[9],pp99[24],pp98[26],pp97[28],pp96[30],pp95[32],pp95[33],pp95[34],pp95[35],pp95[36],pp95[37],pp95[38],pp95[39],pp95[40]};
    CLA_16 KS_57(s57, c57, in57_1, in57_2);
    wire[13:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp114[7],pp114[8],pp114[9],pp99[25],pp98[27],pp97[29],pp96[31],pp96[32],pp96[33],pp96[34],pp96[35],pp96[36],pp96[37],pp96[38]};
    assign in58_2 = {pp115[6],pp115[7],pp115[8],pp115[9],pp99[26],pp98[28],pp97[30],pp97[31],pp97[32],pp97[33],pp97[34],pp97[35],pp97[36],pp97[37]};
    CLA_14 KS_58(s58, c58, in58_1, in58_2);
    wire[11:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp116[6],pp116[7],pp116[8],pp116[9],pp99[27],pp98[29],pp98[30],pp98[31],pp98[32],pp98[33],pp98[34],pp98[35]};
    assign in59_2 = {pp117[5],pp117[6],pp117[7],pp117[8],pp117[9],pp99[28],pp99[29],pp99[30],pp99[31],pp99[32],pp99[33],pp99[34]};
    CLA_12 KS_59(s59, c59, in59_1, in59_2);
    wire[9:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp118[5],pp118[6],pp118[7],pp118[8],pp118[9],pp119[9],pp120[9],pp121[9],pp122[9],pp123[9]};
    assign in60_2 = {pp119[4],pp119[5],pp119[6],pp119[7],pp119[8],pp120[8],pp121[8],pp122[8],pp123[8],pp124[8]};
    CLA_10 KS_60(s60, c60, in60_1, in60_2);
    wire[7:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp120[4],pp120[5],pp120[6],pp120[7],pp121[7],pp122[7],pp123[7],pp124[7]};
    assign in61_2 = {pp121[3],pp121[4],pp121[5],pp121[6],pp122[6],pp123[6],pp124[6],pp125[6]};
    CLA_8 KS_61(s61, c61, in61_1, in61_2);
    wire[5:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp122[3],pp122[4],pp122[5],pp123[5],pp124[5],pp125[5]};
    assign in62_2 = {pp123[2],pp123[3],pp123[4],pp124[4],pp125[4],pp126[4]};
    CLA_6 KS_62(s62, c62, in62_1, in62_2);
    wire[3:0] s63, in63_1, in63_2;
    wire c63;
    assign in63_1 = {pp124[2],pp124[3],pp125[3],pp126[3]};
    assign in63_2 = {pp125[1],pp125[2],pp126[2],pp127[2]};
    CLA_4 KS_63(s63, c63, in63_1, in63_2);
    wire[1:0] s64, in64_1, in64_2;
    wire c64;
    assign in64_1 = {pp126[1],pp127[1]};
    assign in64_2 = {pp127[0],s10[55]};
    CLA_2 KS_64(s64, c64, in64_1, in64_2);

    /*Stage 2*/
    wire[191:0] s65, in65_1, in65_2;
    wire c65;
    assign in65_1 = {pp10[22],pp10[23],pp10[24],pp10[25],pp10[26],pp10[27],pp10[28],pp10[29],pp10[30],pp10[31],pp10[32],pp10[33],pp10[34],pp10[35],pp10[36],pp10[37],pp10[38],pp10[39],pp10[40],pp10[41],pp10[42],pp10[43],pp10[44],pp10[45],pp10[46],pp10[47],pp10[48],pp10[49],pp10[50],pp10[51],pp10[52],pp10[53],pp12[52],pp14[51],pp16[50],pp18[49],pp20[48],pp22[47],pp24[46],pp26[45],pp28[44],pp30[43],pp32[42],pp34[41],pp36[40],pp38[39],pp40[38],pp42[37],pp44[36],pp46[35],pp48[34],pp50[33],pp52[32],pp54[31],pp56[30],pp58[29],pp60[28],pp62[27],pp64[26],pp66[25],pp68[24],pp70[23],pp72[22],pp74[21],pp76[20],pp78[19],pp80[18],pp82[17],pp83[17],pp84[17],pp85[17],pp86[17],pp87[17],pp88[17],pp89[17],pp90[17],pp91[17],pp92[17],pp93[17],pp94[17],pp95[17],pp96[17],pp97[17],pp98[17],pp99[17],pp108[9],pp110[8],pp112[7],pp114[6],pp116[5],pp118[4],pp120[3],pp122[2],pp124[1],pp126[0],s10[54],s11[54],s10[56],pp127[3],pp126[5],pp125[7],pp124[9],pp98[36],pp96[39],pp94[42],pp92[45],pp91[47],pp90[49],pp89[51],pp88[53],pp87[55],pp86[57],pp85[59],pp84[61],pp83[63],pp82[65],pp81[67],pp80[69],pp79[71],pp78[73],pp77[75],pp76[77],pp75[79],pp74[81],pp73[83],pp72[85],pp71[87],pp70[89],pp69[91],pp68[93],pp67[95],pp66[97],pp65[99],pp126[39],pp124[42],pp122[45],pp120[48],pp118[51],pp116[54],pp114[57],pp112[60],pp110[63],pp108[66],pp106[69],pp104[72],pp102[75],pp100[78],pp78[101],pp77[103],pp76[105],pp75[107],pp74[109],pp73[111],pp72[113],pp71[115],pp70[117],pp69[119],pp68[121],pp67[123],pp66[125],pp65[127],pp66[127],pp67[127],pp68[127],pp69[127],pp70[127],pp71[127],pp72[127],pp100[100],pp100[101],pp100[102],pp100[103],pp100[104],pp100[105],pp100[106],pp100[107],pp100[108],pp100[109],pp100[110],pp100[111],pp100[112],pp100[113],pp100[114],pp100[115],pp100[116],pp100[117],pp100[118],pp100[119],pp100[120],pp100[121],pp100[122],pp100[123]};
    assign in65_2 = {pp11[21],pp11[22],pp11[23],pp11[24],pp11[25],pp11[26],pp11[27],pp11[28],pp11[29],pp11[30],pp11[31],pp11[32],pp11[33],pp11[34],pp11[35],pp11[36],pp11[37],pp11[38],pp11[39],pp11[40],pp11[41],pp11[42],pp11[43],pp11[44],pp11[45],pp11[46],pp11[47],pp11[48],pp11[49],pp11[50],pp11[51],pp11[52],pp13[51],pp15[50],pp17[49],pp19[48],pp21[47],pp23[46],pp25[45],pp27[44],pp29[43],pp31[42],pp33[41],pp35[40],pp37[39],pp39[38],pp41[37],pp43[36],pp45[35],pp47[34],pp49[33],pp51[32],pp53[31],pp55[30],pp57[29],pp59[28],pp61[27],pp63[26],pp65[25],pp67[24],pp69[23],pp71[22],pp73[21],pp75[20],pp77[19],pp79[18],pp81[17],pp83[16],pp84[16],pp85[16],pp86[16],pp87[16],pp88[16],pp89[16],pp90[16],pp91[16],pp92[16],pp93[16],pp94[16],pp95[16],pp96[16],pp97[16],pp98[16],pp99[16],pp107[9],pp109[8],pp111[7],pp113[6],pp115[5],pp117[4],pp119[3],pp121[2],pp123[1],pp125[0],s10[53],s11[53],s12[53],s11[55],s10[57],pp127[4],pp126[6],pp125[8],pp99[35],pp97[38],pp95[41],pp93[44],pp92[46],pp91[48],pp90[50],pp89[52],pp88[54],pp87[56],pp86[58],pp85[60],pp84[62],pp83[64],pp82[66],pp81[68],pp80[70],pp79[72],pp78[74],pp77[76],pp76[78],pp75[80],pp74[82],pp73[84],pp72[86],pp71[88],pp70[90],pp69[92],pp68[94],pp67[96],pp66[98],pp127[38],pp125[41],pp123[44],pp121[47],pp119[50],pp117[53],pp115[56],pp113[59],pp111[62],pp109[65],pp107[68],pp105[71],pp103[74],pp101[77],pp79[100],pp78[102],pp77[104],pp76[106],pp75[108],pp74[110],pp73[112],pp72[114],pp71[116],pp70[118],pp69[120],pp68[122],pp67[124],pp66[126],pp67[126],pp68[126],pp69[126],pp70[126],pp71[126],pp72[126],pp73[126],pp73[127],pp101[100],pp101[101],pp101[102],pp101[103],pp101[104],pp101[105],pp101[106],pp101[107],pp101[108],pp101[109],pp101[110],pp101[111],pp101[112],pp101[113],pp101[114],pp101[115],pp101[116],pp101[117],pp101[118],pp101[119],pp101[120],pp101[121],pp101[122]};
    CLA_192 KS_65(s65, c65, in65_1, in65_2);
    wire[189:0] s66, in66_1, in66_2;
    wire c66;
    assign in66_1 = {pp12[21],pp12[22],pp12[23],pp12[24],pp12[25],pp12[26],pp12[27],pp12[28],pp12[29],pp12[30],pp12[31],pp12[32],pp12[33],pp12[34],pp12[35],pp12[36],pp12[37],pp12[38],pp12[39],pp12[40],pp12[41],pp12[42],pp12[43],pp12[44],pp12[45],pp12[46],pp12[47],pp12[48],pp12[49],pp12[50],pp12[51],pp14[50],pp16[49],pp18[48],pp20[47],pp22[46],pp24[45],pp26[44],pp28[43],pp30[42],pp32[41],pp34[40],pp36[39],pp38[38],pp40[37],pp42[36],pp44[35],pp46[34],pp48[33],pp50[32],pp52[31],pp54[30],pp56[29],pp58[28],pp60[27],pp62[26],pp64[25],pp66[24],pp68[23],pp70[22],pp72[21],pp74[20],pp76[19],pp78[18],pp80[17],pp82[16],pp84[15],pp85[15],pp86[15],pp87[15],pp88[15],pp89[15],pp90[15],pp91[15],pp92[15],pp93[15],pp94[15],pp95[15],pp96[15],pp97[15],pp98[15],pp99[15],pp106[9],pp108[8],pp110[7],pp112[6],pp114[5],pp116[4],pp118[3],pp120[2],pp122[1],pp124[0],s10[52],s11[52],s12[52],s13[52],s12[54],s11[56],s10[58],pp127[5],pp126[7],pp125[9],pp98[37],pp96[40],pp94[43],pp93[45],pp92[47],pp91[49],pp90[51],pp89[53],pp88[55],pp87[57],pp86[59],pp85[61],pp84[63],pp83[65],pp82[67],pp81[69],pp80[71],pp79[73],pp78[75],pp77[77],pp76[79],pp75[81],pp74[83],pp73[85],pp72[87],pp71[89],pp70[91],pp69[93],pp68[95],pp67[97],pp66[99],pp126[40],pp124[43],pp122[46],pp120[49],pp118[52],pp116[55],pp114[58],pp112[61],pp110[64],pp108[67],pp106[70],pp104[73],pp102[76],pp100[79],pp79[101],pp78[103],pp77[105],pp76[107],pp75[109],pp74[111],pp73[113],pp72[115],pp71[117],pp70[119],pp69[121],pp68[123],pp67[125],pp68[125],pp69[125],pp70[125],pp71[125],pp72[125],pp73[125],pp74[125],pp74[126],pp74[127],pp102[100],pp102[101],pp102[102],pp102[103],pp102[104],pp102[105],pp102[106],pp102[107],pp102[108],pp102[109],pp102[110],pp102[111],pp102[112],pp102[113],pp102[114],pp102[115],pp102[116],pp102[117],pp102[118],pp102[119],pp102[120]};
    assign in66_2 = {pp13[20],pp13[21],pp13[22],pp13[23],pp13[24],pp13[25],pp13[26],pp13[27],pp13[28],pp13[29],pp13[30],pp13[31],pp13[32],pp13[33],pp13[34],pp13[35],pp13[36],pp13[37],pp13[38],pp13[39],pp13[40],pp13[41],pp13[42],pp13[43],pp13[44],pp13[45],pp13[46],pp13[47],pp13[48],pp13[49],pp13[50],pp15[49],pp17[48],pp19[47],pp21[46],pp23[45],pp25[44],pp27[43],pp29[42],pp31[41],pp33[40],pp35[39],pp37[38],pp39[37],pp41[36],pp43[35],pp45[34],pp47[33],pp49[32],pp51[31],pp53[30],pp55[29],pp57[28],pp59[27],pp61[26],pp63[25],pp65[24],pp67[23],pp69[22],pp71[21],pp73[20],pp75[19],pp77[18],pp79[17],pp81[16],pp83[15],pp85[14],pp86[14],pp87[14],pp88[14],pp89[14],pp90[14],pp91[14],pp92[14],pp93[14],pp94[14],pp95[14],pp96[14],pp97[14],pp98[14],pp99[14],pp105[9],pp107[8],pp109[7],pp111[6],pp113[5],pp115[4],pp117[3],pp119[2],pp121[1],pp123[0],s10[51],s11[51],s12[51],s13[51],s14[51],s13[53],s12[55],s11[57],s65[100],pp127[6],pp126[8],pp99[36],pp97[39],pp95[42],pp94[44],pp93[46],pp92[48],pp91[50],pp90[52],pp89[54],pp88[56],pp87[58],pp86[60],pp85[62],pp84[64],pp83[66],pp82[68],pp81[70],pp80[72],pp79[74],pp78[76],pp77[78],pp76[80],pp75[82],pp74[84],pp73[86],pp72[88],pp71[90],pp70[92],pp69[94],pp68[96],pp67[98],pp127[39],pp125[42],pp123[45],pp121[48],pp119[51],pp117[54],pp115[57],pp113[60],pp111[63],pp109[66],pp107[69],pp105[72],pp103[75],pp101[78],pp80[100],pp79[102],pp78[104],pp77[106],pp76[108],pp75[110],pp74[112],pp73[114],pp72[116],pp71[118],pp70[120],pp69[122],pp68[124],pp69[124],pp70[124],pp71[124],pp72[124],pp73[124],pp74[124],pp75[124],pp75[125],pp75[126],pp75[127],pp103[100],pp103[101],pp103[102],pp103[103],pp103[104],pp103[105],pp103[106],pp103[107],pp103[108],pp103[109],pp103[110],pp103[111],pp103[112],pp103[113],pp103[114],pp103[115],pp103[116],pp103[117],pp103[118],pp103[119]};
    CLA_190 KS_66(s66, c66, in66_1, in66_2);
    wire[187:0] s67, in67_1, in67_2;
    wire c67;
    assign in67_1 = {pp14[20],pp14[21],pp14[22],pp14[23],pp14[24],pp14[25],pp14[26],pp14[27],pp14[28],pp14[29],pp14[30],pp14[31],pp14[32],pp14[33],pp14[34],pp14[35],pp14[36],pp14[37],pp14[38],pp14[39],pp14[40],pp14[41],pp14[42],pp14[43],pp14[44],pp14[45],pp14[46],pp14[47],pp14[48],pp14[49],pp16[48],pp18[47],pp20[46],pp22[45],pp24[44],pp26[43],pp28[42],pp30[41],pp32[40],pp34[39],pp36[38],pp38[37],pp40[36],pp42[35],pp44[34],pp46[33],pp48[32],pp50[31],pp52[30],pp54[29],pp56[28],pp58[27],pp60[26],pp62[25],pp64[24],pp66[23],pp68[22],pp70[21],pp72[20],pp74[19],pp76[18],pp78[17],pp80[16],pp82[15],pp84[14],pp86[13],pp87[13],pp88[13],pp89[13],pp90[13],pp91[13],pp92[13],pp93[13],pp94[13],pp95[13],pp96[13],pp97[13],pp98[13],pp99[13],pp104[9],pp106[8],pp108[7],pp110[6],pp112[5],pp114[4],pp116[3],pp118[2],pp120[1],pp122[0],s10[50],s11[50],s12[50],s13[50],s14[50],s15[50],s14[52],s13[54],s12[56],s10[59],s65[101],pp127[7],pp126[9],pp98[38],pp96[41],pp95[43],pp94[45],pp93[47],pp92[49],pp91[51],pp90[53],pp89[55],pp88[57],pp87[59],pp86[61],pp85[63],pp84[65],pp83[67],pp82[69],pp81[71],pp80[73],pp79[75],pp78[77],pp77[79],pp76[81],pp75[83],pp74[85],pp73[87],pp72[89],pp71[91],pp70[93],pp69[95],pp68[97],pp67[99],pp126[41],pp124[44],pp122[47],pp120[50],pp118[53],pp116[56],pp114[59],pp112[62],pp110[65],pp108[68],pp106[71],pp104[74],pp102[77],pp100[80],pp80[101],pp79[103],pp78[105],pp77[107],pp76[109],pp75[111],pp74[113],pp73[115],pp72[117],pp71[119],pp70[121],pp69[123],pp70[123],pp71[123],pp72[123],pp73[123],pp74[123],pp75[123],pp76[123],pp76[124],pp76[125],pp76[126],pp76[127],pp104[100],pp104[101],pp104[102],pp104[103],pp104[104],pp104[105],pp104[106],pp104[107],pp104[108],pp104[109],pp104[110],pp104[111],pp104[112],pp104[113],pp104[114],pp104[115],pp104[116],pp104[117]};
    assign in67_2 = {pp15[19],pp15[20],pp15[21],pp15[22],pp15[23],pp15[24],pp15[25],pp15[26],pp15[27],pp15[28],pp15[29],pp15[30],pp15[31],pp15[32],pp15[33],pp15[34],pp15[35],pp15[36],pp15[37],pp15[38],pp15[39],pp15[40],pp15[41],pp15[42],pp15[43],pp15[44],pp15[45],pp15[46],pp15[47],pp15[48],pp17[47],pp19[46],pp21[45],pp23[44],pp25[43],pp27[42],pp29[41],pp31[40],pp33[39],pp35[38],pp37[37],pp39[36],pp41[35],pp43[34],pp45[33],pp47[32],pp49[31],pp51[30],pp53[29],pp55[28],pp57[27],pp59[26],pp61[25],pp63[24],pp65[23],pp67[22],pp69[21],pp71[20],pp73[19],pp75[18],pp77[17],pp79[16],pp81[15],pp83[14],pp85[13],pp87[12],pp88[12],pp89[12],pp90[12],pp91[12],pp92[12],pp93[12],pp94[12],pp95[12],pp96[12],pp97[12],pp98[12],pp99[12],pp103[9],pp105[8],pp107[7],pp109[6],pp111[5],pp113[4],pp115[3],pp117[2],pp119[1],pp121[0],s10[49],s11[49],s12[49],s13[49],s14[49],s15[49],s16[49],s15[51],s14[53],s13[55],s11[58],s66[100],s65[102],pp127[8],pp99[37],pp97[40],pp96[42],pp95[44],pp94[46],pp93[48],pp92[50],pp91[52],pp90[54],pp89[56],pp88[58],pp87[60],pp86[62],pp85[64],pp84[66],pp83[68],pp82[70],pp81[72],pp80[74],pp79[76],pp78[78],pp77[80],pp76[82],pp75[84],pp74[86],pp73[88],pp72[90],pp71[92],pp70[94],pp69[96],pp68[98],pp127[40],pp125[43],pp123[46],pp121[49],pp119[52],pp117[55],pp115[58],pp113[61],pp111[64],pp109[67],pp107[70],pp105[73],pp103[76],pp101[79],pp81[100],pp80[102],pp79[104],pp78[106],pp77[108],pp76[110],pp75[112],pp74[114],pp73[116],pp72[118],pp71[120],pp70[122],pp71[122],pp72[122],pp73[122],pp74[122],pp75[122],pp76[122],pp77[122],pp77[123],pp77[124],pp77[125],pp77[126],pp77[127],pp105[100],pp105[101],pp105[102],pp105[103],pp105[104],pp105[105],pp105[106],pp105[107],pp105[108],pp105[109],pp105[110],pp105[111],pp105[112],pp105[113],pp105[114],pp105[115],pp105[116]};
    CLA_188 KS_67(s67, c67, in67_1, in67_2);
    wire[185:0] s68, in68_1, in68_2;
    wire c68;
    assign in68_1 = {pp16[19],pp16[20],pp16[21],pp16[22],pp16[23],pp16[24],pp16[25],pp16[26],pp16[27],pp16[28],pp16[29],pp16[30],pp16[31],pp16[32],pp16[33],pp16[34],pp16[35],pp16[36],pp16[37],pp16[38],pp16[39],pp16[40],pp16[41],pp16[42],pp16[43],pp16[44],pp16[45],pp16[46],pp16[47],pp18[46],pp20[45],pp22[44],pp24[43],pp26[42],pp28[41],pp30[40],pp32[39],pp34[38],pp36[37],pp38[36],pp40[35],pp42[34],pp44[33],pp46[32],pp48[31],pp50[30],pp52[29],pp54[28],pp56[27],pp58[26],pp60[25],pp62[24],pp64[23],pp66[22],pp68[21],pp70[20],pp72[19],pp74[18],pp76[17],pp78[16],pp80[15],pp82[14],pp84[13],pp86[12],pp88[11],pp89[11],pp90[11],pp91[11],pp92[11],pp93[11],pp94[11],pp95[11],pp96[11],pp97[11],pp98[11],pp99[11],pp102[9],pp104[8],pp106[7],pp108[6],pp110[5],pp112[4],pp114[3],pp116[2],pp118[1],pp120[0],s10[48],s11[48],s12[48],s13[48],s14[48],s15[48],s16[48],s17[48],s16[50],s15[52],s14[54],s12[57],s10[60],s66[101],s65[103],pp127[9],pp98[39],pp97[41],pp96[43],pp95[45],pp94[47],pp93[49],pp92[51],pp91[53],pp90[55],pp89[57],pp88[59],pp87[61],pp86[63],pp85[65],pp84[67],pp83[69],pp82[71],pp81[73],pp80[75],pp79[77],pp78[79],pp77[81],pp76[83],pp75[85],pp74[87],pp73[89],pp72[91],pp71[93],pp70[95],pp69[97],pp68[99],pp126[42],pp124[45],pp122[48],pp120[51],pp118[54],pp116[57],pp114[60],pp112[63],pp110[66],pp108[69],pp106[72],pp104[75],pp102[78],pp100[81],pp81[101],pp80[103],pp79[105],pp78[107],pp77[109],pp76[111],pp75[113],pp74[115],pp73[117],pp72[119],pp71[121],pp72[121],pp73[121],pp74[121],pp75[121],pp76[121],pp77[121],pp78[121],pp78[122],pp78[123],pp78[124],pp78[125],pp78[126],pp78[127],pp106[100],pp106[101],pp106[102],pp106[103],pp106[104],pp106[105],pp106[106],pp106[107],pp106[108],pp106[109],pp106[110],pp106[111],pp106[112],pp106[113],pp106[114]};
    assign in68_2 = {pp17[18],pp17[19],pp17[20],pp17[21],pp17[22],pp17[23],pp17[24],pp17[25],pp17[26],pp17[27],pp17[28],pp17[29],pp17[30],pp17[31],pp17[32],pp17[33],pp17[34],pp17[35],pp17[36],pp17[37],pp17[38],pp17[39],pp17[40],pp17[41],pp17[42],pp17[43],pp17[44],pp17[45],pp17[46],pp19[45],pp21[44],pp23[43],pp25[42],pp27[41],pp29[40],pp31[39],pp33[38],pp35[37],pp37[36],pp39[35],pp41[34],pp43[33],pp45[32],pp47[31],pp49[30],pp51[29],pp53[28],pp55[27],pp57[26],pp59[25],pp61[24],pp63[23],pp65[22],pp67[21],pp69[20],pp71[19],pp73[18],pp75[17],pp77[16],pp79[15],pp81[14],pp83[13],pp85[12],pp87[11],pp89[10],pp90[10],pp91[10],pp92[10],pp93[10],pp94[10],pp95[10],pp96[10],pp97[10],pp98[10],pp99[10],pp101[9],pp103[8],pp105[7],pp107[6],pp109[5],pp111[4],pp113[3],pp115[2],pp117[1],pp119[0],s10[47],s11[47],s12[47],s13[47],s14[47],s15[47],s16[47],s17[47],s18[47],s17[49],s16[51],s15[53],s13[56],s11[59],s67[100],s66[102],s65[104],pp99[38],pp98[40],pp97[42],pp96[44],pp95[46],pp94[48],pp93[50],pp92[52],pp91[54],pp90[56],pp89[58],pp88[60],pp87[62],pp86[64],pp85[66],pp84[68],pp83[70],pp82[72],pp81[74],pp80[76],pp79[78],pp78[80],pp77[82],pp76[84],pp75[86],pp74[88],pp73[90],pp72[92],pp71[94],pp70[96],pp69[98],pp127[41],pp125[44],pp123[47],pp121[50],pp119[53],pp117[56],pp115[59],pp113[62],pp111[65],pp109[68],pp107[71],pp105[74],pp103[77],pp101[80],pp82[100],pp81[102],pp80[104],pp79[106],pp78[108],pp77[110],pp76[112],pp75[114],pp74[116],pp73[118],pp72[120],pp73[120],pp74[120],pp75[120],pp76[120],pp77[120],pp78[120],pp79[120],pp79[121],pp79[122],pp79[123],pp79[124],pp79[125],pp79[126],pp79[127],pp107[100],pp107[101],pp107[102],pp107[103],pp107[104],pp107[105],pp107[106],pp107[107],pp107[108],pp107[109],pp107[110],pp107[111],pp107[112],pp107[113]};
    CLA_186 KS_68(s68, c68, in68_1, in68_2);
    wire[183:0] s69, in69_1, in69_2;
    wire c69;
    assign in69_1 = {pp18[18],pp18[19],pp18[20],pp18[21],pp18[22],pp18[23],pp18[24],pp18[25],pp18[26],pp18[27],pp18[28],pp18[29],pp18[30],pp18[31],pp18[32],pp18[33],pp18[34],pp18[35],pp18[36],pp18[37],pp18[38],pp18[39],pp18[40],pp18[41],pp18[42],pp18[43],pp18[44],pp18[45],pp20[44],pp22[43],pp24[42],pp26[41],pp28[40],pp30[39],pp32[38],pp34[37],pp36[36],pp38[35],pp40[34],pp42[33],pp44[32],pp46[31],pp48[30],pp50[29],pp52[28],pp54[27],pp56[26],pp58[25],pp60[24],pp62[23],pp64[22],pp66[21],pp68[20],pp70[19],pp72[18],pp74[17],pp76[16],pp78[15],pp80[14],pp82[13],pp84[12],pp86[11],pp88[10],pp0[99],pp100[0],pp100[1],pp100[2],pp100[3],pp100[4],pp100[5],pp100[6],pp100[7],pp100[8],pp100[9],pp102[8],pp104[7],pp106[6],pp108[5],pp110[4],pp112[3],pp114[2],pp116[1],pp118[0],s10[46],s11[46],s12[46],s13[46],s14[46],s15[46],s16[46],s17[46],s18[46],s19[46],s18[48],s17[50],s16[52],s14[55],s12[58],s10[61],s67[101],s66[103],s65[105],pp99[39],pp98[41],pp97[43],pp96[45],pp95[47],pp94[49],pp93[51],pp92[53],pp91[55],pp90[57],pp89[59],pp88[61],pp87[63],pp86[65],pp85[67],pp84[69],pp83[71],pp82[73],pp81[75],pp80[77],pp79[79],pp78[81],pp77[83],pp76[85],pp75[87],pp74[89],pp73[91],pp72[93],pp71[95],pp70[97],pp69[99],pp126[43],pp124[46],pp122[49],pp120[52],pp118[55],pp116[58],pp114[61],pp112[64],pp110[67],pp108[70],pp106[73],pp104[76],pp102[79],pp100[82],pp82[101],pp81[103],pp80[105],pp79[107],pp78[109],pp77[111],pp76[113],pp75[115],pp74[117],pp73[119],pp74[119],pp75[119],pp76[119],pp77[119],pp78[119],pp79[119],pp80[119],pp80[120],pp80[121],pp80[122],pp80[123],pp80[124],pp80[125],pp80[126],pp80[127],pp108[100],pp108[101],pp108[102],pp108[103],pp108[104],pp108[105],pp108[106],pp108[107],pp108[108],pp108[109],pp108[110],pp108[111]};
    assign in69_2 = {pp19[17],pp19[18],pp19[19],pp19[20],pp19[21],pp19[22],pp19[23],pp19[24],pp19[25],pp19[26],pp19[27],pp19[28],pp19[29],pp19[30],pp19[31],pp19[32],pp19[33],pp19[34],pp19[35],pp19[36],pp19[37],pp19[38],pp19[39],pp19[40],pp19[41],pp19[42],pp19[43],pp19[44],pp21[43],pp23[42],pp25[41],pp27[40],pp29[39],pp31[38],pp33[37],pp35[36],pp37[35],pp39[34],pp41[33],pp43[32],pp45[31],pp47[30],pp49[29],pp51[28],pp53[27],pp55[26],pp57[25],pp59[24],pp61[23],pp63[22],pp65[21],pp67[20],pp69[19],pp71[18],pp73[17],pp75[16],pp77[15],pp79[14],pp81[13],pp83[12],pp85[11],pp87[10],pp0[98],pp1[98],pp1[99],pp101[0],pp101[1],pp101[2],pp101[3],pp101[4],pp101[5],pp101[6],pp101[7],pp101[8],pp103[7],pp105[6],pp107[5],pp109[4],pp111[3],pp113[2],pp115[1],pp117[0],s10[45],s11[45],s12[45],s13[45],s14[45],s15[45],s16[45],s17[45],s18[45],s19[45],s20[45],s19[47],s18[49],s17[51],s15[54],s13[57],s11[60],s68[100],s67[102],s66[104],s65[106],pp99[40],pp98[42],pp97[44],pp96[46],pp95[48],pp94[50],pp93[52],pp92[54],pp91[56],pp90[58],pp89[60],pp88[62],pp87[64],pp86[66],pp85[68],pp84[70],pp83[72],pp82[74],pp81[76],pp80[78],pp79[80],pp78[82],pp77[84],pp76[86],pp75[88],pp74[90],pp73[92],pp72[94],pp71[96],pp70[98],pp127[42],pp125[45],pp123[48],pp121[51],pp119[54],pp117[57],pp115[60],pp113[63],pp111[66],pp109[69],pp107[72],pp105[75],pp103[78],pp101[81],pp83[100],pp82[102],pp81[104],pp80[106],pp79[108],pp78[110],pp77[112],pp76[114],pp75[116],pp74[118],pp75[118],pp76[118],pp77[118],pp78[118],pp79[118],pp80[118],pp81[118],pp81[119],pp81[120],pp81[121],pp81[122],pp81[123],pp81[124],pp81[125],pp81[126],pp81[127],pp109[100],pp109[101],pp109[102],pp109[103],pp109[104],pp109[105],pp109[106],pp109[107],pp109[108],pp109[109],pp109[110]};
    CLA_184 KS_69(s69, c69, in69_1, in69_2);
    wire[181:0] s70, in70_1, in70_2;
    wire c70;
    assign in70_1 = {pp20[17],pp20[18],pp20[19],pp20[20],pp20[21],pp20[22],pp20[23],pp20[24],pp20[25],pp20[26],pp20[27],pp20[28],pp20[29],pp20[30],pp20[31],pp20[32],pp20[33],pp20[34],pp20[35],pp20[36],pp20[37],pp20[38],pp20[39],pp20[40],pp20[41],pp20[42],pp20[43],pp22[42],pp24[41],pp26[40],pp28[39],pp30[38],pp32[37],pp34[36],pp36[35],pp38[34],pp40[33],pp42[32],pp44[31],pp46[30],pp48[29],pp50[28],pp52[27],pp54[26],pp56[25],pp58[24],pp60[23],pp62[22],pp64[21],pp66[20],pp68[19],pp70[18],pp72[17],pp74[16],pp76[15],pp78[14],pp80[13],pp82[12],pp84[11],pp86[10],pp0[97],pp1[97],pp2[97],pp2[98],pp2[99],pp102[0],pp102[1],pp102[2],pp102[3],pp102[4],pp102[5],pp102[6],pp102[7],pp104[6],pp106[5],pp108[4],pp110[3],pp112[2],pp114[1],pp116[0],s10[44],s11[44],s12[44],s13[44],s14[44],s15[44],s16[44],s17[44],s18[44],s19[44],s20[44],s21[44],s20[46],s19[48],s18[50],s16[53],s14[56],s12[59],s10[62],s68[101],s67[103],s66[105],s65[107],pp99[41],pp98[43],pp97[45],pp96[47],pp95[49],pp94[51],pp93[53],pp92[55],pp91[57],pp90[59],pp89[61],pp88[63],pp87[65],pp86[67],pp85[69],pp84[71],pp83[73],pp82[75],pp81[77],pp80[79],pp79[81],pp78[83],pp77[85],pp76[87],pp75[89],pp74[91],pp73[93],pp72[95],pp71[97],pp70[99],pp126[44],pp124[47],pp122[50],pp120[53],pp118[56],pp116[59],pp114[62],pp112[65],pp110[68],pp108[71],pp106[74],pp104[77],pp102[80],pp100[83],pp83[101],pp82[103],pp81[105],pp80[107],pp79[109],pp78[111],pp77[113],pp76[115],pp75[117],pp76[117],pp77[117],pp78[117],pp79[117],pp80[117],pp81[117],pp82[117],pp82[118],pp82[119],pp82[120],pp82[121],pp82[122],pp82[123],pp82[124],pp82[125],pp82[126],pp82[127],pp110[100],pp110[101],pp110[102],pp110[103],pp110[104],pp110[105],pp110[106],pp110[107],pp110[108]};
    assign in70_2 = {pp21[16],pp21[17],pp21[18],pp21[19],pp21[20],pp21[21],pp21[22],pp21[23],pp21[24],pp21[25],pp21[26],pp21[27],pp21[28],pp21[29],pp21[30],pp21[31],pp21[32],pp21[33],pp21[34],pp21[35],pp21[36],pp21[37],pp21[38],pp21[39],pp21[40],pp21[41],pp21[42],pp23[41],pp25[40],pp27[39],pp29[38],pp31[37],pp33[36],pp35[35],pp37[34],pp39[33],pp41[32],pp43[31],pp45[30],pp47[29],pp49[28],pp51[27],pp53[26],pp55[25],pp57[24],pp59[23],pp61[22],pp63[21],pp65[20],pp67[19],pp69[18],pp71[17],pp73[16],pp75[15],pp77[14],pp79[13],pp81[12],pp83[11],pp85[10],pp0[96],pp1[96],pp2[96],pp3[96],pp3[97],pp3[98],pp3[99],pp103[0],pp103[1],pp103[2],pp103[3],pp103[4],pp103[5],pp103[6],pp105[5],pp107[4],pp109[3],pp111[2],pp113[1],pp115[0],s10[43],s11[43],s12[43],s13[43],s14[43],s15[43],s16[43],s17[43],s18[43],s19[43],s20[43],s21[43],s22[43],s21[45],s20[47],s19[49],s17[52],s15[55],s13[58],s11[61],s69[100],s68[102],s67[104],s66[106],s65[108],pp99[42],pp98[44],pp97[46],pp96[48],pp95[50],pp94[52],pp93[54],pp92[56],pp91[58],pp90[60],pp89[62],pp88[64],pp87[66],pp86[68],pp85[70],pp84[72],pp83[74],pp82[76],pp81[78],pp80[80],pp79[82],pp78[84],pp77[86],pp76[88],pp75[90],pp74[92],pp73[94],pp72[96],pp71[98],pp127[43],pp125[46],pp123[49],pp121[52],pp119[55],pp117[58],pp115[61],pp113[64],pp111[67],pp109[70],pp107[73],pp105[76],pp103[79],pp101[82],pp84[100],pp83[102],pp82[104],pp81[106],pp80[108],pp79[110],pp78[112],pp77[114],pp76[116],pp77[116],pp78[116],pp79[116],pp80[116],pp81[116],pp82[116],pp83[116],pp83[117],pp83[118],pp83[119],pp83[120],pp83[121],pp83[122],pp83[123],pp83[124],pp83[125],pp83[126],pp83[127],pp111[100],pp111[101],pp111[102],pp111[103],pp111[104],pp111[105],pp111[106],pp111[107]};
    CLA_182 KS_70(s70, c70, in70_1, in70_2);
    wire[179:0] s71, in71_1, in71_2;
    wire c71;
    assign in71_1 = {pp22[16],pp22[17],pp22[18],pp22[19],pp22[20],pp22[21],pp22[22],pp22[23],pp22[24],pp22[25],pp22[26],pp22[27],pp22[28],pp22[29],pp22[30],pp22[31],pp22[32],pp22[33],pp22[34],pp22[35],pp22[36],pp22[37],pp22[38],pp22[39],pp22[40],pp22[41],pp24[40],pp26[39],pp28[38],pp30[37],pp32[36],pp34[35],pp36[34],pp38[33],pp40[32],pp42[31],pp44[30],pp46[29],pp48[28],pp50[27],pp52[26],pp54[25],pp56[24],pp58[23],pp60[22],pp62[21],pp64[20],pp66[19],pp68[18],pp70[17],pp72[16],pp74[15],pp76[14],pp78[13],pp80[12],pp82[11],pp84[10],pp0[95],pp1[95],pp2[95],pp3[95],pp4[95],pp4[96],pp4[97],pp4[98],pp4[99],pp104[0],pp104[1],pp104[2],pp104[3],pp104[4],pp104[5],pp106[4],pp108[3],pp110[2],pp112[1],pp114[0],s10[42],s11[42],s12[42],s13[42],s14[42],s15[42],s16[42],s17[42],s18[42],s19[42],s20[42],s21[42],s22[42],s23[42],s22[44],s21[46],s20[48],s18[51],s16[54],s14[57],s12[60],s10[63],s69[101],s68[103],s67[105],s66[107],s65[109],pp99[43],pp98[45],pp97[47],pp96[49],pp95[51],pp94[53],pp93[55],pp92[57],pp91[59],pp90[61],pp89[63],pp88[65],pp87[67],pp86[69],pp85[71],pp84[73],pp83[75],pp82[77],pp81[79],pp80[81],pp79[83],pp78[85],pp77[87],pp76[89],pp75[91],pp74[93],pp73[95],pp72[97],pp71[99],pp126[45],pp124[48],pp122[51],pp120[54],pp118[57],pp116[60],pp114[63],pp112[66],pp110[69],pp108[72],pp106[75],pp104[78],pp102[81],pp100[84],pp84[101],pp83[103],pp82[105],pp81[107],pp80[109],pp79[111],pp78[113],pp77[115],pp78[115],pp79[115],pp80[115],pp81[115],pp82[115],pp83[115],pp84[115],pp84[116],pp84[117],pp84[118],pp84[119],pp84[120],pp84[121],pp84[122],pp84[123],pp84[124],pp84[125],pp84[126],pp84[127],pp112[100],pp112[101],pp112[102],pp112[103],pp112[104],pp112[105]};
    assign in71_2 = {pp23[15],pp23[16],pp23[17],pp23[18],pp23[19],pp23[20],pp23[21],pp23[22],pp23[23],pp23[24],pp23[25],pp23[26],pp23[27],pp23[28],pp23[29],pp23[30],pp23[31],pp23[32],pp23[33],pp23[34],pp23[35],pp23[36],pp23[37],pp23[38],pp23[39],pp23[40],pp25[39],pp27[38],pp29[37],pp31[36],pp33[35],pp35[34],pp37[33],pp39[32],pp41[31],pp43[30],pp45[29],pp47[28],pp49[27],pp51[26],pp53[25],pp55[24],pp57[23],pp59[22],pp61[21],pp63[20],pp65[19],pp67[18],pp69[17],pp71[16],pp73[15],pp75[14],pp77[13],pp79[12],pp81[11],pp83[10],pp0[94],pp1[94],pp2[94],pp3[94],pp4[94],pp5[94],pp5[95],pp5[96],pp5[97],pp5[98],pp5[99],pp105[0],pp105[1],pp105[2],pp105[3],pp105[4],pp107[3],pp109[2],pp111[1],pp113[0],s10[41],s11[41],s12[41],s13[41],s14[41],s15[41],s16[41],s17[41],s18[41],s19[41],s20[41],s21[41],s22[41],s23[41],s24[41],s23[43],s22[45],s21[47],s19[50],s17[53],s15[56],s13[59],s11[62],s70[100],s69[102],s68[104],s67[106],s66[108],s65[110],pp99[44],pp98[46],pp97[48],pp96[50],pp95[52],pp94[54],pp93[56],pp92[58],pp91[60],pp90[62],pp89[64],pp88[66],pp87[68],pp86[70],pp85[72],pp84[74],pp83[76],pp82[78],pp81[80],pp80[82],pp79[84],pp78[86],pp77[88],pp76[90],pp75[92],pp74[94],pp73[96],pp72[98],pp127[44],pp125[47],pp123[50],pp121[53],pp119[56],pp117[59],pp115[62],pp113[65],pp111[68],pp109[71],pp107[74],pp105[77],pp103[80],pp101[83],pp85[100],pp84[102],pp83[104],pp82[106],pp81[108],pp80[110],pp79[112],pp78[114],pp79[114],pp80[114],pp81[114],pp82[114],pp83[114],pp84[114],pp85[114],pp85[115],pp85[116],pp85[117],pp85[118],pp85[119],pp85[120],pp85[121],pp85[122],pp85[123],pp85[124],pp85[125],pp85[126],pp85[127],pp113[100],pp113[101],pp113[102],pp113[103],pp113[104]};
    CLA_180 KS_71(s71, c71, in71_1, in71_2);
    wire[177:0] s72, in72_1, in72_2;
    wire c72;
    assign in72_1 = {pp24[15],pp24[16],pp24[17],pp24[18],pp24[19],pp24[20],pp24[21],pp24[22],pp24[23],pp24[24],pp24[25],pp24[26],pp24[27],pp24[28],pp24[29],pp24[30],pp24[31],pp24[32],pp24[33],pp24[34],pp24[35],pp24[36],pp24[37],pp24[38],pp24[39],pp26[38],pp28[37],pp30[36],pp32[35],pp34[34],pp36[33],pp38[32],pp40[31],pp42[30],pp44[29],pp46[28],pp48[27],pp50[26],pp52[25],pp54[24],pp56[23],pp58[22],pp60[21],pp62[20],pp64[19],pp66[18],pp68[17],pp70[16],pp72[15],pp74[14],pp76[13],pp78[12],pp80[11],pp82[10],pp0[93],pp1[93],pp2[93],pp3[93],pp4[93],pp5[93],pp6[93],pp6[94],pp6[95],pp6[96],pp6[97],pp6[98],pp6[99],pp106[0],pp106[1],pp106[2],pp106[3],pp108[2],pp110[1],pp112[0],s10[40],s11[40],s12[40],s13[40],s14[40],s15[40],s16[40],s17[40],s18[40],s19[40],s20[40],s21[40],s22[40],s23[40],s24[40],s25[40],s24[42],s23[44],s22[46],s20[49],s18[52],s16[55],s14[58],s12[61],s10[64],s70[101],s69[103],s68[105],s67[107],s66[109],s65[111],pp99[45],pp98[47],pp97[49],pp96[51],pp95[53],pp94[55],pp93[57],pp92[59],pp91[61],pp90[63],pp89[65],pp88[67],pp87[69],pp86[71],pp85[73],pp84[75],pp83[77],pp82[79],pp81[81],pp80[83],pp79[85],pp78[87],pp77[89],pp76[91],pp75[93],pp74[95],pp73[97],pp72[99],pp126[46],pp124[49],pp122[52],pp120[55],pp118[58],pp116[61],pp114[64],pp112[67],pp110[70],pp108[73],pp106[76],pp104[79],pp102[82],pp100[85],pp85[101],pp84[103],pp83[105],pp82[107],pp81[109],pp80[111],pp79[113],pp80[113],pp81[113],pp82[113],pp83[113],pp84[113],pp85[113],pp86[113],pp86[114],pp86[115],pp86[116],pp86[117],pp86[118],pp86[119],pp86[120],pp86[121],pp86[122],pp86[123],pp86[124],pp86[125],pp86[126],pp86[127],pp114[100],pp114[101],pp114[102]};
    assign in72_2 = {pp25[14],pp25[15],pp25[16],pp25[17],pp25[18],pp25[19],pp25[20],pp25[21],pp25[22],pp25[23],pp25[24],pp25[25],pp25[26],pp25[27],pp25[28],pp25[29],pp25[30],pp25[31],pp25[32],pp25[33],pp25[34],pp25[35],pp25[36],pp25[37],pp25[38],pp27[37],pp29[36],pp31[35],pp33[34],pp35[33],pp37[32],pp39[31],pp41[30],pp43[29],pp45[28],pp47[27],pp49[26],pp51[25],pp53[24],pp55[23],pp57[22],pp59[21],pp61[20],pp63[19],pp65[18],pp67[17],pp69[16],pp71[15],pp73[14],pp75[13],pp77[12],pp79[11],pp81[10],pp0[92],pp1[92],pp2[92],pp3[92],pp4[92],pp5[92],pp6[92],pp7[92],pp7[93],pp7[94],pp7[95],pp7[96],pp7[97],pp7[98],pp7[99],pp107[0],pp107[1],pp107[2],pp109[1],pp111[0],s10[39],s11[39],s12[39],s13[39],s14[39],s15[39],s16[39],s17[39],s18[39],s19[39],s20[39],s21[39],s22[39],s23[39],s24[39],s25[39],s26[39],s25[41],s24[43],s23[45],s21[48],s19[51],s17[54],s15[57],s13[60],s11[63],s71[100],s70[102],s69[104],s68[106],s67[108],s66[110],s65[112],pp99[46],pp98[48],pp97[50],pp96[52],pp95[54],pp94[56],pp93[58],pp92[60],pp91[62],pp90[64],pp89[66],pp88[68],pp87[70],pp86[72],pp85[74],pp84[76],pp83[78],pp82[80],pp81[82],pp80[84],pp79[86],pp78[88],pp77[90],pp76[92],pp75[94],pp74[96],pp73[98],pp127[45],pp125[48],pp123[51],pp121[54],pp119[57],pp117[60],pp115[63],pp113[66],pp111[69],pp109[72],pp107[75],pp105[78],pp103[81],pp101[84],pp86[100],pp85[102],pp84[104],pp83[106],pp82[108],pp81[110],pp80[112],pp81[112],pp82[112],pp83[112],pp84[112],pp85[112],pp86[112],pp87[112],pp87[113],pp87[114],pp87[115],pp87[116],pp87[117],pp87[118],pp87[119],pp87[120],pp87[121],pp87[122],pp87[123],pp87[124],pp87[125],pp87[126],pp87[127],pp115[100],pp115[101]};
    CLA_178 KS_72(s72, c72, in72_1, in72_2);
    wire[175:0] s73, in73_1, in73_2;
    wire c73;
    assign in73_1 = {pp26[14],pp26[15],pp26[16],pp26[17],pp26[18],pp26[19],pp26[20],pp26[21],pp26[22],pp26[23],pp26[24],pp26[25],pp26[26],pp26[27],pp26[28],pp26[29],pp26[30],pp26[31],pp26[32],pp26[33],pp26[34],pp26[35],pp26[36],pp26[37],pp28[36],pp30[35],pp32[34],pp34[33],pp36[32],pp38[31],pp40[30],pp42[29],pp44[28],pp46[27],pp48[26],pp50[25],pp52[24],pp54[23],pp56[22],pp58[21],pp60[20],pp62[19],pp64[18],pp66[17],pp68[16],pp70[15],pp72[14],pp74[13],pp76[12],pp78[11],pp80[10],pp0[91],pp1[91],pp2[91],pp3[91],pp4[91],pp5[91],pp6[91],pp7[91],pp8[91],pp8[92],pp8[93],pp8[94],pp8[95],pp8[96],pp8[97],pp8[98],pp8[99],pp108[0],pp108[1],pp110[0],s10[38],s11[38],s12[38],s13[38],s14[38],s15[38],s16[38],s17[38],s18[38],s19[38],s20[38],s21[38],s22[38],s23[38],s24[38],s25[38],s26[38],s27[38],s26[40],s25[42],s24[44],s22[47],s20[50],s18[53],s16[56],s14[59],s12[62],s10[65],s71[101],s70[103],s69[105],s68[107],s67[109],s66[111],s65[113],pp99[47],pp98[49],pp97[51],pp96[53],pp95[55],pp94[57],pp93[59],pp92[61],pp91[63],pp90[65],pp89[67],pp88[69],pp87[71],pp86[73],pp85[75],pp84[77],pp83[79],pp82[81],pp81[83],pp80[85],pp79[87],pp78[89],pp77[91],pp76[93],pp75[95],pp74[97],pp73[99],pp126[47],pp124[50],pp122[53],pp120[56],pp118[59],pp116[62],pp114[65],pp112[68],pp110[71],pp108[74],pp106[77],pp104[80],pp102[83],pp100[86],pp86[101],pp85[103],pp84[105],pp83[107],pp82[109],pp81[111],pp82[111],pp83[111],pp84[111],pp85[111],pp86[111],pp87[111],pp88[111],pp88[112],pp88[113],pp88[114],pp88[115],pp88[116],pp88[117],pp88[118],pp88[119],pp88[120],pp88[121],pp88[122],pp88[123],pp88[124],pp88[125],pp88[126],pp88[127]};
    assign in73_2 = {pp27[13],pp27[14],pp27[15],pp27[16],pp27[17],pp27[18],pp27[19],pp27[20],pp27[21],pp27[22],pp27[23],pp27[24],pp27[25],pp27[26],pp27[27],pp27[28],pp27[29],pp27[30],pp27[31],pp27[32],pp27[33],pp27[34],pp27[35],pp27[36],pp29[35],pp31[34],pp33[33],pp35[32],pp37[31],pp39[30],pp41[29],pp43[28],pp45[27],pp47[26],pp49[25],pp51[24],pp53[23],pp55[22],pp57[21],pp59[20],pp61[19],pp63[18],pp65[17],pp67[16],pp69[15],pp71[14],pp73[13],pp75[12],pp77[11],pp79[10],pp0[90],pp1[90],pp2[90],pp3[90],pp4[90],pp5[90],pp6[90],pp7[90],pp8[90],pp9[90],pp9[91],pp9[92],pp9[93],pp9[94],pp9[95],pp9[96],pp9[97],pp9[98],pp9[99],pp109[0],s10[37],s11[37],s12[37],s13[37],s14[37],s15[37],s16[37],s17[37],s18[37],s19[37],s20[37],s21[37],s22[37],s23[37],s24[37],s25[37],s26[37],s27[37],s28[37],s27[39],s26[41],s25[43],s23[46],s21[49],s19[52],s17[55],s15[58],s13[61],s11[64],s72[100],s71[102],s70[104],s69[106],s68[108],s67[110],s66[112],s65[114],pp99[48],pp98[50],pp97[52],pp96[54],pp95[56],pp94[58],pp93[60],pp92[62],pp91[64],pp90[66],pp89[68],pp88[70],pp87[72],pp86[74],pp85[76],pp84[78],pp83[80],pp82[82],pp81[84],pp80[86],pp79[88],pp78[90],pp77[92],pp76[94],pp75[96],pp74[98],pp127[46],pp125[49],pp123[52],pp121[55],pp119[58],pp117[61],pp115[64],pp113[67],pp111[70],pp109[73],pp107[76],pp105[79],pp103[82],pp101[85],pp87[100],pp86[102],pp85[104],pp84[106],pp83[108],pp82[110],pp83[110],pp84[110],pp85[110],pp86[110],pp87[110],pp88[110],pp89[110],pp89[111],pp89[112],pp89[113],pp89[114],pp89[115],pp89[116],pp89[117],pp89[118],pp89[119],pp89[120],pp89[121],pp89[122],pp89[123],pp89[124],pp89[125],pp89[126]};
    CLA_176 KS_73(s73, c73, in73_1, in73_2);
    wire[173:0] s74, in74_1, in74_2;
    wire c74;
    assign in74_1 = {pp28[13],pp28[14],pp28[15],pp28[16],pp28[17],pp28[18],pp28[19],pp28[20],pp28[21],pp28[22],pp28[23],pp28[24],pp28[25],pp28[26],pp28[27],pp28[28],pp28[29],pp28[30],pp28[31],pp28[32],pp28[33],pp28[34],pp28[35],pp30[34],pp32[33],pp34[32],pp36[31],pp38[30],pp40[29],pp42[28],pp44[27],pp46[26],pp48[25],pp50[24],pp52[23],pp54[22],pp56[21],pp58[20],pp60[19],pp62[18],pp64[17],pp66[16],pp68[15],pp70[14],pp72[13],pp74[12],pp76[11],pp78[10],pp0[89],pp1[89],pp2[89],pp3[89],pp4[89],pp5[89],pp6[89],pp7[89],pp8[89],pp9[89],pp90[9],pp91[9],pp92[9],pp93[9],pp94[9],pp95[9],pp96[9],pp97[9],pp98[9],pp99[9],s10[36],s11[36],s12[36],s13[36],s14[36],s15[36],s16[36],s17[36],s18[36],s19[36],s20[36],s21[36],s22[36],s23[36],s24[36],s25[36],s26[36],s27[36],s28[36],s29[36],s28[38],s27[40],s26[42],s24[45],s22[48],s20[51],s18[54],s16[57],s14[60],s12[63],s10[66],s72[101],s71[103],s70[105],s69[107],s68[109],s67[111],s66[113],s65[115],pp99[49],pp98[51],pp97[53],pp96[55],pp95[57],pp94[59],pp93[61],pp92[63],pp91[65],pp90[67],pp89[69],pp88[71],pp87[73],pp86[75],pp85[77],pp84[79],pp83[81],pp82[83],pp81[85],pp80[87],pp79[89],pp78[91],pp77[93],pp76[95],pp75[97],pp74[99],pp126[48],pp124[51],pp122[54],pp120[57],pp118[60],pp116[63],pp114[66],pp112[69],pp110[72],pp108[75],pp106[78],pp104[81],pp102[84],pp100[87],pp87[101],pp86[103],pp85[105],pp84[107],pp83[109],pp84[109],pp85[109],pp86[109],pp87[109],pp88[109],pp89[109],pp90[109],pp90[110],pp90[111],pp90[112],pp90[113],pp90[114],pp90[115],pp90[116],pp90[117],pp90[118],pp90[119],pp90[120],pp90[121],pp90[122],pp90[123],pp90[124]};
    assign in74_2 = {pp29[12],pp29[13],pp29[14],pp29[15],pp29[16],pp29[17],pp29[18],pp29[19],pp29[20],pp29[21],pp29[22],pp29[23],pp29[24],pp29[25],pp29[26],pp29[27],pp29[28],pp29[29],pp29[30],pp29[31],pp29[32],pp29[33],pp29[34],pp31[33],pp33[32],pp35[31],pp37[30],pp39[29],pp41[28],pp43[27],pp45[26],pp47[25],pp49[24],pp51[23],pp53[22],pp55[21],pp57[20],pp59[19],pp61[18],pp63[17],pp65[16],pp67[15],pp69[14],pp71[13],pp73[12],pp75[11],pp77[10],pp0[88],pp1[88],pp2[88],pp3[88],pp4[88],pp5[88],pp6[88],pp7[88],pp8[88],pp9[88],pp89[9],pp91[8],pp92[8],pp93[8],pp94[8],pp95[8],pp96[8],pp97[8],pp98[8],pp99[8],s10[35],s11[35],s12[35],s13[35],s14[35],s15[35],s16[35],s17[35],s18[35],s19[35],s20[35],s21[35],s22[35],s23[35],s24[35],s25[35],s26[35],s27[35],s28[35],s29[35],s30[35],s29[37],s28[39],s27[41],s25[44],s23[47],s21[50],s19[53],s17[56],s15[59],s13[62],s11[65],s73[100],s72[102],s71[104],s70[106],s69[108],s68[110],s67[112],s66[114],s65[116],pp99[50],pp98[52],pp97[54],pp96[56],pp95[58],pp94[60],pp93[62],pp92[64],pp91[66],pp90[68],pp89[70],pp88[72],pp87[74],pp86[76],pp85[78],pp84[80],pp83[82],pp82[84],pp81[86],pp80[88],pp79[90],pp78[92],pp77[94],pp76[96],pp75[98],pp127[47],pp125[50],pp123[53],pp121[56],pp119[59],pp117[62],pp115[65],pp113[68],pp111[71],pp109[74],pp107[77],pp105[80],pp103[83],pp101[86],pp88[100],pp87[102],pp86[104],pp85[106],pp84[108],pp85[108],pp86[108],pp87[108],pp88[108],pp89[108],pp90[108],pp91[108],pp91[109],pp91[110],pp91[111],pp91[112],pp91[113],pp91[114],pp91[115],pp91[116],pp91[117],pp91[118],pp91[119],pp91[120],pp91[121],pp91[122],pp91[123]};
    CLA_174 KS_74(s74, c74, in74_1, in74_2);
    wire[171:0] s75, in75_1, in75_2;
    wire c75;
    assign in75_1 = {pp30[12],pp30[13],pp30[14],pp30[15],pp30[16],pp30[17],pp30[18],pp30[19],pp30[20],pp30[21],pp30[22],pp30[23],pp30[24],pp30[25],pp30[26],pp30[27],pp30[28],pp30[29],pp30[30],pp30[31],pp30[32],pp30[33],pp32[32],pp34[31],pp36[30],pp38[29],pp40[28],pp42[27],pp44[26],pp46[25],pp48[24],pp50[23],pp52[22],pp54[21],pp56[20],pp58[19],pp60[18],pp62[17],pp64[16],pp66[15],pp68[14],pp70[13],pp72[12],pp74[11],pp76[10],pp0[87],pp1[87],pp2[87],pp3[87],pp4[87],pp5[87],pp6[87],pp7[87],pp8[87],pp9[87],pp88[9],pp90[8],pp92[7],pp93[7],pp94[7],pp95[7],pp96[7],pp97[7],pp98[7],pp99[7],s10[34],s11[34],s12[34],s13[34],s14[34],s15[34],s16[34],s17[34],s18[34],s19[34],s20[34],s21[34],s22[34],s23[34],s24[34],s25[34],s26[34],s27[34],s28[34],s29[34],s30[34],s31[34],s30[36],s29[38],s28[40],s26[43],s24[46],s22[49],s20[52],s18[55],s16[58],s14[61],s12[64],s10[67],s73[101],s72[103],s71[105],s70[107],s69[109],s68[111],s67[113],s66[115],s65[117],pp99[51],pp98[53],pp97[55],pp96[57],pp95[59],pp94[61],pp93[63],pp92[65],pp91[67],pp90[69],pp89[71],pp88[73],pp87[75],pp86[77],pp85[79],pp84[81],pp83[83],pp82[85],pp81[87],pp80[89],pp79[91],pp78[93],pp77[95],pp76[97],pp75[99],pp126[49],pp124[52],pp122[55],pp120[58],pp118[61],pp116[64],pp114[67],pp112[70],pp110[73],pp108[76],pp106[79],pp104[82],pp102[85],pp100[88],pp88[101],pp87[103],pp86[105],pp85[107],pp86[107],pp87[107],pp88[107],pp89[107],pp90[107],pp91[107],pp92[107],pp92[108],pp92[109],pp92[110],pp92[111],pp92[112],pp92[113],pp92[114],pp92[115],pp92[116],pp92[117],pp92[118],pp92[119],pp92[120],pp92[121]};
    assign in75_2 = {pp31[11],pp31[12],pp31[13],pp31[14],pp31[15],pp31[16],pp31[17],pp31[18],pp31[19],pp31[20],pp31[21],pp31[22],pp31[23],pp31[24],pp31[25],pp31[26],pp31[27],pp31[28],pp31[29],pp31[30],pp31[31],pp31[32],pp33[31],pp35[30],pp37[29],pp39[28],pp41[27],pp43[26],pp45[25],pp47[24],pp49[23],pp51[22],pp53[21],pp55[20],pp57[19],pp59[18],pp61[17],pp63[16],pp65[15],pp67[14],pp69[13],pp71[12],pp73[11],pp75[10],pp0[86],pp1[86],pp2[86],pp3[86],pp4[86],pp5[86],pp6[86],pp7[86],pp8[86],pp9[86],pp87[9],pp89[8],pp91[7],pp93[6],pp94[6],pp95[6],pp96[6],pp97[6],pp98[6],pp99[6],s10[33],s11[33],s12[33],s13[33],s14[33],s15[33],s16[33],s17[33],s18[33],s19[33],s20[33],s21[33],s22[33],s23[33],s24[33],s25[33],s26[33],s27[33],s28[33],s29[33],s30[33],s31[33],s32[33],s31[35],s30[37],s29[39],s27[42],s25[45],s23[48],s21[51],s19[54],s17[57],s15[60],s13[63],s11[66],s74[100],s73[102],s72[104],s71[106],s70[108],s69[110],s68[112],s67[114],s66[116],s65[118],pp99[52],pp98[54],pp97[56],pp96[58],pp95[60],pp94[62],pp93[64],pp92[66],pp91[68],pp90[70],pp89[72],pp88[74],pp87[76],pp86[78],pp85[80],pp84[82],pp83[84],pp82[86],pp81[88],pp80[90],pp79[92],pp78[94],pp77[96],pp76[98],pp127[48],pp125[51],pp123[54],pp121[57],pp119[60],pp117[63],pp115[66],pp113[69],pp111[72],pp109[75],pp107[78],pp105[81],pp103[84],pp101[87],pp89[100],pp88[102],pp87[104],pp86[106],pp87[106],pp88[106],pp89[106],pp90[106],pp91[106],pp92[106],pp93[106],pp93[107],pp93[108],pp93[109],pp93[110],pp93[111],pp93[112],pp93[113],pp93[114],pp93[115],pp93[116],pp93[117],pp93[118],pp93[119],pp93[120]};
    CLA_172 KS_75(s75, c75, in75_1, in75_2);
    wire[169:0] s76, in76_1, in76_2;
    wire c76;
    assign in76_1 = {pp32[11],pp32[12],pp32[13],pp32[14],pp32[15],pp32[16],pp32[17],pp32[18],pp32[19],pp32[20],pp32[21],pp32[22],pp32[23],pp32[24],pp32[25],pp32[26],pp32[27],pp32[28],pp32[29],pp32[30],pp32[31],pp34[30],pp36[29],pp38[28],pp40[27],pp42[26],pp44[25],pp46[24],pp48[23],pp50[22],pp52[21],pp54[20],pp56[19],pp58[18],pp60[17],pp62[16],pp64[15],pp66[14],pp68[13],pp70[12],pp72[11],pp74[10],pp0[85],pp1[85],pp2[85],pp3[85],pp4[85],pp5[85],pp6[85],pp7[85],pp8[85],pp9[85],pp86[9],pp88[8],pp90[7],pp92[6],pp94[5],pp95[5],pp96[5],pp97[5],pp98[5],pp99[5],s10[32],s11[32],s12[32],s13[32],s14[32],s15[32],s16[32],s17[32],s18[32],s19[32],s20[32],s21[32],s22[32],s23[32],s24[32],s25[32],s26[32],s27[32],s28[32],s29[32],s30[32],s31[32],s32[32],s33[32],s32[34],s31[36],s30[38],s28[41],s26[44],s24[47],s22[50],s20[53],s18[56],s16[59],s14[62],s12[65],s10[68],s74[101],s73[103],s72[105],s71[107],s70[109],s69[111],s68[113],s67[115],s66[117],s65[119],pp99[53],pp98[55],pp97[57],pp96[59],pp95[61],pp94[63],pp93[65],pp92[67],pp91[69],pp90[71],pp89[73],pp88[75],pp87[77],pp86[79],pp85[81],pp84[83],pp83[85],pp82[87],pp81[89],pp80[91],pp79[93],pp78[95],pp77[97],pp76[99],pp126[50],pp124[53],pp122[56],pp120[59],pp118[62],pp116[65],pp114[68],pp112[71],pp110[74],pp108[77],pp106[80],pp104[83],pp102[86],pp100[89],pp89[101],pp88[103],pp87[105],pp88[105],pp89[105],pp90[105],pp91[105],pp92[105],pp93[105],pp94[105],pp94[106],pp94[107],pp94[108],pp94[109],pp94[110],pp94[111],pp94[112],pp94[113],pp94[114],pp94[115],pp94[116],pp94[117],pp94[118]};
    assign in76_2 = {pp33[10],pp33[11],pp33[12],pp33[13],pp33[14],pp33[15],pp33[16],pp33[17],pp33[18],pp33[19],pp33[20],pp33[21],pp33[22],pp33[23],pp33[24],pp33[25],pp33[26],pp33[27],pp33[28],pp33[29],pp33[30],pp35[29],pp37[28],pp39[27],pp41[26],pp43[25],pp45[24],pp47[23],pp49[22],pp51[21],pp53[20],pp55[19],pp57[18],pp59[17],pp61[16],pp63[15],pp65[14],pp67[13],pp69[12],pp71[11],pp73[10],pp0[84],pp1[84],pp2[84],pp3[84],pp4[84],pp5[84],pp6[84],pp7[84],pp8[84],pp9[84],pp85[9],pp87[8],pp89[7],pp91[6],pp93[5],pp95[4],pp96[4],pp97[4],pp98[4],pp99[4],s10[31],s11[31],s12[31],s13[31],s14[31],s15[31],s16[31],s17[31],s18[31],s19[31],s20[31],s21[31],s22[31],s23[31],s24[31],s25[31],s26[31],s27[31],s28[31],s29[31],s30[31],s31[31],s32[31],s33[31],s34[31],s33[33],s32[35],s31[37],s29[40],s27[43],s25[46],s23[49],s21[52],s19[55],s17[58],s15[61],s13[64],s11[67],s75[100],s74[102],s73[104],s72[106],s71[108],s70[110],s69[112],s68[114],s67[116],s66[118],s65[120],pp99[54],pp98[56],pp97[58],pp96[60],pp95[62],pp94[64],pp93[66],pp92[68],pp91[70],pp90[72],pp89[74],pp88[76],pp87[78],pp86[80],pp85[82],pp84[84],pp83[86],pp82[88],pp81[90],pp80[92],pp79[94],pp78[96],pp77[98],pp127[49],pp125[52],pp123[55],pp121[58],pp119[61],pp117[64],pp115[67],pp113[70],pp111[73],pp109[76],pp107[79],pp105[82],pp103[85],pp101[88],pp90[100],pp89[102],pp88[104],pp89[104],pp90[104],pp91[104],pp92[104],pp93[104],pp94[104],pp95[104],pp95[105],pp95[106],pp95[107],pp95[108],pp95[109],pp95[110],pp95[111],pp95[112],pp95[113],pp95[114],pp95[115],pp95[116],pp95[117]};
    CLA_170 KS_76(s76, c76, in76_1, in76_2);
    wire[167:0] s77, in77_1, in77_2;
    wire c77;
    assign in77_1 = {pp34[10],pp34[11],pp34[12],pp34[13],pp34[14],pp34[15],pp34[16],pp34[17],pp34[18],pp34[19],pp34[20],pp34[21],pp34[22],pp34[23],pp34[24],pp34[25],pp34[26],pp34[27],pp34[28],pp34[29],pp36[28],pp38[27],pp40[26],pp42[25],pp44[24],pp46[23],pp48[22],pp50[21],pp52[20],pp54[19],pp56[18],pp58[17],pp60[16],pp62[15],pp64[14],pp66[13],pp68[12],pp70[11],pp72[10],pp0[83],pp1[83],pp2[83],pp3[83],pp4[83],pp5[83],pp6[83],pp7[83],pp8[83],pp9[83],pp84[9],pp86[8],pp88[7],pp90[6],pp92[5],pp94[4],pp96[3],pp97[3],pp98[3],pp99[3],s10[30],s11[30],s12[30],s13[30],s14[30],s15[30],s16[30],s17[30],s18[30],s19[30],s20[30],s21[30],s22[30],s23[30],s24[30],s25[30],s26[30],s27[30],s28[30],s29[30],s30[30],s31[30],s32[30],s33[30],s34[30],s35[30],s34[32],s33[34],s32[36],s30[39],s28[42],s26[45],s24[48],s22[51],s20[54],s18[57],s16[60],s14[63],s12[66],s10[69],s75[101],s74[103],s73[105],s72[107],s71[109],s70[111],s69[113],s68[115],s67[117],s66[119],s65[121],pp99[55],pp98[57],pp97[59],pp96[61],pp95[63],pp94[65],pp93[67],pp92[69],pp91[71],pp90[73],pp89[75],pp88[77],pp87[79],pp86[81],pp85[83],pp84[85],pp83[87],pp82[89],pp81[91],pp80[93],pp79[95],pp78[97],pp77[99],pp126[51],pp124[54],pp122[57],pp120[60],pp118[63],pp116[66],pp114[69],pp112[72],pp110[75],pp108[78],pp106[81],pp104[84],pp102[87],pp100[90],pp90[101],pp89[103],pp90[103],pp91[103],pp92[103],pp93[103],pp94[103],pp95[103],pp96[103],pp96[104],pp96[105],pp96[106],pp96[107],pp96[108],pp96[109],pp96[110],pp96[111],pp96[112],pp96[113],pp96[114],pp96[115]};
    assign in77_2 = {pp0[44],pp35[10],pp35[11],pp35[12],pp35[13],pp35[14],pp35[15],pp35[16],pp35[17],pp35[18],pp35[19],pp35[20],pp35[21],pp35[22],pp35[23],pp35[24],pp35[25],pp35[26],pp35[27],pp35[28],pp37[27],pp39[26],pp41[25],pp43[24],pp45[23],pp47[22],pp49[21],pp51[20],pp53[19],pp55[18],pp57[17],pp59[16],pp61[15],pp63[14],pp65[13],pp67[12],pp69[11],pp71[10],pp0[82],pp1[82],pp2[82],pp3[82],pp4[82],pp5[82],pp6[82],pp7[82],pp8[82],pp9[82],pp83[9],pp85[8],pp87[7],pp89[6],pp91[5],pp93[4],pp95[3],pp97[2],pp98[2],pp99[2],s10[29],s11[29],s12[29],s13[29],s14[29],s15[29],s16[29],s17[29],s18[29],s19[29],s20[29],s21[29],s22[29],s23[29],s24[29],s25[29],s26[29],s27[29],s28[29],s29[29],s30[29],s31[29],s32[29],s33[29],s34[29],s35[29],s36[29],s35[31],s34[33],s33[35],s31[38],s29[41],s27[44],s25[47],s23[50],s21[53],s19[56],s17[59],s15[62],s13[65],s11[68],s76[100],s75[102],s74[104],s73[106],s72[108],s71[110],s70[112],s69[114],s68[116],s67[118],s66[120],s65[122],pp99[56],pp98[58],pp97[60],pp96[62],pp95[64],pp94[66],pp93[68],pp92[70],pp91[72],pp90[74],pp89[76],pp88[78],pp87[80],pp86[82],pp85[84],pp84[86],pp83[88],pp82[90],pp81[92],pp80[94],pp79[96],pp78[98],pp127[50],pp125[53],pp123[56],pp121[59],pp119[62],pp117[65],pp115[68],pp113[71],pp111[74],pp109[77],pp107[80],pp105[83],pp103[86],pp101[89],pp91[100],pp90[102],pp91[102],pp92[102],pp93[102],pp94[102],pp95[102],pp96[102],pp97[102],pp97[103],pp97[104],pp97[105],pp97[106],pp97[107],pp97[108],pp97[109],pp97[110],pp97[111],pp97[112],pp97[113],pp97[114]};
    CLA_168 KS_77(s77, c77, in77_1, in77_2);
    wire[165:0] s78, in78_1, in78_2;
    wire c78;
    assign in78_1 = {pp0[45],pp36[10],pp36[11],pp36[12],pp36[13],pp36[14],pp36[15],pp36[16],pp36[17],pp36[18],pp36[19],pp36[20],pp36[21],pp36[22],pp36[23],pp36[24],pp36[25],pp36[26],pp36[27],pp38[26],pp40[25],pp42[24],pp44[23],pp46[22],pp48[21],pp50[20],pp52[19],pp54[18],pp56[17],pp58[16],pp60[15],pp62[14],pp64[13],pp66[12],pp68[11],pp70[10],pp0[81],pp1[81],pp2[81],pp3[81],pp4[81],pp5[81],pp6[81],pp7[81],pp8[81],pp9[81],pp82[9],pp84[8],pp86[7],pp88[6],pp90[5],pp92[4],pp94[3],pp96[2],pp98[1],pp99[1],s10[28],s11[28],s12[28],s13[28],s14[28],s15[28],s16[28],s17[28],s18[28],s19[28],s20[28],s21[28],s22[28],s23[28],s24[28],s25[28],s26[28],s27[28],s28[28],s29[28],s30[28],s31[28],s32[28],s33[28],s34[28],s35[28],s36[28],s37[28],s36[30],s35[32],s34[34],s32[37],s30[40],s28[43],s26[46],s24[49],s22[52],s20[55],s18[58],s16[61],s14[64],s12[67],s10[70],s76[101],s75[103],s74[105],s73[107],s72[109],s71[111],s70[113],s69[115],s68[117],s67[119],s66[121],s65[123],pp99[57],pp98[59],pp97[61],pp96[63],pp95[65],pp94[67],pp93[69],pp92[71],pp91[73],pp90[75],pp89[77],pp88[79],pp87[81],pp86[83],pp85[85],pp84[87],pp83[89],pp82[91],pp81[93],pp80[95],pp79[97],pp78[99],pp126[52],pp124[55],pp122[58],pp120[61],pp118[64],pp116[67],pp114[70],pp112[73],pp110[76],pp108[79],pp106[82],pp104[85],pp102[88],pp100[91],pp91[101],pp92[101],pp93[101],pp94[101],pp95[101],pp96[101],pp97[101],pp98[101],pp98[102],pp98[103],pp98[104],pp98[105],pp98[106],pp98[107],pp98[108],pp98[109],pp98[110],pp98[111],pp98[112]};
    assign in78_2 = {pp1[44],pp0[46],pp37[10],pp37[11],pp37[12],pp37[13],pp37[14],pp37[15],pp37[16],pp37[17],pp37[18],pp37[19],pp37[20],pp37[21],pp37[22],pp37[23],pp37[24],pp37[25],pp37[26],pp39[25],pp41[24],pp43[23],pp45[22],pp47[21],pp49[20],pp51[19],pp53[18],pp55[17],pp57[16],pp59[15],pp61[14],pp63[13],pp65[12],pp67[11],pp69[10],pp0[80],pp1[80],pp2[80],pp3[80],pp4[80],pp5[80],pp6[80],pp7[80],pp8[80],pp9[80],pp81[9],pp83[8],pp85[7],pp87[6],pp89[5],pp91[4],pp93[3],pp95[2],pp97[1],pp99[0],s10[27],s11[27],s12[27],s13[27],s14[27],s15[27],s16[27],s17[27],s18[27],s19[27],s20[27],s21[27],s22[27],s23[27],s24[27],s25[27],s26[27],s27[27],s28[27],s29[27],s30[27],s31[27],s32[27],s33[27],s34[27],s35[27],s36[27],s37[27],s38[27],s37[29],s36[31],s35[33],s33[36],s31[39],s29[42],s27[45],s25[48],s23[51],s21[54],s19[57],s17[60],s15[63],s13[66],s11[69],s77[100],s76[102],s75[104],s74[106],s73[108],s72[110],s71[112],s70[114],s69[116],s68[118],s67[120],s66[122],s65[124],pp99[58],pp98[60],pp97[62],pp96[64],pp95[66],pp94[68],pp93[70],pp92[72],pp91[74],pp90[76],pp89[78],pp88[80],pp87[82],pp86[84],pp85[86],pp84[88],pp83[90],pp82[92],pp81[94],pp80[96],pp79[98],pp127[51],pp125[54],pp123[57],pp121[60],pp119[63],pp117[66],pp115[69],pp113[72],pp111[75],pp109[78],pp107[81],pp105[84],pp103[87],pp101[90],pp92[100],pp93[100],pp94[100],pp95[100],pp96[100],pp97[100],pp98[100],pp99[100],pp99[101],pp99[102],pp99[103],pp99[104],pp99[105],pp99[106],pp99[107],pp99[108],pp99[109],pp99[110],pp99[111]};
    CLA_166 KS_78(s78, c78, in78_1, in78_2);
    wire[163:0] s79, in79_1, in79_2;
    wire c79;
    assign in79_1 = {pp1[45],pp0[47],pp38[10],pp38[11],pp38[12],pp38[13],pp38[14],pp38[15],pp38[16],pp38[17],pp38[18],pp38[19],pp38[20],pp38[21],pp38[22],pp38[23],pp38[24],pp38[25],pp40[24],pp42[23],pp44[22],pp46[21],pp48[20],pp50[19],pp52[18],pp54[17],pp56[16],pp58[15],pp60[14],pp62[13],pp64[12],pp66[11],pp68[10],pp0[79],pp1[79],pp2[79],pp3[79],pp4[79],pp5[79],pp6[79],pp7[79],pp8[79],pp9[79],pp80[9],pp82[8],pp84[7],pp86[6],pp88[5],pp90[4],pp92[3],pp94[2],pp96[1],pp98[0],s10[26],s11[26],s12[26],s13[26],s14[26],s15[26],s16[26],s17[26],s18[26],s19[26],s20[26],s21[26],s22[26],s23[26],s24[26],s25[26],s26[26],s27[26],s28[26],s29[26],s30[26],s31[26],s32[26],s33[26],s34[26],s35[26],s36[26],s37[26],s38[26],s39[26],s38[28],s37[30],s36[32],s34[35],s32[38],s30[41],s28[44],s26[47],s24[50],s22[53],s20[56],s18[59],s16[62],s14[65],s12[68],s10[71],s77[101],s76[103],s75[105],s74[107],s73[109],s72[111],s71[113],s70[115],s69[117],s68[119],s67[121],s66[123],s65[125],pp99[59],pp98[61],pp97[63],pp96[65],pp95[67],pp94[69],pp93[71],pp92[73],pp91[75],pp90[77],pp89[79],pp88[81],pp87[83],pp86[85],pp85[87],pp84[89],pp83[91],pp82[93],pp81[95],pp80[97],pp79[99],pp126[53],pp124[56],pp122[59],pp120[62],pp118[65],pp116[68],pp114[71],pp112[74],pp110[77],pp108[80],pp106[83],pp104[86],pp102[89],pp100[92],pp100[93],pp100[94],pp100[95],pp100[96],pp100[97],pp100[98],pp100[99],pp101[99],pp102[99],pp103[99],pp104[99],pp105[99],pp106[99],pp107[99],pp108[99],pp109[99],pp110[99]};
    assign in79_2 = {pp2[44],pp1[46],pp0[48],pp39[10],pp39[11],pp39[12],pp39[13],pp39[14],pp39[15],pp39[16],pp39[17],pp39[18],pp39[19],pp39[20],pp39[21],pp39[22],pp39[23],pp39[24],pp41[23],pp43[22],pp45[21],pp47[20],pp49[19],pp51[18],pp53[17],pp55[16],pp57[15],pp59[14],pp61[13],pp63[12],pp65[11],pp67[10],pp0[78],pp1[78],pp2[78],pp3[78],pp4[78],pp5[78],pp6[78],pp7[78],pp8[78],pp9[78],pp79[9],pp81[8],pp83[7],pp85[6],pp87[5],pp89[4],pp91[3],pp93[2],pp95[1],pp97[0],s10[25],s11[25],s12[25],s13[25],s14[25],s15[25],s16[25],s17[25],s18[25],s19[25],s20[25],s21[25],s22[25],s23[25],s24[25],s25[25],s26[25],s27[25],s28[25],s29[25],s30[25],s31[25],s32[25],s33[25],s34[25],s35[25],s36[25],s37[25],s38[25],s39[25],s40[25],s39[27],s38[29],s37[31],s35[34],s33[37],s31[40],s29[43],s27[46],s25[49],s23[52],s21[55],s19[58],s17[61],s15[64],s13[67],s11[70],s78[100],s77[102],s76[104],s75[106],s74[108],s73[110],s72[112],s71[114],s70[116],s69[118],s68[120],s67[122],s66[124],s65[126],pp99[60],pp98[62],pp97[64],pp96[66],pp95[68],pp94[70],pp93[72],pp92[74],pp91[76],pp90[78],pp89[80],pp88[82],pp87[84],pp86[86],pp85[88],pp84[90],pp83[92],pp82[94],pp81[96],pp80[98],pp127[52],pp125[55],pp123[58],pp121[61],pp119[64],pp117[67],pp115[70],pp113[73],pp111[76],pp109[79],pp107[82],pp105[85],pp103[88],pp101[91],pp101[92],pp101[93],pp101[94],pp101[95],pp101[96],pp101[97],pp101[98],pp102[98],pp103[98],pp104[98],pp105[98],pp106[98],pp107[98],pp108[98],pp109[98],pp110[98],pp111[98]};
    CLA_164 KS_79(s79, c79, in79_1, in79_2);
    wire[161:0] s80, in80_1, in80_2;
    wire c80;
    assign in80_1 = {pp2[45],pp1[47],pp0[49],pp40[10],pp40[11],pp40[12],pp40[13],pp40[14],pp40[15],pp40[16],pp40[17],pp40[18],pp40[19],pp40[20],pp40[21],pp40[22],pp40[23],pp42[22],pp44[21],pp46[20],pp48[19],pp50[18],pp52[17],pp54[16],pp56[15],pp58[14],pp60[13],pp62[12],pp64[11],pp66[10],pp0[77],pp1[77],pp2[77],pp3[77],pp4[77],pp5[77],pp6[77],pp7[77],pp8[77],pp9[77],pp78[9],pp80[8],pp82[7],pp84[6],pp86[5],pp88[4],pp90[3],pp92[2],pp94[1],pp96[0],s10[24],s11[24],s12[24],s13[24],s14[24],s15[24],s16[24],s17[24],s18[24],s19[24],s20[24],s21[24],s22[24],s23[24],s24[24],s25[24],s26[24],s27[24],s28[24],s29[24],s30[24],s31[24],s32[24],s33[24],s34[24],s35[24],s36[24],s37[24],s38[24],s39[24],s40[24],s41[24],s40[26],s39[28],s38[30],s36[33],s34[36],s32[39],s30[42],s28[45],s26[48],s24[51],s22[54],s20[57],s18[60],s16[63],s14[66],s12[69],s10[72],s78[101],s77[103],s76[105],s75[107],s74[109],s73[111],s72[113],s71[115],s70[117],s69[119],s68[121],s67[123],s66[125],s65[127],pp99[61],pp98[63],pp97[65],pp96[67],pp95[69],pp94[71],pp93[73],pp92[75],pp91[77],pp90[79],pp89[81],pp88[83],pp87[85],pp86[87],pp85[89],pp84[91],pp83[93],pp82[95],pp81[97],pp80[99],pp126[54],pp124[57],pp122[60],pp120[63],pp118[66],pp116[69],pp114[72],pp112[75],pp110[78],pp108[81],pp106[84],pp104[87],pp102[90],pp102[91],pp102[92],pp102[93],pp102[94],pp102[95],pp102[96],pp102[97],pp103[97],pp104[97],pp105[97],pp106[97],pp107[97],pp108[97],pp109[97],pp110[97],pp111[97]};
    assign in80_2 = {pp3[44],pp2[46],pp1[48],pp0[50],pp41[10],pp41[11],pp41[12],pp41[13],pp41[14],pp41[15],pp41[16],pp41[17],pp41[18],pp41[19],pp41[20],pp41[21],pp41[22],pp43[21],pp45[20],pp47[19],pp49[18],pp51[17],pp53[16],pp55[15],pp57[14],pp59[13],pp61[12],pp63[11],pp65[10],pp0[76],pp1[76],pp2[76],pp3[76],pp4[76],pp5[76],pp6[76],pp7[76],pp8[76],pp9[76],pp77[9],pp79[8],pp81[7],pp83[6],pp85[5],pp87[4],pp89[3],pp91[2],pp93[1],pp95[0],s10[23],s11[23],s12[23],s13[23],s14[23],s15[23],s16[23],s17[23],s18[23],s19[23],s20[23],s21[23],s22[23],s23[23],s24[23],s25[23],s26[23],s27[23],s28[23],s29[23],s30[23],s31[23],s32[23],s33[23],s34[23],s35[23],s36[23],s37[23],s38[23],s39[23],s40[23],s41[23],s42[23],s41[25],s40[27],s39[29],s37[32],s35[35],s33[38],s31[41],s29[44],s27[47],s25[50],s23[53],s21[56],s19[59],s17[62],s15[65],s13[68],s11[71],s79[100],s78[102],s77[104],s76[106],s75[108],s74[110],s73[112],s72[114],s71[116],s70[118],s69[120],s68[122],s67[124],s66[126],s65[128],pp99[62],pp98[64],pp97[66],pp96[68],pp95[70],pp94[72],pp93[74],pp92[76],pp91[78],pp90[80],pp89[82],pp88[84],pp87[86],pp86[88],pp85[90],pp84[92],pp83[94],pp82[96],pp81[98],pp127[53],pp125[56],pp123[59],pp121[62],pp119[65],pp117[68],pp115[71],pp113[74],pp111[77],pp109[80],pp107[83],pp105[86],pp103[89],pp103[90],pp103[91],pp103[92],pp103[93],pp103[94],pp103[95],pp103[96],pp104[96],pp105[96],pp106[96],pp107[96],pp108[96],pp109[96],pp110[96],pp111[96],pp112[96]};
    CLA_162 KS_80(s80, c80, in80_1, in80_2);
    wire[159:0] s81, in81_1, in81_2;
    wire c81;
    assign in81_1 = {pp3[45],pp2[47],pp1[49],pp0[51],pp42[10],pp42[11],pp42[12],pp42[13],pp42[14],pp42[15],pp42[16],pp42[17],pp42[18],pp42[19],pp42[20],pp42[21],pp44[20],pp46[19],pp48[18],pp50[17],pp52[16],pp54[15],pp56[14],pp58[13],pp60[12],pp62[11],pp64[10],pp0[75],pp1[75],pp2[75],pp3[75],pp4[75],pp5[75],pp6[75],pp7[75],pp8[75],pp9[75],pp76[9],pp78[8],pp80[7],pp82[6],pp84[5],pp86[4],pp88[3],pp90[2],pp92[1],pp94[0],s10[22],s11[22],s12[22],s13[22],s14[22],s15[22],s16[22],s17[22],s18[22],s19[22],s20[22],s21[22],s22[22],s23[22],s24[22],s25[22],s26[22],s27[22],s28[22],s29[22],s30[22],s31[22],s32[22],s33[22],s34[22],s35[22],s36[22],s37[22],s38[22],s39[22],s40[22],s41[22],s42[22],s43[22],s42[24],s41[26],s40[28],s38[31],s36[34],s34[37],s32[40],s30[43],s28[46],s26[49],s24[52],s22[55],s20[58],s18[61],s16[64],s14[67],s12[70],s10[73],s79[101],s78[103],s77[105],s76[107],s75[109],s74[111],s73[113],s72[115],s71[117],s70[119],s69[121],s68[123],s67[125],s66[127],s65[129],pp99[63],pp98[65],pp97[67],pp96[69],pp95[71],pp94[73],pp93[75],pp92[77],pp91[79],pp90[81],pp89[83],pp88[85],pp87[87],pp86[89],pp85[91],pp84[93],pp83[95],pp82[97],pp81[99],pp126[55],pp124[58],pp122[61],pp120[64],pp118[67],pp116[70],pp114[73],pp112[76],pp110[79],pp108[82],pp106[85],pp104[88],pp104[89],pp104[90],pp104[91],pp104[92],pp104[93],pp104[94],pp104[95],pp105[95],pp106[95],pp107[95],pp108[95],pp109[95],pp110[95],pp111[95],pp112[95]};
    assign in81_2 = {pp4[44],pp3[46],pp2[48],pp1[50],pp0[52],pp43[10],pp43[11],pp43[12],pp43[13],pp43[14],pp43[15],pp43[16],pp43[17],pp43[18],pp43[19],pp43[20],pp45[19],pp47[18],pp49[17],pp51[16],pp53[15],pp55[14],pp57[13],pp59[12],pp61[11],pp63[10],pp0[74],pp1[74],pp2[74],pp3[74],pp4[74],pp5[74],pp6[74],pp7[74],pp8[74],pp9[74],pp75[9],pp77[8],pp79[7],pp81[6],pp83[5],pp85[4],pp87[3],pp89[2],pp91[1],pp93[0],s10[21],s11[21],s12[21],s13[21],s14[21],s15[21],s16[21],s17[21],s18[21],s19[21],s20[21],s21[21],s22[21],s23[21],s24[21],s25[21],s26[21],s27[21],s28[21],s29[21],s30[21],s31[21],s32[21],s33[21],s34[21],s35[21],s36[21],s37[21],s38[21],s39[21],s40[21],s41[21],s42[21],s43[21],s44[21],s43[23],s42[25],s41[27],s39[30],s37[33],s35[36],s33[39],s31[42],s29[45],s27[48],s25[51],s23[54],s21[57],s19[60],s17[63],s15[66],s13[69],s11[72],s80[100],s79[102],s78[104],s77[106],s76[108],s75[110],s74[112],s73[114],s72[116],s71[118],s70[120],s69[122],s68[124],s67[126],s66[128],s65[130],pp99[64],pp98[66],pp97[68],pp96[70],pp95[72],pp94[74],pp93[76],pp92[78],pp91[80],pp90[82],pp89[84],pp88[86],pp87[88],pp86[90],pp85[92],pp84[94],pp83[96],pp82[98],pp127[54],pp125[57],pp123[60],pp121[63],pp119[66],pp117[69],pp115[72],pp113[75],pp111[78],pp109[81],pp107[84],pp105[87],pp105[88],pp105[89],pp105[90],pp105[91],pp105[92],pp105[93],pp105[94],pp106[94],pp107[94],pp108[94],pp109[94],pp110[94],pp111[94],pp112[94],pp113[94]};
    CLA_160 KS_81(s81, c81, in81_1, in81_2);
    wire[157:0] s82, in82_1, in82_2;
    wire c82;
    assign in82_1 = {pp4[45],pp3[47],pp2[49],pp1[51],pp0[53],pp44[10],pp44[11],pp44[12],pp44[13],pp44[14],pp44[15],pp44[16],pp44[17],pp44[18],pp44[19],pp46[18],pp48[17],pp50[16],pp52[15],pp54[14],pp56[13],pp58[12],pp60[11],pp62[10],pp0[73],pp1[73],pp2[73],pp3[73],pp4[73],pp5[73],pp6[73],pp7[73],pp8[73],pp9[73],pp74[9],pp76[8],pp78[7],pp80[6],pp82[5],pp84[4],pp86[3],pp88[2],pp90[1],pp92[0],s10[20],s11[20],s12[20],s13[20],s14[20],s15[20],s16[20],s17[20],s18[20],s19[20],s20[20],s21[20],s22[20],s23[20],s24[20],s25[20],s26[20],s27[20],s28[20],s29[20],s30[20],s31[20],s32[20],s33[20],s34[20],s35[20],s36[20],s37[20],s38[20],s39[20],s40[20],s41[20],s42[20],s43[20],s44[20],s45[20],s44[22],s43[24],s42[26],s40[29],s38[32],s36[35],s34[38],s32[41],s30[44],s28[47],s26[50],s24[53],s22[56],s20[59],s18[62],s16[65],s14[68],s12[71],s10[74],s80[101],s79[103],s78[105],s77[107],s76[109],s75[111],s74[113],s73[115],s72[117],s71[119],s70[121],s69[123],s68[125],s67[127],s66[129],s65[131],pp99[65],pp98[67],pp97[69],pp96[71],pp95[73],pp94[75],pp93[77],pp92[79],pp91[81],pp90[83],pp89[85],pp88[87],pp87[89],pp86[91],pp85[93],pp84[95],pp83[97],pp82[99],pp126[56],pp124[59],pp122[62],pp120[65],pp118[68],pp116[71],pp114[74],pp112[77],pp110[80],pp108[83],pp106[86],pp106[87],pp106[88],pp106[89],pp106[90],pp106[91],pp106[92],pp106[93],pp107[93],pp108[93],pp109[93],pp110[93],pp111[93],pp112[93],pp113[93]};
    assign in82_2 = {pp5[44],pp4[46],pp3[48],pp2[50],pp1[52],pp0[54],pp45[10],pp45[11],pp45[12],pp45[13],pp45[14],pp45[15],pp45[16],pp45[17],pp45[18],pp47[17],pp49[16],pp51[15],pp53[14],pp55[13],pp57[12],pp59[11],pp61[10],pp0[72],pp1[72],pp2[72],pp3[72],pp4[72],pp5[72],pp6[72],pp7[72],pp8[72],pp9[72],pp73[9],pp75[8],pp77[7],pp79[6],pp81[5],pp83[4],pp85[3],pp87[2],pp89[1],pp91[0],s10[19],s11[19],s12[19],s13[19],s14[19],s15[19],s16[19],s17[19],s18[19],s19[19],s20[19],s21[19],s22[19],s23[19],s24[19],s25[19],s26[19],s27[19],s28[19],s29[19],s30[19],s31[19],s32[19],s33[19],s34[19],s35[19],s36[19],s37[19],s38[19],s39[19],s40[19],s41[19],s42[19],s43[19],s44[19],s45[19],s46[19],s45[21],s44[23],s43[25],s41[28],s39[31],s37[34],s35[37],s33[40],s31[43],s29[46],s27[49],s25[52],s23[55],s21[58],s19[61],s17[64],s15[67],s13[70],s11[73],s81[100],s80[102],s79[104],s78[106],s77[108],s76[110],s75[112],s74[114],s73[116],s72[118],s71[120],s70[122],s69[124],s68[126],s67[128],s66[130],s65[132],pp99[66],pp98[68],pp97[70],pp96[72],pp95[74],pp94[76],pp93[78],pp92[80],pp91[82],pp90[84],pp89[86],pp88[88],pp87[90],pp86[92],pp85[94],pp84[96],pp83[98],pp127[55],pp125[58],pp123[61],pp121[64],pp119[67],pp117[70],pp115[73],pp113[76],pp111[79],pp109[82],pp107[85],pp107[86],pp107[87],pp107[88],pp107[89],pp107[90],pp107[91],pp107[92],pp108[92],pp109[92],pp110[92],pp111[92],pp112[92],pp113[92],pp114[92]};
    CLA_158 KS_82(s82, c82, in82_1, in82_2);
    wire[155:0] s83, in83_1, in83_2;
    wire c83;
    assign in83_1 = {pp5[45],pp4[47],pp3[49],pp2[51],pp1[53],pp0[55],pp46[10],pp46[11],pp46[12],pp46[13],pp46[14],pp46[15],pp46[16],pp46[17],pp48[16],pp50[15],pp52[14],pp54[13],pp56[12],pp58[11],pp60[10],pp0[71],pp1[71],pp2[71],pp3[71],pp4[71],pp5[71],pp6[71],pp7[71],pp8[71],pp9[71],pp72[9],pp74[8],pp76[7],pp78[6],pp80[5],pp82[4],pp84[3],pp86[2],pp88[1],pp90[0],s10[18],s11[18],s12[18],s13[18],s14[18],s15[18],s16[18],s17[18],s18[18],s19[18],s20[18],s21[18],s22[18],s23[18],s24[18],s25[18],s26[18],s27[18],s28[18],s29[18],s30[18],s31[18],s32[18],s33[18],s34[18],s35[18],s36[18],s37[18],s38[18],s39[18],s40[18],s41[18],s42[18],s43[18],s44[18],s45[18],s46[18],s47[18],s46[20],s45[22],s44[24],s42[27],s40[30],s38[33],s36[36],s34[39],s32[42],s30[45],s28[48],s26[51],s24[54],s22[57],s20[60],s18[63],s16[66],s14[69],s12[72],s10[75],s81[101],s80[103],s79[105],s78[107],s77[109],s76[111],s75[113],s74[115],s73[117],s72[119],s71[121],s70[123],s69[125],s68[127],s67[129],s66[131],s65[133],pp99[67],pp98[69],pp97[71],pp96[73],pp95[75],pp94[77],pp93[79],pp92[81],pp91[83],pp90[85],pp89[87],pp88[89],pp87[91],pp86[93],pp85[95],pp84[97],pp83[99],pp126[57],pp124[60],pp122[63],pp120[66],pp118[69],pp116[72],pp114[75],pp112[78],pp110[81],pp108[84],pp108[85],pp108[86],pp108[87],pp108[88],pp108[89],pp108[90],pp108[91],pp109[91],pp110[91],pp111[91],pp112[91],pp113[91],pp114[91]};
    assign in83_2 = {pp6[44],pp5[46],pp4[48],pp3[50],pp2[52],pp1[54],pp0[56],pp47[10],pp47[11],pp47[12],pp47[13],pp47[14],pp47[15],pp47[16],pp49[15],pp51[14],pp53[13],pp55[12],pp57[11],pp59[10],pp0[70],pp1[70],pp2[70],pp3[70],pp4[70],pp5[70],pp6[70],pp7[70],pp8[70],pp9[70],pp71[9],pp73[8],pp75[7],pp77[6],pp79[5],pp81[4],pp83[3],pp85[2],pp87[1],pp89[0],s10[17],s11[17],s12[17],s13[17],s14[17],s15[17],s16[17],s17[17],s18[17],s19[17],s20[17],s21[17],s22[17],s23[17],s24[17],s25[17],s26[17],s27[17],s28[17],s29[17],s30[17],s31[17],s32[17],s33[17],s34[17],s35[17],s36[17],s37[17],s38[17],s39[17],s40[17],s41[17],s42[17],s43[17],s44[17],s45[17],s46[17],s47[17],s48[17],s47[19],s46[21],s45[23],s43[26],s41[29],s39[32],s37[35],s35[38],s33[41],s31[44],s29[47],s27[50],s25[53],s23[56],s21[59],s19[62],s17[65],s15[68],s13[71],s11[74],s82[100],s81[102],s80[104],s79[106],s78[108],s77[110],s76[112],s75[114],s74[116],s73[118],s72[120],s71[122],s70[124],s69[126],s68[128],s67[130],s66[132],s65[134],pp99[68],pp98[70],pp97[72],pp96[74],pp95[76],pp94[78],pp93[80],pp92[82],pp91[84],pp90[86],pp89[88],pp88[90],pp87[92],pp86[94],pp85[96],pp84[98],pp127[56],pp125[59],pp123[62],pp121[65],pp119[68],pp117[71],pp115[74],pp113[77],pp111[80],pp109[83],pp109[84],pp109[85],pp109[86],pp109[87],pp109[88],pp109[89],pp109[90],pp110[90],pp111[90],pp112[90],pp113[90],pp114[90],pp115[90]};
    CLA_156 KS_83(s83, c83, in83_1, in83_2);
    wire[153:0] s84, in84_1, in84_2;
    wire c84;
    assign in84_1 = {pp6[45],pp5[47],pp4[49],pp3[51],pp2[53],pp1[55],pp0[57],pp48[10],pp48[11],pp48[12],pp48[13],pp48[14],pp48[15],pp50[14],pp52[13],pp54[12],pp56[11],pp58[10],pp0[69],pp1[69],pp2[69],pp3[69],pp4[69],pp5[69],pp6[69],pp7[69],pp8[69],pp9[69],pp70[9],pp72[8],pp74[7],pp76[6],pp78[5],pp80[4],pp82[3],pp84[2],pp86[1],pp88[0],s10[16],s11[16],s12[16],s13[16],s14[16],s15[16],s16[16],s17[16],s18[16],s19[16],s20[16],s21[16],s22[16],s23[16],s24[16],s25[16],s26[16],s27[16],s28[16],s29[16],s30[16],s31[16],s32[16],s33[16],s34[16],s35[16],s36[16],s37[16],s38[16],s39[16],s40[16],s41[16],s42[16],s43[16],s44[16],s45[16],s46[16],s47[16],s48[16],s49[16],s48[18],s47[20],s46[22],s44[25],s42[28],s40[31],s38[34],s36[37],s34[40],s32[43],s30[46],s28[49],s26[52],s24[55],s22[58],s20[61],s18[64],s16[67],s14[70],s12[73],s10[76],s82[101],s81[103],s80[105],s79[107],s78[109],s77[111],s76[113],s75[115],s74[117],s73[119],s72[121],s71[123],s70[125],s69[127],s68[129],s67[131],s66[133],s65[135],pp99[69],pp98[71],pp97[73],pp96[75],pp95[77],pp94[79],pp93[81],pp92[83],pp91[85],pp90[87],pp89[89],pp88[91],pp87[93],pp86[95],pp85[97],pp84[99],pp126[58],pp124[61],pp122[64],pp120[67],pp118[70],pp116[73],pp114[76],pp112[79],pp110[82],pp110[83],pp110[84],pp110[85],pp110[86],pp110[87],pp110[88],pp110[89],pp111[89],pp112[89],pp113[89],pp114[89],pp115[89]};
    assign in84_2 = {pp7[44],pp6[46],pp5[48],pp4[50],pp3[52],pp2[54],pp1[56],pp0[58],pp49[10],pp49[11],pp49[12],pp49[13],pp49[14],pp51[13],pp53[12],pp55[11],pp57[10],pp0[68],pp1[68],pp2[68],pp3[68],pp4[68],pp5[68],pp6[68],pp7[68],pp8[68],pp9[68],pp69[9],pp71[8],pp73[7],pp75[6],pp77[5],pp79[4],pp81[3],pp83[2],pp85[1],pp87[0],s10[15],s11[15],s12[15],s13[15],s14[15],s15[15],s16[15],s17[15],s18[15],s19[15],s20[15],s21[15],s22[15],s23[15],s24[15],s25[15],s26[15],s27[15],s28[15],s29[15],s30[15],s31[15],s32[15],s33[15],s34[15],s35[15],s36[15],s37[15],s38[15],s39[15],s40[15],s41[15],s42[15],s43[15],s44[15],s45[15],s46[15],s47[15],s48[15],s49[15],s50[15],s49[17],s48[19],s47[21],s45[24],s43[27],s41[30],s39[33],s37[36],s35[39],s33[42],s31[45],s29[48],s27[51],s25[54],s23[57],s21[60],s19[63],s17[66],s15[69],s13[72],s11[75],s83[100],s82[102],s81[104],s80[106],s79[108],s78[110],s77[112],s76[114],s75[116],s74[118],s73[120],s72[122],s71[124],s70[126],s69[128],s68[130],s67[132],s66[134],s65[136],pp99[70],pp98[72],pp97[74],pp96[76],pp95[78],pp94[80],pp93[82],pp92[84],pp91[86],pp90[88],pp89[90],pp88[92],pp87[94],pp86[96],pp85[98],pp127[57],pp125[60],pp123[63],pp121[66],pp119[69],pp117[72],pp115[75],pp113[78],pp111[81],pp111[82],pp111[83],pp111[84],pp111[85],pp111[86],pp111[87],pp111[88],pp112[88],pp113[88],pp114[88],pp115[88],pp116[88]};
    CLA_154 KS_84(s84, c84, in84_1, in84_2);
    wire[151:0] s85, in85_1, in85_2;
    wire c85;
    assign in85_1 = {pp7[45],pp6[47],pp5[49],pp4[51],pp3[53],pp2[55],pp1[57],pp0[59],pp50[10],pp50[11],pp50[12],pp50[13],pp52[12],pp54[11],pp56[10],pp0[67],pp1[67],pp2[67],pp3[67],pp4[67],pp5[67],pp6[67],pp7[67],pp8[67],pp9[67],pp68[9],pp70[8],pp72[7],pp74[6],pp76[5],pp78[4],pp80[3],pp82[2],pp84[1],pp86[0],s10[14],s11[14],s12[14],s13[14],s14[14],s15[14],s16[14],s17[14],s18[14],s19[14],s20[14],s21[14],s22[14],s23[14],s24[14],s25[14],s26[14],s27[14],s28[14],s29[14],s30[14],s31[14],s32[14],s33[14],s34[14],s35[14],s36[14],s37[14],s38[14],s39[14],s40[14],s41[14],s42[14],s43[14],s44[14],s45[14],s46[14],s47[14],s48[14],s49[14],s50[14],s51[14],s50[16],s49[18],s48[20],s46[23],s44[26],s42[29],s40[32],s38[35],s36[38],s34[41],s32[44],s30[47],s28[50],s26[53],s24[56],s22[59],s20[62],s18[65],s16[68],s14[71],s12[74],s10[77],s83[101],s82[103],s81[105],s80[107],s79[109],s78[111],s77[113],s76[115],s75[117],s74[119],s73[121],s72[123],s71[125],s70[127],s69[129],s68[131],s67[133],s66[135],s65[137],pp99[71],pp98[73],pp97[75],pp96[77],pp95[79],pp94[81],pp93[83],pp92[85],pp91[87],pp90[89],pp89[91],pp88[93],pp87[95],pp86[97],pp85[99],pp126[59],pp124[62],pp122[65],pp120[68],pp118[71],pp116[74],pp114[77],pp112[80],pp112[81],pp112[82],pp112[83],pp112[84],pp112[85],pp112[86],pp112[87],pp113[87],pp114[87],pp115[87],pp116[87]};
    assign in85_2 = {pp8[44],pp7[46],pp6[48],pp5[50],pp4[52],pp3[54],pp2[56],pp1[58],pp0[60],pp51[10],pp51[11],pp51[12],pp53[11],pp55[10],pp0[66],pp1[66],pp2[66],pp3[66],pp4[66],pp5[66],pp6[66],pp7[66],pp8[66],pp9[66],pp67[9],pp69[8],pp71[7],pp73[6],pp75[5],pp77[4],pp79[3],pp81[2],pp83[1],pp85[0],s10[13],s11[13],s12[13],s13[13],s14[13],s15[13],s16[13],s17[13],s18[13],s19[13],s20[13],s21[13],s22[13],s23[13],s24[13],s25[13],s26[13],s27[13],s28[13],s29[13],s30[13],s31[13],s32[13],s33[13],s34[13],s35[13],s36[13],s37[13],s38[13],s39[13],s40[13],s41[13],s42[13],s43[13],s44[13],s45[13],s46[13],s47[13],s48[13],s49[13],s50[13],s51[13],s52[13],s51[15],s50[17],s49[19],s47[22],s45[25],s43[28],s41[31],s39[34],s37[37],s35[40],s33[43],s31[46],s29[49],s27[52],s25[55],s23[58],s21[61],s19[64],s17[67],s15[70],s13[73],s11[76],s84[100],s83[102],s82[104],s81[106],s80[108],s79[110],s78[112],s77[114],s76[116],s75[118],s74[120],s73[122],s72[124],s71[126],s70[128],s69[130],s68[132],s67[134],s66[136],s65[138],pp99[72],pp98[74],pp97[76],pp96[78],pp95[80],pp94[82],pp93[84],pp92[86],pp91[88],pp90[90],pp89[92],pp88[94],pp87[96],pp86[98],pp127[58],pp125[61],pp123[64],pp121[67],pp119[70],pp117[73],pp115[76],pp113[79],pp113[80],pp113[81],pp113[82],pp113[83],pp113[84],pp113[85],pp113[86],pp114[86],pp115[86],pp116[86],pp117[86]};
    CLA_152 KS_85(s85, c85, in85_1, in85_2);
    wire[149:0] s86, in86_1, in86_2;
    wire c86;
    assign in86_1 = {pp8[45],pp7[47],pp6[49],pp5[51],pp4[53],pp3[55],pp2[57],pp1[59],pp0[61],pp52[10],pp52[11],pp54[10],pp0[65],pp1[65],pp2[65],pp3[65],pp4[65],pp5[65],pp6[65],pp7[65],pp8[65],pp9[65],pp66[9],pp68[8],pp70[7],pp72[6],pp74[5],pp76[4],pp78[3],pp80[2],pp82[1],pp84[0],s10[12],s11[12],s12[12],s13[12],s14[12],s15[12],s16[12],s17[12],s18[12],s19[12],s20[12],s21[12],s22[12],s23[12],s24[12],s25[12],s26[12],s27[12],s28[12],s29[12],s30[12],s31[12],s32[12],s33[12],s34[12],s35[12],s36[12],s37[12],s38[12],s39[12],s40[12],s41[12],s42[12],s43[12],s44[12],s45[12],s46[12],s47[12],s48[12],s49[12],s50[12],s51[12],s52[12],s53[12],s52[14],s51[16],s50[18],s48[21],s46[24],s44[27],s42[30],s40[33],s38[36],s36[39],s34[42],s32[45],s30[48],s28[51],s26[54],s24[57],s22[60],s20[63],s18[66],s16[69],s14[72],s12[75],s10[78],s84[101],s83[103],s82[105],s81[107],s80[109],s79[111],s78[113],s77[115],s76[117],s75[119],s74[121],s73[123],s72[125],s71[127],s70[129],s69[131],s68[133],s67[135],s66[137],s65[139],pp99[73],pp98[75],pp97[77],pp96[79],pp95[81],pp94[83],pp93[85],pp92[87],pp91[89],pp90[91],pp89[93],pp88[95],pp87[97],pp86[99],pp126[60],pp124[63],pp122[66],pp120[69],pp118[72],pp116[75],pp114[78],pp114[79],pp114[80],pp114[81],pp114[82],pp114[83],pp114[84],pp114[85],pp115[85],pp116[85],pp117[85]};
    assign in86_2 = {pp9[44],pp8[46],pp7[48],pp6[50],pp5[52],pp4[54],pp3[56],pp2[58],pp1[60],pp0[62],pp53[10],pp0[64],pp1[64],pp2[64],pp3[64],pp4[64],pp5[64],pp6[64],pp7[64],pp8[64],pp9[64],pp65[9],pp67[8],pp69[7],pp71[6],pp73[5],pp75[4],pp77[3],pp79[2],pp81[1],pp83[0],s10[11],s11[11],s12[11],s13[11],s14[11],s15[11],s16[11],s17[11],s18[11],s19[11],s20[11],s21[11],s22[11],s23[11],s24[11],s25[11],s26[11],s27[11],s28[11],s29[11],s30[11],s31[11],s32[11],s33[11],s34[11],s35[11],s36[11],s37[11],s38[11],s39[11],s40[11],s41[11],s42[11],s43[11],s44[11],s45[11],s46[11],s47[11],s48[11],s49[11],s50[11],s51[11],s52[11],s53[11],s54[11],s53[13],s52[15],s51[17],s49[20],s47[23],s45[26],s43[29],s41[32],s39[35],s37[38],s35[41],s33[44],s31[47],s29[50],s27[53],s25[56],s23[59],s21[62],s19[65],s17[68],s15[71],s13[74],s11[77],s85[100],s84[102],s83[104],s82[106],s81[108],s80[110],s79[112],s78[114],s77[116],s76[118],s75[120],s74[122],s73[124],s72[126],s71[128],s70[130],s69[132],s68[134],s67[136],s66[138],s65[140],pp99[74],pp98[76],pp97[78],pp96[80],pp95[82],pp94[84],pp93[86],pp92[88],pp91[90],pp90[92],pp89[94],pp88[96],pp87[98],pp127[59],pp125[62],pp123[65],pp121[68],pp119[71],pp117[74],pp115[77],pp115[78],pp115[79],pp115[80],pp115[81],pp115[82],pp115[83],pp115[84],pp116[84],pp117[84],pp118[84]};
    CLA_150 KS_86(s86, c86, in86_1, in86_2);
    wire[147:0] s87, in87_1, in87_2;
    wire c87;
    assign in87_1 = {pp9[45],pp8[47],pp7[49],pp6[51],pp5[53],pp4[55],pp3[57],pp2[59],pp1[61],pp0[63],pp1[63],pp2[63],pp3[63],pp4[63],pp5[63],pp6[63],pp7[63],pp8[63],pp9[63],pp64[9],pp66[8],pp68[7],pp70[6],pp72[5],pp74[4],pp76[3],pp78[2],pp80[1],pp82[0],s10[10],s11[10],s12[10],s13[10],s14[10],s15[10],s16[10],s17[10],s18[10],s19[10],s20[10],s21[10],s22[10],s23[10],s24[10],s25[10],s26[10],s27[10],s28[10],s29[10],s30[10],s31[10],s32[10],s33[10],s34[10],s35[10],s36[10],s37[10],s38[10],s39[10],s40[10],s41[10],s42[10],s43[10],s44[10],s45[10],s46[10],s47[10],s48[10],s49[10],s50[10],s51[10],s52[10],s53[10],s54[10],s55[10],s54[12],s53[14],s52[16],s50[19],s48[22],s46[25],s44[28],s42[31],s40[34],s38[37],s36[40],s34[43],s32[46],s30[49],s28[52],s26[55],s24[58],s22[61],s20[64],s18[67],s16[70],s14[73],s12[76],s10[79],s85[101],s84[103],s83[105],s82[107],s81[109],s80[111],s79[113],s78[115],s77[117],s76[119],s75[121],s74[123],s73[125],s72[127],s71[129],s70[131],s69[133],s68[135],s67[137],s66[139],s10[100],pp99[75],pp98[77],pp97[79],pp96[81],pp95[83],pp94[85],pp93[87],pp92[89],pp91[91],pp90[93],pp89[95],pp88[97],pp87[99],pp126[61],pp124[64],pp122[67],pp120[70],pp118[73],pp116[76],pp116[77],pp116[78],pp116[79],pp116[80],pp116[81],pp116[82],pp116[83],pp117[83],pp118[83]};
    assign in87_2 = {pp45[9],pp9[46],pp8[48],pp7[50],pp6[52],pp5[54],pp4[56],pp3[58],pp2[60],pp1[62],pp2[62],pp3[62],pp4[62],pp5[62],pp6[62],pp7[62],pp8[62],pp9[62],pp63[9],pp65[8],pp67[7],pp69[6],pp71[5],pp73[4],pp75[3],pp77[2],pp79[1],pp81[0],s65[50],s65[51],s65[52],s65[53],s65[54],s65[55],s65[56],s65[57],s65[58],s65[59],s65[60],s65[61],s65[62],s65[63],s65[64],s65[65],s65[66],s65[67],s65[68],s65[69],s65[70],s65[71],s65[72],s65[73],s65[74],s65[75],s65[76],s65[77],s65[78],s65[79],s65[80],s65[81],s65[82],s65[83],s65[84],s65[85],s65[86],s65[87],s65[88],s65[89],s65[90],s65[91],s65[92],s65[93],s65[94],s65[95],s65[96],s55[11],s54[13],s53[15],s51[18],s49[21],s47[24],s45[27],s43[30],s41[33],s39[36],s37[39],s35[42],s33[45],s31[48],s29[51],s27[54],s25[57],s23[60],s21[63],s19[66],s17[69],s15[72],s13[75],s11[78],s86[100],s85[102],s84[104],s83[106],s82[108],s81[110],s80[112],s79[114],s78[116],s77[118],s76[120],s75[122],s74[124],s73[126],s72[128],s71[130],s70[132],s69[134],s68[136],s67[138],s65[141],s10[101],pp99[76],pp98[78],pp97[80],pp96[82],pp95[84],pp94[86],pp93[88],pp92[90],pp91[92],pp90[94],pp89[96],pp88[98],pp127[60],pp125[63],pp123[66],pp121[69],pp119[72],pp117[75],pp117[76],pp117[77],pp117[78],pp117[79],pp117[80],pp117[81],pp117[82],pp118[82],pp119[82]};
    CLA_148 KS_87(s87, c87, in87_1, in87_2);
    wire[145:0] s88, in88_1, in88_2;
    wire c88;
    assign in88_1 = {pp46[9],pp9[47],pp8[49],pp7[51],pp6[53],pp5[55],pp4[57],pp3[59],pp2[61],pp3[61],pp4[61],pp5[61],pp6[61],pp7[61],pp8[61],pp9[61],pp62[9],pp64[8],pp66[7],pp68[6],pp70[5],pp72[4],pp74[3],pp76[2],pp78[1],pp80[0],s65[49],s66[49],s66[50],s66[51],s66[52],s66[53],s66[54],s66[55],s66[56],s66[57],s66[58],s66[59],s66[60],s66[61],s66[62],s66[63],s66[64],s66[65],s66[66],s66[67],s66[68],s66[69],s66[70],s66[71],s66[72],s66[73],s66[74],s66[75],s66[76],s66[77],s66[78],s66[79],s66[80],s66[81],s66[82],s66[83],s66[84],s66[85],s66[86],s66[87],s66[88],s66[89],s66[90],s66[91],s66[92],s66[93],s66[94],s66[95],s56[10],s55[12],s54[14],s52[17],s50[20],s48[23],s46[26],s44[29],s42[32],s40[35],s38[38],s36[41],s34[44],s32[47],s30[50],s28[53],s26[56],s24[59],s22[62],s20[65],s18[68],s16[71],s14[74],s12[77],s10[80],s86[101],s85[103],s84[105],s83[107],s82[109],s81[111],s80[113],s79[115],s78[117],s77[119],s76[121],s75[123],s74[125],s73[127],s72[129],s71[131],s70[133],s69[135],s68[137],s66[140],s11[100],s10[102],pp99[77],pp98[79],pp97[81],pp96[83],pp95[85],pp94[87],pp93[89],pp92[91],pp91[93],pp90[95],pp89[97],pp88[99],pp126[62],pp124[65],pp122[68],pp120[71],pp118[74],pp118[75],pp118[76],pp118[77],pp118[78],pp118[79],pp118[80],pp118[81],pp119[81]};
    assign in88_2 = {pp47[8],pp47[9],pp9[48],pp8[50],pp7[52],pp6[54],pp5[56],pp4[58],pp3[60],pp4[60],pp5[60],pp6[60],pp7[60],pp8[60],pp9[60],pp61[9],pp63[8],pp65[7],pp67[6],pp69[5],pp71[4],pp73[3],pp75[2],pp77[1],pp79[0],s65[48],s66[48],s67[48],s67[49],s67[50],s67[51],s67[52],s67[53],s67[54],s67[55],s67[56],s67[57],s67[58],s67[59],s67[60],s67[61],s67[62],s67[63],s67[64],s67[65],s67[66],s67[67],s67[68],s67[69],s67[70],s67[71],s67[72],s67[73],s67[74],s67[75],s67[76],s67[77],s67[78],s67[79],s67[80],s67[81],s67[82],s67[83],s67[84],s67[85],s67[86],s67[87],s67[88],s67[89],s67[90],s67[91],s67[92],s67[93],s67[94],s65[97],s56[11],s55[13],s53[16],s51[19],s49[22],s47[25],s45[28],s43[31],s41[34],s39[37],s37[40],s35[43],s33[46],s31[49],s29[52],s27[55],s25[58],s23[61],s21[64],s19[67],s17[70],s15[73],s13[76],s11[79],s87[100],s86[102],s85[104],s84[106],s83[108],s82[110],s81[112],s80[114],s79[116],s78[118],s77[120],s76[122],s75[124],s74[126],s73[128],s72[130],s71[132],s70[134],s69[136],s67[139],s65[142],s11[101],s10[103],pp99[78],pp98[80],pp97[82],pp96[84],pp95[86],pp94[88],pp93[90],pp92[92],pp91[94],pp90[96],pp89[98],pp127[61],pp125[64],pp123[67],pp121[70],pp119[73],pp119[74],pp119[75],pp119[76],pp119[77],pp119[78],pp119[79],pp119[80],pp120[80]};
    CLA_146 KS_88(s88, c88, in88_1, in88_2);
    wire[143:0] s89, in89_1, in89_2;
    wire c89;
    assign in89_1 = {pp48[8],pp48[9],pp9[49],pp8[51],pp7[53],pp6[55],pp5[57],pp4[59],pp5[59],pp6[59],pp7[59],pp8[59],pp9[59],pp60[9],pp62[8],pp64[7],pp66[6],pp68[5],pp70[4],pp72[3],pp74[2],pp76[1],pp78[0],s65[47],s66[47],s67[47],s68[47],s68[48],s68[49],s68[50],s68[51],s68[52],s68[53],s68[54],s68[55],s68[56],s68[57],s68[58],s68[59],s68[60],s68[61],s68[62],s68[63],s68[64],s68[65],s68[66],s68[67],s68[68],s68[69],s68[70],s68[71],s68[72],s68[73],s68[74],s68[75],s68[76],s68[77],s68[78],s68[79],s68[80],s68[81],s68[82],s68[83],s68[84],s68[85],s68[86],s68[87],s68[88],s68[89],s68[90],s68[91],s68[92],s68[93],s66[96],s57[10],s56[12],s54[15],s52[18],s50[21],s48[24],s46[27],s44[30],s42[33],s40[36],s38[39],s36[42],s34[45],s32[48],s30[51],s28[54],s26[57],s24[60],s22[63],s20[66],s18[69],s16[72],s14[75],s12[78],s10[81],s87[101],s86[103],s85[105],s84[107],s83[109],s82[111],s81[113],s80[115],s79[117],s78[119],s77[121],s76[123],s75[125],s74[127],s73[129],s72[131],s71[133],s70[135],s68[138],s66[141],s12[100],s11[102],s10[104],pp99[79],pp98[81],pp97[83],pp96[85],pp95[87],pp94[89],pp93[91],pp92[93],pp91[95],pp90[97],pp89[99],pp126[63],pp124[66],pp122[69],pp120[72],pp120[73],pp120[74],pp120[75],pp120[76],pp120[77],pp120[78],pp120[79]};
    assign in89_2 = {pp49[7],pp49[8],pp49[9],pp9[50],pp8[52],pp7[54],pp6[56],pp5[58],pp6[58],pp7[58],pp8[58],pp9[58],pp59[9],pp61[8],pp63[7],pp65[6],pp67[5],pp69[4],pp71[3],pp73[2],pp75[1],pp77[0],s65[46],s66[46],s67[46],s68[46],s69[46],s69[47],s69[48],s69[49],s69[50],s69[51],s69[52],s69[53],s69[54],s69[55],s69[56],s69[57],s69[58],s69[59],s69[60],s69[61],s69[62],s69[63],s69[64],s69[65],s69[66],s69[67],s69[68],s69[69],s69[70],s69[71],s69[72],s69[73],s69[74],s69[75],s69[76],s69[77],s69[78],s69[79],s69[80],s69[81],s69[82],s69[83],s69[84],s69[85],s69[86],s69[87],s69[88],s69[89],s69[90],s69[91],s69[92],s67[95],s65[98],s57[11],s55[14],s53[17],s51[20],s49[23],s47[26],s45[29],s43[32],s41[35],s39[38],s37[41],s35[44],s33[47],s31[50],s29[53],s27[56],s25[59],s23[62],s21[65],s19[68],s17[71],s15[74],s13[77],s11[80],s88[100],s87[102],s86[104],s85[106],s84[108],s83[110],s82[112],s81[114],s80[116],s79[118],s78[120],s77[122],s76[124],s75[126],s74[128],s73[130],s72[132],s71[134],s69[137],s67[140],s65[143],s12[101],s11[103],s10[105],pp99[80],pp98[82],pp97[84],pp96[86],pp95[88],pp94[90],pp93[92],pp92[94],pp91[96],pp90[98],pp127[62],pp125[65],pp123[68],pp121[71],pp121[72],pp121[73],pp121[74],pp121[75],pp121[76],pp121[77],pp121[78]};
    CLA_144 KS_89(s89, c89, in89_1, in89_2);
    wire[141:0] s90, in90_1, in90_2;
    wire c90;
    assign in90_1 = {pp50[7],pp50[8],pp50[9],pp9[51],pp8[53],pp7[55],pp6[57],pp7[57],pp8[57],pp9[57],pp58[9],pp60[8],pp62[7],pp64[6],pp66[5],pp68[4],pp70[3],pp72[2],pp74[1],pp76[0],s65[45],s66[45],s67[45],s68[45],s69[45],s70[45],s70[46],s70[47],s70[48],s70[49],s70[50],s70[51],s70[52],s70[53],s70[54],s70[55],s70[56],s70[57],s70[58],s70[59],s70[60],s70[61],s70[62],s70[63],s70[64],s70[65],s70[66],s70[67],s70[68],s70[69],s70[70],s70[71],s70[72],s70[73],s70[74],s70[75],s70[76],s70[77],s70[78],s70[79],s70[80],s70[81],s70[82],s70[83],s70[84],s70[85],s70[86],s70[87],s70[88],s70[89],s70[90],s70[91],s68[94],s66[97],s58[10],s56[13],s54[16],s52[19],s50[22],s48[25],s46[28],s44[31],s42[34],s40[37],s38[40],s36[43],s34[46],s32[49],s30[52],s28[55],s26[58],s24[61],s22[64],s20[67],s18[70],s16[73],s14[76],s12[79],s10[82],s88[101],s87[103],s86[105],s85[107],s84[109],s83[111],s82[113],s81[115],s80[117],s79[119],s78[121],s77[123],s76[125],s75[127],s74[129],s73[131],s72[133],s70[136],s68[139],s66[142],s13[100],s12[102],s11[104],s10[106],pp99[81],pp98[83],pp97[85],pp96[87],pp95[89],pp94[91],pp93[93],pp92[95],pp91[97],pp90[99],pp126[64],pp124[67],pp122[70],pp122[71],pp122[72],pp122[73],pp122[74],pp122[75],pp122[76]};
    assign in90_2 = {pp51[6],pp51[7],pp51[8],pp51[9],pp9[52],pp8[54],pp7[56],pp8[56],pp9[56],pp57[9],pp59[8],pp61[7],pp63[6],pp65[5],pp67[4],pp69[3],pp71[2],pp73[1],pp75[0],s65[44],s66[44],s67[44],s68[44],s69[44],s70[44],s71[44],s71[45],s71[46],s71[47],s71[48],s71[49],s71[50],s71[51],s71[52],s71[53],s71[54],s71[55],s71[56],s71[57],s71[58],s71[59],s71[60],s71[61],s71[62],s71[63],s71[64],s71[65],s71[66],s71[67],s71[68],s71[69],s71[70],s71[71],s71[72],s71[73],s71[74],s71[75],s71[76],s71[77],s71[78],s71[79],s71[80],s71[81],s71[82],s71[83],s71[84],s71[85],s71[86],s71[87],s71[88],s71[89],s71[90],s69[93],s67[96],s65[99],s57[12],s55[15],s53[18],s51[21],s49[24],s47[27],s45[30],s43[33],s41[36],s39[39],s37[42],s35[45],s33[48],s31[51],s29[54],s27[57],s25[60],s23[63],s21[66],s19[69],s17[72],s15[75],s13[78],s11[81],s89[100],s88[102],s87[104],s86[106],s85[108],s84[110],s83[112],s82[114],s81[116],s80[118],s79[120],s78[122],s77[124],s76[126],s75[128],s74[130],s73[132],s71[135],s69[138],s67[141],s65[144],s13[101],s12[103],s11[105],s10[107],pp99[82],pp98[84],pp97[86],pp96[88],pp95[90],pp94[92],pp93[94],pp92[96],pp91[98],pp127[63],pp125[66],pp123[69],pp123[70],pp123[71],pp123[72],pp123[73],pp123[74],pp123[75]};
    CLA_142 KS_90(s90, c90, in90_1, in90_2);
    wire[139:0] s91, in91_1, in91_2;
    wire c91;
    assign in91_1 = {pp52[6],pp52[7],pp52[8],pp52[9],pp9[53],pp8[55],pp9[55],pp56[9],pp58[8],pp60[7],pp62[6],pp64[5],pp66[4],pp68[3],pp70[2],pp72[1],pp74[0],s65[43],s66[43],s67[43],s68[43],s69[43],s70[43],s71[43],s72[43],s72[44],s72[45],s72[46],s72[47],s72[48],s72[49],s72[50],s72[51],s72[52],s72[53],s72[54],s72[55],s72[56],s72[57],s72[58],s72[59],s72[60],s72[61],s72[62],s72[63],s72[64],s72[65],s72[66],s72[67],s72[68],s72[69],s72[70],s72[71],s72[72],s72[73],s72[74],s72[75],s72[76],s72[77],s72[78],s72[79],s72[80],s72[81],s72[82],s72[83],s72[84],s72[85],s72[86],s72[87],s72[88],s72[89],s70[92],s68[95],s66[98],s58[11],s56[14],s54[17],s52[20],s50[23],s48[26],s46[29],s44[32],s42[35],s40[38],s38[41],s36[44],s34[47],s32[50],s30[53],s28[56],s26[59],s24[62],s22[65],s20[68],s18[71],s16[74],s14[77],s12[80],s10[83],s89[101],s88[103],s87[105],s86[107],s85[109],s84[111],s83[113],s82[115],s81[117],s80[119],s79[121],s78[123],s77[125],s76[127],s75[129],s74[131],s72[134],s70[137],s68[140],s66[143],s14[100],s13[102],s12[104],s11[106],s10[108],pp99[83],pp98[85],pp97[87],pp96[89],pp95[91],pp94[93],pp93[95],pp92[97],pp91[99],pp126[65],pp124[68],pp124[69],pp124[70],pp124[71],pp124[72],pp124[73]};
    assign in91_2 = {pp53[5],pp53[6],pp53[7],pp53[8],pp53[9],pp9[54],pp55[9],pp57[8],pp59[7],pp61[6],pp63[5],pp65[4],pp67[3],pp69[2],pp71[1],pp73[0],s65[42],s66[42],s67[42],s68[42],s69[42],s70[42],s71[42],s72[42],s73[42],s73[43],s73[44],s73[45],s73[46],s73[47],s73[48],s73[49],s73[50],s73[51],s73[52],s73[53],s73[54],s73[55],s73[56],s73[57],s73[58],s73[59],s73[60],s73[61],s73[62],s73[63],s73[64],s73[65],s73[66],s73[67],s73[68],s73[69],s73[70],s73[71],s73[72],s73[73],s73[74],s73[75],s73[76],s73[77],s73[78],s73[79],s73[80],s73[81],s73[82],s73[83],s73[84],s73[85],s73[86],s73[87],s73[88],s71[91],s69[94],s67[97],s59[10],s57[13],s55[16],s53[19],s51[22],s49[25],s47[28],s45[31],s43[34],s41[37],s39[40],s37[43],s35[46],s33[49],s31[52],s29[55],s27[58],s25[61],s23[64],s21[67],s19[70],s17[73],s15[76],s13[79],s11[82],s90[100],s89[102],s88[104],s87[106],s86[108],s85[110],s84[112],s83[114],s82[116],s81[118],s80[120],s79[122],s78[124],s77[126],s76[128],s75[130],s73[133],s71[136],s69[139],s67[142],s65[145],s14[101],s13[103],s12[105],s11[107],s10[109],pp99[84],pp98[86],pp97[88],pp96[90],pp95[92],pp94[94],pp93[96],pp92[98],pp127[64],pp125[67],pp125[68],pp125[69],pp125[70],pp125[71],pp125[72]};
    CLA_140 KS_91(s91, c91, in91_1, in91_2);
    wire[137:0] s92, in92_1, in92_2;
    wire c92;
    assign in92_1 = {pp54[5],pp54[6],pp54[7],pp54[8],pp54[9],pp56[8],pp58[7],pp60[6],pp62[5],pp64[4],pp66[3],pp68[2],pp70[1],pp72[0],s65[41],s66[41],s67[41],s68[41],s69[41],s70[41],s71[41],s72[41],s73[41],s74[41],s74[42],s74[43],s74[44],s74[45],s74[46],s74[47],s74[48],s74[49],s74[50],s74[51],s74[52],s74[53],s74[54],s74[55],s74[56],s74[57],s74[58],s74[59],s74[60],s74[61],s74[62],s74[63],s74[64],s74[65],s74[66],s74[67],s74[68],s74[69],s74[70],s74[71],s74[72],s74[73],s74[74],s74[75],s74[76],s74[77],s74[78],s74[79],s74[80],s74[81],s74[82],s74[83],s74[84],s74[85],s74[86],s74[87],s72[90],s70[93],s68[96],s66[99],s58[12],s56[15],s54[18],s52[21],s50[24],s48[27],s46[30],s44[33],s42[36],s40[39],s38[42],s36[45],s34[48],s32[51],s30[54],s28[57],s26[60],s24[63],s22[66],s20[69],s18[72],s16[75],s14[78],s12[81],s10[84],s90[101],s89[103],s88[105],s87[107],s86[109],s85[111],s84[113],s83[115],s82[117],s81[119],s80[121],s79[123],s78[125],s77[127],s76[129],s74[132],s72[135],s70[138],s68[141],s66[144],s65[146],s65[147],s65[148],s65[149],s65[150],s65[151],pp99[85],pp98[87],pp97[89],pp96[91],pp95[93],pp94[95],pp93[97],pp92[99],pp126[66],pp126[67],pp126[68],pp126[69],pp126[70]};
    assign in92_2 = {pp55[4],pp55[5],pp55[6],pp55[7],pp55[8],pp57[7],pp59[6],pp61[5],pp63[4],pp65[3],pp67[2],pp69[1],pp71[0],s65[40],s66[40],s67[40],s68[40],s69[40],s70[40],s71[40],s72[40],s73[40],s74[40],s75[40],s75[41],s75[42],s75[43],s75[44],s75[45],s75[46],s75[47],s75[48],s75[49],s75[50],s75[51],s75[52],s75[53],s75[54],s75[55],s75[56],s75[57],s75[58],s75[59],s75[60],s75[61],s75[62],s75[63],s75[64],s75[65],s75[66],s75[67],s75[68],s75[69],s75[70],s75[71],s75[72],s75[73],s75[74],s75[75],s75[76],s75[77],s75[78],s75[79],s75[80],s75[81],s75[82],s75[83],s75[84],s75[85],s75[86],s73[89],s71[92],s69[95],s67[98],s59[11],s57[14],s55[17],s53[20],s51[23],s49[26],s47[29],s45[32],s43[35],s41[38],s39[41],s37[44],s35[47],s33[50],s31[53],s29[56],s27[59],s25[62],s23[65],s21[68],s19[71],s17[74],s15[77],s13[80],s11[83],s91[100],s90[102],s89[104],s88[106],s87[108],s86[110],s85[112],s84[114],s83[116],s82[118],s81[120],s80[122],s79[124],s78[126],s77[128],s75[131],s73[134],s71[137],s69[140],s67[143],s66[145],s66[146],s66[147],s66[148],s66[149],s66[150],s65[152],pp99[86],pp98[88],pp97[90],pp96[92],pp95[94],pp94[96],pp93[98],pp127[65],pp127[66],pp127[67],pp127[68],pp127[69]};
    CLA_138 KS_92(s92, c92, in92_1, in92_2);
    wire[135:0] s93, in93_1, in93_2;
    wire c93;
    assign in93_1 = {pp56[4],pp56[5],pp56[6],pp56[7],pp58[6],pp60[5],pp62[4],pp64[3],pp66[2],pp68[1],pp70[0],s65[39],s66[39],s67[39],s68[39],s69[39],s70[39],s71[39],s72[39],s73[39],s74[39],s75[39],s76[39],s76[40],s76[41],s76[42],s76[43],s76[44],s76[45],s76[46],s76[47],s76[48],s76[49],s76[50],s76[51],s76[52],s76[53],s76[54],s76[55],s76[56],s76[57],s76[58],s76[59],s76[60],s76[61],s76[62],s76[63],s76[64],s76[65],s76[66],s76[67],s76[68],s76[69],s76[70],s76[71],s76[72],s76[73],s76[74],s76[75],s76[76],s76[77],s76[78],s76[79],s76[80],s76[81],s76[82],s76[83],s76[84],s76[85],s74[88],s72[91],s70[94],s68[97],s67[99],s58[13],s56[16],s54[19],s52[22],s50[25],s48[28],s46[31],s44[34],s42[37],s40[40],s38[43],s36[46],s34[49],s32[52],s30[55],s28[58],s26[61],s24[64],s22[67],s20[70],s18[73],s16[76],s14[79],s12[82],s10[85],s91[101],s90[103],s89[105],s88[107],s87[109],s86[111],s85[113],s84[115],s83[117],s82[119],s81[121],s80[123],s79[125],s78[127],s76[130],s74[133],s72[136],s70[139],s68[142],s67[144],s67[145],s67[146],s67[147],s67[148],s67[149],s66[151],s65[153],pp99[87],pp98[89],pp97[91],pp96[93],pp95[95],pp94[97],pp93[99],pp94[99],pp95[99],pp96[99]};
    assign in93_2 = {pp57[3],pp57[4],pp57[5],pp57[6],pp59[5],pp61[4],pp63[3],pp65[2],pp67[1],pp69[0],s65[38],s66[38],s67[38],s68[38],s69[38],s70[38],s71[38],s72[38],s73[38],s74[38],s75[38],s76[38],s77[38],s77[39],s77[40],s77[41],s77[42],s77[43],s77[44],s77[45],s77[46],s77[47],s77[48],s77[49],s77[50],s77[51],s77[52],s77[53],s77[54],s77[55],s77[56],s77[57],s77[58],s77[59],s77[60],s77[61],s77[62],s77[63],s77[64],s77[65],s77[66],s77[67],s77[68],s77[69],s77[70],s77[71],s77[72],s77[73],s77[74],s77[75],s77[76],s77[77],s77[78],s77[79],s77[80],s77[81],s77[82],s77[83],s77[84],s75[87],s73[90],s71[93],s69[96],s68[98],s68[99],s57[15],s55[18],s53[21],s51[24],s49[27],s47[30],s45[33],s43[36],s41[39],s39[42],s37[45],s35[48],s33[51],s31[54],s29[57],s27[60],s25[63],s23[66],s21[69],s19[72],s17[75],s15[78],s13[81],s11[84],s92[100],s91[102],s90[104],s89[106],s88[108],s87[110],s86[112],s85[114],s84[116],s83[118],s82[120],s81[122],s80[124],s79[126],s77[129],s75[132],s73[135],s71[138],s69[141],s68[143],s68[144],s68[145],s68[146],s68[147],s68[148],s67[150],s66[152],s65[154],pp99[88],pp98[90],pp97[92],pp96[94],pp95[96],pp94[98],pp95[98],pp96[98],pp97[98]};
    CLA_136 KS_93(s93, c93, in93_1, in93_2);
    wire[133:0] s94, in94_1, in94_2;
    wire c94;
    assign in94_1 = {pp58[3],pp58[4],pp58[5],pp60[4],pp62[3],pp64[2],pp66[1],pp68[0],s65[37],s66[37],s67[37],s68[37],s69[37],s70[37],s71[37],s72[37],s73[37],s74[37],s75[37],s76[37],s77[37],s78[37],s78[38],s78[39],s78[40],s78[41],s78[42],s78[43],s78[44],s78[45],s78[46],s78[47],s78[48],s78[49],s78[50],s78[51],s78[52],s78[53],s78[54],s78[55],s78[56],s78[57],s78[58],s78[59],s78[60],s78[61],s78[62],s78[63],s78[64],s78[65],s78[66],s78[67],s78[68],s78[69],s78[70],s78[71],s78[72],s78[73],s78[74],s78[75],s78[76],s78[77],s78[78],s78[79],s78[80],s78[81],s78[82],s78[83],s76[86],s74[89],s72[92],s70[95],s69[97],s69[98],s69[99],s56[17],s54[20],s52[23],s50[26],s48[29],s46[32],s44[35],s42[38],s40[41],s38[44],s36[47],s34[50],s32[53],s30[56],s28[59],s26[62],s24[65],s22[68],s20[71],s18[74],s16[77],s14[80],s12[83],s10[86],s92[101],s91[103],s90[105],s89[107],s88[109],s87[111],s86[113],s85[115],s84[117],s83[119],s82[121],s81[123],s80[125],s78[128],s76[131],s74[134],s72[137],s70[140],s69[142],s69[143],s69[144],s69[145],s69[146],s69[147],s68[149],s67[151],s66[153],s65[155],pp99[89],pp98[91],pp97[93],pp96[95],pp95[97],pp96[97],pp97[97]};
    assign in94_2 = {pp59[2],pp59[3],pp59[4],pp61[3],pp63[2],pp65[1],pp67[0],s65[36],s66[36],s67[36],s68[36],s69[36],s70[36],s71[36],s72[36],s73[36],s74[36],s75[36],s76[36],s77[36],s78[36],s79[36],s79[37],s79[38],s79[39],s79[40],s79[41],s79[42],s79[43],s79[44],s79[45],s79[46],s79[47],s79[48],s79[49],s79[50],s79[51],s79[52],s79[53],s79[54],s79[55],s79[56],s79[57],s79[58],s79[59],s79[60],s79[61],s79[62],s79[63],s79[64],s79[65],s79[66],s79[67],s79[68],s79[69],s79[70],s79[71],s79[72],s79[73],s79[74],s79[75],s79[76],s79[77],s79[78],s79[79],s79[80],s79[81],s79[82],s77[85],s75[88],s73[91],s71[94],s70[96],s70[97],s70[98],s70[99],s55[19],s53[22],s51[25],s49[28],s47[31],s45[34],s43[37],s41[40],s39[43],s37[46],s35[49],s33[52],s31[55],s29[58],s27[61],s25[64],s23[67],s21[70],s19[73],s17[76],s15[79],s13[82],s11[85],s93[100],s92[102],s91[104],s90[106],s89[108],s88[110],s87[112],s86[114],s85[116],s84[118],s83[120],s82[122],s81[124],s79[127],s77[130],s75[133],s73[136],s71[139],s70[141],s70[142],s70[143],s70[144],s70[145],s70[146],s69[148],s68[150],s67[152],s66[154],s65[156],pp99[90],pp98[92],pp97[94],pp96[96],pp97[96],pp98[96]};
    CLA_134 KS_94(s94, c94, in94_1, in94_2);
    wire[131:0] s95, in95_1, in95_2;
    wire c95;
    assign in95_1 = {pp60[2],pp60[3],pp62[2],pp64[1],pp66[0],s65[35],s66[35],s67[35],s68[35],s69[35],s70[35],s71[35],s72[35],s73[35],s74[35],s75[35],s76[35],s77[35],s78[35],s79[35],s80[35],s80[36],s80[37],s80[38],s80[39],s80[40],s80[41],s80[42],s80[43],s80[44],s80[45],s80[46],s80[47],s80[48],s80[49],s80[50],s80[51],s80[52],s80[53],s80[54],s80[55],s80[56],s80[57],s80[58],s80[59],s80[60],s80[61],s80[62],s80[63],s80[64],s80[65],s80[66],s80[67],s80[68],s80[69],s80[70],s80[71],s80[72],s80[73],s80[74],s80[75],s80[76],s80[77],s80[78],s80[79],s80[80],s80[81],s78[84],s76[87],s74[90],s72[93],s71[95],s71[96],s71[97],s71[98],s71[99],s54[21],s52[24],s50[27],s48[30],s46[33],s44[36],s42[39],s40[42],s38[45],s36[48],s34[51],s32[54],s30[57],s28[60],s26[63],s24[66],s22[69],s20[72],s18[75],s16[78],s14[81],s12[84],s10[87],s93[101],s92[103],s91[105],s90[107],s89[109],s88[111],s87[113],s86[115],s85[117],s84[119],s83[121],s82[123],s80[126],s78[129],s76[132],s74[135],s72[138],s71[140],s71[141],s71[142],s71[143],s71[144],s71[145],s70[147],s69[149],s68[151],s67[153],s66[155],s65[157],pp99[91],pp98[93],pp97[95],pp98[95]};
    assign in95_2 = {pp61[1],pp61[2],pp63[1],pp65[0],s65[34],s66[34],s67[34],s68[34],s69[34],s70[34],s71[34],s72[34],s73[34],s74[34],s75[34],s76[34],s77[34],s78[34],s79[34],s80[34],s81[34],s81[35],s81[36],s81[37],s81[38],s81[39],s81[40],s81[41],s81[42],s81[43],s81[44],s81[45],s81[46],s81[47],s81[48],s81[49],s81[50],s81[51],s81[52],s81[53],s81[54],s81[55],s81[56],s81[57],s81[58],s81[59],s81[60],s81[61],s81[62],s81[63],s81[64],s81[65],s81[66],s81[67],s81[68],s81[69],s81[70],s81[71],s81[72],s81[73],s81[74],s81[75],s81[76],s81[77],s81[78],s81[79],s81[80],s79[83],s77[86],s75[89],s73[92],s72[94],s72[95],s72[96],s72[97],s72[98],s72[99],s53[23],s51[26],s49[29],s47[32],s45[35],s43[38],s41[41],s39[44],s37[47],s35[50],s33[53],s31[56],s29[59],s27[62],s25[65],s23[68],s21[71],s19[74],s17[77],s15[80],s13[83],s11[86],s94[100],s93[102],s92[104],s91[106],s90[108],s89[110],s88[112],s87[114],s86[116],s85[118],s84[120],s83[122],s81[125],s79[128],s77[131],s75[134],s73[137],s72[139],s72[140],s72[141],s72[142],s72[143],s72[144],s71[146],s70[148],s69[150],s68[152],s67[154],s66[156],s65[158],pp99[92],pp98[94],pp99[94]};
    CLA_132 KS_95(s95, c95, in95_1, in95_2);
    wire[129:0] s96, in96_1, in96_2;
    wire c96;
    assign in96_1 = {pp62[1],pp64[0],s65[33],s66[33],s67[33],s68[33],s69[33],s70[33],s71[33],s72[33],s73[33],s74[33],s75[33],s76[33],s77[33],s78[33],s79[33],s80[33],s81[33],s82[33],s82[34],s82[35],s82[36],s82[37],s82[38],s82[39],s82[40],s82[41],s82[42],s82[43],s82[44],s82[45],s82[46],s82[47],s82[48],s82[49],s82[50],s82[51],s82[52],s82[53],s82[54],s82[55],s82[56],s82[57],s82[58],s82[59],s82[60],s82[61],s82[62],s82[63],s82[64],s82[65],s82[66],s82[67],s82[68],s82[69],s82[70],s82[71],s82[72],s82[73],s82[74],s82[75],s82[76],s82[77],s82[78],s82[79],s80[82],s78[85],s76[88],s74[91],s73[93],s73[94],s73[95],s73[96],s73[97],s73[98],s73[99],s52[25],s50[28],s48[31],s46[34],s44[37],s42[40],s40[43],s38[46],s36[49],s34[52],s32[55],s30[58],s28[61],s26[64],s24[67],s22[70],s20[73],s18[76],s16[79],s14[82],s12[85],s10[88],s94[101],s93[103],s92[105],s91[107],s90[109],s89[111],s88[113],s87[115],s86[117],s85[119],s84[121],s82[124],s80[127],s78[130],s76[133],s74[136],s73[138],s73[139],s73[140],s73[141],s73[142],s73[143],s72[145],s71[147],s70[149],s69[151],s68[153],s67[155],s66[157],s65[159],pp99[93]};
    assign in96_2 = {pp63[0],s65[32],s66[32],s67[32],s68[32],s69[32],s70[32],s71[32],s72[32],s73[32],s74[32],s75[32],s76[32],s77[32],s78[32],s79[32],s80[32],s81[32],s82[32],s83[32],s83[33],s83[34],s83[35],s83[36],s83[37],s83[38],s83[39],s83[40],s83[41],s83[42],s83[43],s83[44],s83[45],s83[46],s83[47],s83[48],s83[49],s83[50],s83[51],s83[52],s83[53],s83[54],s83[55],s83[56],s83[57],s83[58],s83[59],s83[60],s83[61],s83[62],s83[63],s83[64],s83[65],s83[66],s83[67],s83[68],s83[69],s83[70],s83[71],s83[72],s83[73],s83[74],s83[75],s83[76],s83[77],s83[78],s81[81],s79[84],s77[87],s75[90],s74[92],s74[93],s74[94],s74[95],s74[96],s74[97],s74[98],s74[99],s51[27],s49[30],s47[33],s45[36],s43[39],s41[42],s39[45],s37[48],s35[51],s33[54],s31[57],s29[60],s27[63],s25[66],s23[69],s21[72],s19[75],s17[78],s15[81],s13[84],s11[87],s95[100],s94[102],s93[104],s92[106],s91[108],s90[110],s89[112],s88[114],s87[116],s86[118],s85[120],s83[123],s81[126],s79[129],s77[132],s75[135],s74[137],s74[138],s74[139],s74[140],s74[141],s74[142],s73[144],s72[146],s71[148],s70[150],s69[152],s68[154],s67[156],s66[158],s65[160]};
    CLA_130 KS_96(s96, c96, in96_1, in96_2);

    /*Stage 3*/
    wire[223:0] s97, in97_1, in97_2;
    wire c97;
    assign in97_1 = {pp0[16],pp0[17],pp0[18],pp0[19],pp10[10],pp10[11],pp10[12],pp10[13],pp10[14],pp10[15],pp10[16],pp10[17],pp10[18],pp10[19],pp10[20],pp10[21],pp12[20],pp14[19],pp16[18],pp18[17],pp20[16],pp22[15],pp24[14],pp26[13],pp28[12],pp30[11],pp32[10],pp0[43],pp1[43],pp2[43],pp3[43],pp4[43],pp5[43],pp6[43],pp7[43],pp8[43],pp9[43],pp44[9],pp46[8],pp48[7],pp50[6],pp52[5],pp54[4],pp56[3],pp58[2],pp60[1],pp62[0],s65[31],s66[31],s67[31],s68[31],s69[31],s70[31],s71[31],s72[31],s73[31],s74[31],s75[31],s76[31],s77[31],s78[31],s79[31],s80[31],s81[31],s82[31],s83[31],s84[31],s84[32],s84[33],s84[34],s84[35],s84[36],s84[37],s84[38],s84[39],s84[40],s84[41],s84[42],s84[43],s84[44],s84[45],s84[46],s84[47],s84[48],s84[49],s84[50],s84[51],s84[52],s84[53],s84[54],s84[55],s84[56],s84[57],s84[58],s84[59],s84[60],s84[61],s84[62],s84[63],s84[64],s84[65],s84[66],s84[67],s84[68],s84[69],s84[70],s84[71],s84[72],s84[73],s84[74],s84[75],s84[76],s84[77],s82[80],s80[83],s78[86],s76[89],s75[91],s75[92],s75[93],s75[94],s75[95],s75[96],s75[97],s75[98],s75[99],s50[29],s48[32],s46[35],s44[38],s42[41],s40[44],s38[47],s36[50],s34[53],s32[56],s30[59],s28[62],s26[65],s24[68],s22[71],s20[74],s18[77],s16[80],s14[83],s12[86],s10[89],s95[101],s94[103],s93[105],s92[107],s91[109],s90[111],s89[113],s88[115],s87[117],s86[119],s84[122],s82[125],s80[128],s78[131],s76[134],s75[136],s75[137],s75[138],s75[139],s75[140],s75[141],s74[143],s73[145],s72[147],s71[149],s70[151],s69[153],s68[155],s67[157],s66[159],s65[161],pp99[95],pp98[97],pp97[99],pp126[71],pp124[74],pp122[77],pp121[79],pp120[81],pp119[83],pp118[85],pp117[87],pp116[89],pp115[91],pp114[93],pp113[95],pp112[97],pp111[99],pp98[113],pp96[116],pp94[119],pp92[122],pp90[125],pp116[100],pp114[103],pp112[106],pp110[109],pp108[112],pp106[115],pp104[118],pp102[121],pp100[124],pp100[125],pp100[126],pp100[127],pp101[127],pp102[127],pp103[127],pp104[127],pp105[127],pp106[127],pp107[127],pp108[127],pp109[127],pp110[127],pp111[127],pp112[127]};
    assign in97_2 = {pp1[15],pp1[16],pp1[17],pp1[18],pp0[20],pp11[10],pp11[11],pp11[12],pp11[13],pp11[14],pp11[15],pp11[16],pp11[17],pp11[18],pp11[19],pp11[20],pp13[19],pp15[18],pp17[17],pp19[16],pp21[15],pp23[14],pp25[13],pp27[12],pp29[11],pp31[10],pp0[42],pp1[42],pp2[42],pp3[42],pp4[42],pp5[42],pp6[42],pp7[42],pp8[42],pp9[42],pp43[9],pp45[8],pp47[7],pp49[6],pp51[5],pp53[4],pp55[3],pp57[2],pp59[1],pp61[0],s65[30],s66[30],s67[30],s68[30],s69[30],s70[30],s71[30],s72[30],s73[30],s74[30],s75[30],s76[30],s77[30],s78[30],s79[30],s80[30],s81[30],s82[30],s83[30],s84[30],s85[30],s85[31],s85[32],s85[33],s85[34],s85[35],s85[36],s85[37],s85[38],s85[39],s85[40],s85[41],s85[42],s85[43],s85[44],s85[45],s85[46],s85[47],s85[48],s85[49],s85[50],s85[51],s85[52],s85[53],s85[54],s85[55],s85[56],s85[57],s85[58],s85[59],s85[60],s85[61],s85[62],s85[63],s85[64],s85[65],s85[66],s85[67],s85[68],s85[69],s85[70],s85[71],s85[72],s85[73],s85[74],s85[75],s85[76],s83[79],s81[82],s79[85],s77[88],s76[90],s76[91],s76[92],s76[93],s76[94],s76[95],s76[96],s76[97],s76[98],s76[99],s49[31],s47[34],s45[37],s43[40],s41[43],s39[46],s37[49],s35[52],s33[55],s31[58],s29[61],s27[64],s25[67],s23[70],s21[73],s19[76],s17[79],s15[82],s13[85],s11[88],s96[100],s95[102],s94[104],s93[106],s92[108],s91[110],s90[112],s89[114],s88[116],s87[118],s85[121],s83[124],s81[127],s79[130],s77[133],s76[135],s76[136],s76[137],s76[138],s76[139],s76[140],s75[142],s74[144],s73[146],s72[148],s71[150],s70[152],s69[154],s68[156],s67[158],s66[160],s65[162],pp99[96],pp98[98],pp127[70],pp125[73],pp123[76],pp122[78],pp121[80],pp120[82],pp119[84],pp118[86],pp117[88],pp116[90],pp115[92],pp114[94],pp113[96],pp112[98],pp99[112],pp97[115],pp95[118],pp93[121],pp91[124],pp89[127],pp115[102],pp113[105],pp111[108],pp109[111],pp107[114],pp105[117],pp103[120],pp101[123],pp101[124],pp101[125],pp101[126],pp102[126],pp103[126],pp104[126],pp105[126],pp106[126],pp107[126],pp108[126],pp109[126],pp110[126],pp111[126],pp112[126],pp113[126]};
    CLA_224 KS_97(s97, c97, in97_1, in97_2);
    wire[221:0] s98, in98_1, in98_2;
    wire c98;
    assign in98_1 = {pp2[15],pp2[16],pp2[17],pp1[19],pp0[21],pp12[10],pp12[11],pp12[12],pp12[13],pp12[14],pp12[15],pp12[16],pp12[17],pp12[18],pp12[19],pp14[18],pp16[17],pp18[16],pp20[15],pp22[14],pp24[13],pp26[12],pp28[11],pp30[10],pp0[41],pp1[41],pp2[41],pp3[41],pp4[41],pp5[41],pp6[41],pp7[41],pp8[41],pp9[41],pp42[9],pp44[8],pp46[7],pp48[6],pp50[5],pp52[4],pp54[3],pp56[2],pp58[1],pp60[0],s65[29],s66[29],s67[29],s68[29],s69[29],s70[29],s71[29],s72[29],s73[29],s74[29],s75[29],s76[29],s77[29],s78[29],s79[29],s80[29],s81[29],s82[29],s83[29],s84[29],s85[29],s86[29],s86[30],s86[31],s86[32],s86[33],s86[34],s86[35],s86[36],s86[37],s86[38],s86[39],s86[40],s86[41],s86[42],s86[43],s86[44],s86[45],s86[46],s86[47],s86[48],s86[49],s86[50],s86[51],s86[52],s86[53],s86[54],s86[55],s86[56],s86[57],s86[58],s86[59],s86[60],s86[61],s86[62],s97[100],s97[101],s97[102],s97[103],s97[104],s97[105],s97[106],s97[107],s97[108],s97[109],s97[110],s97[111],s97[112],s97[113],s97[114],s97[115],s97[116],s97[117],s97[118],s97[119],s97[120],s97[121],s97[122],s97[123],s97[124],s97[125],s97[126],s97[127],s97[128],s97[129],s97[130],s97[131],s97[132],s97[133],s97[134],s97[135],s97[136],s97[137],s97[138],s97[139],s97[140],s97[141],s97[142],s97[143],s97[144],s97[145],s97[146],s97[147],s96[101],s95[103],s94[105],s93[107],s92[109],s91[111],s90[113],s89[115],s88[117],s86[120],s84[123],s82[126],s80[129],s78[132],s77[134],s77[135],s77[136],s77[137],s77[138],s77[139],s76[141],s75[143],s74[145],s73[147],s72[149],s71[151],s70[153],s69[155],s68[157],s67[159],s66[161],s65[163],pp99[97],pp98[99],pp126[72],pp124[75],pp123[77],pp122[79],pp121[81],pp120[83],pp119[85],pp118[87],pp117[89],pp116[91],pp115[93],pp114[95],pp113[97],pp112[99],pp98[114],pp96[117],pp94[120],pp92[123],pp90[126],pp116[101],pp114[104],pp112[107],pp110[110],pp108[113],pp106[116],pp104[119],pp102[122],pp102[123],pp102[124],pp102[125],pp103[125],pp104[125],pp105[125],pp106[125],pp107[125],pp108[125],pp109[125],pp110[125],pp111[125],pp112[125],pp113[125]};
    assign in98_2 = {pp3[14],pp3[15],pp3[16],pp2[18],pp1[20],pp0[22],pp13[10],pp13[11],pp13[12],pp13[13],pp13[14],pp13[15],pp13[16],pp13[17],pp13[18],pp15[17],pp17[16],pp19[15],pp21[14],pp23[13],pp25[12],pp27[11],pp29[10],pp0[40],pp1[40],pp2[40],pp3[40],pp4[40],pp5[40],pp6[40],pp7[40],pp8[40],pp9[40],pp41[9],pp43[8],pp45[7],pp47[6],pp49[5],pp51[4],pp53[3],pp55[2],pp57[1],pp59[0],s65[28],s66[28],s67[28],s68[28],s69[28],s70[28],s71[28],s72[28],s73[28],s74[28],s75[28],s76[28],s77[28],s78[28],s79[28],s80[28],s81[28],s82[28],s83[28],s84[28],s85[28],s86[28],s87[28],s87[29],s87[30],s87[31],s87[32],s87[33],s87[34],s87[35],s87[36],s87[37],s87[38],s87[39],s87[40],s87[41],s87[42],s87[43],s87[44],s87[45],s87[46],s87[47],s87[48],s87[49],s87[50],s87[51],s87[52],s87[53],s87[54],s87[55],s87[56],s87[57],s87[58],s87[59],s87[60],s87[61],s86[63],s86[64],s86[65],s86[66],s86[67],s86[68],s86[69],s86[70],s86[71],s86[72],s86[73],s86[74],s86[75],s84[78],s82[81],s80[84],s78[87],s77[89],s77[90],s77[91],s77[92],s77[93],s77[94],s77[95],s77[96],s77[97],s77[98],s77[99],s48[33],s46[36],s44[39],s42[42],s40[45],s38[48],s36[51],s34[54],s32[57],s30[60],s28[63],s26[66],s24[69],s22[72],s20[75],s18[78],s16[81],s14[84],s12[87],s10[90],s97[148],s96[102],s95[104],s94[106],s93[108],s92[110],s91[112],s90[114],s89[116],s87[119],s85[122],s83[125],s81[128],s79[131],s78[133],s78[134],s78[135],s78[136],s78[137],s78[138],s77[140],s76[142],s75[144],s74[146],s73[148],s72[150],s71[152],s70[154],s69[156],s68[158],s67[160],s66[162],s65[164],pp99[98],pp127[71],pp125[74],pp124[76],pp123[78],pp122[80],pp121[82],pp120[84],pp119[86],pp118[88],pp117[90],pp116[92],pp115[94],pp114[96],pp113[98],pp99[113],pp97[116],pp95[119],pp93[122],pp91[125],pp117[100],pp115[103],pp113[106],pp111[109],pp109[112],pp107[115],pp105[118],pp103[121],pp103[122],pp103[123],pp103[124],pp104[124],pp105[124],pp106[124],pp107[124],pp108[124],pp109[124],pp110[124],pp111[124],pp112[124],pp113[124],pp114[124]};
    CLA_222 KS_98(s98, c98, in98_1, in98_2);
    wire[219:0] s99, in99_1, in99_2;
    wire c99;
    assign in99_1 = {pp4[14],pp4[15],pp3[17],pp2[19],pp1[21],pp0[23],pp14[10],pp14[11],pp14[12],pp14[13],pp14[14],pp14[15],pp14[16],pp14[17],pp16[16],pp18[15],pp20[14],pp22[13],pp24[12],pp26[11],pp28[10],pp0[39],pp1[39],pp2[39],pp3[39],pp4[39],pp5[39],pp6[39],pp7[39],pp8[39],pp9[39],pp40[9],pp42[8],pp44[7],pp46[6],pp48[5],pp50[4],pp52[3],pp54[2],pp56[1],pp58[0],s65[27],s66[27],s67[27],s68[27],s69[27],s70[27],s71[27],s72[27],s73[27],s74[27],s75[27],s76[27],s77[27],s78[27],s79[27],s80[27],s81[27],s82[27],s83[27],s84[27],s85[27],s86[27],s87[27],s88[27],s88[28],s88[29],s88[30],s88[31],s88[32],s88[33],s88[34],s88[35],s88[36],s88[37],s88[38],s88[39],s88[40],s88[41],s88[42],s88[43],s88[44],s88[45],s88[46],s88[47],s88[48],s88[49],s88[50],s88[51],s88[52],s88[53],s88[54],s88[55],s88[56],s88[57],s88[58],s88[59],s88[60],s87[62],s98[100],s98[101],s98[102],s98[103],s98[104],s98[105],s98[106],s98[107],s98[108],s98[109],s98[110],s98[111],s98[112],s98[113],s98[114],s98[115],s98[116],s98[117],s98[118],s98[119],s98[120],s98[121],s98[122],s98[123],s98[124],s98[125],s98[126],s98[127],s98[128],s98[129],s98[130],s98[131],s98[132],s98[133],s98[134],s98[135],s98[136],s98[137],s98[138],s98[139],s98[140],s98[141],s98[142],s98[143],s98[144],s98[145],s98[146],s98[147],s97[149],s96[103],s95[105],s94[107],s93[109],s92[111],s91[113],s90[115],s88[118],s86[121],s84[124],s82[127],s80[130],s79[132],s79[133],s79[134],s79[135],s79[136],s79[137],s78[139],s77[141],s76[143],s75[145],s74[147],s73[149],s72[151],s71[153],s70[155],s69[157],s68[159],s67[161],s66[163],s65[165],pp99[99],pp126[73],pp125[75],pp124[77],pp123[79],pp122[81],pp121[83],pp120[85],pp119[87],pp118[89],pp117[91],pp116[93],pp115[95],pp114[97],pp113[99],pp98[115],pp96[118],pp94[121],pp92[124],pp90[127],pp116[102],pp114[105],pp112[108],pp110[111],pp108[114],pp106[117],pp104[120],pp104[121],pp104[122],pp104[123],pp105[123],pp106[123],pp107[123],pp108[123],pp109[123],pp110[123],pp111[123],pp112[123],pp113[123],pp114[123]};
    assign in99_2 = {pp5[13],pp5[14],pp4[16],pp3[18],pp2[20],pp1[22],pp0[24],pp15[10],pp15[11],pp15[12],pp15[13],pp15[14],pp15[15],pp15[16],pp17[15],pp19[14],pp21[13],pp23[12],pp25[11],pp27[10],pp0[38],pp1[38],pp2[38],pp3[38],pp4[38],pp5[38],pp6[38],pp7[38],pp8[38],pp9[38],pp39[9],pp41[8],pp43[7],pp45[6],pp47[5],pp49[4],pp51[3],pp53[2],pp55[1],pp57[0],s65[26],s66[26],s67[26],s68[26],s69[26],s70[26],s71[26],s72[26],s73[26],s74[26],s75[26],s76[26],s77[26],s78[26],s79[26],s80[26],s81[26],s82[26],s83[26],s84[26],s85[26],s86[26],s87[26],s88[26],s89[26],s89[27],s89[28],s89[29],s89[30],s89[31],s89[32],s89[33],s89[34],s89[35],s89[36],s89[37],s89[38],s89[39],s89[40],s89[41],s89[42],s89[43],s89[44],s89[45],s89[46],s89[47],s89[48],s89[49],s89[50],s89[51],s89[52],s89[53],s89[54],s89[55],s89[56],s89[57],s89[58],s89[59],s88[61],s87[63],s87[64],s87[65],s87[66],s87[67],s87[68],s87[69],s87[70],s87[71],s87[72],s87[73],s87[74],s85[77],s83[80],s81[83],s79[86],s78[88],s78[89],s78[90],s78[91],s78[92],s78[93],s78[94],s78[95],s78[96],s78[97],s78[98],s78[99],s47[35],s45[38],s43[41],s41[44],s39[47],s37[50],s35[53],s33[56],s31[59],s29[62],s27[65],s25[68],s23[71],s21[74],s19[77],s17[80],s15[83],s13[86],s11[89],s1[100],s98[148],s97[150],s96[104],s95[106],s94[108],s93[110],s92[112],s91[114],s89[117],s87[120],s85[123],s83[126],s81[129],s80[131],s80[132],s80[133],s80[134],s80[135],s80[136],s79[138],s78[140],s77[142],s76[144],s75[146],s74[148],s73[150],s72[152],s71[154],s70[156],s69[158],s68[160],s67[162],s66[164],s65[166],pp127[72],pp126[74],pp125[76],pp124[78],pp123[80],pp122[82],pp121[84],pp120[86],pp119[88],pp118[90],pp117[92],pp116[94],pp115[96],pp114[98],pp99[114],pp97[117],pp95[120],pp93[123],pp91[126],pp117[101],pp115[104],pp113[107],pp111[110],pp109[113],pp107[116],pp105[119],pp105[120],pp105[121],pp105[122],pp106[122],pp107[122],pp108[122],pp109[122],pp110[122],pp111[122],pp112[122],pp113[122],pp114[122],pp115[122]};
    CLA_220 KS_99(s99, c99, in99_1, in99_2);
    wire[217:0] s100, in100_1, in100_2;
    wire c100;
    assign in100_1 = {pp6[13],pp5[15],pp4[17],pp3[19],pp2[21],pp1[23],pp0[25],pp16[10],pp16[11],pp16[12],pp16[13],pp16[14],pp16[15],pp18[14],pp20[13],pp22[12],pp24[11],pp26[10],pp0[37],pp1[37],pp2[37],pp3[37],pp4[37],pp5[37],pp6[37],pp7[37],pp8[37],pp9[37],pp38[9],pp40[8],pp42[7],pp44[6],pp46[5],pp48[4],pp50[3],pp52[2],pp54[1],pp56[0],s65[25],s66[25],s67[25],s68[25],s69[25],s70[25],s71[25],s72[25],s73[25],s74[25],s75[25],s76[25],s77[25],s78[25],s79[25],s80[25],s81[25],s82[25],s83[25],s84[25],s85[25],s86[25],s87[25],s88[25],s89[25],s90[25],s90[26],s90[27],s90[28],s90[29],s90[30],s90[31],s90[32],s90[33],s90[34],s90[35],s90[36],s90[37],s90[38],s90[39],s90[40],s90[41],s90[42],s90[43],s90[44],s90[45],s90[46],s90[47],s90[48],s90[49],s90[50],s90[51],s90[52],s90[53],s90[54],s90[55],s90[56],s90[57],s90[58],s89[60],s88[62],s99[100],s99[101],s99[102],s99[103],s99[104],s99[105],s99[106],s99[107],s99[108],s99[109],s99[110],s99[111],s99[112],s99[113],s99[114],s99[115],s99[116],s99[117],s99[118],s99[119],s99[120],s99[121],s99[122],s99[123],s99[124],s99[125],s99[126],s99[127],s99[128],s99[129],s99[130],s99[131],s99[132],s99[133],s99[134],s99[135],s99[136],s99[137],s99[138],s99[139],s99[140],s99[141],s99[142],s99[143],s99[144],s99[145],s99[146],s99[147],s98[149],s97[151],s96[105],s95[107],s94[109],s93[111],s92[113],s90[116],s88[119],s86[122],s84[125],s82[128],s81[130],s81[131],s81[132],s81[133],s81[134],s81[135],s80[137],s79[139],s78[141],s77[143],s76[145],s75[147],s74[149],s73[151],s72[153],s71[155],s70[157],s69[159],s68[161],s67[163],s66[165],s65[167],pp127[73],pp126[75],pp125[77],pp124[79],pp123[81],pp122[83],pp121[85],pp120[87],pp119[89],pp118[91],pp117[93],pp116[95],pp115[97],pp114[99],pp98[116],pp96[119],pp94[122],pp92[125],pp118[100],pp116[103],pp114[106],pp112[109],pp110[112],pp108[115],pp106[118],pp106[119],pp106[120],pp106[121],pp107[121],pp108[121],pp109[121],pp110[121],pp111[121],pp112[121],pp113[121],pp114[121],pp115[121]};
    assign in100_2 = {pp7[12],pp6[14],pp5[16],pp4[18],pp3[20],pp2[22],pp1[24],pp0[26],pp17[10],pp17[11],pp17[12],pp17[13],pp17[14],pp19[13],pp21[12],pp23[11],pp25[10],pp0[36],pp1[36],pp2[36],pp3[36],pp4[36],pp5[36],pp6[36],pp7[36],pp8[36],pp9[36],pp37[9],pp39[8],pp41[7],pp43[6],pp45[5],pp47[4],pp49[3],pp51[2],pp53[1],pp55[0],s65[24],s66[24],s67[24],s68[24],s69[24],s70[24],s71[24],s72[24],s73[24],s74[24],s75[24],s76[24],s77[24],s78[24],s79[24],s80[24],s81[24],s82[24],s83[24],s84[24],s85[24],s86[24],s87[24],s88[24],s89[24],s90[24],s91[24],s91[25],s91[26],s91[27],s91[28],s91[29],s91[30],s91[31],s91[32],s91[33],s91[34],s91[35],s91[36],s91[37],s91[38],s91[39],s91[40],s91[41],s91[42],s91[43],s91[44],s91[45],s91[46],s91[47],s91[48],s91[49],s91[50],s91[51],s91[52],s91[53],s91[54],s91[55],s91[56],s91[57],s90[59],s89[61],s88[63],s88[64],s88[65],s88[66],s88[67],s88[68],s88[69],s88[70],s88[71],s88[72],s88[73],s86[76],s84[79],s82[82],s80[85],s79[87],s79[88],s79[89],s79[90],s79[91],s79[92],s79[93],s79[94],s79[95],s79[96],s79[97],s79[98],s79[99],s46[37],s44[40],s42[43],s40[46],s38[49],s36[52],s34[55],s32[58],s30[61],s28[64],s26[67],s24[70],s22[73],s20[76],s18[79],s16[82],s14[85],s12[88],s10[91],s1[101],s99[148],s98[150],s97[152],s96[106],s95[108],s94[110],s93[112],s91[115],s89[118],s87[121],s85[124],s83[127],s82[129],s82[130],s82[131],s82[132],s82[133],s82[134],s81[136],s80[138],s79[140],s78[142],s77[144],s76[146],s75[148],s74[150],s73[152],s72[154],s71[156],s70[158],s69[160],s68[162],s67[164],s66[166],s65[168],pp127[74],pp126[76],pp125[78],pp124[80],pp123[82],pp122[84],pp121[86],pp120[88],pp119[90],pp118[92],pp117[94],pp116[96],pp115[98],pp99[115],pp97[118],pp95[121],pp93[124],pp91[127],pp117[102],pp115[105],pp113[108],pp111[111],pp109[114],pp107[117],pp107[118],pp107[119],pp107[120],pp108[120],pp109[120],pp110[120],pp111[120],pp112[120],pp113[120],pp114[120],pp115[120],pp116[120]};
    CLA_218 KS_100(s100, c100, in100_1, in100_2);
    wire[215:0] s101, in101_1, in101_2;
    wire c101;
    assign in101_1 = {pp7[13],pp6[15],pp5[17],pp4[19],pp3[21],pp2[23],pp1[25],pp0[27],pp18[10],pp18[11],pp18[12],pp18[13],pp20[12],pp22[11],pp24[10],s100[16],s100[17],s100[18],s100[19],s100[20],s100[21],s100[22],s100[23],s100[24],s100[25],s100[26],s100[27],s100[28],s100[29],s100[30],s100[31],s100[32],s100[33],s100[34],s100[35],s100[36],s100[37],s100[38],s100[39],s100[40],s100[41],s100[42],s100[43],s100[44],s100[45],s100[46],s100[47],s100[48],s100[49],s100[50],s100[51],s100[52],s100[53],s100[54],s100[55],s100[56],s100[57],s100[58],s100[59],s100[60],s100[61],s100[62],s100[63],s100[64],s100[65],s100[66],s100[67],s100[68],s100[69],s100[70],s100[71],s100[72],s100[73],s100[74],s100[75],s100[76],s100[77],s100[78],s100[79],s100[80],s100[81],s100[82],s100[83],s100[84],s100[85],s100[86],s100[87],s100[88],s100[89],s100[90],s100[91],s100[92],s100[93],s100[94],s100[95],s100[96],s100[97],s100[98],s100[99],s100[100],s100[101],s100[102],s100[103],s100[104],s100[105],s100[106],s100[107],s100[108],s100[109],s100[110],s100[111],s100[112],s100[113],s100[114],s100[115],s100[116],s100[117],s100[118],s100[119],s100[120],s100[121],s100[122],s100[123],s100[124],s100[125],s100[126],s100[127],s100[128],s100[129],s100[130],s100[131],s100[132],s100[133],s100[134],s100[135],s100[136],s100[137],s100[138],s100[139],s100[140],s100[141],s100[142],s100[143],s100[144],s100[145],s100[146],s100[147],s100[148],s100[149],s100[150],s100[151],s100[152],s100[153],s100[154],s100[155],s100[156],s100[157],s100[158],s100[159],s100[160],s100[161],s100[162],s100[163],s100[164],s100[165],s100[166],s100[167],s100[168],s100[169],s100[170],s100[171],s100[172],s100[173],s100[174],s100[175],s100[176],s100[177],s100[178],s100[179],s100[180],s100[181],s100[182],pp127[75],pp126[77],pp125[79],pp124[81],pp123[83],pp122[85],pp121[87],pp120[89],pp119[91],pp118[93],pp117[95],pp116[97],pp115[99],pp98[117],pp96[120],pp94[123],pp92[126],pp118[101],pp116[104],pp114[107],pp112[110],pp110[113],pp108[116],pp108[117],pp108[118],pp108[119],pp109[119],pp110[119],pp111[119],pp112[119],pp113[119],pp114[119],pp115[119],pp116[119]};
    assign in101_2 = {pp8[12],pp7[14],pp6[16],pp5[18],pp4[20],pp3[22],pp2[24],pp1[26],pp0[28],pp19[10],pp19[11],pp19[12],pp21[11],pp23[10],s100[15],pp0[35],pp1[35],pp2[35],pp3[35],pp4[35],pp5[35],pp6[35],pp7[35],pp8[35],pp9[35],pp36[9],pp38[8],pp40[7],pp42[6],pp44[5],pp46[4],pp48[3],pp50[2],pp52[1],pp54[0],s65[23],s66[23],s67[23],s68[23],s69[23],s70[23],s71[23],s72[23],s73[23],s74[23],s75[23],s76[23],s77[23],s78[23],s79[23],s80[23],s81[23],s82[23],s83[23],s84[23],s85[23],s86[23],s87[23],s88[23],s89[23],s90[23],s91[23],s92[23],s92[24],s92[25],s92[26],s92[27],s92[28],s92[29],s92[30],s92[31],s92[32],s92[33],s92[34],s92[35],s92[36],s92[37],s92[38],s92[39],s92[40],s92[41],s92[42],s92[43],s92[44],s92[45],s92[46],s92[47],s92[48],s92[49],s92[50],s92[51],s92[52],s92[53],s92[54],s92[55],s92[56],s91[58],s90[60],s89[62],s89[63],s89[64],s89[65],s89[66],s89[67],s89[68],s89[69],s89[70],s89[71],s89[72],s87[75],s85[78],s83[81],s81[84],s80[86],s80[87],s80[88],s80[89],s80[90],s80[91],s80[92],s80[93],s80[94],s80[95],s80[96],s80[97],s80[98],s80[99],s45[39],s43[42],s41[45],s39[48],s37[51],s35[54],s33[57],s31[60],s29[63],s27[66],s25[69],s23[72],s21[75],s19[78],s17[81],s15[84],s13[87],s11[90],s2[100],s1[102],s99[149],s98[151],s97[153],s96[107],s95[109],s94[111],s92[114],s90[117],s88[120],s86[123],s84[126],s83[128],s83[129],s83[130],s83[131],s83[132],s83[133],s82[135],s81[137],s80[139],s79[141],s78[143],s77[145],s76[147],s75[149],s74[151],s73[153],s72[155],s71[157],s70[159],s69[161],s68[163],s67[165],s66[167],s65[169],s100[183],pp127[76],pp126[78],pp125[80],pp124[82],pp123[84],pp122[86],pp121[88],pp120[90],pp119[92],pp118[94],pp117[96],pp116[98],pp99[116],pp97[119],pp95[122],pp93[125],pp119[100],pp117[103],pp115[106],pp113[109],pp111[112],pp109[115],pp109[116],pp109[117],pp109[118],pp110[118],pp111[118],pp112[118],pp113[118],pp114[118],pp115[118],pp116[118],pp117[118]};
    CLA_216 KS_101(s101, c101, in101_1, in101_2);
    wire[213:0] s102, in102_1, in102_2;
    wire c102;
    assign in102_1 = {pp8[13],pp7[15],pp6[17],pp5[19],pp4[21],pp3[23],pp2[25],pp1[27],s100[10],pp20[10],pp20[11],pp22[10],s100[14],s101[14],s101[15],s101[16],s101[17],s101[18],s101[19],s101[20],s101[21],s101[22],s101[23],s101[24],s101[25],s101[26],s101[27],s101[28],s101[29],s101[30],s101[31],s101[32],s101[33],s101[34],s101[35],s101[36],s101[37],s101[38],s101[39],s101[40],s101[41],s101[42],s101[43],s101[44],s101[45],s101[46],s101[47],s101[48],s101[49],s101[50],s101[51],s101[52],s101[53],s101[54],s101[55],s101[56],s101[57],s101[58],s101[59],s101[60],s101[61],s101[62],s101[63],s101[64],s101[65],s101[66],s101[67],s101[68],s101[69],s101[70],s101[71],s101[72],s101[73],s101[74],s101[75],s101[76],s101[77],s101[78],s101[79],s101[80],s101[81],s101[82],s101[83],s101[84],s101[85],s101[86],s101[87],s101[88],s101[89],s101[90],s101[91],s101[92],s101[93],s101[94],s101[95],s101[96],s101[97],s101[98],s101[99],s101[100],s101[101],s101[102],s101[103],s101[104],s101[105],s101[106],s101[107],s101[108],s101[109],s101[110],s101[111],s101[112],s101[113],s101[114],s101[115],s101[116],s101[117],s101[118],s101[119],s101[120],s101[121],s101[122],s101[123],s101[124],s101[125],s101[126],s101[127],s101[128],s101[129],s101[130],s101[131],s101[132],s101[133],s101[134],s101[135],s101[136],s101[137],s101[138],s101[139],s101[140],s101[141],s101[142],s101[143],s101[144],s101[145],s101[146],s101[147],s101[148],s101[149],s101[150],s101[151],s101[152],s101[153],s101[154],s101[155],s101[156],s101[157],s101[158],s101[159],s101[160],s101[161],s101[162],s101[163],s101[164],s101[165],s101[166],s101[167],s101[168],s101[169],s101[170],s101[171],s101[172],s101[173],s101[174],s101[175],s101[176],s101[177],s101[178],s101[179],s101[180],s101[181],s101[182],s100[184],pp127[77],pp126[79],pp125[81],pp124[83],pp123[85],pp122[87],pp121[89],pp120[91],pp119[93],pp118[95],pp117[97],pp116[99],pp98[118],pp96[121],pp94[124],pp92[127],pp118[102],pp116[105],pp114[108],pp112[111],pp110[114],pp110[115],pp110[116],pp110[117],pp111[117],pp112[117],pp113[117],pp114[117],pp115[117],pp116[117],pp117[117]};
    assign in102_2 = {pp9[12],pp8[14],pp7[16],pp6[18],pp5[20],pp4[22],pp3[24],pp2[26],pp0[29],s100[11],pp21[10],s100[13],s101[13],pp0[34],pp1[34],pp2[34],pp3[34],pp4[34],pp5[34],pp6[34],pp7[34],pp8[34],pp9[34],pp35[9],pp37[8],pp39[7],pp41[6],pp43[5],pp45[4],pp47[3],pp49[2],pp51[1],pp53[0],s65[22],s66[22],s67[22],s68[22],s69[22],s70[22],s71[22],s72[22],s73[22],s74[22],s75[22],s76[22],s77[22],s78[22],s79[22],s80[22],s81[22],s82[22],s83[22],s84[22],s85[22],s86[22],s87[22],s88[22],s89[22],s90[22],s91[22],s92[22],s93[22],s93[23],s93[24],s93[25],s93[26],s93[27],s93[28],s93[29],s93[30],s93[31],s93[32],s93[33],s93[34],s93[35],s93[36],s93[37],s93[38],s93[39],s93[40],s93[41],s93[42],s93[43],s93[44],s93[45],s93[46],s93[47],s93[48],s93[49],s93[50],s93[51],s93[52],s93[53],s93[54],s93[55],s92[57],s91[59],s90[61],s90[62],s90[63],s90[64],s90[65],s90[66],s90[67],s90[68],s90[69],s90[70],s90[71],s88[74],s86[77],s84[80],s82[83],s81[85],s81[86],s81[87],s81[88],s81[89],s81[90],s81[91],s81[92],s81[93],s81[94],s81[95],s81[96],s81[97],s81[98],s81[99],s44[41],s42[44],s40[47],s38[50],s36[53],s34[56],s32[59],s30[62],s28[65],s26[68],s24[71],s22[74],s20[77],s18[80],s16[83],s14[86],s12[89],s10[92],s2[101],s1[103],s99[150],s98[152],s97[154],s96[108],s95[110],s93[113],s91[116],s89[119],s87[122],s85[125],s84[127],s84[128],s84[129],s84[130],s84[131],s84[132],s83[134],s82[136],s81[138],s80[140],s79[142],s78[144],s77[146],s76[148],s75[150],s74[152],s73[154],s72[156],s71[158],s70[160],s69[162],s68[164],s67[166],s66[168],s65[170],s101[183],s100[185],pp127[78],pp126[80],pp125[82],pp124[84],pp123[86],pp122[88],pp121[90],pp120[92],pp119[94],pp118[96],pp117[98],pp99[117],pp97[120],pp95[123],pp93[126],pp119[101],pp117[104],pp115[107],pp113[110],pp111[113],pp111[114],pp111[115],pp111[116],pp112[116],pp113[116],pp114[116],pp115[116],pp116[116],pp117[116],pp118[116]};
    CLA_214 KS_102(s102, c102, in102_1, in102_2);
    wire[211:0] s103, in103_1, in103_2;
    wire c103;
    assign in103_1 = {pp9[13],pp8[15],pp7[17],pp6[19],pp5[21],pp4[23],pp3[25],pp1[28],s101[10],s100[12],s101[12],s102[12],s102[13],s102[14],s102[15],s102[16],s102[17],s102[18],s102[19],s102[20],s102[21],s102[22],s102[23],s102[24],s102[25],s102[26],s102[27],s102[28],s102[29],s102[30],s102[31],s102[32],s102[33],s102[34],s102[35],s102[36],s102[37],s102[38],s102[39],s102[40],s102[41],s102[42],s102[43],s102[44],s102[45],s102[46],s102[47],s102[48],s102[49],s102[50],s102[51],s102[52],s102[53],s102[54],s102[55],s102[56],s102[57],s102[58],s102[59],s102[60],s102[61],s102[62],s102[63],s102[64],s102[65],s102[66],s102[67],s102[68],s102[69],s102[70],s102[71],s102[72],s102[73],s102[74],s102[75],s102[76],s102[77],s102[78],s102[79],s102[80],s102[81],s102[82],s102[83],s102[84],s102[85],s102[86],s102[87],s102[88],s102[89],s102[90],s102[91],s102[92],s102[93],s102[94],s102[95],s102[96],s102[97],s102[98],s102[99],s102[100],s102[101],s102[102],s102[103],s102[104],s102[105],s102[106],s102[107],s102[108],s102[109],s102[110],s102[111],s102[112],s102[113],s102[114],s102[115],s102[116],s102[117],s102[118],s102[119],s102[120],s102[121],s102[122],s102[123],s102[124],s102[125],s102[126],s102[127],s102[128],s102[129],s102[130],s102[131],s102[132],s102[133],s102[134],s102[135],s102[136],s102[137],s102[138],s102[139],s102[140],s102[141],s102[142],s102[143],s102[144],s102[145],s102[146],s102[147],s102[148],s102[149],s102[150],s102[151],s102[152],s102[153],s102[154],s102[155],s102[156],s102[157],s102[158],s102[159],s102[160],s102[161],s102[162],s102[163],s102[164],s102[165],s102[166],s102[167],s102[168],s102[169],s102[170],s102[171],s102[172],s102[173],s102[174],s102[175],s102[176],s102[177],s102[178],s102[179],s102[180],s102[181],s102[182],s101[184],s100[186],pp127[79],pp126[81],pp125[83],pp124[85],pp123[87],pp122[89],pp121[91],pp120[93],pp119[95],pp118[97],pp117[99],pp98[119],pp96[122],pp94[125],pp120[100],pp118[103],pp116[106],pp114[109],pp112[112],pp112[113],pp112[114],pp112[115],pp113[115],pp114[115],pp115[115],pp116[115],pp117[115],pp118[115]};
    assign in103_2 = {pp13[9],pp9[14],pp8[16],pp7[18],pp6[20],pp5[22],pp4[24],pp2[27],pp0[30],s101[11],s102[11],pp0[33],pp1[33],pp2[33],pp3[33],pp4[33],pp5[33],pp6[33],pp7[33],pp8[33],pp9[33],pp34[9],pp36[8],pp38[7],pp40[6],pp42[5],pp44[4],pp46[3],pp48[2],pp50[1],pp52[0],s65[21],s66[21],s67[21],s68[21],s69[21],s70[21],s71[21],s72[21],s73[21],s74[21],s75[21],s76[21],s77[21],s78[21],s79[21],s80[21],s81[21],s82[21],s83[21],s84[21],s85[21],s86[21],s87[21],s88[21],s89[21],s90[21],s91[21],s92[21],s93[21],s94[21],s94[22],s94[23],s94[24],s94[25],s94[26],s94[27],s94[28],s94[29],s94[30],s94[31],s94[32],s94[33],s94[34],s94[35],s94[36],s94[37],s94[38],s94[39],s94[40],s94[41],s94[42],s94[43],s94[44],s94[45],s94[46],s94[47],s94[48],s94[49],s94[50],s94[51],s94[52],s94[53],s94[54],s93[56],s92[58],s91[60],s91[61],s91[62],s91[63],s91[64],s91[65],s91[66],s91[67],s91[68],s91[69],s91[70],s89[73],s87[76],s85[79],s83[82],s82[84],s82[85],s82[86],s82[87],s82[88],s82[89],s82[90],s82[91],s82[92],s82[93],s82[94],s82[95],s82[96],s82[97],s82[98],s82[99],s43[43],s41[46],s39[49],s37[52],s35[55],s33[58],s31[61],s29[64],s27[67],s25[70],s23[73],s21[76],s19[79],s17[82],s15[85],s13[88],s11[91],s3[100],s2[102],s1[104],s99[151],s98[153],s97[155],s96[109],s94[112],s92[115],s90[118],s88[121],s86[124],s85[126],s85[127],s85[128],s85[129],s85[130],s85[131],s84[133],s83[135],s82[137],s81[139],s80[141],s79[143],s78[145],s77[147],s76[149],s75[151],s74[153],s73[155],s72[157],s71[159],s70[161],s69[163],s68[165],s67[167],s66[169],s65[171],s102[183],s101[185],s100[187],pp127[80],pp126[82],pp125[84],pp124[86],pp123[88],pp122[90],pp121[92],pp120[94],pp119[96],pp118[98],pp99[118],pp97[121],pp95[124],pp93[127],pp119[102],pp117[105],pp115[108],pp113[111],pp113[112],pp113[113],pp113[114],pp114[114],pp115[114],pp116[114],pp117[114],pp118[114],pp119[114]};
    CLA_212 KS_103(s103, c103, in103_1, in103_2);
    wire[209:0] s104, in104_1, in104_2;
    wire c104;
    assign in104_1 = {pp14[9],pp9[15],pp8[17],pp7[19],pp6[21],pp5[23],pp3[26],pp1[29],s102[10],s103[10],s103[11],s103[12],s103[13],s103[14],s103[15],s103[16],s103[17],s103[18],s103[19],s103[20],s103[21],s103[22],s103[23],s103[24],s103[25],s103[26],s103[27],s103[28],s103[29],s103[30],s103[31],s103[32],s103[33],s103[34],s103[35],s103[36],s103[37],s103[38],s103[39],s103[40],s103[41],s103[42],s103[43],s103[44],s103[45],s103[46],s103[47],s103[48],s103[49],s103[50],s103[51],s103[52],s103[53],s103[54],s103[55],s103[56],s103[57],s103[58],s103[59],s103[60],s103[61],s103[62],s103[63],s103[64],s103[65],s103[66],s103[67],s103[68],s103[69],s103[70],s103[71],s103[72],s103[73],s103[74],s103[75],s103[76],s103[77],s103[78],s103[79],s103[80],s103[81],s103[82],s103[83],s103[84],s103[85],s103[86],s103[87],s103[88],s103[89],s103[90],s103[91],s103[92],s103[93],s103[94],s103[95],s103[96],s103[97],s103[98],s103[99],s103[100],s103[101],s103[102],s103[103],s103[104],s103[105],s103[106],s103[107],s103[108],s103[109],s103[110],s103[111],s103[112],s103[113],s103[114],s103[115],s103[116],s103[117],s103[118],s103[119],s103[120],s103[121],s103[122],s103[123],s103[124],s103[125],s103[126],s103[127],s103[128],s103[129],s103[130],s103[131],s103[132],s103[133],s103[134],s103[135],s103[136],s103[137],s103[138],s103[139],s103[140],s103[141],s103[142],s103[143],s103[144],s103[145],s103[146],s103[147],s103[148],s103[149],s103[150],s103[151],s103[152],s103[153],s103[154],s103[155],s103[156],s103[157],s103[158],s103[159],s103[160],s103[161],s103[162],s103[163],s103[164],s103[165],s103[166],s103[167],s103[168],s103[169],s103[170],s103[171],s103[172],s103[173],s103[174],s103[175],s103[176],s103[177],s103[178],s103[179],s103[180],s103[181],s103[182],s102[184],s101[186],s100[188],pp127[81],pp126[83],pp125[85],pp124[87],pp123[89],pp122[91],pp121[93],pp120[95],pp119[97],pp118[99],pp98[120],pp96[123],pp94[126],pp120[101],pp118[104],pp116[107],pp114[110],pp114[111],pp114[112],pp114[113],pp115[113],pp116[113],pp117[113],pp118[113],pp119[113]};
    assign in104_2 = {pp15[8],pp15[9],pp9[16],pp8[18],pp7[20],pp6[22],pp4[25],pp2[28],pp0[31],pp0[32],pp1[32],pp2[32],pp3[32],pp4[32],pp5[32],pp6[32],pp7[32],pp8[32],pp9[32],pp33[9],pp35[8],pp37[7],pp39[6],pp41[5],pp43[4],pp45[3],pp47[2],pp49[1],pp51[0],s65[20],s66[20],s67[20],s68[20],s69[20],s70[20],s71[20],s72[20],s73[20],s74[20],s75[20],s76[20],s77[20],s78[20],s79[20],s80[20],s81[20],s82[20],s83[20],s84[20],s85[20],s86[20],s87[20],s88[20],s89[20],s90[20],s91[20],s92[20],s93[20],s94[20],s95[20],s95[21],s95[22],s95[23],s95[24],s95[25],s95[26],s95[27],s95[28],s95[29],s95[30],s95[31],s95[32],s95[33],s95[34],s95[35],s95[36],s95[37],s95[38],s95[39],s95[40],s95[41],s95[42],s95[43],s95[44],s95[45],s95[46],s95[47],s95[48],s95[49],s95[50],s95[51],s95[52],s95[53],s94[55],s93[57],s92[59],s92[60],s92[61],s92[62],s92[63],s92[64],s92[65],s92[66],s92[67],s92[68],s92[69],s90[72],s88[75],s86[78],s84[81],s83[83],s83[84],s83[85],s83[86],s83[87],s83[88],s83[89],s83[90],s83[91],s83[92],s83[93],s83[94],s83[95],s83[96],s83[97],s83[98],s83[99],s42[45],s40[48],s38[51],s36[54],s34[57],s32[60],s30[63],s28[66],s26[69],s24[72],s22[75],s20[78],s18[81],s16[84],s14[87],s12[90],s10[93],s3[101],s2[103],s1[105],s99[152],s98[154],s97[156],s95[111],s93[114],s91[117],s89[120],s87[123],s86[125],s86[126],s86[127],s86[128],s86[129],s86[130],s85[132],s84[134],s83[136],s82[138],s81[140],s80[142],s79[144],s78[146],s77[148],s76[150],s75[152],s74[154],s73[156],s72[158],s71[160],s70[162],s69[164],s68[166],s67[168],s66[170],s65[172],s103[183],s102[185],s101[187],s100[189],pp127[82],pp126[84],pp125[86],pp124[88],pp123[90],pp122[92],pp121[94],pp120[96],pp119[98],pp99[119],pp97[122],pp95[125],pp121[100],pp119[103],pp117[106],pp115[109],pp115[110],pp115[111],pp115[112],pp116[112],pp117[112],pp118[112],pp119[112],pp120[112]};
    CLA_210 KS_104(s104, c104, in104_1, in104_2);
    wire[207:0] s105, in105_1, in105_2;
    wire c105;
    assign in105_1 = {pp16[8],pp16[9],pp9[17],pp8[19],pp7[21],pp5[24],pp3[27],pp1[30],pp1[31],s104[10],s104[11],s104[12],s104[13],s104[14],s104[15],s104[16],s104[17],s104[18],s104[19],s104[20],s104[21],s104[22],s104[23],s104[24],s104[25],s104[26],s104[27],s104[28],s104[29],s104[30],s104[31],s104[32],s104[33],s104[34],s104[35],s104[36],s104[37],s104[38],s104[39],s104[40],s104[41],s104[42],s104[43],s104[44],s104[45],s104[46],s104[47],s104[48],s104[49],s104[50],s104[51],s104[52],s104[53],s104[54],s104[55],s104[56],s104[57],s104[58],s104[59],s104[60],s104[61],s104[62],s104[63],s104[64],s104[65],s104[66],s104[67],s104[68],s104[69],s104[70],s104[71],s104[72],s104[73],s104[74],s104[75],s104[76],s104[77],s104[78],s104[79],s104[80],s104[81],s104[82],s104[83],s104[84],s104[85],s104[86],s104[87],s104[88],s104[89],s104[90],s104[91],s104[92],s104[93],s104[94],s104[95],s104[96],s104[97],s104[98],s104[99],s104[100],s104[101],s104[102],s104[103],s104[104],s104[105],s104[106],s104[107],s104[108],s104[109],s104[110],s104[111],s104[112],s104[113],s104[114],s104[115],s104[116],s104[117],s104[118],s104[119],s104[120],s104[121],s104[122],s104[123],s104[124],s104[125],s104[126],s104[127],s104[128],s104[129],s104[130],s104[131],s104[132],s104[133],s104[134],s104[135],s104[136],s104[137],s104[138],s104[139],s104[140],s104[141],s104[142],s104[143],s104[144],s104[145],s104[146],s104[147],s104[148],s104[149],s104[150],s104[151],s104[152],s104[153],s104[154],s104[155],s104[156],s104[157],s104[158],s104[159],s104[160],s104[161],s104[162],s104[163],s104[164],s104[165],s104[166],s104[167],s104[168],s104[169],s104[170],s104[171],s104[172],s104[173],s104[174],s104[175],s104[176],s104[177],s104[178],s104[179],s104[180],s104[181],s104[182],s103[184],s102[186],s101[188],s100[190],pp127[83],pp126[85],pp125[87],pp124[89],pp123[91],pp122[93],pp121[95],pp120[97],pp119[99],pp98[121],pp96[124],pp94[127],pp120[102],pp118[105],pp116[108],pp116[109],pp116[110],pp116[111],pp117[111],pp118[111],pp119[111],pp120[111]};
    assign in105_2 = {pp17[7],pp17[8],pp17[9],pp9[18],pp8[20],pp6[23],pp4[26],pp2[29],pp2[30],pp2[31],pp3[31],pp4[31],pp5[31],pp6[31],pp7[31],pp8[31],pp9[31],pp32[9],pp34[8],pp36[7],pp38[6],pp40[5],pp42[4],pp44[3],pp46[2],pp48[1],pp50[0],s65[19],s66[19],s67[19],s68[19],s69[19],s70[19],s71[19],s72[19],s73[19],s74[19],s75[19],s76[19],s77[19],s78[19],s79[19],s80[19],s81[19],s82[19],s83[19],s84[19],s85[19],s86[19],s87[19],s88[19],s89[19],s90[19],s91[19],s92[19],s93[19],s94[19],s95[19],s96[19],s96[20],s96[21],s96[22],s96[23],s96[24],s96[25],s96[26],s96[27],s96[28],s96[29],s96[30],s96[31],s96[32],s96[33],s96[34],s96[35],s96[36],s96[37],s96[38],s96[39],s96[40],s96[41],s96[42],s96[43],s96[44],s96[45],s96[46],s96[47],s96[48],s96[49],s96[50],s96[51],s96[52],s95[54],s94[56],s93[58],s93[59],s93[60],s93[61],s93[62],s93[63],s93[64],s93[65],s93[66],s93[67],s93[68],s91[71],s89[74],s87[77],s85[80],s84[82],s84[83],s84[84],s84[85],s84[86],s84[87],s84[88],s84[89],s84[90],s84[91],s84[92],s84[93],s84[94],s84[95],s84[96],s84[97],s84[98],s84[99],s41[47],s39[50],s37[53],s35[56],s33[59],s31[62],s29[65],s27[68],s25[71],s23[74],s21[77],s19[80],s17[83],s15[86],s13[89],s11[92],s4[100],s3[102],s2[104],s1[106],s99[153],s98[155],s96[110],s94[113],s92[116],s90[119],s88[122],s87[124],s87[125],s87[126],s87[127],s87[128],s87[129],s86[131],s85[133],s84[135],s83[137],s82[139],s81[141],s80[143],s79[145],s78[147],s77[149],s76[151],s75[153],s74[155],s73[157],s72[159],s71[161],s70[163],s69[165],s68[167],s67[169],s66[171],s65[173],s104[183],s103[185],s102[187],s101[189],s100[191],pp127[84],pp126[86],pp125[88],pp124[90],pp123[92],pp122[94],pp121[96],pp120[98],pp99[120],pp97[123],pp95[126],pp121[101],pp119[104],pp117[107],pp117[108],pp117[109],pp117[110],pp118[110],pp119[110],pp120[110],pp121[110]};
    CLA_208 KS_105(s105, c105, in105_1, in105_2);
    wire[205:0] s106, in106_1, in106_2;
    wire c106;
    assign in106_1 = {pp18[7],pp18[8],pp18[9],pp9[19],pp7[22],pp5[25],pp3[28],pp3[29],pp3[30],s105[10],s105[11],s105[12],s105[13],s105[14],s105[15],s105[16],s105[17],s105[18],s105[19],s105[20],s105[21],s105[22],s105[23],s105[24],s105[25],s105[26],s105[27],s105[28],s105[29],s105[30],s105[31],s105[32],s105[33],s105[34],s105[35],s105[36],s105[37],s105[38],s105[39],s105[40],s105[41],s105[42],s105[43],s105[44],s105[45],s105[46],s105[47],s105[48],s105[49],s105[50],s105[51],s105[52],s105[53],s105[54],s105[55],s105[56],s105[57],s105[58],s105[59],s105[60],s105[61],s105[62],s105[63],s105[64],s105[65],s105[66],s105[67],s105[68],s105[69],s105[70],s105[71],s105[72],s105[73],s105[74],s105[75],s105[76],s105[77],s105[78],s105[79],s105[80],s105[81],s105[82],s105[83],s105[84],s105[85],s105[86],s105[87],s105[88],s105[89],s105[90],s105[91],s105[92],s105[93],s105[94],s105[95],s105[96],s105[97],s105[98],s105[99],s105[100],s105[101],s105[102],s105[103],s105[104],s105[105],s105[106],s105[107],s105[108],s105[109],s105[110],s105[111],s105[112],s105[113],s105[114],s105[115],s105[116],s105[117],s105[118],s105[119],s105[120],s105[121],s105[122],s105[123],s105[124],s105[125],s105[126],s105[127],s105[128],s105[129],s105[130],s105[131],s105[132],s105[133],s105[134],s105[135],s105[136],s105[137],s105[138],s105[139],s105[140],s105[141],s105[142],s105[143],s105[144],s105[145],s105[146],s105[147],s105[148],s105[149],s105[150],s105[151],s105[152],s105[153],s105[154],s105[155],s105[156],s105[157],s105[158],s105[159],s105[160],s105[161],s105[162],s105[163],s105[164],s105[165],s105[166],s105[167],s105[168],s105[169],s105[170],s105[171],s105[172],s105[173],s105[174],s105[175],s105[176],s105[177],s105[178],s105[179],s105[180],s105[181],s105[182],s104[184],s103[186],s102[188],s101[190],s100[192],pp127[85],pp126[87],pp125[89],pp124[91],pp123[93],pp122[95],pp121[97],pp120[99],pp98[122],pp96[125],pp122[100],pp120[103],pp118[106],pp118[107],pp118[108],pp118[109],pp119[109],pp120[109],pp121[109]};
    assign in106_2 = {pp19[6],pp19[7],pp19[8],pp19[9],pp8[21],pp6[24],pp4[27],pp4[28],pp4[29],pp4[30],pp5[30],pp6[30],pp7[30],pp8[30],pp9[30],pp31[9],pp33[8],pp35[7],pp37[6],pp39[5],pp41[4],pp43[3],pp45[2],pp47[1],pp49[0],s65[18],s66[18],s67[18],s68[18],s69[18],s70[18],s71[18],s72[18],s73[18],s74[18],s75[18],s76[18],s77[18],s78[18],s79[18],s80[18],s81[18],s82[18],s83[18],s84[18],s85[18],s86[18],s87[18],s88[18],s89[18],s90[18],s91[18],s92[18],s93[18],s94[18],s95[18],s96[18],s97[66],s97[67],s97[68],s97[69],s97[70],s97[71],s97[72],s97[73],s97[74],s97[75],s97[76],s97[77],s97[78],s97[79],s97[80],s97[81],s97[82],s97[83],s97[84],s97[85],s97[86],s97[87],s97[88],s97[89],s97[90],s97[91],s97[92],s97[93],s97[94],s97[95],s97[96],s97[97],s97[98],s97[99],s96[53],s95[55],s94[57],s94[58],s94[59],s94[60],s94[61],s94[62],s94[63],s94[64],s94[65],s94[66],s94[67],s92[70],s90[73],s88[76],s86[79],s85[81],s85[82],s85[83],s85[84],s85[85],s85[86],s85[87],s85[88],s85[89],s85[90],s85[91],s85[92],s85[93],s85[94],s85[95],s85[96],s85[97],s85[98],s85[99],s40[49],s38[52],s36[55],s34[58],s32[61],s30[64],s28[67],s26[70],s24[73],s22[76],s20[79],s18[82],s16[85],s14[88],s12[91],s10[94],s4[101],s3[103],s2[105],s1[107],s99[154],s97[157],s95[112],s93[115],s91[118],s89[121],s88[123],s88[124],s88[125],s88[126],s88[127],s88[128],s87[130],s86[132],s85[134],s84[136],s83[138],s82[140],s81[142],s80[144],s79[146],s78[148],s77[150],s76[152],s75[154],s74[156],s73[158],s72[160],s71[162],s70[164],s69[166],s68[168],s67[170],s66[172],s65[174],s105[183],s104[185],s103[187],s102[189],s101[191],s100[193],pp127[86],pp126[88],pp125[90],pp124[92],pp123[94],pp122[96],pp121[98],pp99[121],pp97[124],pp95[127],pp121[102],pp119[105],pp119[106],pp119[107],pp119[108],pp120[108],pp121[108],pp122[108]};
    CLA_206 KS_106(s106, c106, in106_1, in106_2);
    wire[203:0] s107, in107_1, in107_2;
    wire c107;
    assign in107_1 = {pp20[6],pp20[7],pp20[8],pp9[20],pp7[23],pp5[26],pp5[27],pp5[28],pp5[29],s106[10],s106[11],s106[12],s106[13],s106[14],s106[15],s106[16],s106[17],s106[18],s106[19],s106[20],s106[21],s106[22],s106[23],s106[24],s106[25],s106[26],s106[27],s106[28],s106[29],s106[30],s106[31],s106[32],s106[33],s106[34],s106[35],s106[36],s106[37],s106[38],s106[39],s106[40],s106[41],s106[42],s106[43],s106[44],s106[45],s106[46],s106[47],s106[48],s106[49],s106[50],s106[51],s106[52],s106[53],s106[54],s106[55],s106[56],s106[57],s106[58],s106[59],s106[60],s106[61],s106[62],s106[63],s106[64],s106[65],s106[66],s106[67],s106[68],s106[69],s106[70],s106[71],s106[72],s106[73],s106[74],s106[75],s106[76],s106[77],s106[78],s106[79],s106[80],s106[81],s106[82],s106[83],s106[84],s106[85],s106[86],s106[87],s106[88],s106[89],s106[90],s106[91],s106[92],s106[93],s106[94],s106[95],s106[96],s106[97],s106[98],s106[99],s106[100],s106[101],s106[102],s106[103],s106[104],s106[105],s106[106],s106[107],s106[108],s106[109],s106[110],s106[111],s106[112],s106[113],s106[114],s106[115],s106[116],s106[117],s106[118],s106[119],s106[120],s106[121],s106[122],s106[123],s106[124],s106[125],s106[126],s106[127],s106[128],s106[129],s106[130],s106[131],s106[132],s106[133],s106[134],s106[135],s106[136],s106[137],s106[138],s106[139],s106[140],s106[141],s106[142],s106[143],s106[144],s106[145],s106[146],s106[147],s106[148],s106[149],s106[150],s106[151],s106[152],s106[153],s106[154],s106[155],s106[156],s106[157],s106[158],s106[159],s106[160],s106[161],s106[162],s106[163],s106[164],s106[165],s106[166],s106[167],s106[168],s106[169],s106[170],s106[171],s106[172],s106[173],s106[174],s106[175],s106[176],s106[177],s106[178],s106[179],s106[180],s106[181],s106[182],s105[184],s104[186],s103[188],s102[190],s101[192],s100[194],pp127[87],pp126[89],pp125[91],pp124[93],pp123[95],pp122[97],pp121[99],pp98[123],pp96[126],pp122[101],pp120[104],pp120[105],pp120[106],pp120[107],pp121[107],pp122[107]};
    assign in107_2 = {pp21[5],pp21[6],pp21[7],pp20[9],pp8[22],pp6[25],pp6[26],pp6[27],pp6[28],pp6[29],pp7[29],pp8[29],pp9[29],pp30[9],pp32[8],pp34[7],pp36[6],pp38[5],pp40[4],pp42[3],pp44[2],pp46[1],pp48[0],s65[17],s66[17],s67[17],s68[17],s69[17],s70[17],s71[17],s72[17],s73[17],s74[17],s75[17],s76[17],s77[17],s78[17],s79[17],s80[17],s81[17],s82[17],s83[17],s84[17],s85[17],s86[17],s87[17],s88[17],s89[17],s90[17],s91[17],s92[17],s93[17],s94[17],s95[17],s96[17],s97[65],s98[65],s98[66],s98[67],s98[68],s98[69],s98[70],s98[71],s98[72],s98[73],s98[74],s98[75],s98[76],s98[77],s98[78],s98[79],s98[80],s98[81],s98[82],s98[83],s98[84],s98[85],s98[86],s98[87],s98[88],s98[89],s98[90],s98[91],s98[92],s98[93],s98[94],s98[95],s98[96],s98[97],s98[98],s98[99],s96[54],s95[56],s95[57],s95[58],s95[59],s95[60],s95[61],s95[62],s95[63],s95[64],s95[65],s95[66],s93[69],s91[72],s89[75],s87[78],s86[80],s86[81],s86[82],s86[83],s86[84],s86[85],s86[86],s86[87],s86[88],s86[89],s86[90],s86[91],s86[92],s86[93],s86[94],s86[95],s86[96],s86[97],s86[98],s86[99],s39[51],s37[54],s35[57],s33[60],s31[63],s29[66],s27[69],s25[72],s23[75],s21[78],s19[81],s17[84],s15[87],s13[90],s11[93],s5[100],s4[102],s3[104],s2[106],s1[108],s98[156],s96[111],s94[114],s92[117],s90[120],s89[122],s89[123],s89[124],s89[125],s89[126],s89[127],s88[129],s87[131],s86[133],s85[135],s84[137],s83[139],s82[141],s81[143],s80[145],s79[147],s78[149],s77[151],s76[153],s75[155],s74[157],s73[159],s72[161],s71[163],s70[165],s69[167],s68[169],s67[171],s66[173],s65[175],s106[183],s105[185],s104[187],s103[189],s102[191],s101[193],s100[195],pp127[88],pp126[90],pp125[92],pp124[94],pp123[96],pp122[98],pp99[122],pp97[125],pp123[100],pp121[103],pp121[104],pp121[105],pp121[106],pp122[106],pp123[106]};
    CLA_204 KS_107(s107, c107, in107_1, in107_2);
    wire[201:0] s108, in108_1, in108_2;
    wire c108;
    assign in108_1 = {pp22[5],pp22[6],pp21[8],pp9[21],pp7[24],pp7[25],pp7[26],pp7[27],pp7[28],s107[10],s107[11],s107[12],s107[13],s107[14],s107[15],s107[16],s107[17],s107[18],s107[19],s107[20],s107[21],s107[22],s107[23],s107[24],s107[25],s107[26],s107[27],s107[28],s107[29],s107[30],s107[31],s107[32],s107[33],s107[34],s107[35],s107[36],s107[37],s107[38],s107[39],s107[40],s107[41],s107[42],s107[43],s107[44],s107[45],s107[46],s107[47],s107[48],s107[49],s107[50],s107[51],s107[52],s107[53],s107[54],s107[55],s107[56],s107[57],s107[58],s107[59],s107[60],s107[61],s107[62],s107[63],s107[64],s107[65],s107[66],s107[67],s107[68],s107[69],s107[70],s107[71],s107[72],s107[73],s107[74],s107[75],s107[76],s107[77],s107[78],s107[79],s107[80],s107[81],s107[82],s107[83],s107[84],s107[85],s107[86],s107[87],s107[88],s107[89],s107[90],s107[91],s107[92],s107[93],s107[94],s107[95],s107[96],s107[97],s107[98],s107[99],s107[100],s107[101],s107[102],s107[103],s107[104],s107[105],s107[106],s107[107],s107[108],s107[109],s107[110],s107[111],s107[112],s107[113],s107[114],s107[115],s107[116],s107[117],s107[118],s107[119],s107[120],s107[121],s107[122],s107[123],s107[124],s107[125],s107[126],s107[127],s107[128],s107[129],s107[130],s107[131],s107[132],s107[133],s107[134],s107[135],s107[136],s107[137],s107[138],s107[139],s107[140],s107[141],s107[142],s107[143],s107[144],s107[145],s107[146],s107[147],s107[148],s107[149],s107[150],s107[151],s107[152],s107[153],s107[154],s107[155],s107[156],s107[157],s107[158],s107[159],s107[160],s107[161],s107[162],s107[163],s107[164],s107[165],s107[166],s107[167],s107[168],s107[169],s107[170],s107[171],s107[172],s107[173],s107[174],s107[175],s107[176],s107[177],s107[178],s107[179],s107[180],s107[181],s107[182],s106[184],s105[186],s104[188],s103[190],s102[192],s101[194],s100[196],pp127[89],pp126[91],pp125[93],pp124[95],pp123[97],pp122[99],pp98[124],pp96[127],pp122[102],pp122[103],pp122[104],pp122[105],pp123[105]};
    assign in108_2 = {pp23[4],pp23[5],pp22[7],pp21[9],pp8[23],pp8[24],pp8[25],pp8[26],pp8[27],pp8[28],pp9[28],pp29[9],pp31[8],pp33[7],pp35[6],pp37[5],pp39[4],pp41[3],pp43[2],pp45[1],pp47[0],s65[16],s66[16],s67[16],s68[16],s69[16],s70[16],s71[16],s72[16],s73[16],s74[16],s75[16],s76[16],s77[16],s78[16],s79[16],s80[16],s81[16],s82[16],s83[16],s84[16],s85[16],s86[16],s87[16],s88[16],s89[16],s90[16],s91[16],s92[16],s93[16],s94[16],s95[16],s96[16],s97[64],s98[64],s99[64],s99[65],s99[66],s99[67],s99[68],s99[69],s99[70],s99[71],s99[72],s99[73],s99[74],s99[75],s99[76],s99[77],s99[78],s99[79],s99[80],s99[81],s99[82],s99[83],s99[84],s99[85],s99[86],s99[87],s99[88],s99[89],s99[90],s99[91],s99[92],s99[93],s99[94],s99[95],s99[96],s99[97],s99[98],s99[99],s96[55],s96[56],s96[57],s96[58],s96[59],s96[60],s96[61],s96[62],s96[63],s96[64],s96[65],s94[68],s92[71],s90[74],s88[77],s87[79],s87[80],s87[81],s87[82],s87[83],s87[84],s87[85],s87[86],s87[87],s87[88],s87[89],s87[90],s87[91],s87[92],s87[93],s87[94],s87[95],s87[96],s87[97],s87[98],s87[99],s38[53],s36[56],s34[59],s32[62],s30[65],s28[68],s26[71],s24[74],s22[77],s20[80],s18[83],s16[86],s14[89],s12[92],s10[95],s5[101],s4[103],s3[105],s2[107],s99[155],s97[158],s95[113],s93[116],s91[119],s90[121],s90[122],s90[123],s90[124],s90[125],s90[126],s89[128],s88[130],s87[132],s86[134],s85[136],s84[138],s83[140],s82[142],s81[144],s80[146],s79[148],s78[150],s77[152],s76[154],s75[156],s74[158],s73[160],s72[162],s71[164],s70[166],s69[168],s68[170],s67[172],s66[174],s65[176],s107[183],s106[185],s105[187],s104[189],s103[191],s102[193],s101[195],s100[197],pp127[90],pp126[92],pp125[94],pp124[96],pp123[98],pp99[123],pp97[126],pp123[101],pp123[102],pp123[103],pp123[104],pp124[104]};
    CLA_202 KS_108(s108, c108, in108_1, in108_2);
    wire[199:0] s109, in109_1, in109_2;
    wire c109;
    assign in109_1 = {pp24[4],pp23[6],pp22[8],pp9[22],pp9[23],pp9[24],pp9[25],pp9[26],pp9[27],s108[10],s108[11],s108[12],s108[13],s108[14],s108[15],s108[16],s108[17],s108[18],s108[19],s108[20],s108[21],s108[22],s108[23],s108[24],s108[25],s108[26],s108[27],s108[28],s108[29],s108[30],s108[31],s108[32],s108[33],s108[34],s108[35],s108[36],s108[37],s108[38],s108[39],s108[40],s108[41],s108[42],s108[43],s108[44],s108[45],s108[46],s108[47],s108[48],s108[49],s108[50],s108[51],s108[52],s108[53],s108[54],s108[55],s108[56],s108[57],s108[58],s108[59],s108[60],s108[61],s108[62],s108[63],s108[64],s108[65],s108[66],s108[67],s108[68],s108[69],s108[70],s108[71],s108[72],s108[73],s108[74],s108[75],s108[76],s108[77],s108[78],s108[79],s108[80],s108[81],s108[82],s108[83],s108[84],s108[85],s108[86],s108[87],s108[88],s108[89],s108[90],s108[91],s108[92],s108[93],s108[94],s108[95],s108[96],s108[97],s108[98],s108[99],s108[100],s108[101],s108[102],s108[103],s108[104],s108[105],s108[106],s108[107],s108[108],s108[109],s108[110],s108[111],s108[112],s108[113],s108[114],s108[115],s108[116],s108[117],s108[118],s108[119],s108[120],s108[121],s108[122],s108[123],s108[124],s108[125],s108[126],s108[127],s108[128],s108[129],s108[130],s108[131],s108[132],s108[133],s108[134],s108[135],s108[136],s108[137],s108[138],s108[139],s108[140],s108[141],s108[142],s108[143],s108[144],s108[145],s108[146],s108[147],s108[148],s108[149],s108[150],s108[151],s108[152],s108[153],s108[154],s108[155],s108[156],s108[157],s108[158],s108[159],s108[160],s108[161],s108[162],s108[163],s108[164],s108[165],s108[166],s108[167],s108[168],s108[169],s108[170],s108[171],s108[172],s108[173],s108[174],s108[175],s108[176],s108[177],s108[178],s108[179],s108[180],s108[181],s108[182],s107[184],s106[186],s105[188],s104[190],s103[192],s102[194],s101[196],s100[198],pp127[91],pp126[93],pp125[95],pp124[97],pp123[99],pp98[125],pp124[100],pp124[101],pp124[102],pp124[103]};
    assign in109_2 = {pp25[3],pp24[5],pp23[7],pp22[9],pp23[9],pp24[9],pp25[9],pp26[9],pp27[9],pp28[9],pp30[8],pp32[7],pp34[6],pp36[5],pp38[4],pp40[3],pp42[2],pp44[1],pp46[0],s65[15],s66[15],s67[15],s68[15],s69[15],s70[15],s71[15],s72[15],s73[15],s74[15],s75[15],s76[15],s77[15],s78[15],s79[15],s80[15],s81[15],s82[15],s83[15],s84[15],s85[15],s86[15],s87[15],s88[15],s89[15],s90[15],s91[15],s92[15],s93[15],s94[15],s95[15],s96[15],s97[63],s98[63],s99[63],s1[18],s1[19],s1[20],s1[21],s1[22],s1[23],s1[24],s1[25],s1[26],s1[27],s1[28],s1[29],s1[30],s1[31],s1[32],s1[33],s1[34],s1[35],s1[36],s1[37],s1[38],s1[39],s1[40],s1[41],s1[42],s1[43],s1[44],s1[45],s1[46],s1[47],s1[48],s1[49],s1[50],s1[51],s1[52],s1[53],s1[54],s1[55],s1[56],s1[57],s1[58],s1[59],s1[60],s1[61],s1[62],s1[63],s1[64],s95[67],s93[70],s91[73],s89[76],s88[78],s88[79],s88[80],s88[81],s88[82],s88[83],s88[84],s88[85],s88[86],s88[87],s88[88],s88[89],s88[90],s88[91],s88[92],s88[93],s88[94],s88[95],s88[96],s88[97],s88[98],s88[99],s37[55],s35[58],s33[61],s31[64],s29[67],s27[70],s25[73],s23[76],s21[79],s19[82],s17[85],s15[88],s13[91],s11[94],s6[100],s5[102],s4[104],s3[106],s1[109],s98[157],s96[112],s94[115],s92[118],s91[120],s91[121],s91[122],s91[123],s91[124],s91[125],s90[127],s89[129],s88[131],s87[133],s86[135],s85[137],s84[139],s83[141],s82[143],s81[145],s80[147],s79[149],s78[151],s77[153],s76[155],s75[157],s74[159],s73[161],s72[163],s71[165],s70[167],s69[169],s68[171],s67[173],s66[175],s65[177],s108[183],s107[185],s106[187],s105[189],s104[191],s103[193],s102[195],s101[197],s100[199],pp127[92],pp126[94],pp125[96],pp124[98],pp99[124],pp97[127],pp125[100],pp125[101],pp125[102]};
    CLA_200 KS_109(s109, c109, in109_1, in109_2);
    wire[197:0] s110, in110_1, in110_2;
    wire c110;
    assign in110_1 = {pp25[4],pp24[6],pp23[8],pp24[8],pp25[8],pp26[8],pp27[8],pp28[8],pp29[8],s109[10],s109[11],s109[12],s109[13],s109[14],s109[15],s109[16],s109[17],s109[18],s109[19],s109[20],s109[21],s109[22],s109[23],s109[24],s109[25],s109[26],s109[27],s109[28],s109[29],s109[30],s109[31],s109[32],s109[33],s109[34],s109[35],s109[36],s109[37],s109[38],s109[39],s109[40],s109[41],s109[42],s109[43],s109[44],s109[45],s109[46],s109[47],s109[48],s109[49],s109[50],s109[51],s109[52],s109[53],s109[54],s109[55],s109[56],s109[57],s109[58],s109[59],s109[60],s109[61],s109[62],s109[63],s109[64],s109[65],s109[66],s109[67],s109[68],s109[69],s109[70],s109[71],s109[72],s109[73],s109[74],s109[75],s109[76],s109[77],s109[78],s109[79],s109[80],s109[81],s109[82],s109[83],s109[84],s109[85],s109[86],s109[87],s109[88],s109[89],s109[90],s109[91],s109[92],s109[93],s109[94],s109[95],s109[96],s109[97],s109[98],s109[99],s109[100],s109[101],s109[102],s109[103],s109[104],s109[105],s109[106],s109[107],s109[108],s109[109],s109[110],s109[111],s109[112],s109[113],s109[114],s109[115],s109[116],s109[117],s109[118],s109[119],s109[120],s109[121],s109[122],s109[123],s109[124],s109[125],s109[126],s109[127],s109[128],s109[129],s109[130],s109[131],s109[132],s109[133],s109[134],s109[135],s109[136],s109[137],s109[138],s109[139],s109[140],s109[141],s109[142],s109[143],s109[144],s109[145],s109[146],s109[147],s109[148],s109[149],s109[150],s109[151],s109[152],s109[153],s109[154],s109[155],s109[156],s109[157],s109[158],s109[159],s109[160],s109[161],s109[162],s109[163],s109[164],s109[165],s109[166],s109[167],s109[168],s109[169],s109[170],s109[171],s109[172],s109[173],s109[174],s109[175],s109[176],s109[177],s109[178],s109[179],s109[180],s109[181],s109[182],s108[184],s107[186],s106[188],s105[190],s104[192],s103[194],s102[196],s101[198],s100[200],pp127[93],pp126[95],pp125[97],pp124[99],pp98[126],pp98[127],pp126[100]};
    assign in110_2 = {pp26[3],pp25[5],pp24[7],pp25[7],pp26[7],pp27[7],pp28[7],pp29[7],pp30[7],pp31[7],pp33[6],pp35[5],pp37[4],pp39[3],pp41[2],pp43[1],pp45[0],s65[14],s66[14],s67[14],s68[14],s69[14],s70[14],s71[14],s72[14],s73[14],s74[14],s75[14],s76[14],s77[14],s78[14],s79[14],s80[14],s81[14],s82[14],s83[14],s84[14],s85[14],s86[14],s87[14],s88[14],s89[14],s90[14],s91[14],s92[14],s93[14],s94[14],s95[14],s96[14],s97[62],s98[62],s99[62],s1[17],s2[17],s2[18],s2[19],s2[20],s2[21],s2[22],s2[23],s2[24],s2[25],s2[26],s2[27],s2[28],s2[29],s2[30],s2[31],s2[32],s2[33],s2[34],s2[35],s2[36],s2[37],s2[38],s2[39],s2[40],s2[41],s2[42],s2[43],s2[44],s2[45],s2[46],s2[47],s2[48],s2[49],s2[50],s2[51],s2[52],s2[53],s2[54],s2[55],s2[56],s2[57],s2[58],s2[59],s2[60],s2[61],s2[62],s2[63],s96[66],s94[69],s92[72],s90[75],s89[77],s89[78],s89[79],s89[80],s89[81],s89[82],s89[83],s89[84],s89[85],s89[86],s89[87],s89[88],s89[89],s89[90],s89[91],s89[92],s89[93],s89[94],s89[95],s89[96],s89[97],s89[98],s89[99],s36[57],s34[60],s32[63],s30[66],s28[69],s26[72],s24[75],s22[78],s20[81],s18[84],s16[87],s14[90],s12[93],s10[96],s6[101],s5[103],s4[105],s2[108],s99[156],s97[159],s95[114],s93[117],s92[119],s92[120],s92[121],s92[122],s92[123],s92[124],s91[126],s90[128],s89[130],s88[132],s87[134],s86[136],s85[138],s84[140],s83[142],s82[144],s81[146],s80[148],s79[150],s78[152],s77[154],s76[156],s75[158],s74[160],s73[162],s72[164],s71[166],s70[168],s69[170],s68[172],s67[174],s66[176],s65[178],s109[183],s108[185],s107[187],s106[189],s105[191],s104[193],s103[195],s102[197],s101[199],s100[201],pp127[94],pp126[96],pp125[98],pp99[125],pp99[126],pp99[127]};
    CLA_198 KS_110(s110, c110, in110_1, in110_2);
    wire[195:0] s111, in111_1, in111_2;
    wire c111;
    assign in111_1 = {pp26[4],pp25[6],pp26[6],pp27[6],pp28[6],pp29[6],pp30[6],pp31[6],pp32[6],s110[10],s110[11],s110[12],s110[13],s110[14],s110[15],s110[16],s110[17],s110[18],s110[19],s110[20],s110[21],s110[22],s110[23],s110[24],s110[25],s110[26],s110[27],s110[28],s110[29],s110[30],s110[31],s110[32],s110[33],s110[34],s110[35],s110[36],s110[37],s110[38],s110[39],s110[40],s110[41],s110[42],s110[43],s110[44],s110[45],s110[46],s110[47],s110[48],s110[49],s110[50],s110[51],s110[52],s110[53],s110[54],s110[55],s110[56],s110[57],s110[58],s110[59],s110[60],s110[61],s110[62],s110[63],s110[64],s110[65],s110[66],s110[67],s110[68],s110[69],s110[70],s110[71],s110[72],s110[73],s110[74],s110[75],s110[76],s110[77],s110[78],s110[79],s110[80],s110[81],s110[82],s110[83],s110[84],s110[85],s110[86],s110[87],s110[88],s110[89],s110[90],s110[91],s110[92],s110[93],s110[94],s110[95],s110[96],s110[97],s110[98],s110[99],s110[100],s110[101],s110[102],s110[103],s110[104],s110[105],s110[106],s110[107],s110[108],s110[109],s110[110],s110[111],s110[112],s110[113],s110[114],s110[115],s110[116],s110[117],s110[118],s110[119],s110[120],s110[121],s110[122],s110[123],s110[124],s110[125],s110[126],s110[127],s110[128],s110[129],s110[130],s110[131],s110[132],s110[133],s110[134],s110[135],s110[136],s110[137],s110[138],s110[139],s110[140],s110[141],s110[142],s110[143],s110[144],s110[145],s110[146],s110[147],s110[148],s110[149],s110[150],s110[151],s110[152],s110[153],s110[154],s110[155],s110[156],s110[157],s110[158],s110[159],s110[160],s110[161],s110[162],s110[163],s110[164],s110[165],s110[166],s110[167],s110[168],s110[169],s110[170],s110[171],s110[172],s110[173],s110[174],s110[175],s110[176],s110[177],s110[178],s110[179],s110[180],s110[181],s110[182],s109[184],s108[186],s107[188],s106[190],s105[192],s104[194],s103[196],s102[198],s101[200],s100[202],pp127[95],pp126[97],pp125[99],pp126[99]};
    assign in111_2 = {pp27[3],pp26[5],pp27[5],pp28[5],pp29[5],pp30[5],pp31[5],pp32[5],pp33[5],pp34[5],pp36[4],pp38[3],pp40[2],pp42[1],pp44[0],s65[13],s66[13],s67[13],s68[13],s69[13],s70[13],s71[13],s72[13],s73[13],s74[13],s75[13],s76[13],s77[13],s78[13],s79[13],s80[13],s81[13],s82[13],s83[13],s84[13],s85[13],s86[13],s87[13],s88[13],s89[13],s90[13],s91[13],s92[13],s93[13],s94[13],s95[13],s96[13],s97[61],s98[61],s99[61],s1[16],s2[16],s3[16],s3[17],s3[18],s3[19],s3[20],s3[21],s3[22],s3[23],s3[24],s3[25],s3[26],s3[27],s3[28],s3[29],s3[30],s3[31],s3[32],s3[33],s3[34],s3[35],s3[36],s3[37],s3[38],s3[39],s3[40],s3[41],s3[42],s3[43],s3[44],s3[45],s3[46],s3[47],s3[48],s3[49],s3[50],s3[51],s3[52],s3[53],s3[54],s3[55],s3[56],s3[57],s3[58],s3[59],s3[60],s3[61],s3[62],s1[65],s95[68],s93[71],s91[74],s90[76],s90[77],s90[78],s90[79],s90[80],s90[81],s90[82],s90[83],s90[84],s90[85],s90[86],s90[87],s90[88],s90[89],s90[90],s90[91],s90[92],s90[93],s90[94],s90[95],s90[96],s90[97],s90[98],s90[99],s35[59],s33[62],s31[65],s29[68],s27[71],s25[74],s23[77],s21[80],s19[83],s17[86],s15[89],s13[92],s11[95],s7[100],s6[102],s5[104],s3[107],s1[110],s98[158],s96[113],s94[116],s93[118],s93[119],s93[120],s93[121],s93[122],s93[123],s92[125],s91[127],s90[129],s89[131],s88[133],s87[135],s86[137],s85[139],s84[141],s83[143],s82[145],s81[147],s80[149],s79[151],s78[153],s77[155],s76[157],s75[159],s74[161],s73[163],s72[165],s71[167],s70[169],s69[171],s68[173],s67[175],s66[177],s65[179],s110[183],s109[185],s108[187],s107[189],s106[191],s105[193],s104[195],s103[197],s102[199],s101[201],s100[203],pp127[96],pp126[98],pp127[98]};
    CLA_196 KS_111(s111, c111, in111_1, in111_2);
    wire[193:0] s112, in112_1, in112_2;
    wire c112;
    assign in112_1 = {pp27[4],pp28[4],pp29[4],pp30[4],pp31[4],pp32[4],pp33[4],pp34[4],pp35[4],s111[10],s111[11],s111[12],s111[13],s111[14],s111[15],s111[16],s111[17],s111[18],s111[19],s111[20],s111[21],s111[22],s111[23],s111[24],s111[25],s111[26],s111[27],s111[28],s111[29],s111[30],s111[31],s111[32],s111[33],s111[34],s111[35],s111[36],s111[37],s111[38],s111[39],s111[40],s111[41],s111[42],s111[43],s111[44],s111[45],s111[46],s111[47],s111[48],s111[49],s111[50],s111[51],s111[52],s111[53],s111[54],s111[55],s111[56],s111[57],s111[58],s111[59],s111[60],s111[61],s111[62],s111[63],s111[64],s111[65],s111[66],s111[67],s111[68],s111[69],s111[70],s111[71],s111[72],s111[73],s111[74],s111[75],s111[76],s111[77],s111[78],s111[79],s111[80],s111[81],s111[82],s111[83],s111[84],s111[85],s111[86],s111[87],s111[88],s111[89],s111[90],s111[91],s111[92],s111[93],s111[94],s111[95],s111[96],s111[97],s111[98],s111[99],s111[100],s111[101],s111[102],s111[103],s111[104],s111[105],s111[106],s111[107],s111[108],s111[109],s111[110],s111[111],s111[112],s111[113],s111[114],s111[115],s111[116],s111[117],s111[118],s111[119],s111[120],s111[121],s111[122],s111[123],s111[124],s111[125],s111[126],s111[127],s111[128],s111[129],s111[130],s111[131],s111[132],s111[133],s111[134],s111[135],s111[136],s111[137],s111[138],s111[139],s111[140],s111[141],s111[142],s111[143],s111[144],s111[145],s111[146],s111[147],s111[148],s111[149],s111[150],s111[151],s111[152],s111[153],s111[154],s111[155],s111[156],s111[157],s111[158],s111[159],s111[160],s111[161],s111[162],s111[163],s111[164],s111[165],s111[166],s111[167],s111[168],s111[169],s111[170],s111[171],s111[172],s111[173],s111[174],s111[175],s111[176],s111[177],s111[178],s111[179],s111[180],s111[181],s111[182],s110[184],s109[186],s108[188],s107[190],s106[192],s105[194],s104[196],s103[198],s102[200],s101[202],s100[204],pp127[97]};
    assign in112_2 = {pp28[3],pp29[3],pp30[3],pp31[3],pp32[3],pp33[3],pp34[3],pp35[3],pp36[3],pp37[3],pp39[2],pp41[1],pp43[0],s65[12],s66[12],s67[12],s68[12],s69[12],s70[12],s71[12],s72[12],s73[12],s74[12],s75[12],s76[12],s77[12],s78[12],s79[12],s80[12],s81[12],s82[12],s83[12],s84[12],s85[12],s86[12],s87[12],s88[12],s89[12],s90[12],s91[12],s92[12],s93[12],s94[12],s95[12],s96[12],s97[60],s98[60],s99[60],s1[15],s2[15],s3[15],s4[15],s4[16],s4[17],s4[18],s4[19],s4[20],s4[21],s4[22],s4[23],s4[24],s4[25],s4[26],s4[27],s4[28],s4[29],s4[30],s4[31],s4[32],s4[33],s4[34],s4[35],s4[36],s4[37],s4[38],s4[39],s4[40],s4[41],s4[42],s4[43],s4[44],s4[45],s4[46],s4[47],s4[48],s4[49],s4[50],s4[51],s4[52],s4[53],s4[54],s4[55],s4[56],s4[57],s4[58],s4[59],s4[60],s4[61],s2[64],s96[67],s94[70],s92[73],s91[75],s91[76],s91[77],s91[78],s91[79],s91[80],s91[81],s91[82],s91[83],s91[84],s91[85],s91[86],s91[87],s91[88],s91[89],s91[90],s91[91],s91[92],s91[93],s91[94],s91[95],s91[96],s91[97],s91[98],s91[99],s34[61],s32[64],s30[67],s28[70],s26[73],s24[76],s22[79],s20[82],s18[85],s16[88],s14[91],s12[94],s10[97],s7[101],s6[103],s4[106],s2[109],s99[157],s97[160],s95[115],s94[117],s94[118],s94[119],s94[120],s94[121],s94[122],s93[124],s92[126],s91[128],s90[130],s89[132],s88[134],s87[136],s86[138],s85[140],s84[142],s83[144],s82[146],s81[148],s80[150],s79[152],s78[154],s77[156],s76[158],s75[160],s74[162],s73[164],s72[166],s71[168],s70[170],s69[172],s68[174],s67[176],s66[178],s65[180],s111[183],s110[185],s109[187],s108[189],s107[191],s106[193],s105[195],s104[197],s103[199],s102[201],s101[203],s100[205]};
    CLA_194 KS_112(s112, c112, in112_1, in112_2);

    /*Stage 4*/
    wire[239:0] s113, in113_1, in113_2;
    wire c113;
    assign in113_1 = {pp0[8],pp0[9],pp0[10],pp0[11],pp0[12],pp0[13],pp0[14],pp0[15],pp2[14],pp4[13],pp6[12],pp8[11],pp9[11],pp12[9],pp14[8],pp16[7],pp18[6],pp20[5],pp22[4],pp24[3],pp26[2],pp27[2],pp28[2],pp29[2],pp30[2],pp31[2],pp32[2],pp33[2],pp34[2],pp35[2],pp36[2],pp37[2],pp38[2],s112[10],s112[11],s112[12],s112[13],s112[14],s112[15],s112[16],s112[17],s112[18],s112[19],s112[20],s112[21],s112[22],s112[23],s112[24],s112[25],s112[26],s112[27],s112[28],s112[29],s112[30],s112[31],s112[32],s112[33],s112[34],s112[35],s112[36],s112[37],s112[38],s112[39],s112[40],s112[41],s112[42],s112[43],s112[44],s112[45],s112[46],s112[47],s112[48],s112[49],s112[50],s112[51],s112[52],s112[53],s112[54],s112[55],s112[56],s112[57],s112[58],s112[59],s112[60],s112[61],s112[62],s112[63],s112[64],s112[65],s112[66],s112[67],s112[68],s112[69],s112[70],s112[71],s112[72],s112[73],s112[74],s112[75],s112[76],s112[77],s112[78],s112[79],s112[80],s112[81],s112[82],s112[83],s112[84],s112[85],s112[86],s112[87],s112[88],s112[89],s112[90],s112[91],s112[92],s112[93],s112[94],s112[95],s112[96],s112[97],s112[98],s112[99],s112[100],s112[101],s112[102],s112[103],s112[104],s112[105],s112[106],s112[107],s112[108],s112[109],s112[110],s112[111],s112[112],s112[113],s112[114],s112[115],s112[116],s112[117],s112[118],s112[119],s112[120],s112[121],s112[122],s112[123],s112[124],s112[125],s112[126],s112[127],s112[128],s112[129],s112[130],s112[131],s112[132],s112[133],s112[134],s112[135],s112[136],s112[137],s112[138],s112[139],s112[140],s112[141],s112[142],s112[143],s112[144],s112[145],s112[146],s112[147],s112[148],s112[149],s112[150],s112[151],s112[152],s112[153],s112[154],s112[155],s112[156],s112[157],s112[158],s112[159],s112[160],s112[161],s112[162],s112[163],s112[164],s112[165],s112[166],s112[167],s112[168],s112[169],s112[170],s112[171],s112[172],s112[173],s112[174],s112[175],s112[176],s112[177],s112[178],s112[179],s112[180],s112[181],s112[182],s111[184],s110[186],s109[188],s108[190],s107[192],s106[194],s105[196],s104[198],s103[200],s102[202],s101[204],s100[206],pp127[99],pp126[101],pp125[103],pp124[105],pp123[107],pp122[109],pp121[111],pp120[113],pp119[115],pp118[117],pp117[119],pp116[121],pp115[123],pp114[125],pp113[127],pp114[127],pp115[127],pp116[127],pp117[127],pp118[127],pp119[127],pp120[127]};
    assign in113_2 = {pp1[7],pp1[8],pp10[0],pp1[10],pp1[11],pp1[12],pp1[13],pp1[14],pp3[13],pp5[12],pp7[11],pp9[10],pp11[9],pp13[8],pp15[7],pp17[6],pp19[5],pp21[4],pp23[3],pp25[2],pp27[1],pp28[1],pp29[1],pp30[1],pp31[1],pp32[1],pp33[1],pp34[1],pp35[1],pp36[1],pp37[1],pp38[1],pp39[1],pp40[1],pp42[0],s65[11],s66[11],s67[11],s68[11],s69[11],s70[11],s71[11],s72[11],s73[11],s74[11],s75[11],s76[11],s77[11],s78[11],s79[11],s80[11],s81[11],s82[11],s83[11],s84[11],s85[11],s86[11],s87[11],s88[11],s89[11],s90[11],s91[11],s92[11],s93[11],s94[11],s95[11],s96[11],s97[59],s98[59],s99[59],s1[14],s2[14],s3[14],s4[14],s5[14],s5[15],s5[16],s5[17],s5[18],s5[19],s5[20],s5[21],s5[22],s5[23],s5[24],s5[25],s5[26],s5[27],s5[28],s5[29],s5[30],s5[31],s5[32],s5[33],s5[34],s5[35],s5[36],s5[37],s5[38],s5[39],s5[40],s5[41],s5[42],s5[43],s5[44],s5[45],s5[46],s5[47],s5[48],s5[49],s5[50],s5[51],s5[52],s5[53],s5[54],s5[55],s5[56],s5[57],s5[58],s5[59],s5[60],s3[63],s1[66],s95[69],s93[72],s92[74],s92[75],s92[76],s92[77],s92[78],s92[79],s92[80],s92[81],s92[82],s92[83],s92[84],s92[85],s92[86],s92[87],s92[88],s92[89],s92[90],s92[91],s92[92],s92[93],s92[94],s92[95],s92[96],s92[97],s92[98],s92[99],s33[63],s31[66],s29[69],s27[72],s25[75],s23[78],s21[81],s19[84],s17[87],s15[90],s13[93],s11[96],s8[100],s7[102],s5[105],s3[108],s1[111],s98[159],s96[114],s95[116],s95[117],s95[118],s95[119],s95[120],s95[121],s94[123],s93[125],s92[127],s91[129],s90[131],s89[133],s88[135],s87[137],s86[139],s85[141],s84[143],s83[145],s82[147],s81[149],s80[151],s79[153],s78[155],s77[157],s76[159],s75[161],s74[163],s73[165],s72[167],s71[169],s70[171],s69[173],s68[175],s67[177],s66[179],s65[181],s112[183],s111[185],s110[187],s109[189],s108[191],s107[193],s106[195],s105[197],s104[199],s103[201],s102[203],s101[205],s100[207],pp127[100],pp126[102],pp125[104],pp124[106],pp123[108],pp122[110],pp121[112],pp120[114],pp119[116],pp118[118],pp117[120],pp116[122],pp115[124],pp114[126],pp115[126],pp116[126],pp117[126],pp118[126],pp119[126],pp120[126],pp121[126]};
    CLA_240 KS_113(s113, c113, in113_1, in113_2);
    wire[237:0] s114, in114_1, in114_2;
    wire c114;
    assign in114_1 = {pp2[7],s113[2],pp10[1],pp2[10],pp2[11],pp2[12],pp2[13],pp4[12],pp6[11],s113[10],s113[11],s113[12],s113[13],s113[14],s113[15],s113[16],s113[17],s113[18],s113[19],s113[20],s113[21],s113[22],s113[23],s113[24],s113[25],s113[26],s113[27],s113[28],s113[29],s113[30],s113[31],s113[32],s113[33],s113[34],s113[35],s113[36],s113[37],s113[38],s113[39],s113[40],s113[41],s113[42],s113[43],s113[44],s113[45],s113[46],s113[47],s113[48],s113[49],s113[50],s113[51],s113[52],s113[53],s113[54],s113[55],s113[56],s113[57],s113[58],s113[59],s113[60],s113[61],s113[62],s113[63],s113[64],s113[65],s113[66],s113[67],s113[68],s113[69],s113[70],s113[71],s113[72],s113[73],s113[74],s113[75],s113[76],s113[77],s113[78],s113[79],s113[80],s113[81],s113[82],s113[83],s113[84],s113[85],s113[86],s113[87],s113[88],s113[89],s113[90],s113[91],s113[92],s113[93],s113[94],s113[95],s113[96],s113[97],s113[98],s113[99],s113[100],s113[101],s113[102],s113[103],s113[104],s113[105],s113[106],s113[107],s113[108],s113[109],s113[110],s113[111],s113[112],s113[113],s113[114],s113[115],s113[116],s113[117],s113[118],s113[119],s113[120],s113[121],s113[122],s113[123],s113[124],s113[125],s113[126],s113[127],s113[128],s113[129],s113[130],s113[131],s113[132],s113[133],s113[134],s113[135],s113[136],s113[137],s113[138],s113[139],s113[140],s113[141],s113[142],s113[143],s113[144],s113[145],s113[146],s113[147],s113[148],s113[149],s113[150],s113[151],s113[152],s113[153],s113[154],s113[155],s113[156],s113[157],s113[158],s113[159],s113[160],s113[161],s113[162],s113[163],s113[164],s113[165],s113[166],s113[167],s113[168],s113[169],s113[170],s113[171],s113[172],s113[173],s113[174],s113[175],s113[176],s113[177],s113[178],s113[179],s113[180],s113[181],s113[182],s113[183],s113[184],s113[185],s113[186],s113[187],s113[188],s113[189],s113[190],s113[191],s113[192],s113[193],s113[194],s113[195],s113[196],s113[197],s113[198],s113[199],s113[200],s113[201],s113[202],s113[203],s113[204],s113[205],s113[206],s112[184],s111[186],s110[188],s109[190],s108[192],s107[194],s106[196],s105[198],s104[200],s103[202],s102[204],s101[206],s100[208],pp127[101],pp126[103],pp125[105],pp124[107],pp123[109],pp122[111],pp121[113],pp120[115],pp119[117],pp118[119],pp117[121],pp116[123],pp115[125],pp116[125],pp117[125],pp118[125],pp119[125],pp120[125],pp121[125]};
    assign in114_2 = {pp3[6],pp1[9],pp11[0],pp10[2],pp3[10],pp3[11],pp3[12],pp5[11],pp7[10],pp8[10],pp10[9],pp12[8],pp14[7],pp16[6],pp18[5],pp20[4],pp22[3],pp24[2],pp26[1],pp28[0],pp29[0],pp30[0],pp31[0],pp32[0],pp33[0],pp34[0],pp35[0],pp36[0],pp37[0],pp38[0],pp39[0],pp40[0],pp41[0],s65[10],s66[10],s67[10],s68[10],s69[10],s70[10],s71[10],s72[10],s73[10],s74[10],s75[10],s76[10],s77[10],s78[10],s79[10],s80[10],s81[10],s82[10],s83[10],s84[10],s85[10],s86[10],s87[10],s88[10],s89[10],s90[10],s91[10],s92[10],s93[10],s94[10],s95[10],s96[10],s97[58],s98[58],s99[58],s1[13],s2[13],s3[13],s4[13],s5[13],s6[13],s6[14],s6[15],s6[16],s6[17],s6[18],s6[19],s6[20],s6[21],s6[22],s6[23],s6[24],s6[25],s6[26],s6[27],s6[28],s6[29],s6[30],s6[31],s6[32],s6[33],s6[34],s6[35],s6[36],s6[37],s6[38],s6[39],s6[40],s6[41],s6[42],s6[43],s6[44],s6[45],s6[46],s6[47],s6[48],s6[49],s6[50],s6[51],s6[52],s6[53],s6[54],s6[55],s6[56],s6[57],s6[58],s6[59],s4[62],s2[65],s96[68],s94[71],s93[73],s93[74],s93[75],s93[76],s93[77],s93[78],s93[79],s93[80],s93[81],s93[82],s93[83],s93[84],s93[85],s93[86],s93[87],s93[88],s93[89],s93[90],s93[91],s93[92],s93[93],s93[94],s93[95],s93[96],s93[97],s93[98],s93[99],s32[65],s30[68],s28[71],s26[74],s24[77],s22[80],s20[83],s18[86],s16[89],s14[92],s12[95],s10[98],s8[101],s6[104],s4[107],s2[110],s99[158],s97[161],s96[115],s96[116],s96[117],s96[118],s96[119],s96[120],s95[122],s94[124],s93[126],s92[128],s91[130],s90[132],s89[134],s88[136],s87[138],s86[140],s85[142],s84[144],s83[146],s82[148],s81[150],s80[152],s79[154],s78[156],s77[158],s76[160],s75[162],s74[164],s73[166],s72[168],s71[170],s70[172],s69[174],s68[176],s67[178],s66[180],s65[182],s113[207],s112[185],s111[187],s110[189],s109[191],s108[193],s107[195],s106[197],s105[199],s104[201],s103[203],s102[205],s101[207],s100[209],pp127[102],pp126[104],pp125[106],pp124[108],pp123[110],pp122[112],pp121[114],pp120[116],pp119[118],pp118[120],pp117[122],pp116[124],pp117[124],pp118[124],pp119[124],pp120[124],pp121[124],pp122[124]};
    CLA_238 KS_114(s114, c114, in114_1, in114_2);
    wire[235:0] s115, in115_1, in115_2;
    wire c115;
    assign in115_1 = {pp2[8],s113[3],pp11[1],pp10[3],pp4[10],pp4[11],pp6[10],pp10[7],pp10[8],s114[10],s114[11],s114[12],s114[13],s114[14],s114[15],s114[16],s114[17],s114[18],s114[19],s114[20],s114[21],s114[22],s114[23],s114[24],s114[25],s114[26],s114[27],s114[28],s114[29],s114[30],s114[31],s114[32],s114[33],s114[34],s114[35],s114[36],s114[37],s114[38],s114[39],s114[40],s114[41],s114[42],s114[43],s114[44],s114[45],s114[46],s114[47],s114[48],s114[49],s114[50],s114[51],s114[52],s114[53],s114[54],s114[55],s114[56],s114[57],s114[58],s114[59],s114[60],s114[61],s114[62],s114[63],s114[64],s114[65],s114[66],s114[67],s114[68],s114[69],s114[70],s114[71],s114[72],s114[73],s114[74],s114[75],s114[76],s114[77],s114[78],s114[79],s114[80],s114[81],s114[82],s114[83],s114[84],s114[85],s114[86],s114[87],s114[88],s114[89],s114[90],s114[91],s114[92],s114[93],s114[94],s114[95],s114[96],s114[97],s114[98],s114[99],s114[100],s114[101],s114[102],s114[103],s114[104],s114[105],s114[106],s114[107],s114[108],s114[109],s114[110],s114[111],s114[112],s114[113],s114[114],s114[115],s114[116],s114[117],s114[118],s114[119],s114[120],s114[121],s114[122],s114[123],s114[124],s114[125],s114[126],s114[127],s114[128],s114[129],s114[130],s114[131],s114[132],s114[133],s114[134],s114[135],s114[136],s114[137],s114[138],s114[139],s114[140],s114[141],s114[142],s114[143],s114[144],s114[145],s114[146],s114[147],s114[148],s114[149],s114[150],s114[151],s114[152],s114[153],s114[154],s114[155],s114[156],s114[157],s114[158],s114[159],s114[160],s114[161],s114[162],s114[163],s114[164],s114[165],s114[166],s114[167],s114[168],s114[169],s114[170],s114[171],s114[172],s114[173],s114[174],s114[175],s114[176],s114[177],s114[178],s114[179],s114[180],s114[181],s114[182],s114[183],s114[184],s114[185],s114[186],s114[187],s114[188],s114[189],s114[190],s114[191],s114[192],s114[193],s114[194],s114[195],s114[196],s114[197],s114[198],s114[199],s114[200],s114[201],s114[202],s114[203],s114[204],s114[205],s114[206],s113[208],s112[186],s111[188],s110[190],s109[192],s108[194],s107[196],s106[198],s105[200],s104[202],s103[204],s102[206],s101[208],s100[210],pp127[103],pp126[105],pp125[107],pp124[109],pp123[111],pp122[113],pp121[115],pp120[117],pp119[119],pp118[121],pp117[123],pp118[123],pp119[123],pp120[123],pp121[123],pp122[123]};
    assign in115_2 = {pp3[7],s114[2],pp12[0],pp11[2],pp10[4],pp5[10],pp10[6],pp11[6],pp11[7],pp11[8],pp13[7],pp15[6],pp17[5],pp19[4],pp21[3],pp23[2],pp25[1],pp27[0],s97[12],s97[13],s97[14],s97[15],s97[16],s97[17],s97[18],s97[19],s97[20],s97[21],s97[22],s97[23],s97[24],s97[25],s97[26],s97[27],s97[28],s97[29],s97[30],s97[31],s97[32],s97[33],s97[34],s97[35],s97[36],s97[37],s97[38],s97[39],s97[40],s97[41],s97[42],s97[43],s97[44],s97[45],s97[46],s97[47],s97[48],s97[49],s97[50],s97[51],s97[52],s97[53],s97[54],s97[55],s97[56],s97[57],s98[57],s99[57],s1[12],s2[12],s3[12],s4[12],s5[12],s6[12],s7[12],s7[13],s7[14],s7[15],s7[16],s7[17],s7[18],s7[19],s7[20],s7[21],s7[22],s7[23],s7[24],s7[25],s7[26],s7[27],s7[28],s7[29],s7[30],s7[31],s7[32],s7[33],s7[34],s7[35],s7[36],s7[37],s7[38],s7[39],s7[40],s7[41],s7[42],s7[43],s7[44],s7[45],s7[46],s7[47],s7[48],s7[49],s7[50],s7[51],s7[52],s7[53],s7[54],s7[55],s7[56],s7[57],s7[58],s5[61],s3[64],s1[67],s95[70],s94[72],s94[73],s94[74],s94[75],s94[76],s94[77],s94[78],s94[79],s94[80],s94[81],s94[82],s94[83],s94[84],s94[85],s94[86],s94[87],s94[88],s94[89],s94[90],s94[91],s94[92],s94[93],s94[94],s94[95],s94[96],s94[97],s94[98],s94[99],s31[67],s29[70],s27[73],s25[76],s23[79],s21[82],s19[85],s17[88],s15[91],s13[94],s11[97],s9[100],s7[103],s5[106],s3[109],s1[112],s98[160],s97[162],s97[163],s97[164],s97[165],s97[166],s97[167],s96[121],s95[123],s94[125],s93[127],s92[129],s91[131],s90[133],s89[135],s88[137],s87[139],s86[141],s85[143],s84[145],s83[147],s82[149],s81[151],s80[153],s79[155],s78[157],s77[159],s76[161],s75[163],s74[165],s73[167],s72[169],s71[171],s70[173],s69[175],s68[177],s67[179],s66[181],s65[183],s114[207],s113[209],s112[187],s111[189],s110[191],s109[193],s108[195],s107[197],s106[199],s105[201],s104[203],s103[205],s102[207],s101[209],s100[211],pp127[104],pp126[106],pp125[108],pp124[110],pp123[112],pp122[114],pp121[116],pp120[118],pp119[120],pp118[122],pp119[122],pp120[122],pp121[122],pp122[122],pp123[122]};
    CLA_236 KS_115(s115, c115, in115_1, in115_2);
    wire[233:0] s116, in116_1, in116_2;
    wire c116;
    assign in116_1 = {pp2[9],s113[4],pp12[1],pp11[3],pp10[5],pp11[5],pp12[5],pp12[6],pp12[7],s115[10],s115[11],s115[12],s115[13],s115[14],s115[15],s115[16],s115[17],s115[18],s115[19],s115[20],s115[21],s115[22],s115[23],s115[24],s115[25],s115[26],s115[27],s115[28],s115[29],s115[30],s115[31],s115[32],s115[33],s115[34],s115[35],s115[36],s115[37],s115[38],s115[39],s115[40],s115[41],s115[42],s115[43],s115[44],s115[45],s115[46],s115[47],s115[48],s115[49],s115[50],s115[51],s115[52],s115[53],s115[54],s115[55],s115[56],s115[57],s115[58],s115[59],s115[60],s115[61],s115[62],s115[63],s115[64],s115[65],s115[66],s115[67],s115[68],s115[69],s115[70],s115[71],s115[72],s115[73],s115[74],s115[75],s115[76],s115[77],s115[78],s115[79],s115[80],s115[81],s115[82],s115[83],s115[84],s115[85],s115[86],s115[87],s115[88],s115[89],s115[90],s115[91],s115[92],s115[93],s115[94],s115[95],s115[96],s115[97],s115[98],s115[99],s115[100],s115[101],s115[102],s115[103],s115[104],s115[105],s115[106],s115[107],s115[108],s115[109],s115[110],s115[111],s115[112],s115[113],s115[114],s115[115],s115[116],s115[117],s115[118],s115[119],s115[120],s115[121],s115[122],s115[123],s115[124],s115[125],s115[126],s115[127],s115[128],s115[129],s115[130],s115[131],s115[132],s115[133],s115[134],s115[135],s115[136],s115[137],s115[138],s115[139],s115[140],s115[141],s115[142],s115[143],s115[144],s115[145],s115[146],s115[147],s115[148],s115[149],s115[150],s115[151],s115[152],s115[153],s115[154],s115[155],s115[156],s115[157],s115[158],s115[159],s115[160],s115[161],s115[162],s115[163],s115[164],s115[165],s115[166],s115[167],s115[168],s115[169],s115[170],s115[171],s115[172],s115[173],s115[174],s115[175],s115[176],s115[177],s115[178],s115[179],s115[180],s115[181],s115[182],s115[183],s115[184],s115[185],s115[186],s115[187],s115[188],s115[189],s115[190],s115[191],s115[192],s115[193],s115[194],s115[195],s115[196],s115[197],s115[198],s115[199],s115[200],s115[201],s115[202],s115[203],s115[204],s115[205],s115[206],s114[208],s113[210],s112[188],s111[190],s110[192],s109[194],s108[196],s107[198],s106[200],s105[202],s104[204],s103[206],s102[208],s101[210],s100[212],pp127[105],pp126[107],pp125[109],pp124[111],pp123[113],pp122[115],pp121[117],pp120[119],pp119[121],pp120[121],pp121[121],pp122[121],pp123[121]};
    assign in116_2 = {pp3[8],s114[3],pp13[0],pp12[2],pp11[4],pp12[4],pp13[4],pp13[5],pp13[6],pp14[6],pp16[5],pp18[4],pp20[3],pp22[2],pp24[1],pp26[0],s97[11],s98[11],s98[12],s98[13],s98[14],s98[15],s98[16],s98[17],s98[18],s98[19],s98[20],s98[21],s98[22],s98[23],s98[24],s98[25],s98[26],s98[27],s98[28],s98[29],s98[30],s98[31],s98[32],s98[33],s98[34],s98[35],s98[36],s98[37],s98[38],s98[39],s98[40],s98[41],s98[42],s98[43],s98[44],s98[45],s98[46],s98[47],s98[48],s98[49],s98[50],s98[51],s98[52],s98[53],s98[54],s98[55],s98[56],s99[56],s1[11],s2[11],s3[11],s4[11],s5[11],s6[11],s7[11],s8[11],s8[12],s8[13],s8[14],s8[15],s8[16],s8[17],s8[18],s8[19],s8[20],s8[21],s8[22],s8[23],s8[24],s8[25],s8[26],s8[27],s8[28],s8[29],s8[30],s8[31],s8[32],s8[33],s8[34],s8[35],s8[36],s8[37],s8[38],s8[39],s8[40],s8[41],s8[42],s8[43],s8[44],s8[45],s8[46],s8[47],s8[48],s8[49],s8[50],s8[51],s8[52],s8[53],s8[54],s8[55],s8[56],s8[57],s6[60],s4[63],s2[66],s96[69],s95[71],s95[72],s95[73],s95[74],s95[75],s95[76],s95[77],s95[78],s95[79],s95[80],s95[81],s95[82],s95[83],s95[84],s95[85],s95[86],s95[87],s95[88],s95[89],s95[90],s95[91],s95[92],s95[93],s95[94],s95[95],s95[96],s95[97],s95[98],s95[99],s30[69],s28[72],s26[75],s24[78],s22[81],s20[84],s18[87],s16[90],s14[93],s12[96],s10[99],s8[102],s6[105],s4[108],s2[111],s99[159],s98[161],s98[162],s98[163],s98[164],s98[165],s98[166],s97[168],s96[122],s95[124],s94[126],s93[128],s92[130],s91[132],s90[134],s89[136],s88[138],s87[140],s86[142],s85[144],s84[146],s83[148],s82[150],s81[152],s80[154],s79[156],s78[158],s77[160],s76[162],s75[164],s74[166],s73[168],s72[170],s71[172],s70[174],s69[176],s68[178],s67[180],s66[182],s65[184],s115[207],s114[209],s113[211],s112[189],s111[191],s110[193],s109[195],s108[197],s107[199],s106[201],s105[203],s104[205],s103[207],s102[209],s101[211],s100[213],pp127[106],pp126[108],pp125[110],pp124[112],pp123[114],pp122[116],pp121[118],pp120[120],pp121[120],pp122[120],pp123[120],pp124[120]};
    CLA_234 KS_116(s116, c116, in116_1, in116_2);
    wire[231:0] s117, in117_1, in117_2;
    wire c117;
    assign in117_1 = {s115[2],s113[5],pp13[1],pp12[3],pp13[3],pp14[3],pp14[4],pp14[5],pp15[5],s116[10],s116[11],s116[12],s116[13],s116[14],s116[15],s116[16],s116[17],s116[18],s116[19],s116[20],s116[21],s116[22],s116[23],s116[24],s116[25],s116[26],s116[27],s116[28],s116[29],s116[30],s116[31],s116[32],s116[33],s116[34],s116[35],s116[36],s116[37],s116[38],s116[39],s116[40],s116[41],s116[42],s116[43],s116[44],s116[45],s116[46],s116[47],s116[48],s116[49],s116[50],s116[51],s116[52],s116[53],s116[54],s116[55],s116[56],s116[57],s116[58],s116[59],s116[60],s116[61],s116[62],s116[63],s116[64],s116[65],s116[66],s116[67],s116[68],s116[69],s116[70],s116[71],s116[72],s116[73],s116[74],s116[75],s116[76],s116[77],s116[78],s116[79],s116[80],s116[81],s116[82],s116[83],s116[84],s116[85],s116[86],s116[87],s116[88],s116[89],s116[90],s116[91],s116[92],s116[93],s116[94],s116[95],s116[96],s116[97],s116[98],s116[99],s116[100],s116[101],s116[102],s116[103],s116[104],s116[105],s116[106],s116[107],s116[108],s116[109],s116[110],s116[111],s116[112],s116[113],s116[114],s116[115],s116[116],s116[117],s116[118],s116[119],s116[120],s116[121],s116[122],s116[123],s116[124],s116[125],s116[126],s116[127],s116[128],s116[129],s116[130],s116[131],s116[132],s116[133],s116[134],s116[135],s116[136],s116[137],s116[138],s116[139],s116[140],s116[141],s116[142],s116[143],s116[144],s116[145],s116[146],s116[147],s116[148],s116[149],s116[150],s116[151],s116[152],s116[153],s116[154],s116[155],s116[156],s116[157],s116[158],s116[159],s116[160],s116[161],s116[162],s116[163],s116[164],s116[165],s116[166],s116[167],s116[168],s116[169],s116[170],s116[171],s116[172],s116[173],s116[174],s116[175],s116[176],s116[177],s116[178],s116[179],s116[180],s116[181],s116[182],s116[183],s116[184],s116[185],s116[186],s116[187],s116[188],s116[189],s116[190],s116[191],s116[192],s116[193],s116[194],s116[195],s116[196],s116[197],s116[198],s116[199],s116[200],s116[201],s116[202],s116[203],s116[204],s116[205],s116[206],s115[208],s114[210],s113[212],s112[190],s111[192],s110[194],s109[196],s108[198],s107[200],s106[202],s105[204],s104[206],s103[208],s102[210],s101[212],s100[214],pp127[107],pp126[109],pp125[111],pp124[113],pp123[115],pp122[117],pp121[119],pp122[119],pp123[119],pp124[119]};
    assign in117_2 = {pp3[9],s114[4],pp14[0],pp13[2],pp14[2],pp15[2],pp15[3],pp15[4],pp16[4],pp17[4],pp19[3],pp21[2],pp23[1],pp25[0],s97[10],s98[10],s99[10],s99[11],s99[12],s99[13],s99[14],s99[15],s99[16],s99[17],s99[18],s99[19],s99[20],s99[21],s99[22],s99[23],s99[24],s99[25],s99[26],s99[27],s99[28],s99[29],s99[30],s99[31],s99[32],s99[33],s99[34],s99[35],s99[36],s99[37],s99[38],s99[39],s99[40],s99[41],s99[42],s99[43],s99[44],s99[45],s99[46],s99[47],s99[48],s99[49],s99[50],s99[51],s99[52],s99[53],s99[54],s99[55],s1[10],s2[10],s3[10],s4[10],s5[10],s6[10],s7[10],s8[10],s9[10],s9[11],s9[12],s9[13],s9[14],s9[15],s9[16],s9[17],s9[18],s9[19],s9[20],s9[21],s9[22],s9[23],s9[24],s9[25],s9[26],s9[27],s9[28],s9[29],s9[30],s9[31],s9[32],s9[33],s9[34],s9[35],s9[36],s9[37],s9[38],s9[39],s9[40],s9[41],s9[42],s9[43],s9[44],s9[45],s9[46],s9[47],s9[48],s9[49],s9[50],s9[51],s9[52],s9[53],s9[54],s9[55],s9[56],s7[59],s5[62],s3[65],s1[68],s96[70],s96[71],s96[72],s96[73],s96[74],s96[75],s96[76],s96[77],s96[78],s96[79],s96[80],s96[81],s96[82],s96[83],s96[84],s96[85],s96[86],s96[87],s96[88],s96[89],s96[90],s96[91],s96[92],s96[93],s96[94],s96[95],s96[96],s96[97],s96[98],s96[99],s29[71],s27[74],s25[77],s23[80],s21[83],s19[86],s17[89],s15[92],s13[95],s11[98],s9[101],s7[104],s5[107],s3[110],s1[113],s99[160],s99[161],s99[162],s99[163],s99[164],s99[165],s98[167],s97[169],s96[123],s95[125],s94[127],s93[129],s92[131],s91[133],s90[135],s89[137],s88[139],s87[141],s86[143],s85[145],s84[147],s83[149],s82[151],s81[153],s80[155],s79[157],s78[159],s77[161],s76[163],s75[165],s74[167],s73[169],s72[171],s71[173],s70[175],s69[177],s68[179],s67[181],s66[183],s65[185],s116[207],s115[209],s114[211],s113[213],s112[191],s111[193],s110[195],s109[197],s108[199],s107[201],s106[203],s105[205],s104[207],s103[209],s102[211],s101[213],s100[215],pp127[108],pp126[110],pp125[112],pp124[114],pp123[116],pp122[118],pp123[118],pp124[118],pp125[118]};
    CLA_232 KS_117(s117, c117, in117_1, in117_2);
    wire[229:0] s118, in118_1, in118_2;
    wire c118;
    assign in118_1 = {s115[3],s113[6],pp14[1],pp15[1],pp16[1],pp16[2],pp16[3],pp17[3],pp18[3],s117[10],s117[11],s117[12],s117[13],s117[14],s117[15],s117[16],s117[17],s117[18],s117[19],s117[20],s117[21],s117[22],s117[23],s117[24],s117[25],s117[26],s117[27],s117[28],s117[29],s117[30],s117[31],s117[32],s117[33],s117[34],s117[35],s117[36],s117[37],s117[38],s117[39],s117[40],s117[41],s117[42],s117[43],s117[44],s117[45],s117[46],s117[47],s117[48],s117[49],s117[50],s117[51],s117[52],s117[53],s117[54],s117[55],s117[56],s117[57],s117[58],s117[59],s117[60],s117[61],s117[62],s117[63],s117[64],s117[65],s117[66],s117[67],s117[68],s117[69],s117[70],s117[71],s117[72],s117[73],s117[74],s117[75],s117[76],s117[77],s117[78],s117[79],s117[80],s117[81],s117[82],s117[83],s117[84],s117[85],s117[86],s117[87],s117[88],s117[89],s117[90],s117[91],s117[92],s117[93],s117[94],s117[95],s117[96],s117[97],s117[98],s117[99],s117[100],s117[101],s117[102],s117[103],s117[104],s117[105],s117[106],s117[107],s117[108],s117[109],s117[110],s117[111],s117[112],s117[113],s117[114],s117[115],s117[116],s117[117],s117[118],s117[119],s117[120],s117[121],s117[122],s117[123],s117[124],s117[125],s117[126],s117[127],s117[128],s117[129],s117[130],s117[131],s117[132],s117[133],s117[134],s117[135],s117[136],s117[137],s117[138],s117[139],s117[140],s117[141],s117[142],s117[143],s117[144],s117[145],s117[146],s117[147],s117[148],s117[149],s117[150],s117[151],s117[152],s117[153],s117[154],s117[155],s117[156],s117[157],s117[158],s117[159],s117[160],s117[161],s117[162],s117[163],s117[164],s117[165],s117[166],s117[167],s117[168],s117[169],s117[170],s117[171],s117[172],s117[173],s117[174],s117[175],s117[176],s117[177],s117[178],s117[179],s117[180],s117[181],s117[182],s117[183],s117[184],s117[185],s117[186],s117[187],s117[188],s117[189],s117[190],s117[191],s117[192],s117[193],s117[194],s117[195],s117[196],s117[197],s117[198],s117[199],s117[200],s117[201],s117[202],s117[203],s117[204],s117[205],s117[206],s116[208],s115[210],s114[212],s113[214],s112[192],s111[194],s110[196],s109[198],s108[200],s107[202],s106[204],s105[206],s104[208],s103[210],s102[212],s101[214],s100[216],pp127[109],pp126[111],pp125[113],pp124[115],pp123[117],pp124[117],pp125[117]};
    assign in118_2 = {s116[2],s114[5],pp15[0],pp16[0],pp17[0],pp17[1],pp17[2],pp18[2],pp19[2],pp20[2],pp22[1],pp24[0],s100[6],s100[7],s100[8],s100[9],s101[9],s102[9],s103[9],s104[9],s105[9],s106[9],s107[9],s108[9],s109[9],s110[9],s111[9],s112[9],s65[9],s66[9],s67[9],s68[9],s69[9],s70[9],s71[9],s72[9],s73[9],s74[9],s75[9],s76[9],s77[9],s78[9],s79[9],s80[9],s81[9],s82[9],s83[9],s84[9],s85[9],s86[9],s87[9],s88[9],s89[9],s90[9],s91[9],s92[9],s93[9],s94[9],s95[9],s96[9],s10[0],s10[1],s10[2],s10[3],s10[4],s10[5],s10[6],s10[7],s10[8],s10[9],s11[9],s12[9],s13[9],s14[9],s15[9],s16[9],s17[9],s18[9],s19[9],s20[9],s21[9],s22[9],s23[9],s24[9],s25[9],s26[9],s27[9],s28[9],s29[9],s30[9],s31[9],s32[9],s33[9],s34[9],s35[9],s36[9],s37[9],s38[9],s39[9],s40[9],s41[9],s42[9],s43[9],s44[9],s45[9],s46[9],s47[9],s48[9],s49[9],s50[9],s51[9],s52[9],s53[9],s54[9],s55[9],s56[9],s8[58],s6[61],s4[64],s2[67],s1[69],s1[70],s1[71],s1[72],s1[73],s1[74],s1[75],s1[76],s1[77],s1[78],s1[79],s1[80],s1[81],s1[82],s1[83],s1[84],s1[85],s1[86],s1[87],s1[88],s1[89],s1[90],s1[91],s1[92],s1[93],s1[94],s1[95],s1[96],s1[97],s1[98],s1[99],s28[73],s26[76],s24[79],s22[82],s20[85],s18[88],s16[91],s14[94],s12[97],s11[99],s8[103],s6[106],s4[109],s2[112],s1[114],s1[115],s1[116],s1[117],s1[118],s1[119],s99[166],s98[168],s97[170],s96[124],s95[126],s94[128],s93[130],s92[132],s91[134],s90[136],s89[138],s88[140],s87[142],s86[144],s85[146],s84[148],s83[150],s82[152],s81[154],s80[156],s79[158],s78[160],s77[162],s76[164],s75[166],s74[168],s73[170],s72[172],s71[174],s70[176],s69[178],s68[180],s67[182],s66[184],s65[186],s117[207],s116[209],s115[211],s114[213],s113[215],s112[193],s111[195],s110[197],s109[199],s108[201],s107[203],s106[205],s105[207],s104[209],s103[211],s102[213],s101[215],s100[217],pp127[110],pp126[112],pp125[114],pp124[116],pp125[116],pp126[116]};
    CLA_230 KS_118(s118, c118, in118_1, in118_2);
    wire[227:0] s119, in119_1, in119_2;
    wire c119;
    assign in119_1 = {s115[4],s113[7],s113[8],s113[9],pp18[0],pp18[1],pp19[1],pp20[1],pp21[1],s118[10],s118[11],s118[12],s118[13],s118[14],s118[15],s118[16],s118[17],s118[18],s118[19],s118[20],s118[21],s118[22],s118[23],s118[24],s118[25],s118[26],s118[27],s118[28],s118[29],s118[30],s118[31],s118[32],s118[33],s118[34],s118[35],s118[36],s118[37],s118[38],s118[39],s118[40],s118[41],s118[42],s118[43],s118[44],s118[45],s118[46],s118[47],s118[48],s118[49],s118[50],s118[51],s118[52],s118[53],s118[54],s118[55],s118[56],s118[57],s118[58],s118[59],s118[60],s118[61],s118[62],s118[63],s118[64],s118[65],s118[66],s118[67],s118[68],s118[69],s118[70],s118[71],s118[72],s118[73],s118[74],s118[75],s118[76],s118[77],s118[78],s118[79],s118[80],s118[81],s118[82],s118[83],s118[84],s118[85],s118[86],s118[87],s118[88],s118[89],s118[90],s118[91],s118[92],s118[93],s118[94],s118[95],s118[96],s118[97],s118[98],s118[99],s118[100],s118[101],s118[102],s118[103],s118[104],s118[105],s118[106],s118[107],s118[108],s118[109],s118[110],s118[111],s118[112],s118[113],s118[114],s118[115],s118[116],s118[117],s118[118],s118[119],s118[120],s118[121],s118[122],s118[123],s118[124],s118[125],s118[126],s118[127],s118[128],s118[129],s118[130],s118[131],s118[132],s118[133],s118[134],s118[135],s118[136],s118[137],s118[138],s118[139],s118[140],s118[141],s118[142],s118[143],s118[144],s118[145],s118[146],s118[147],s118[148],s118[149],s118[150],s118[151],s118[152],s118[153],s118[154],s118[155],s118[156],s118[157],s118[158],s118[159],s118[160],s118[161],s118[162],s118[163],s118[164],s118[165],s118[166],s118[167],s118[168],s118[169],s118[170],s118[171],s118[172],s118[173],s118[174],s118[175],s118[176],s118[177],s118[178],s118[179],s118[180],s118[181],s118[182],s118[183],s118[184],s118[185],s118[186],s118[187],s118[188],s118[189],s118[190],s118[191],s118[192],s118[193],s118[194],s118[195],s118[196],s118[197],s118[198],s118[199],s118[200],s118[201],s118[202],s118[203],s118[204],s118[205],s118[206],s117[208],s116[210],s115[212],s114[214],s113[216],s113[217],s113[218],s113[219],s113[220],s113[221],s113[222],s113[223],s113[224],s113[225],s113[226],s113[227],s113[228],s113[229],pp127[111],pp126[113],pp125[115],pp126[115]};
    assign in119_2 = {s116[3],s114[6],s114[7],s114[8],s114[9],pp19[0],pp20[0],pp21[0],pp22[0],pp23[0],s100[5],s101[5],s101[6],s101[7],s101[8],s102[8],s103[8],s104[8],s105[8],s106[8],s107[8],s108[8],s109[8],s110[8],s111[8],s112[8],s65[8],s66[8],s67[8],s68[8],s69[8],s70[8],s71[8],s72[8],s73[8],s74[8],s75[8],s76[8],s77[8],s78[8],s79[8],s80[8],s81[8],s82[8],s83[8],s84[8],s85[8],s86[8],s87[8],s88[8],s89[8],s90[8],s91[8],s92[8],s93[8],s94[8],s95[8],s96[8],s1[8],s1[9],s11[0],s11[1],s11[2],s11[3],s11[4],s11[5],s11[6],s11[7],s11[8],s12[8],s13[8],s14[8],s15[8],s16[8],s17[8],s18[8],s19[8],s20[8],s21[8],s22[8],s23[8],s24[8],s25[8],s26[8],s27[8],s28[8],s29[8],s30[8],s31[8],s32[8],s33[8],s34[8],s35[8],s36[8],s37[8],s38[8],s39[8],s40[8],s41[8],s42[8],s43[8],s44[8],s45[8],s46[8],s47[8],s48[8],s49[8],s50[8],s51[8],s52[8],s53[8],s54[8],s55[8],s56[8],s57[8],s9[57],s7[60],s5[63],s3[66],s2[68],s2[69],s2[70],s2[71],s2[72],s2[73],s2[74],s2[75],s2[76],s2[77],s2[78],s2[79],s2[80],s2[81],s2[82],s2[83],s2[84],s2[85],s2[86],s2[87],s2[88],s2[89],s2[90],s2[91],s2[92],s2[93],s2[94],s2[95],s2[96],s2[97],s2[98],s2[99],s27[75],s25[78],s23[81],s21[84],s19[87],s17[90],s15[93],s13[96],s12[98],s9[102],s7[105],s5[108],s3[111],s2[113],s2[114],s2[115],s2[116],s2[117],s2[118],s1[120],s99[167],s98[169],s97[171],s96[125],s95[127],s94[129],s93[131],s92[133],s91[135],s90[137],s89[139],s88[141],s87[143],s86[145],s85[147],s84[149],s83[151],s82[153],s81[155],s80[157],s79[159],s78[161],s77[163],s76[165],s75[167],s74[169],s73[171],s72[173],s71[175],s70[177],s69[179],s68[181],s67[183],s66[185],s65[187],s118[207],s117[209],s116[211],s115[213],s114[215],s114[216],s114[217],s114[218],s114[219],s114[220],s114[221],s114[222],s114[223],s114[224],s114[225],s114[226],s114[227],s114[228],s113[230],pp127[112],pp126[114],pp127[114]};
    CLA_228 KS_119(s119, c119, in119_1, in119_2);
    wire[225:0] s120, in120_1, in120_2;
    wire c120;
    assign in120_1 = {s115[5],s115[6],s115[7],s115[8],s100[0],s100[1],s100[2],s100[3],s100[4],s119[10],s119[11],s119[12],s119[13],s119[14],s119[15],s119[16],s119[17],s119[18],s119[19],s119[20],s119[21],s119[22],s119[23],s119[24],s119[25],s119[26],s119[27],s119[28],s119[29],s119[30],s119[31],s119[32],s119[33],s119[34],s119[35],s119[36],s119[37],s119[38],s119[39],s119[40],s119[41],s119[42],s119[43],s119[44],s119[45],s119[46],s119[47],s119[48],s119[49],s119[50],s119[51],s119[52],s119[53],s119[54],s119[55],s119[56],s119[57],s119[58],s119[59],s119[60],s119[61],s119[62],s119[63],s119[64],s119[65],s119[66],s119[67],s119[68],s119[69],s119[70],s119[71],s119[72],s119[73],s119[74],s119[75],s119[76],s119[77],s119[78],s119[79],s119[80],s119[81],s119[82],s119[83],s119[84],s119[85],s119[86],s119[87],s119[88],s119[89],s119[90],s119[91],s119[92],s119[93],s119[94],s119[95],s119[96],s119[97],s119[98],s119[99],s119[100],s119[101],s119[102],s119[103],s119[104],s119[105],s119[106],s119[107],s119[108],s119[109],s119[110],s119[111],s119[112],s119[113],s119[114],s119[115],s119[116],s119[117],s119[118],s119[119],s119[120],s119[121],s119[122],s119[123],s119[124],s119[125],s119[126],s119[127],s119[128],s119[129],s119[130],s119[131],s119[132],s119[133],s119[134],s119[135],s119[136],s119[137],s119[138],s119[139],s119[140],s119[141],s119[142],s119[143],s119[144],s119[145],s119[146],s119[147],s119[148],s119[149],s119[150],s119[151],s119[152],s119[153],s119[154],s119[155],s119[156],s119[157],s119[158],s119[159],s119[160],s119[161],s119[162],s119[163],s119[164],s119[165],s119[166],s119[167],s119[168],s119[169],s119[170],s119[171],s119[172],s119[173],s119[174],s119[175],s119[176],s119[177],s119[178],s119[179],s119[180],s119[181],s119[182],s119[183],s119[184],s119[185],s119[186],s119[187],s119[188],s119[189],s119[190],s119[191],s119[192],s119[193],s119[194],s119[195],s119[196],s119[197],s119[198],s119[199],s119[200],s119[201],s119[202],s119[203],s119[204],s119[205],s119[206],s118[208],s117[210],s116[212],s115[214],s115[215],s115[216],s115[217],s115[218],s115[219],s115[220],s115[221],s115[222],s115[223],s115[224],s115[225],s115[226],s115[227],s114[229],s113[231],pp127[113]};
    assign in120_2 = {s116[4],s116[5],s116[6],s116[7],s115[9],s101[0],s101[1],s101[2],s101[3],s101[4],s102[4],s102[5],s102[6],s102[7],s103[7],s104[7],s105[7],s106[7],s107[7],s108[7],s109[7],s110[7],s111[7],s112[7],s65[7],s66[7],s67[7],s68[7],s69[7],s70[7],s71[7],s72[7],s73[7],s74[7],s75[7],s76[7],s77[7],s78[7],s79[7],s80[7],s81[7],s82[7],s83[7],s84[7],s85[7],s86[7],s87[7],s88[7],s89[7],s90[7],s91[7],s92[7],s93[7],s94[7],s95[7],s96[7],s1[7],s2[7],s2[8],s2[9],s12[0],s12[1],s12[2],s12[3],s12[4],s12[5],s12[6],s12[7],s13[7],s14[7],s15[7],s16[7],s17[7],s18[7],s19[7],s20[7],s21[7],s22[7],s23[7],s24[7],s25[7],s26[7],s27[7],s28[7],s29[7],s30[7],s31[7],s32[7],s33[7],s34[7],s35[7],s36[7],s37[7],s38[7],s39[7],s40[7],s41[7],s42[7],s43[7],s44[7],s45[7],s46[7],s47[7],s48[7],s49[7],s50[7],s51[7],s52[7],s53[7],s54[7],s55[7],s56[7],s57[7],s58[7],s57[9],s8[59],s6[62],s4[65],s3[67],s3[68],s3[69],s3[70],s3[71],s3[72],s3[73],s3[74],s3[75],s3[76],s3[77],s3[78],s3[79],s3[80],s3[81],s3[82],s3[83],s3[84],s3[85],s3[86],s3[87],s3[88],s3[89],s3[90],s3[91],s3[92],s3[93],s3[94],s3[95],s3[96],s3[97],s3[98],s3[99],s26[77],s24[80],s22[83],s20[86],s18[89],s16[92],s14[95],s13[97],s12[99],s8[104],s6[107],s4[110],s3[112],s3[113],s3[114],s3[115],s3[116],s3[117],s2[119],s1[121],s99[168],s98[170],s97[172],s96[126],s95[128],s94[130],s93[132],s92[134],s91[136],s90[138],s89[140],s88[142],s87[144],s86[146],s85[148],s84[150],s83[152],s82[154],s81[156],s80[158],s79[160],s78[162],s77[164],s76[166],s75[168],s74[170],s73[172],s72[174],s71[176],s70[178],s69[180],s68[182],s67[184],s66[186],s65[188],s119[207],s118[209],s117[211],s116[213],s116[214],s116[215],s116[216],s116[217],s116[218],s116[219],s116[220],s116[221],s116[222],s116[223],s116[224],s116[225],s116[226],s115[228],s114[230],s113[232]};
    CLA_226 KS_120(s120, c120, in120_1, in120_2);

    /*Stage 5*/
    wire[247:0] s121, in121_1, in121_2;
    wire c121;
    assign in121_1 = {pp0[4],pp0[5],pp0[6],pp0[7],s113[0],s113[1],s114[1],s115[1],s116[1],s117[1],s117[2],s117[3],s117[4],s117[5],s117[6],s116[8],s116[9],s102[0],s102[1],s102[2],s102[3],s120[10],s120[11],s120[12],s120[13],s120[14],s120[15],s120[16],s120[17],s120[18],s120[19],s120[20],s120[21],s120[22],s120[23],s120[24],s120[25],s120[26],s120[27],s120[28],s120[29],s120[30],s120[31],s120[32],s120[33],s120[34],s120[35],s120[36],s120[37],s120[38],s120[39],s120[40],s120[41],s120[42],s120[43],s120[44],s120[45],s120[46],s120[47],s120[48],s120[49],s120[50],s120[51],s120[52],s120[53],s120[54],s120[55],s120[56],s120[57],s120[58],s120[59],s120[60],s120[61],s120[62],s120[63],s120[64],s120[65],s120[66],s120[67],s120[68],s120[69],s120[70],s120[71],s120[72],s120[73],s120[74],s120[75],s120[76],s120[77],s120[78],s120[79],s120[80],s120[81],s120[82],s120[83],s120[84],s120[85],s120[86],s120[87],s120[88],s120[89],s120[90],s120[91],s120[92],s120[93],s120[94],s120[95],s120[96],s120[97],s120[98],s120[99],s120[100],s120[101],s120[102],s120[103],s120[104],s120[105],s120[106],s120[107],s120[108],s120[109],s120[110],s120[111],s120[112],s120[113],s120[114],s120[115],s120[116],s120[117],s120[118],s120[119],s120[120],s120[121],s120[122],s120[123],s120[124],s120[125],s120[126],s120[127],s120[128],s120[129],s120[130],s120[131],s120[132],s120[133],s120[134],s120[135],s120[136],s120[137],s120[138],s120[139],s120[140],s120[141],s120[142],s120[143],s120[144],s120[145],s120[146],s120[147],s120[148],s120[149],s120[150],s120[151],s120[152],s120[153],s120[154],s120[155],s120[156],s120[157],s120[158],s120[159],s120[160],s120[161],s120[162],s120[163],s120[164],s120[165],s120[166],s120[167],s120[168],s120[169],s120[170],s120[171],s120[172],s120[173],s120[174],s120[175],s120[176],s120[177],s120[178],s120[179],s120[180],s120[181],s120[182],s120[183],s120[184],s120[185],s120[186],s120[187],s120[188],s120[189],s120[190],s120[191],s120[192],s120[193],s120[194],s120[195],s120[196],s120[197],s120[198],s120[199],s120[200],s120[201],s120[202],s120[203],s120[204],s120[205],s120[206],s119[208],s118[210],s117[212],s117[213],s117[214],s117[215],s117[216],s117[217],s117[218],s117[219],s117[220],s117[221],s117[222],s117[223],s117[224],s117[225],s116[227],s115[229],s114[231],s113[233],pp127[115],pp126[117],pp125[119],pp124[121],pp123[123],pp122[125],pp121[127],pp122[127],pp123[127],pp124[127]};
    assign in121_2 = {pp1[3],pp1[4],pp1[5],pp1[6],pp2[6],s114[0],s115[0],s116[0],s117[0],s118[0],s118[1],s118[2],s118[3],s118[4],s118[5],s117[7],s117[8],s117[9],s103[0],s103[1],s103[2],s103[3],s103[4],s103[5],s103[6],s104[6],s105[6],s106[6],s107[6],s108[6],s109[6],s110[6],s111[6],s112[6],s65[6],s66[6],s67[6],s68[6],s69[6],s70[6],s71[6],s72[6],s73[6],s74[6],s75[6],s76[6],s77[6],s78[6],s79[6],s80[6],s81[6],s82[6],s83[6],s84[6],s85[6],s86[6],s87[6],s88[6],s89[6],s90[6],s91[6],s92[6],s93[6],s94[6],s95[6],s96[6],s1[6],s2[6],s3[6],s3[7],s3[8],s3[9],s13[0],s13[1],s13[2],s13[3],s13[4],s13[5],s13[6],s14[6],s15[6],s16[6],s17[6],s18[6],s19[6],s20[6],s21[6],s22[6],s23[6],s24[6],s25[6],s26[6],s27[6],s28[6],s29[6],s30[6],s31[6],s32[6],s33[6],s34[6],s35[6],s36[6],s37[6],s38[6],s39[6],s40[6],s41[6],s42[6],s43[6],s44[6],s45[6],s46[6],s47[6],s48[6],s49[6],s50[6],s51[6],s52[6],s53[6],s54[6],s55[6],s56[6],s57[6],s58[6],s59[6],s58[8],s9[58],s7[61],s5[64],s4[66],s4[67],s4[68],s4[69],s4[70],s4[71],s4[72],s4[73],s4[74],s4[75],s4[76],s4[77],s4[78],s4[79],s4[80],s4[81],s4[82],s4[83],s4[84],s4[85],s4[86],s4[87],s4[88],s4[89],s4[90],s4[91],s4[92],s4[93],s4[94],s4[95],s4[96],s4[97],s4[98],s4[99],s25[79],s23[82],s21[85],s19[88],s17[91],s15[94],s14[96],s13[98],s9[103],s7[106],s5[109],s4[111],s4[112],s4[113],s4[114],s4[115],s4[116],s3[118],s2[120],s1[122],s99[169],s98[171],s97[173],s96[127],s95[129],s94[131],s93[133],s92[135],s91[137],s90[139],s89[141],s88[143],s87[145],s86[147],s85[149],s84[151],s83[153],s82[155],s81[157],s80[159],s79[161],s78[163],s77[165],s76[167],s75[169],s74[171],s73[173],s72[175],s71[177],s70[179],s69[181],s68[183],s67[185],s66[187],s65[189],s120[207],s119[209],s118[211],s118[212],s118[213],s118[214],s118[215],s118[216],s118[217],s118[218],s118[219],s118[220],s118[221],s118[222],s118[223],s118[224],s117[226],s116[228],s115[230],s114[232],s113[234],pp127[116],pp126[118],pp125[120],pp124[122],pp123[124],pp122[126],pp123[126],pp124[126],pp125[126]};
    CLA_248 KS_121(s121, c121, in121_1, in121_2);
    wire[245:0] s122, in122_1, in122_2;
    wire c122;
    assign in122_1 = {pp2[3],s121[2],s121[3],s121[4],s121[5],s121[6],s121[7],s121[8],s121[9],s121[10],s121[11],s121[12],s121[13],s121[14],s121[15],s121[16],s121[17],s121[18],s121[19],s121[20],s121[21],s121[22],s121[23],s121[24],s121[25],s121[26],s121[27],s121[28],s121[29],s121[30],s121[31],s121[32],s121[33],s121[34],s121[35],s121[36],s121[37],s121[38],s121[39],s121[40],s121[41],s121[42],s121[43],s121[44],s121[45],s121[46],s121[47],s121[48],s121[49],s121[50],s121[51],s121[52],s121[53],s121[54],s121[55],s121[56],s121[57],s121[58],s121[59],s121[60],s121[61],s121[62],s121[63],s121[64],s121[65],s121[66],s121[67],s121[68],s121[69],s121[70],s121[71],s121[72],s121[73],s121[74],s121[75],s121[76],s121[77],s121[78],s121[79],s121[80],s121[81],s121[82],s121[83],s121[84],s121[85],s121[86],s121[87],s121[88],s121[89],s121[90],s121[91],s121[92],s121[93],s121[94],s121[95],s121[96],s121[97],s121[98],s121[99],s121[100],s121[101],s121[102],s121[103],s121[104],s121[105],s121[106],s121[107],s121[108],s121[109],s121[110],s121[111],s121[112],s121[113],s121[114],s121[115],s121[116],s121[117],s121[118],s121[119],s121[120],s121[121],s121[122],s121[123],s121[124],s121[125],s121[126],s121[127],s121[128],s121[129],s121[130],s121[131],s121[132],s121[133],s121[134],s121[135],s121[136],s121[137],s121[138],s121[139],s121[140],s121[141],s121[142],s121[143],s121[144],s121[145],s121[146],s121[147],s121[148],s121[149],s121[150],s121[151],s121[152],s121[153],s121[154],s121[155],s121[156],s121[157],s121[158],s121[159],s121[160],s121[161],s121[162],s121[163],s121[164],s121[165],s121[166],s121[167],s121[168],s121[169],s121[170],s121[171],s121[172],s121[173],s121[174],s121[175],s121[176],s121[177],s121[178],s121[179],s121[180],s121[181],s121[182],s121[183],s121[184],s121[185],s121[186],s121[187],s121[188],s121[189],s121[190],s121[191],s121[192],s121[193],s121[194],s121[195],s121[196],s121[197],s121[198],s121[199],s121[200],s121[201],s121[202],s121[203],s121[204],s121[205],s121[206],s121[207],s121[208],s121[209],s121[210],s121[211],s121[212],s121[213],s121[214],s121[215],s121[216],s121[217],s121[218],s120[208],s119[210],s119[211],s119[212],s119[213],s119[214],s119[215],s119[216],s119[217],s119[218],s119[219],s119[220],s119[221],s119[222],s119[223],s118[225],s117[227],s116[229],s115[231],s114[233],s113[235],pp127[117],pp126[119],pp125[121],pp124[123],pp123[125],pp124[125],pp125[125]};
    assign in122_2 = {pp3[2],pp2[4],pp2[5],pp3[5],pp4[5],pp4[6],pp4[7],pp4[8],pp4[9],s119[0],s119[1],s119[2],s119[3],s119[4],s118[6],s118[7],s118[8],s118[9],s104[0],s104[1],s104[2],s104[3],s104[4],s104[5],s105[5],s106[5],s107[5],s108[5],s109[5],s110[5],s111[5],s112[5],s65[5],s66[5],s67[5],s68[5],s69[5],s70[5],s71[5],s72[5],s73[5],s74[5],s75[5],s76[5],s77[5],s78[5],s79[5],s80[5],s81[5],s82[5],s83[5],s84[5],s85[5],s86[5],s87[5],s88[5],s89[5],s90[5],s91[5],s92[5],s93[5],s94[5],s95[5],s96[5],s1[5],s2[5],s3[5],s4[5],s4[6],s4[7],s4[8],s4[9],s14[0],s14[1],s14[2],s14[3],s14[4],s14[5],s15[5],s16[5],s17[5],s18[5],s19[5],s20[5],s21[5],s22[5],s23[5],s24[5],s25[5],s26[5],s27[5],s28[5],s29[5],s30[5],s31[5],s32[5],s33[5],s34[5],s35[5],s36[5],s37[5],s38[5],s39[5],s40[5],s41[5],s42[5],s43[5],s44[5],s45[5],s46[5],s47[5],s48[5],s49[5],s50[5],s51[5],s52[5],s53[5],s54[5],s55[5],s56[5],s57[5],s58[5],s59[5],s60[5],s59[7],s58[9],s8[60],s6[63],s5[65],s5[66],s5[67],s5[68],s5[69],s5[70],s5[71],s5[72],s5[73],s5[74],s5[75],s5[76],s5[77],s5[78],s5[79],s5[80],s5[81],s5[82],s5[83],s5[84],s5[85],s5[86],s5[87],s5[88],s5[89],s5[90],s5[91],s5[92],s5[93],s5[94],s5[95],s5[96],s5[97],s5[98],s5[99],s24[81],s22[84],s20[87],s18[90],s16[93],s15[95],s14[97],s13[99],s8[105],s6[108],s5[110],s5[111],s5[112],s5[113],s5[114],s5[115],s4[117],s3[119],s2[121],s1[123],s99[170],s98[172],s97[174],s96[128],s95[130],s94[132],s93[134],s92[136],s91[138],s90[140],s89[142],s88[144],s87[146],s86[148],s85[150],s84[152],s83[154],s82[156],s81[158],s80[160],s79[162],s78[164],s77[166],s76[168],s75[170],s74[172],s73[174],s72[176],s71[178],s70[180],s69[182],s68[184],s67[186],s66[188],s65[190],s121[219],s120[209],s120[210],s120[211],s120[212],s120[213],s120[214],s120[215],s120[216],s120[217],s120[218],s120[219],s120[220],s120[221],s120[222],s119[224],s118[226],s117[228],s116[230],s115[232],s114[234],s113[236],pp127[118],pp126[120],pp125[122],pp124[124],pp125[124],pp126[124]};
    CLA_246 KS_122(s122, c122, in122_1, in122_2);
    wire[243:0] s123, in123_1, in123_2;
    wire c123;
    assign in123_1 = {pp3[3],s122[2],s122[3],s122[4],s122[5],s122[6],s122[7],s122[8],s122[9],s122[10],s122[11],s122[12],s122[13],s122[14],s122[15],s122[16],s122[17],s122[18],s122[19],s122[20],s122[21],s122[22],s122[23],s122[24],s122[25],s122[26],s122[27],s122[28],s122[29],s122[30],s122[31],s122[32],s122[33],s122[34],s122[35],s122[36],s122[37],s122[38],s122[39],s122[40],s122[41],s122[42],s122[43],s122[44],s122[45],s122[46],s122[47],s122[48],s122[49],s122[50],s122[51],s122[52],s122[53],s122[54],s122[55],s122[56],s122[57],s122[58],s122[59],s122[60],s122[61],s122[62],s122[63],s122[64],s122[65],s122[66],s122[67],s122[68],s122[69],s122[70],s122[71],s122[72],s122[73],s122[74],s122[75],s122[76],s122[77],s122[78],s122[79],s122[80],s122[81],s122[82],s122[83],s122[84],s122[85],s122[86],s122[87],s122[88],s122[89],s122[90],s122[91],s122[92],s122[93],s122[94],s122[95],s122[96],s122[97],s122[98],s122[99],s122[100],s122[101],s122[102],s122[103],s122[104],s122[105],s122[106],s122[107],s122[108],s122[109],s122[110],s122[111],s122[112],s122[113],s122[114],s122[115],s122[116],s122[117],s122[118],s122[119],s122[120],s122[121],s122[122],s122[123],s122[124],s122[125],s122[126],s122[127],s122[128],s122[129],s122[130],s122[131],s122[132],s122[133],s122[134],s122[135],s122[136],s122[137],s122[138],s122[139],s122[140],s122[141],s122[142],s122[143],s122[144],s122[145],s122[146],s122[147],s122[148],s122[149],s122[150],s122[151],s122[152],s122[153],s122[154],s122[155],s122[156],s122[157],s122[158],s122[159],s122[160],s122[161],s122[162],s122[163],s122[164],s122[165],s122[166],s122[167],s122[168],s122[169],s122[170],s122[171],s122[172],s122[173],s122[174],s122[175],s122[176],s122[177],s122[178],s122[179],s122[180],s122[181],s122[182],s122[183],s122[184],s122[185],s122[186],s122[187],s122[188],s122[189],s122[190],s122[191],s122[192],s122[193],s122[194],s122[195],s122[196],s122[197],s122[198],s122[199],s122[200],s122[201],s122[202],s122[203],s122[204],s122[205],s122[206],s122[207],s122[208],s122[209],s122[210],s122[211],s122[212],s122[213],s122[214],s122[215],s122[216],s122[217],s122[218],s121[220],s121[221],s121[222],s121[223],s121[224],s121[225],s121[226],s121[227],s121[228],s121[229],s121[230],s121[231],s121[232],s121[233],s120[223],s119[225],s118[227],s117[229],s116[231],s115[233],s114[235],s113[237],pp127[119],pp126[121],pp125[123],pp126[123]};
    assign in123_2 = {pp4[2],pp3[4],pp4[4],pp5[4],pp5[5],pp5[6],pp5[7],pp5[8],pp5[9],s120[0],s120[1],s120[2],s120[3],s119[5],s119[6],s119[7],s119[8],s119[9],s105[0],s105[1],s105[2],s105[3],s105[4],s106[4],s107[4],s108[4],s109[4],s110[4],s111[4],s112[4],s65[4],s66[4],s67[4],s68[4],s69[4],s70[4],s71[4],s72[4],s73[4],s74[4],s75[4],s76[4],s77[4],s78[4],s79[4],s80[4],s81[4],s82[4],s83[4],s84[4],s85[4],s86[4],s87[4],s88[4],s89[4],s90[4],s91[4],s92[4],s93[4],s94[4],s95[4],s96[4],s1[4],s2[4],s3[4],s4[4],s5[4],s5[5],s5[6],s5[7],s5[8],s5[9],s15[0],s15[1],s15[2],s15[3],s15[4],s16[4],s17[4],s18[4],s19[4],s20[4],s21[4],s22[4],s23[4],s24[4],s25[4],s26[4],s27[4],s28[4],s29[4],s30[4],s31[4],s32[4],s33[4],s34[4],s35[4],s36[4],s37[4],s38[4],s39[4],s40[4],s41[4],s42[4],s43[4],s44[4],s45[4],s46[4],s47[4],s48[4],s49[4],s50[4],s51[4],s52[4],s53[4],s54[4],s55[4],s56[4],s57[4],s58[4],s59[4],s60[4],s61[4],s60[6],s59[8],s9[59],s7[62],s6[64],s6[65],s6[66],s6[67],s6[68],s6[69],s6[70],s6[71],s6[72],s6[73],s6[74],s6[75],s6[76],s6[77],s6[78],s6[79],s6[80],s6[81],s6[82],s6[83],s6[84],s6[85],s6[86],s6[87],s6[88],s6[89],s6[90],s6[91],s6[92],s6[93],s6[94],s6[95],s6[96],s6[97],s6[98],s6[99],s23[83],s21[86],s19[89],s17[92],s16[94],s15[96],s14[98],s9[104],s7[107],s6[109],s6[110],s6[111],s6[112],s6[113],s6[114],s5[116],s4[118],s3[120],s2[122],s1[124],s99[171],s98[173],s97[175],s96[129],s95[131],s94[133],s93[135],s92[137],s91[139],s90[141],s89[143],s88[145],s87[147],s86[149],s85[151],s84[153],s83[155],s82[157],s81[159],s80[161],s79[163],s78[165],s77[167],s76[169],s75[171],s74[173],s73[175],s72[177],s71[179],s70[181],s69[183],s68[185],s67[187],s66[189],s65[191],s122[219],s122[220],s122[221],s122[222],s122[223],s122[224],s122[225],s122[226],s122[227],s122[228],s122[229],s122[230],s122[231],s122[232],s121[234],s120[224],s119[226],s118[228],s117[230],s116[232],s115[234],s114[236],s113[238],pp127[120],pp126[122],pp127[122]};
    CLA_244 KS_123(s123, c123, in123_1, in123_2);
    wire[241:0] s124, in124_1, in124_2;
    wire c124;
    assign in124_1 = {pp4[3],s123[2],s123[3],s123[4],s123[5],s123[6],s123[7],s123[8],s123[9],s123[10],s123[11],s123[12],s123[13],s123[14],s123[15],s123[16],s123[17],s123[18],s123[19],s123[20],s123[21],s123[22],s123[23],s123[24],s123[25],s123[26],s123[27],s123[28],s123[29],s123[30],s123[31],s123[32],s123[33],s123[34],s123[35],s123[36],s123[37],s123[38],s123[39],s123[40],s123[41],s123[42],s123[43],s123[44],s123[45],s123[46],s123[47],s123[48],s123[49],s123[50],s123[51],s123[52],s123[53],s123[54],s123[55],s123[56],s123[57],s123[58],s123[59],s123[60],s123[61],s123[62],s123[63],s123[64],s123[65],s123[66],s123[67],s123[68],s123[69],s123[70],s123[71],s123[72],s123[73],s123[74],s123[75],s123[76],s123[77],s123[78],s123[79],s123[80],s123[81],s123[82],s123[83],s123[84],s123[85],s123[86],s123[87],s123[88],s123[89],s123[90],s123[91],s123[92],s123[93],s123[94],s123[95],s123[96],s123[97],s123[98],s123[99],s123[100],s123[101],s123[102],s123[103],s123[104],s123[105],s123[106],s123[107],s123[108],s123[109],s123[110],s123[111],s123[112],s123[113],s123[114],s123[115],s123[116],s123[117],s123[118],s123[119],s123[120],s123[121],s123[122],s123[123],s123[124],s123[125],s123[126],s123[127],s123[128],s123[129],s123[130],s123[131],s123[132],s123[133],s123[134],s123[135],s123[136],s123[137],s123[138],s123[139],s123[140],s123[141],s123[142],s123[143],s123[144],s123[145],s123[146],s123[147],s123[148],s123[149],s123[150],s123[151],s123[152],s123[153],s123[154],s123[155],s123[156],s123[157],s123[158],s123[159],s123[160],s123[161],s123[162],s123[163],s123[164],s123[165],s123[166],s123[167],s123[168],s123[169],s123[170],s123[171],s123[172],s123[173],s123[174],s123[175],s123[176],s123[177],s123[178],s123[179],s123[180],s123[181],s123[182],s123[183],s123[184],s123[185],s123[186],s123[187],s123[188],s123[189],s123[190],s123[191],s123[192],s123[193],s123[194],s123[195],s123[196],s123[197],s123[198],s123[199],s123[200],s123[201],s123[202],s123[203],s123[204],s123[205],s123[206],s123[207],s123[208],s123[209],s123[210],s123[211],s123[212],s123[213],s123[214],s123[215],s123[216],s123[217],s123[218],s123[219],s123[220],s123[221],s123[222],s123[223],s123[224],s123[225],s123[226],s123[227],s123[228],s123[229],s123[230],s123[231],s122[233],s121[235],s120[225],s119[227],s118[229],s117[231],s116[233],s115[235],s114[237],s113[239],pp127[121]};
    assign in124_2 = {pp5[2],pp5[3],pp6[3],pp6[4],pp6[5],pp6[6],pp6[7],pp6[8],pp6[9],pp7[9],pp8[9],pp9[9],s120[4],s120[5],s120[6],s120[7],s120[8],s120[9],s106[0],s106[1],s106[2],s106[3],s107[3],s108[3],s109[3],s110[3],s111[3],s112[3],s65[3],s66[3],s67[3],s68[3],s69[3],s70[3],s71[3],s72[3],s73[3],s74[3],s75[3],s76[3],s77[3],s78[3],s79[3],s80[3],s81[3],s82[3],s83[3],s84[3],s85[3],s86[3],s87[3],s88[3],s89[3],s90[3],s91[3],s92[3],s93[3],s94[3],s95[3],s96[3],s1[3],s2[3],s3[3],s4[3],s5[3],s6[3],s6[4],s6[5],s6[6],s6[7],s6[8],s6[9],s16[0],s16[1],s16[2],s16[3],s17[3],s18[3],s19[3],s20[3],s21[3],s22[3],s23[3],s24[3],s25[3],s26[3],s27[3],s28[3],s29[3],s30[3],s31[3],s32[3],s33[3],s34[3],s35[3],s36[3],s37[3],s38[3],s39[3],s40[3],s41[3],s42[3],s43[3],s44[3],s45[3],s46[3],s47[3],s48[3],s49[3],s50[3],s51[3],s52[3],s53[3],s54[3],s55[3],s56[3],s57[3],s58[3],s59[3],s60[3],s61[3],s62[3],s61[5],s60[7],s59[9],s8[61],s7[63],s7[64],s7[65],s7[66],s7[67],s7[68],s7[69],s7[70],s7[71],s7[72],s7[73],s7[74],s7[75],s7[76],s7[77],s7[78],s7[79],s7[80],s7[81],s7[82],s7[83],s7[84],s7[85],s7[86],s7[87],s7[88],s7[89],s7[90],s7[91],s7[92],s7[93],s7[94],s7[95],s7[96],s7[97],s7[98],s7[99],s22[85],s20[88],s18[91],s17[93],s16[95],s15[97],s14[99],s8[106],s7[108],s7[109],s7[110],s7[111],s7[112],s7[113],s6[115],s5[117],s4[119],s3[121],s2[123],s1[125],s99[172],s98[174],s97[176],s97[177],s97[178],s97[179],s97[180],s97[181],s97[182],s97[183],s97[184],s97[185],s97[186],s97[187],s97[188],s97[189],s97[190],s97[191],s97[192],s97[193],s97[194],s97[195],s97[196],s97[197],s97[198],s97[199],s97[200],s97[201],s97[202],s97[203],s97[204],s97[205],s97[206],s97[207],s97[208],s97[209],s97[210],s97[211],s97[212],s97[213],s97[214],s97[215],s97[216],s97[217],s97[218],s97[219],s97[220],s97[221],s123[232],s122[234],s121[236],s121[237],s121[238],s121[239],s121[240],s121[241],s121[242],s121[243],s121[244]};
    CLA_242 KS_124(s124, c124, in124_1, in124_2);

    /*Stage 6*/
    wire[251:0] s125, in125_1, in125_2;
    wire c125;
    assign in125_1 = {pp0[2],pp0[3],s121[0],s121[1],s122[1],s123[1],s124[1],s124[2],s124[3],s124[4],s124[5],s124[6],s124[7],s124[8],s124[9],s124[10],s124[11],s124[12],s124[13],s124[14],s124[15],s124[16],s124[17],s124[18],s124[19],s124[20],s124[21],s124[22],s124[23],s124[24],s124[25],s124[26],s124[27],s124[28],s124[29],s124[30],s124[31],s124[32],s124[33],s124[34],s124[35],s124[36],s124[37],s124[38],s124[39],s124[40],s124[41],s124[42],s124[43],s124[44],s124[45],s124[46],s124[47],s124[48],s124[49],s124[50],s124[51],s124[52],s124[53],s124[54],s124[55],s124[56],s124[57],s124[58],s124[59],s124[60],s124[61],s124[62],s124[63],s124[64],s124[65],s124[66],s124[67],s124[68],s124[69],s124[70],s124[71],s124[72],s124[73],s124[74],s124[75],s124[76],s124[77],s124[78],s124[79],s124[80],s124[81],s124[82],s124[83],s124[84],s124[85],s124[86],s124[87],s124[88],s124[89],s124[90],s124[91],s124[92],s124[93],s124[94],s124[95],s124[96],s124[97],s124[98],s124[99],s124[100],s124[101],s124[102],s124[103],s124[104],s124[105],s124[106],s124[107],s124[108],s124[109],s124[110],s124[111],s124[112],s124[113],s124[114],s124[115],s124[116],s124[117],s124[118],s124[119],s124[120],s124[121],s124[122],s124[123],s124[124],s124[125],s124[126],s124[127],s124[128],s124[129],s124[130],s124[131],s124[132],s124[133],s124[134],s124[135],s124[136],s124[137],s124[138],s124[139],s124[140],s124[141],s124[142],s124[143],s124[144],s124[145],s124[146],s124[147],s124[148],s124[149],s124[150],s124[151],s124[152],s124[153],s124[154],s124[155],s124[156],s124[157],s124[158],s124[159],s124[160],s124[161],s124[162],s124[163],s124[164],s124[165],s124[166],s124[167],s124[168],s124[169],s124[170],s124[171],s124[172],s124[173],s124[174],s124[175],s124[176],s124[177],s124[178],s124[179],s124[180],s124[181],s124[182],s124[183],s124[184],s124[185],s124[186],s124[187],s124[188],s124[189],s124[190],s124[191],s124[192],s124[193],s124[194],s124[195],s124[196],s124[197],s124[198],s124[199],s124[200],s124[201],s124[202],s124[203],s124[204],s124[205],s124[206],s124[207],s124[208],s124[209],s124[210],s124[211],s124[212],s124[213],s124[214],s124[215],s124[216],s124[217],s124[218],s124[219],s124[220],s124[221],s124[222],s124[223],s124[224],s124[225],s124[226],s124[227],s124[228],s124[229],s124[230],s124[231],s123[233],s122[235],s122[236],s122[237],s122[238],s122[239],s122[240],s122[241],s122[242],s122[243],s121[245],pp127[123],pp126[125],pp125[127],pp126[127]};
    assign in125_2 = {pp1[1],pp1[2],pp2[2],s122[0],s123[0],s124[0],pp6[2],pp7[2],pp7[3],pp7[4],pp7[5],pp7[6],pp7[7],pp7[8],pp8[8],pp9[8],s97[2],s97[3],s97[4],s97[5],s97[6],s97[7],s97[8],s97[9],s107[0],s107[1],s107[2],s108[2],s109[2],s110[2],s111[2],s112[2],s65[2],s66[2],s67[2],s68[2],s69[2],s70[2],s71[2],s72[2],s73[2],s74[2],s75[2],s76[2],s77[2],s78[2],s79[2],s80[2],s81[2],s82[2],s83[2],s84[2],s85[2],s86[2],s87[2],s88[2],s89[2],s90[2],s91[2],s92[2],s93[2],s94[2],s95[2],s96[2],s1[2],s2[2],s3[2],s4[2],s5[2],s6[2],s7[2],s7[3],s7[4],s7[5],s7[6],s7[7],s7[8],s7[9],s17[0],s17[1],s17[2],s18[2],s19[2],s20[2],s21[2],s22[2],s23[2],s24[2],s25[2],s26[2],s27[2],s28[2],s29[2],s30[2],s31[2],s32[2],s33[2],s34[2],s35[2],s36[2],s37[2],s38[2],s39[2],s40[2],s41[2],s42[2],s43[2],s44[2],s45[2],s46[2],s47[2],s48[2],s49[2],s50[2],s51[2],s52[2],s53[2],s54[2],s55[2],s56[2],s57[2],s58[2],s59[2],s60[2],s61[2],s62[2],s63[2],s62[4],s61[6],s60[8],s9[60],s8[62],s8[63],s8[64],s8[65],s8[66],s8[67],s8[68],s8[69],s8[70],s8[71],s8[72],s8[73],s8[74],s8[75],s8[76],s8[77],s8[78],s8[79],s8[80],s8[81],s8[82],s8[83],s8[84],s8[85],s8[86],s8[87],s8[88],s8[89],s8[90],s8[91],s8[92],s8[93],s8[94],s8[95],s8[96],s8[97],s8[98],s8[99],s21[87],s19[90],s18[92],s17[94],s16[96],s15[98],s9[105],s8[107],s8[108],s8[109],s8[110],s8[111],s8[112],s7[114],s6[116],s5[118],s4[120],s3[122],s2[124],s1[126],s99[173],s98[175],s98[176],s98[177],s98[178],s98[179],s98[180],s98[181],s98[182],s98[183],s98[184],s98[185],s98[186],s98[187],s98[188],s98[189],s98[190],s98[191],s98[192],s98[193],s98[194],s98[195],s98[196],s98[197],s98[198],s98[199],s98[200],s98[201],s98[202],s98[203],s98[204],s98[205],s98[206],s98[207],s98[208],s98[209],s98[210],s98[211],s98[212],s98[213],s98[214],s98[215],s98[216],s98[217],s98[218],s98[219],s98[220],s97[222],s124[232],s123[234],s123[235],s123[236],s123[237],s123[238],s123[239],s123[240],s123[241],s123[242],s122[244],s121[246],pp127[124],pp126[126],pp127[126]};
    CLA_252 KS_125(s125, c125, in125_1, in125_2);
    wire[249:0] s126, in126_1, in126_2;
    wire c126;
    assign in126_1 = {pp2[1],s125[2],s125[3],s125[4],s125[5],s125[6],s125[7],s125[8],s125[9],s125[10],s125[11],s125[12],s125[13],s125[14],s125[15],s125[16],s125[17],s125[18],s125[19],s125[20],s125[21],s125[22],s125[23],s125[24],s125[25],s125[26],s125[27],s125[28],s125[29],s125[30],s125[31],s125[32],s125[33],s125[34],s125[35],s125[36],s125[37],s125[38],s125[39],s125[40],s125[41],s125[42],s125[43],s125[44],s125[45],s125[46],s125[47],s125[48],s125[49],s125[50],s125[51],s125[52],s125[53],s125[54],s125[55],s125[56],s125[57],s125[58],s125[59],s125[60],s125[61],s125[62],s125[63],s125[64],s125[65],s125[66],s125[67],s125[68],s125[69],s125[70],s125[71],s125[72],s125[73],s125[74],s125[75],s125[76],s125[77],s125[78],s125[79],s125[80],s125[81],s125[82],s125[83],s125[84],s125[85],s125[86],s125[87],s125[88],s125[89],s125[90],s125[91],s125[92],s125[93],s125[94],s125[95],s125[96],s125[97],s125[98],s125[99],s125[100],s125[101],s125[102],s125[103],s125[104],s125[105],s125[106],s125[107],s125[108],s125[109],s125[110],s125[111],s125[112],s125[113],s125[114],s125[115],s125[116],s125[117],s125[118],s125[119],s125[120],s125[121],s125[122],s125[123],s125[124],s125[125],s125[126],s125[127],s125[128],s125[129],s125[130],s125[131],s125[132],s125[133],s125[134],s125[135],s125[136],s125[137],s125[138],s125[139],s125[140],s125[141],s125[142],s125[143],s125[144],s125[145],s125[146],s125[147],s125[148],s125[149],s125[150],s125[151],s125[152],s125[153],s125[154],s125[155],s125[156],s125[157],s125[158],s125[159],s125[160],s125[161],s125[162],s125[163],s125[164],s125[165],s125[166],s125[167],s125[168],s125[169],s125[170],s125[171],s125[172],s125[173],s125[174],s125[175],s125[176],s125[177],s125[178],s125[179],s125[180],s125[181],s125[182],s125[183],s125[184],s125[185],s125[186],s125[187],s125[188],s125[189],s125[190],s125[191],s125[192],s125[193],s125[194],s125[195],s125[196],s125[197],s125[198],s125[199],s125[200],s125[201],s125[202],s125[203],s125[204],s125[205],s125[206],s125[207],s125[208],s125[209],s125[210],s125[211],s125[212],s125[213],s125[214],s125[215],s125[216],s125[217],s125[218],s125[219],s125[220],s125[221],s125[222],s125[223],s125[224],s125[225],s125[226],s125[227],s125[228],s125[229],s125[230],s125[231],s125[232],s125[233],s125[234],s125[235],s125[236],s125[237],s124[233],s124[234],s124[235],s124[236],s124[237],s124[238],s124[239],s124[240],s124[241],s123[243],s122[245],s121[247],pp127[125]};
    assign in126_2 = {pp3[0],pp3[1],pp4[1],pp5[1],pp6[1],pp7[1],pp8[1],pp8[2],pp8[3],pp8[4],pp8[5],pp8[6],pp8[7],pp9[7],s97[1],s98[1],s98[2],s98[3],s98[4],s98[5],s98[6],s98[7],s98[8],s98[9],s108[0],s108[1],s109[1],s110[1],s111[1],s112[1],s65[1],s66[1],s67[1],s68[1],s69[1],s70[1],s71[1],s72[1],s73[1],s74[1],s75[1],s76[1],s77[1],s78[1],s79[1],s80[1],s81[1],s82[1],s83[1],s84[1],s85[1],s86[1],s87[1],s88[1],s89[1],s90[1],s91[1],s92[1],s93[1],s94[1],s95[1],s96[1],s1[1],s2[1],s3[1],s4[1],s5[1],s6[1],s7[1],s8[1],s8[2],s8[3],s8[4],s8[5],s8[6],s8[7],s8[8],s8[9],s18[0],s18[1],s19[1],s20[1],s21[1],s22[1],s23[1],s24[1],s25[1],s26[1],s27[1],s28[1],s29[1],s30[1],s31[1],s32[1],s33[1],s34[1],s35[1],s36[1],s37[1],s38[1],s39[1],s40[1],s41[1],s42[1],s43[1],s44[1],s45[1],s46[1],s47[1],s48[1],s49[1],s50[1],s51[1],s52[1],s53[1],s54[1],s55[1],s56[1],s57[1],s58[1],s59[1],s60[1],s61[1],s62[1],s63[1],s64[1],s63[3],s62[5],s61[7],s60[9],s9[61],s9[62],s9[63],s9[64],s9[65],s9[66],s9[67],s9[68],s9[69],s9[70],s9[71],s9[72],s9[73],s9[74],s9[75],s9[76],s9[77],s9[78],s9[79],s9[80],s9[81],s9[82],s9[83],s9[84],s9[85],s9[86],s9[87],s9[88],s9[89],s9[90],s9[91],s9[92],s9[93],s9[94],s9[95],s9[96],s9[97],s9[98],s9[99],s20[89],s19[91],s18[93],s17[95],s16[97],s15[99],s9[106],s9[107],s9[108],s9[109],s9[110],s9[111],s8[113],s7[115],s6[117],s5[119],s4[121],s3[123],s2[125],s1[127],s99[174],s99[175],s99[176],s99[177],s99[178],s99[179],s99[180],s99[181],s99[182],s99[183],s99[184],s99[185],s99[186],s99[187],s99[188],s99[189],s99[190],s99[191],s99[192],s99[193],s99[194],s99[195],s99[196],s99[197],s99[198],s99[199],s99[200],s99[201],s99[202],s99[203],s99[204],s99[205],s99[206],s99[207],s99[208],s99[209],s99[210],s99[211],s99[212],s99[213],s99[214],s99[215],s99[216],s99[217],s99[218],s99[219],s98[221],s97[223],s125[238],s125[239],s125[240],s125[241],s125[242],s125[243],s125[244],s125[245],s125[246],s125[247],s125[248],s125[249],s125[250]};
    CLA_250 KS_126(s126, c126, in126_1, in126_2);


    /*Final Stage 6*/
    wire[253:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],s125[0],s125[1],pp4[0],pp5[0],pp6[0],pp7[0],pp8[0],pp9[0],pp9[1],pp9[2],pp9[3],pp9[4],pp9[5],pp9[6],s97[0],s98[0],s99[0],s99[1],s99[2],s99[3],s99[4],s99[5],s99[6],s99[7],s99[8],s99[9],s109[0],s110[0],s111[0],s112[0],s65[0],s66[0],s67[0],s68[0],s69[0],s70[0],s71[0],s72[0],s73[0],s74[0],s75[0],s76[0],s77[0],s78[0],s79[0],s80[0],s81[0],s82[0],s83[0],s84[0],s85[0],s86[0],s87[0],s88[0],s89[0],s90[0],s91[0],s92[0],s93[0],s94[0],s95[0],s96[0],s1[0],s2[0],s3[0],s4[0],s5[0],s6[0],s7[0],s8[0],s9[0],s9[1],s9[2],s9[3],s9[4],s9[5],s9[6],s9[7],s9[8],s9[9],s19[0],s20[0],s21[0],s22[0],s23[0],s24[0],s25[0],s26[0],s27[0],s28[0],s29[0],s30[0],s31[0],s32[0],s33[0],s34[0],s35[0],s36[0],s37[0],s38[0],s39[0],s40[0],s41[0],s42[0],s43[0],s44[0],s45[0],s46[0],s47[0],s48[0],s49[0],s50[0],s51[0],s52[0],s53[0],s54[0],s55[0],s56[0],s57[0],s58[0],s59[0],s60[0],s61[0],s62[0],s63[0],s64[0],p1'b0,c64,c63,c62,c61,c60,c59,c58,c57,c56,c55,c54,c53,c52,c51,c50,c49,c48,c47,c46,c45,c44,c43,c42,c41,c40,c39,c38,c37,c36,c35,c34,c33,c32,c31,c30,c29,c28,c27,c26,c25,c24,c23,c22,c21,c20,c19,c18,c17,c16,c15,c14,c13,c12,c11,c10,c9,c8,c7,c6,c5,c4,c3,c2,c1,c96,c95,c94,c93,c92,c91,c90,c89,c88,c87,c86,c85,c84,c83,c82,c81,c80,c79,c78,c77,c76,c75,c74,c73,c72,c71,c70,c69,c68,c67,c66,c65,c112,c111,c110,c109,c108,c107,c106,c105,c104,c103,c102,c101,c100,c99,c98,c97,c120,c119,c118,c117,c116,c115,c114,c113,c124,c123,c122,c121,s125[251],pp127[127]};
    assign in_2 = {pp1[0],pp2[0],s126[0],s126[1],s126[2],s126[3],s126[4],s126[5],s126[6],s126[7],s126[8],s126[9],s126[10],s126[11],s126[12],s126[13],s126[14],s126[15],s126[16],s126[17],s126[18],s126[19],s126[20],s126[21],s126[22],s126[23],s126[24],s126[25],s126[26],s126[27],s126[28],s126[29],s126[30],s126[31],s126[32],s126[33],s126[34],s126[35],s126[36],s126[37],s126[38],s126[39],s126[40],s126[41],s126[42],s126[43],s126[44],s126[45],s126[46],s126[47],s126[48],s126[49],s126[50],s126[51],s126[52],s126[53],s126[54],s126[55],s126[56],s126[57],s126[58],s126[59],s126[60],s126[61],s126[62],s126[63],s126[64],s126[65],s126[66],s126[67],s126[68],s126[69],s126[70],s126[71],s126[72],s126[73],s126[74],s126[75],s126[76],s126[77],s126[78],s126[79],s126[80],s126[81],s126[82],s126[83],s126[84],s126[85],s126[86],s126[87],s126[88],s126[89],s126[90],s126[91],s126[92],s126[93],s126[94],s126[95],s126[96],s126[97],s126[98],s126[99],s126[100],s126[101],s126[102],s126[103],s126[104],s126[105],s126[106],s126[107],s126[108],s126[109],s126[110],s126[111],s126[112],s126[113],s126[114],s126[115],s126[116],s126[117],s126[118],s126[119],s126[120],s126[121],s126[122],s126[123],s126[124],s126[125],s126[126],s126[127],s126[128],s126[129],s126[130],s126[131],s126[132],s126[133],s126[134],s126[135],s126[136],s126[137],s126[138],s126[139],s126[140],s126[141],s126[142],s126[143],s126[144],s126[145],s126[146],s126[147],s126[148],s126[149],s126[150],s126[151],s126[152],s126[153],s126[154],s126[155],s126[156],s126[157],s126[158],s126[159],s126[160],s126[161],s126[162],s126[163],s126[164],s126[165],s126[166],s126[167],s126[168],s126[169],s126[170],s126[171],s126[172],s126[173],s126[174],s126[175],s126[176],s126[177],s126[178],s126[179],s126[180],s126[181],s126[182],s126[183],s126[184],s126[185],s126[186],s126[187],s126[188],s126[189],s126[190],s126[191],s126[192],s126[193],s126[194],s126[195],s126[196],s126[197],s126[198],s126[199],s126[200],s126[201],s126[202],s126[203],s126[204],s126[205],s126[206],s126[207],s126[208],s126[209],s126[210],s126[211],s126[212],s126[213],s126[214],s126[215],s126[216],s126[217],s126[218],s126[219],s126[220],s126[221],s126[222],s126[223],s126[224],s126[225],s126[226],s126[227],s126[228],s126[229],s126[230],s126[231],s126[232],s126[233],s126[234],s126[235],s126[236],s126[237],s126[238],s126[239],s126[240],s126[241],s126[242],s126[243],s126[244],s126[245],s126[246],s126[247],s126[248],s126[249],c126,c125};
    CLA_254(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = s[126];
    assign product[128] = s[127];
    assign product[129] = s[128];
    assign product[130] = s[129];
    assign product[131] = s[130];
    assign product[132] = s[131];
    assign product[133] = s[132];
    assign product[134] = s[133];
    assign product[135] = s[134];
    assign product[136] = s[135];
    assign product[137] = s[136];
    assign product[138] = s[137];
    assign product[139] = s[138];
    assign product[140] = s[139];
    assign product[141] = s[140];
    assign product[142] = s[141];
    assign product[143] = s[142];
    assign product[144] = s[143];
    assign product[145] = s[144];
    assign product[146] = s[145];
    assign product[147] = s[146];
    assign product[148] = s[147];
    assign product[149] = s[148];
    assign product[150] = s[149];
    assign product[151] = s[150];
    assign product[152] = s[151];
    assign product[153] = s[152];
    assign product[154] = s[153];
    assign product[155] = s[154];
    assign product[156] = s[155];
    assign product[157] = s[156];
    assign product[158] = s[157];
    assign product[159] = s[158];
    assign product[160] = s[159];
    assign product[161] = s[160];
    assign product[162] = s[161];
    assign product[163] = s[162];
    assign product[164] = s[163];
    assign product[165] = s[164];
    assign product[166] = s[165];
    assign product[167] = s[166];
    assign product[168] = s[167];
    assign product[169] = s[168];
    assign product[170] = s[169];
    assign product[171] = s[170];
    assign product[172] = s[171];
    assign product[173] = s[172];
    assign product[174] = s[173];
    assign product[175] = s[174];
    assign product[176] = s[175];
    assign product[177] = s[176];
    assign product[178] = s[177];
    assign product[179] = s[178];
    assign product[180] = s[179];
    assign product[181] = s[180];
    assign product[182] = s[181];
    assign product[183] = s[182];
    assign product[184] = s[183];
    assign product[185] = s[184];
    assign product[186] = s[185];
    assign product[187] = s[186];
    assign product[188] = s[187];
    assign product[189] = s[188];
    assign product[190] = s[189];
    assign product[191] = s[190];
    assign product[192] = s[191];
    assign product[193] = s[192];
    assign product[194] = s[193];
    assign product[195] = s[194];
    assign product[196] = s[195];
    assign product[197] = s[196];
    assign product[198] = s[197];
    assign product[199] = s[198];
    assign product[200] = s[199];
    assign product[201] = s[200];
    assign product[202] = s[201];
    assign product[203] = s[202];
    assign product[204] = s[203];
    assign product[205] = s[204];
    assign product[206] = s[205];
    assign product[207] = s[206];
    assign product[208] = s[207];
    assign product[209] = s[208];
    assign product[210] = s[209];
    assign product[211] = s[210];
    assign product[212] = s[211];
    assign product[213] = s[212];
    assign product[214] = s[213];
    assign product[215] = s[214];
    assign product[216] = s[215];
    assign product[217] = s[216];
    assign product[218] = s[217];
    assign product[219] = s[218];
    assign product[220] = s[219];
    assign product[221] = s[220];
    assign product[222] = s[221];
    assign product[223] = s[222];
    assign product[224] = s[223];
    assign product[225] = s[224];
    assign product[226] = s[225];
    assign product[227] = s[226];
    assign product[228] = s[227];
    assign product[229] = s[228];
    assign product[230] = s[229];
    assign product[231] = s[230];
    assign product[232] = s[231];
    assign product[233] = s[232];
    assign product[234] = s[233];
    assign product[235] = s[234];
    assign product[236] = s[235];
    assign product[237] = s[236];
    assign product[238] = s[237];
    assign product[239] = s[238];
    assign product[240] = s[239];
    assign product[241] = s[240];
    assign product[242] = s[241];
    assign product[243] = s[242];
    assign product[244] = s[243];
    assign product[245] = s[244];
    assign product[246] = s[245];
    assign product[247] = s[246];
    assign product[248] = s[247];
    assign product[249] = s[248];
    assign product[250] = s[249];
    assign product[251] = s[250];
    assign product[252] = s[251];
    assign product[253] = s[252];
    assign product[254] = s[253];
    assign product[255] = c;
endmodule

