module multiplier_64bits_version11(product, A, B);

    output [127:0] product;
    input [63:0] A, B;

    wire [63:0] pp0;
    wire [63:0] pp1;
    wire [63:0] pp2;
    wire [63:0] pp3;
    wire [63:0] pp4;
    wire [63:0] pp5;
    wire [63:0] pp6;
    wire [63:0] pp7;
    wire [63:0] pp8;
    wire [63:0] pp9;
    wire [63:0] pp10;
    wire [63:0] pp11;
    wire [63:0] pp12;
    wire [63:0] pp13;
    wire [63:0] pp14;
    wire [63:0] pp15;
    wire [63:0] pp16;
    wire [63:0] pp17;
    wire [63:0] pp18;
    wire [63:0] pp19;
    wire [63:0] pp20;
    wire [63:0] pp21;
    wire [63:0] pp22;
    wire [63:0] pp23;
    wire [63:0] pp24;
    wire [63:0] pp25;
    wire [63:0] pp26;
    wire [63:0] pp27;
    wire [63:0] pp28;
    wire [63:0] pp29;
    wire [63:0] pp30;
    wire [63:0] pp31;
    wire [63:0] pp32;
    wire [63:0] pp33;
    wire [63:0] pp34;
    wire [63:0] pp35;
    wire [63:0] pp36;
    wire [63:0] pp37;
    wire [63:0] pp38;
    wire [63:0] pp39;
    wire [63:0] pp40;
    wire [63:0] pp41;
    wire [63:0] pp42;
    wire [63:0] pp43;
    wire [63:0] pp44;
    wire [63:0] pp45;
    wire [63:0] pp46;
    wire [63:0] pp47;
    wire [63:0] pp48;
    wire [63:0] pp49;
    wire [63:0] pp50;
    wire [63:0] pp51;
    wire [63:0] pp52;
    wire [63:0] pp53;
    wire [63:0] pp54;
    wire [63:0] pp55;
    wire [63:0] pp56;
    wire [63:0] pp57;
    wire [63:0] pp58;
    wire [63:0] pp59;
    wire [63:0] pp60;
    wire [63:0] pp61;
    wire [63:0] pp62;
    wire [63:0] pp63;


    assign pp0 = A[0] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[63:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[32],pp0[33],pp0[34],pp0[35],pp0[36],pp0[37],pp0[38],pp0[39],pp0[40],pp0[41],pp0[42],pp0[43],pp0[44],pp0[45],pp0[46],pp0[47],pp0[48],pp0[49],pp0[50],pp0[51],pp0[52],pp0[53],pp0[54],pp0[55],pp0[56],pp0[57],pp0[58],pp0[59],pp0[60],pp0[61],pp0[62],pp0[63],pp1[63],pp2[63],pp3[63],pp4[63],pp5[63],pp6[63],pp7[63],pp8[63],pp9[63],pp10[63],pp11[63],pp12[63],pp13[63],pp14[63],pp15[63],pp16[63],pp17[63],pp18[63],pp19[63],pp20[63],pp21[63],pp22[63],pp23[63],pp24[63],pp25[63],pp26[63],pp27[63],pp28[63],pp29[63],pp30[63],pp31[63],pp32[63]};
    assign in1_2 = {pp1[31],pp1[32],pp1[33],pp1[34],pp1[35],pp1[36],pp1[37],pp1[38],pp1[39],pp1[40],pp1[41],pp1[42],pp1[43],pp1[44],pp1[45],pp1[46],pp1[47],pp1[48],pp1[49],pp1[50],pp1[51],pp1[52],pp1[53],pp1[54],pp1[55],pp1[56],pp1[57],pp1[58],pp1[59],pp1[60],pp1[61],pp1[62],pp2[62],pp3[62],pp4[62],pp5[62],pp6[62],pp7[62],pp8[62],pp9[62],pp10[62],pp11[62],pp12[62],pp13[62],pp14[62],pp15[62],pp16[62],pp17[62],pp18[62],pp19[62],pp20[62],pp21[62],pp22[62],pp23[62],pp24[62],pp25[62],pp26[62],pp27[62],pp28[62],pp29[62],pp30[62],pp31[62],pp32[62],pp33[62]};
    CLA_64 KS_1(s1, c1, in1_1, in1_2);
    wire[61:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp2[31],pp2[32],pp2[33],pp2[34],pp2[35],pp2[36],pp2[37],pp2[38],pp2[39],pp2[40],pp2[41],pp2[42],pp2[43],pp2[44],pp2[45],pp2[46],pp2[47],pp2[48],pp2[49],pp2[50],pp2[51],pp2[52],pp2[53],pp2[54],pp2[55],pp2[56],pp2[57],pp2[58],pp2[59],pp2[60],pp2[61],pp3[61],pp4[61],pp5[61],pp6[61],pp7[61],pp8[61],pp9[61],pp10[61],pp11[61],pp12[61],pp13[61],pp14[61],pp15[61],pp16[61],pp17[61],pp18[61],pp19[61],pp20[61],pp21[61],pp22[61],pp23[61],pp24[61],pp25[61],pp26[61],pp27[61],pp28[61],pp29[61],pp30[61],pp31[61],pp32[61],pp33[61]};
    assign in2_2 = {pp3[30],pp3[31],pp3[32],pp3[33],pp3[34],pp3[35],pp3[36],pp3[37],pp3[38],pp3[39],pp3[40],pp3[41],pp3[42],pp3[43],pp3[44],pp3[45],pp3[46],pp3[47],pp3[48],pp3[49],pp3[50],pp3[51],pp3[52],pp3[53],pp3[54],pp3[55],pp3[56],pp3[57],pp3[58],pp3[59],pp3[60],pp4[60],pp5[60],pp6[60],pp7[60],pp8[60],pp9[60],pp10[60],pp11[60],pp12[60],pp13[60],pp14[60],pp15[60],pp16[60],pp17[60],pp18[60],pp19[60],pp20[60],pp21[60],pp22[60],pp23[60],pp24[60],pp25[60],pp26[60],pp27[60],pp28[60],pp29[60],pp30[60],pp31[60],pp32[60],pp33[60],pp34[60]};
    CLA_62 KS_2(s2, c2, in2_1, in2_2);
    wire[59:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp4[30],pp4[31],pp4[32],pp4[33],pp4[34],pp4[35],pp4[36],pp4[37],pp4[38],pp4[39],pp4[40],pp4[41],pp4[42],pp4[43],pp4[44],pp4[45],pp4[46],pp4[47],pp4[48],pp4[49],pp4[50],pp4[51],pp4[52],pp4[53],pp4[54],pp4[55],pp4[56],pp4[57],pp4[58],pp4[59],pp5[59],pp6[59],pp7[59],pp8[59],pp9[59],pp10[59],pp11[59],pp12[59],pp13[59],pp14[59],pp15[59],pp16[59],pp17[59],pp18[59],pp19[59],pp20[59],pp21[59],pp22[59],pp23[59],pp24[59],pp25[59],pp26[59],pp27[59],pp28[59],pp29[59],pp30[59],pp31[59],pp32[59],pp33[59],pp34[59]};
    assign in3_2 = {pp5[29],pp5[30],pp5[31],pp5[32],pp5[33],pp5[34],pp5[35],pp5[36],pp5[37],pp5[38],pp5[39],pp5[40],pp5[41],pp5[42],pp5[43],pp5[44],pp5[45],pp5[46],pp5[47],pp5[48],pp5[49],pp5[50],pp5[51],pp5[52],pp5[53],pp5[54],pp5[55],pp5[56],pp5[57],pp5[58],pp6[58],pp7[58],pp8[58],pp9[58],pp10[58],pp11[58],pp12[58],pp13[58],pp14[58],pp15[58],pp16[58],pp17[58],pp18[58],pp19[58],pp20[58],pp21[58],pp22[58],pp23[58],pp24[58],pp25[58],pp26[58],pp27[58],pp28[58],pp29[58],pp30[58],pp31[58],pp32[58],pp33[58],pp34[58],pp35[58]};
    CLA_60 KS_3(s3, c3, in3_1, in3_2);
    wire[57:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp6[29],pp6[30],pp6[31],pp6[32],pp6[33],pp6[34],pp6[35],pp6[36],pp6[37],pp6[38],pp6[39],pp6[40],pp6[41],pp6[42],pp6[43],pp6[44],pp6[45],pp6[46],pp6[47],pp6[48],pp6[49],pp6[50],pp6[51],pp6[52],pp6[53],pp6[54],pp6[55],pp6[56],pp6[57],pp7[57],pp8[57],pp9[57],pp10[57],pp11[57],pp12[57],pp13[57],pp14[57],pp15[57],pp16[57],pp17[57],pp18[57],pp19[57],pp20[57],pp21[57],pp22[57],pp23[57],pp24[57],pp25[57],pp26[57],pp27[57],pp28[57],pp29[57],pp30[57],pp31[57],pp32[57],pp33[57],pp34[57],pp35[57]};
    assign in4_2 = {pp7[28],pp7[29],pp7[30],pp7[31],pp7[32],pp7[33],pp7[34],pp7[35],pp7[36],pp7[37],pp7[38],pp7[39],pp7[40],pp7[41],pp7[42],pp7[43],pp7[44],pp7[45],pp7[46],pp7[47],pp7[48],pp7[49],pp7[50],pp7[51],pp7[52],pp7[53],pp7[54],pp7[55],pp7[56],pp8[56],pp9[56],pp10[56],pp11[56],pp12[56],pp13[56],pp14[56],pp15[56],pp16[56],pp17[56],pp18[56],pp19[56],pp20[56],pp21[56],pp22[56],pp23[56],pp24[56],pp25[56],pp26[56],pp27[56],pp28[56],pp29[56],pp30[56],pp31[56],pp32[56],pp33[56],pp34[56],pp35[56],pp36[56]};
    CLA_58 KS_4(s4, c4, in4_1, in4_2);
    wire[55:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp8[28],pp8[29],pp8[30],pp8[31],pp8[32],pp8[33],pp8[34],pp8[35],pp8[36],pp8[37],pp8[38],pp8[39],pp8[40],pp8[41],pp8[42],pp8[43],pp8[44],pp8[45],pp8[46],pp8[47],pp8[48],pp8[49],pp8[50],pp8[51],pp8[52],pp8[53],pp8[54],pp8[55],pp9[55],pp10[55],pp11[55],pp12[55],pp13[55],pp14[55],pp15[55],pp16[55],pp17[55],pp18[55],pp19[55],pp20[55],pp21[55],pp22[55],pp23[55],pp24[55],pp25[55],pp26[55],pp27[55],pp28[55],pp29[55],pp30[55],pp31[55],pp32[55],pp33[55],pp34[55],pp35[55],pp36[55]};
    assign in5_2 = {pp9[27],pp9[28],pp9[29],pp9[30],pp9[31],pp9[32],pp9[33],pp9[34],pp9[35],pp9[36],pp9[37],pp9[38],pp9[39],pp9[40],pp9[41],pp9[42],pp9[43],pp9[44],pp9[45],pp9[46],pp9[47],pp9[48],pp9[49],pp9[50],pp9[51],pp9[52],pp9[53],pp9[54],pp10[54],pp11[54],pp12[54],pp13[54],pp14[54],pp15[54],pp16[54],pp17[54],pp18[54],pp19[54],pp20[54],pp21[54],pp22[54],pp23[54],pp24[54],pp25[54],pp26[54],pp27[54],pp28[54],pp29[54],pp30[54],pp31[54],pp32[54],pp33[54],pp34[54],pp35[54],pp36[54],pp37[54]};
    CLA_56 KS_5(s5, c5, in5_1, in5_2);
    wire[53:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp10[27],pp10[28],pp10[29],pp10[30],pp10[31],pp10[32],pp10[33],pp10[34],pp10[35],pp10[36],pp10[37],pp10[38],pp10[39],pp10[40],pp10[41],pp10[42],pp10[43],pp10[44],pp10[45],pp10[46],pp10[47],pp10[48],pp10[49],pp10[50],pp10[51],pp10[52],pp10[53],pp11[53],pp12[53],pp13[53],pp14[53],pp15[53],pp16[53],pp17[53],pp18[53],pp19[53],pp20[53],pp21[53],pp22[53],pp23[53],pp24[53],pp25[53],pp26[53],pp27[53],pp28[53],pp29[53],pp30[53],pp31[53],pp32[53],pp33[53],pp34[53],pp35[53],pp36[53],pp37[53]};
    assign in6_2 = {pp11[26],pp11[27],pp11[28],pp11[29],pp11[30],pp11[31],pp11[32],pp11[33],pp11[34],pp11[35],pp11[36],pp11[37],pp11[38],pp11[39],pp11[40],pp11[41],pp11[42],pp11[43],pp11[44],pp11[45],pp11[46],pp11[47],pp11[48],pp11[49],pp11[50],pp11[51],pp11[52],pp12[52],pp13[52],pp14[52],pp15[52],pp16[52],pp17[52],pp18[52],pp19[52],pp20[52],pp21[52],pp22[52],pp23[52],pp24[52],pp25[52],pp26[52],pp27[52],pp28[52],pp29[52],pp30[52],pp31[52],pp32[52],pp33[52],pp34[52],pp35[52],pp36[52],pp37[52],pp38[52]};
    CLA_54 KS_6(s6, c6, in6_1, in6_2);
    wire[51:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp12[26],pp12[27],pp12[28],pp12[29],pp12[30],pp12[31],pp12[32],pp12[33],pp12[34],pp12[35],pp12[36],pp12[37],pp12[38],pp12[39],pp12[40],pp12[41],pp12[42],pp12[43],pp12[44],pp12[45],pp12[46],pp12[47],pp12[48],pp12[49],pp12[50],pp12[51],pp13[51],pp14[51],pp15[51],pp16[51],pp17[51],pp18[51],pp19[51],pp20[51],pp21[51],pp22[51],pp23[51],pp24[51],pp25[51],pp26[51],pp27[51],pp28[51],pp29[51],pp30[51],pp31[51],pp32[51],pp33[51],pp34[51],pp35[51],pp36[51],pp37[51],pp38[51]};
    assign in7_2 = {pp13[25],pp13[26],pp13[27],pp13[28],pp13[29],pp13[30],pp13[31],pp13[32],pp13[33],pp13[34],pp13[35],pp13[36],pp13[37],pp13[38],pp13[39],pp13[40],pp13[41],pp13[42],pp13[43],pp13[44],pp13[45],pp13[46],pp13[47],pp13[48],pp13[49],pp13[50],pp14[50],pp15[50],pp16[50],pp17[50],pp18[50],pp19[50],pp20[50],pp21[50],pp22[50],pp23[50],pp24[50],pp25[50],pp26[50],pp27[50],pp28[50],pp29[50],pp30[50],pp31[50],pp32[50],pp33[50],pp34[50],pp35[50],pp36[50],pp37[50],pp38[50],pp39[50]};
    CLA_52 KS_7(s7, c7, in7_1, in7_2);
    wire[49:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp14[25],pp14[26],pp14[27],pp14[28],pp14[29],pp14[30],pp14[31],pp14[32],pp14[33],pp14[34],pp14[35],pp14[36],pp14[37],pp14[38],pp14[39],pp14[40],pp14[41],pp14[42],pp14[43],pp14[44],pp14[45],pp14[46],pp14[47],pp14[48],pp14[49],pp15[49],pp16[49],pp17[49],pp18[49],pp19[49],pp20[49],pp21[49],pp22[49],pp23[49],pp24[49],pp25[49],pp26[49],pp27[49],pp28[49],pp29[49],pp30[49],pp31[49],pp32[49],pp33[49],pp34[49],pp35[49],pp36[49],pp37[49],pp38[49],pp39[49]};
    assign in8_2 = {pp15[24],pp15[25],pp15[26],pp15[27],pp15[28],pp15[29],pp15[30],pp15[31],pp15[32],pp15[33],pp15[34],pp15[35],pp15[36],pp15[37],pp15[38],pp15[39],pp15[40],pp15[41],pp15[42],pp15[43],pp15[44],pp15[45],pp15[46],pp15[47],pp15[48],pp16[48],pp17[48],pp18[48],pp19[48],pp20[48],pp21[48],pp22[48],pp23[48],pp24[48],pp25[48],pp26[48],pp27[48],pp28[48],pp29[48],pp30[48],pp31[48],pp32[48],pp33[48],pp34[48],pp35[48],pp36[48],pp37[48],pp38[48],pp39[48],pp40[48]};
    CLA_50 KS_8(s8, c8, in8_1, in8_2);
    wire[47:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp16[24],pp16[25],pp16[26],pp16[27],pp16[28],pp16[29],pp16[30],pp16[31],pp16[32],pp16[33],pp16[34],pp16[35],pp16[36],pp16[37],pp16[38],pp16[39],pp16[40],pp16[41],pp16[42],pp16[43],pp16[44],pp16[45],pp16[46],pp16[47],pp17[47],pp18[47],pp19[47],pp20[47],pp21[47],pp22[47],pp23[47],pp24[47],pp25[47],pp26[47],pp27[47],pp28[47],pp29[47],pp30[47],pp31[47],pp32[47],pp33[47],pp34[47],pp35[47],pp36[47],pp37[47],pp38[47],pp39[47],pp40[47]};
    assign in9_2 = {pp17[23],pp17[24],pp17[25],pp17[26],pp17[27],pp17[28],pp17[29],pp17[30],pp17[31],pp17[32],pp17[33],pp17[34],pp17[35],pp17[36],pp17[37],pp17[38],pp17[39],pp17[40],pp17[41],pp17[42],pp17[43],pp17[44],pp17[45],pp17[46],pp18[46],pp19[46],pp20[46],pp21[46],pp22[46],pp23[46],pp24[46],pp25[46],pp26[46],pp27[46],pp28[46],pp29[46],pp30[46],pp31[46],pp32[46],pp33[46],pp34[46],pp35[46],pp36[46],pp37[46],pp38[46],pp39[46],pp40[46],pp41[46]};
    CLA_48 KS_9(s9, c9, in9_1, in9_2);
    wire[45:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp18[23],pp18[24],pp18[25],pp18[26],pp18[27],pp18[28],pp18[29],pp18[30],pp18[31],pp18[32],pp18[33],pp18[34],pp18[35],pp18[36],pp18[37],pp18[38],pp18[39],pp18[40],pp18[41],pp18[42],pp18[43],pp18[44],pp18[45],pp19[45],pp20[45],pp21[45],pp22[45],pp23[45],pp24[45],pp25[45],pp26[45],pp27[45],pp28[45],pp29[45],pp30[45],pp31[45],pp32[45],pp33[45],pp34[45],pp35[45],pp36[45],pp37[45],pp38[45],pp39[45],pp40[45],pp41[45]};
    assign in10_2 = {pp19[22],pp19[23],pp19[24],pp19[25],pp19[26],pp19[27],pp19[28],pp19[29],pp19[30],pp19[31],pp19[32],pp19[33],pp19[34],pp19[35],pp19[36],pp19[37],pp19[38],pp19[39],pp19[40],pp19[41],pp19[42],pp19[43],pp19[44],pp20[44],pp21[44],pp22[44],pp23[44],pp24[44],pp25[44],pp26[44],pp27[44],pp28[44],pp29[44],pp30[44],pp31[44],pp32[44],pp33[44],pp34[44],pp35[44],pp36[44],pp37[44],pp38[44],pp39[44],pp40[44],pp41[44],pp42[44]};
    CLA_46 KS_10(s10, c10, in10_1, in10_2);
    wire[43:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp20[22],pp20[23],pp20[24],pp20[25],pp20[26],pp20[27],pp20[28],pp20[29],pp20[30],pp20[31],pp20[32],pp20[33],pp20[34],pp20[35],pp20[36],pp20[37],pp20[38],pp20[39],pp20[40],pp20[41],pp20[42],pp20[43],pp21[43],pp22[43],pp23[43],pp24[43],pp25[43],pp26[43],pp27[43],pp28[43],pp29[43],pp30[43],pp31[43],pp32[43],pp33[43],pp34[43],pp35[43],pp36[43],pp37[43],pp38[43],pp39[43],pp40[43],pp41[43],pp42[43]};
    assign in11_2 = {pp21[21],pp21[22],pp21[23],pp21[24],pp21[25],pp21[26],pp21[27],pp21[28],pp21[29],pp21[30],pp21[31],pp21[32],pp21[33],pp21[34],pp21[35],pp21[36],pp21[37],pp21[38],pp21[39],pp21[40],pp21[41],pp21[42],pp22[42],pp23[42],pp24[42],pp25[42],pp26[42],pp27[42],pp28[42],pp29[42],pp30[42],pp31[42],pp32[42],pp33[42],pp34[42],pp35[42],pp36[42],pp37[42],pp38[42],pp39[42],pp40[42],pp41[42],pp42[42],pp43[42]};
    CLA_44 KS_11(s11, c11, in11_1, in11_2);
    wire[41:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp22[21],pp22[22],pp22[23],pp22[24],pp22[25],pp22[26],pp22[27],pp22[28],pp22[29],pp22[30],pp22[31],pp22[32],pp22[33],pp22[34],pp22[35],pp22[36],pp22[37],pp22[38],pp22[39],pp22[40],pp22[41],pp23[41],pp24[41],pp25[41],pp26[41],pp27[41],pp28[41],pp29[41],pp30[41],pp31[41],pp32[41],pp33[41],pp34[41],pp35[41],pp36[41],pp37[41],pp38[41],pp39[41],pp40[41],pp41[41],pp42[41],pp43[41]};
    assign in12_2 = {pp23[20],pp23[21],pp23[22],pp23[23],pp23[24],pp23[25],pp23[26],pp23[27],pp23[28],pp23[29],pp23[30],pp23[31],pp23[32],pp23[33],pp23[34],pp23[35],pp23[36],pp23[37],pp23[38],pp23[39],pp23[40],pp24[40],pp25[40],pp26[40],pp27[40],pp28[40],pp29[40],pp30[40],pp31[40],pp32[40],pp33[40],pp34[40],pp35[40],pp36[40],pp37[40],pp38[40],pp39[40],pp40[40],pp41[40],pp42[40],pp43[40],pp44[40]};
    CLA_42 KS_12(s12, c12, in12_1, in12_2);
    wire[39:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp24[20],pp24[21],pp24[22],pp24[23],pp24[24],pp24[25],pp24[26],pp24[27],pp24[28],pp24[29],pp24[30],pp24[31],pp24[32],pp24[33],pp24[34],pp24[35],pp24[36],pp24[37],pp24[38],pp24[39],pp25[39],pp26[39],pp27[39],pp28[39],pp29[39],pp30[39],pp31[39],pp32[39],pp33[39],pp34[39],pp35[39],pp36[39],pp37[39],pp38[39],pp39[39],pp40[39],pp41[39],pp42[39],pp43[39],pp44[39]};
    assign in13_2 = {pp25[19],pp25[20],pp25[21],pp25[22],pp25[23],pp25[24],pp25[25],pp25[26],pp25[27],pp25[28],pp25[29],pp25[30],pp25[31],pp25[32],pp25[33],pp25[34],pp25[35],pp25[36],pp25[37],pp25[38],pp26[38],pp27[38],pp28[38],pp29[38],pp30[38],pp31[38],pp32[38],pp33[38],pp34[38],pp35[38],pp36[38],pp37[38],pp38[38],pp39[38],pp40[38],pp41[38],pp42[38],pp43[38],pp44[38],pp45[38]};
    CLA_40 KS_13(s13, c13, in13_1, in13_2);
    wire[37:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp26[19],pp26[20],pp26[21],pp26[22],pp26[23],pp26[24],pp26[25],pp26[26],pp26[27],pp26[28],pp26[29],pp26[30],pp26[31],pp26[32],pp26[33],pp26[34],pp26[35],pp26[36],pp26[37],pp27[37],pp28[37],pp29[37],pp30[37],pp31[37],pp32[37],pp33[37],pp34[37],pp35[37],pp36[37],pp37[37],pp38[37],pp39[37],pp40[37],pp41[37],pp42[37],pp43[37],pp44[37],pp45[37]};
    assign in14_2 = {pp27[18],pp27[19],pp27[20],pp27[21],pp27[22],pp27[23],pp27[24],pp27[25],pp27[26],pp27[27],pp27[28],pp27[29],pp27[30],pp27[31],pp27[32],pp27[33],pp27[34],pp27[35],pp27[36],pp28[36],pp29[36],pp30[36],pp31[36],pp32[36],pp33[36],pp34[36],pp35[36],pp36[36],pp37[36],pp38[36],pp39[36],pp40[36],pp41[36],pp42[36],pp43[36],pp44[36],pp45[36],pp46[36]};
    CLA_38 KS_14(s14, c14, in14_1, in14_2);
    wire[35:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp28[18],pp28[19],pp28[20],pp28[21],pp28[22],pp28[23],pp28[24],pp28[25],pp28[26],pp28[27],pp28[28],pp28[29],pp28[30],pp28[31],pp28[32],pp28[33],pp28[34],pp28[35],pp29[35],pp30[35],pp31[35],pp32[35],pp33[35],pp34[35],pp35[35],pp36[35],pp37[35],pp38[35],pp39[35],pp40[35],pp41[35],pp42[35],pp43[35],pp44[35],pp45[35],pp46[35]};
    assign in15_2 = {pp29[17],pp29[18],pp29[19],pp29[20],pp29[21],pp29[22],pp29[23],pp29[24],pp29[25],pp29[26],pp29[27],pp29[28],pp29[29],pp29[30],pp29[31],pp29[32],pp29[33],pp29[34],pp30[34],pp31[34],pp32[34],pp33[34],pp34[34],pp35[34],pp36[34],pp37[34],pp38[34],pp39[34],pp40[34],pp41[34],pp42[34],pp43[34],pp44[34],pp45[34],pp46[34],pp47[34]};
    CLA_36 KS_15(s15, c15, in15_1, in15_2);
    wire[33:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp30[17],pp30[18],pp30[19],pp30[20],pp30[21],pp30[22],pp30[23],pp30[24],pp30[25],pp30[26],pp30[27],pp30[28],pp30[29],pp30[30],pp30[31],pp30[32],pp30[33],pp31[33],pp32[33],pp33[33],pp34[33],pp35[33],pp36[33],pp37[33],pp38[33],pp39[33],pp40[33],pp41[33],pp42[33],pp43[33],pp44[33],pp45[33],pp46[33],pp47[33]};
    assign in16_2 = {pp31[16],pp31[17],pp31[18],pp31[19],pp31[20],pp31[21],pp31[22],pp31[23],pp31[24],pp31[25],pp31[26],pp31[27],pp31[28],pp31[29],pp31[30],pp31[31],pp31[32],pp32[32],pp33[32],pp34[32],pp35[32],pp36[32],pp37[32],pp38[32],pp39[32],pp40[32],pp41[32],pp42[32],pp43[32],pp44[32],pp45[32],pp46[32],pp47[32],pp48[32]};
    CLA_34 KS_16(s16, c16, in16_1, in16_2);
    wire[31:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp32[16],pp32[17],pp32[18],pp32[19],pp32[20],pp32[21],pp32[22],pp32[23],pp32[24],pp32[25],pp32[26],pp32[27],pp32[28],pp32[29],pp32[30],pp32[31],pp33[31],pp34[31],pp35[31],pp36[31],pp37[31],pp38[31],pp39[31],pp40[31],pp41[31],pp42[31],pp43[31],pp44[31],pp45[31],pp46[31],pp47[31],pp48[31]};
    assign in17_2 = {pp33[15],pp33[16],pp33[17],pp33[18],pp33[19],pp33[20],pp33[21],pp33[22],pp33[23],pp33[24],pp33[25],pp33[26],pp33[27],pp33[28],pp33[29],pp33[30],pp34[30],pp35[30],pp36[30],pp37[30],pp38[30],pp39[30],pp40[30],pp41[30],pp42[30],pp43[30],pp44[30],pp45[30],pp46[30],pp47[30],pp48[30],pp49[30]};
    CLA_32 KS_17(s17, c17, in17_1, in17_2);
    wire[29:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp34[15],pp34[16],pp34[17],pp34[18],pp34[19],pp34[20],pp34[21],pp34[22],pp34[23],pp34[24],pp34[25],pp34[26],pp34[27],pp34[28],pp34[29],pp35[29],pp36[29],pp37[29],pp38[29],pp39[29],pp40[29],pp41[29],pp42[29],pp43[29],pp44[29],pp45[29],pp46[29],pp47[29],pp48[29],pp49[29]};
    assign in18_2 = {pp35[14],pp35[15],pp35[16],pp35[17],pp35[18],pp35[19],pp35[20],pp35[21],pp35[22],pp35[23],pp35[24],pp35[25],pp35[26],pp35[27],pp35[28],pp36[28],pp37[28],pp38[28],pp39[28],pp40[28],pp41[28],pp42[28],pp43[28],pp44[28],pp45[28],pp46[28],pp47[28],pp48[28],pp49[28],pp50[28]};
    CLA_30 KS_18(s18, c18, in18_1, in18_2);
    wire[27:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp36[14],pp36[15],pp36[16],pp36[17],pp36[18],pp36[19],pp36[20],pp36[21],pp36[22],pp36[23],pp36[24],pp36[25],pp36[26],pp36[27],pp37[27],pp38[27],pp39[27],pp40[27],pp41[27],pp42[27],pp43[27],pp44[27],pp45[27],pp46[27],pp47[27],pp48[27],pp49[27],pp50[27]};
    assign in19_2 = {pp37[13],pp37[14],pp37[15],pp37[16],pp37[17],pp37[18],pp37[19],pp37[20],pp37[21],pp37[22],pp37[23],pp37[24],pp37[25],pp37[26],pp38[26],pp39[26],pp40[26],pp41[26],pp42[26],pp43[26],pp44[26],pp45[26],pp46[26],pp47[26],pp48[26],pp49[26],pp50[26],pp51[26]};
    CLA_28 KS_19(s19, c19, in19_1, in19_2);
    wire[25:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp38[13],pp38[14],pp38[15],pp38[16],pp38[17],pp38[18],pp38[19],pp38[20],pp38[21],pp38[22],pp38[23],pp38[24],pp38[25],pp39[25],pp40[25],pp41[25],pp42[25],pp43[25],pp44[25],pp45[25],pp46[25],pp47[25],pp48[25],pp49[25],pp50[25],pp51[25]};
    assign in20_2 = {pp39[12],pp39[13],pp39[14],pp39[15],pp39[16],pp39[17],pp39[18],pp39[19],pp39[20],pp39[21],pp39[22],pp39[23],pp39[24],pp40[24],pp41[24],pp42[24],pp43[24],pp44[24],pp45[24],pp46[24],pp47[24],pp48[24],pp49[24],pp50[24],pp51[24],pp52[24]};
    CLA_26 KS_20(s20, c20, in20_1, in20_2);
    wire[23:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp40[12],pp40[13],pp40[14],pp40[15],pp40[16],pp40[17],pp40[18],pp40[19],pp40[20],pp40[21],pp40[22],pp40[23],pp41[23],pp42[23],pp43[23],pp44[23],pp45[23],pp46[23],pp47[23],pp48[23],pp49[23],pp50[23],pp51[23],pp52[23]};
    assign in21_2 = {pp41[11],pp41[12],pp41[13],pp41[14],pp41[15],pp41[16],pp41[17],pp41[18],pp41[19],pp41[20],pp41[21],pp41[22],pp42[22],pp43[22],pp44[22],pp45[22],pp46[22],pp47[22],pp48[22],pp49[22],pp50[22],pp51[22],pp52[22],pp53[22]};
    CLA_24 KS_21(s21, c21, in21_1, in21_2);
    wire[21:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp42[11],pp42[12],pp42[13],pp42[14],pp42[15],pp42[16],pp42[17],pp42[18],pp42[19],pp42[20],pp42[21],pp43[21],pp44[21],pp45[21],pp46[21],pp47[21],pp48[21],pp49[21],pp50[21],pp51[21],pp52[21],pp53[21]};
    assign in22_2 = {pp43[10],pp43[11],pp43[12],pp43[13],pp43[14],pp43[15],pp43[16],pp43[17],pp43[18],pp43[19],pp43[20],pp44[20],pp45[20],pp46[20],pp47[20],pp48[20],pp49[20],pp50[20],pp51[20],pp52[20],pp53[20],pp54[20]};
    CLA_22 KS_22(s22, c22, in22_1, in22_2);
    wire[19:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp44[10],pp44[11],pp44[12],pp44[13],pp44[14],pp44[15],pp44[16],pp44[17],pp44[18],pp44[19],pp45[19],pp46[19],pp47[19],pp48[19],pp49[19],pp50[19],pp51[19],pp52[19],pp53[19],pp54[19]};
    assign in23_2 = {pp45[9],pp45[10],pp45[11],pp45[12],pp45[13],pp45[14],pp45[15],pp45[16],pp45[17],pp45[18],pp46[18],pp47[18],pp48[18],pp49[18],pp50[18],pp51[18],pp52[18],pp53[18],pp54[18],pp55[18]};
    CLA_20 KS_23(s23, c23, in23_1, in23_2);
    wire[17:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp46[9],pp46[10],pp46[11],pp46[12],pp46[13],pp46[14],pp46[15],pp46[16],pp46[17],pp47[17],pp48[17],pp49[17],pp50[17],pp51[17],pp52[17],pp53[17],pp54[17],pp55[17]};
    assign in24_2 = {pp47[8],pp47[9],pp47[10],pp47[11],pp47[12],pp47[13],pp47[14],pp47[15],pp47[16],pp48[16],pp49[16],pp50[16],pp51[16],pp52[16],pp53[16],pp54[16],pp55[16],pp56[16]};
    CLA_18 KS_24(s24, c24, in24_1, in24_2);
    wire[15:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp48[8],pp48[9],pp48[10],pp48[11],pp48[12],pp48[13],pp48[14],pp48[15],pp49[15],pp50[15],pp51[15],pp52[15],pp53[15],pp54[15],pp55[15],pp56[15]};
    assign in25_2 = {pp49[7],pp49[8],pp49[9],pp49[10],pp49[11],pp49[12],pp49[13],pp49[14],pp50[14],pp51[14],pp52[14],pp53[14],pp54[14],pp55[14],pp56[14],pp57[14]};
    CLA_16 KS_25(s25, c25, in25_1, in25_2);
    wire[13:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp50[7],pp50[8],pp50[9],pp50[10],pp50[11],pp50[12],pp50[13],pp51[13],pp52[13],pp53[13],pp54[13],pp55[13],pp56[13],pp57[13]};
    assign in26_2 = {pp51[6],pp51[7],pp51[8],pp51[9],pp51[10],pp51[11],pp51[12],pp52[12],pp53[12],pp54[12],pp55[12],pp56[12],pp57[12],pp58[12]};
    CLA_14 KS_26(s26, c26, in26_1, in26_2);
    wire[11:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp52[6],pp52[7],pp52[8],pp52[9],pp52[10],pp52[11],pp53[11],pp54[11],pp55[11],pp56[11],pp57[11],pp58[11]};
    assign in27_2 = {pp53[5],pp53[6],pp53[7],pp53[8],pp53[9],pp53[10],pp54[10],pp55[10],pp56[10],pp57[10],pp58[10],pp59[10]};
    CLA_12 KS_27(s27, c27, in27_1, in27_2);
    wire[9:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp54[5],pp54[6],pp54[7],pp54[8],pp54[9],pp55[9],pp56[9],pp57[9],pp58[9],pp59[9]};
    assign in28_2 = {pp55[4],pp55[5],pp55[6],pp55[7],pp55[8],pp56[8],pp57[8],pp58[8],pp59[8],pp60[8]};
    CLA_10 KS_28(s28, c28, in28_1, in28_2);
    wire[7:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp56[4],pp56[5],pp56[6],pp56[7],pp57[7],pp58[7],pp59[7],pp60[7]};
    assign in29_2 = {pp57[3],pp57[4],pp57[5],pp57[6],pp58[6],pp59[6],pp60[6],pp61[6]};
    CLA_8 KS_29(s29, c29, in29_1, in29_2);
    wire[5:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp58[3],pp58[4],pp58[5],pp59[5],pp60[5],pp61[5]};
    assign in30_2 = {pp59[2],pp59[3],pp59[4],pp60[4],pp61[4],pp62[4]};
    CLA_6 KS_30(s30, c30, in30_1, in30_2);
    wire[3:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp60[2],pp60[3],pp61[3],pp62[3]};
    assign in31_2 = {pp61[1],pp61[2],pp62[2],pp63[2]};
    CLA_4 KS_31(s31, c31, in31_1, in31_2);
    wire[1:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp62[1],pp63[1]};
    assign in32_2 = {pp63[0],1'b0};
    CLA_2 KS_32(s32, c32, in32_1, in32_2);

    /*Stage 2*/
    wire[95:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp0[16],pp0[17],pp0[18],pp0[19],pp0[20],pp0[21],pp0[22],pp0[23],pp0[24],pp0[25],pp0[26],pp0[27],pp0[28],pp0[29],pp0[30],pp0[31],pp2[30],pp4[29],pp6[28],pp8[27],pp10[26],pp12[25],pp14[24],pp16[23],pp18[22],pp20[21],pp22[20],pp24[19],pp26[18],pp28[17],pp30[16],pp32[15],pp34[14],pp36[13],pp38[12],pp40[11],pp42[10],pp44[9],pp46[8],pp48[7],pp50[6],pp52[5],pp54[4],pp56[3],pp58[2],pp60[1],pp62[0],s1[31],s1[32],s1[33],pp63[3],pp62[5],pp61[7],pp60[9],pp59[11],pp58[13],pp57[15],pp56[17],pp55[19],pp54[21],pp53[23],pp52[25],pp51[27],pp50[29],pp49[31],pp48[33],pp47[35],pp46[37],pp45[39],pp44[41],pp43[43],pp42[45],pp41[47],pp40[49],pp39[51],pp38[53],pp37[55],pp36[57],pp35[59],pp34[61],pp33[63],pp34[63],pp35[63],pp36[63],pp37[63],pp38[63],pp39[63],pp40[63],pp41[63],pp42[63],pp43[63],pp44[63],pp45[63],pp46[63],pp47[63],pp48[63]};
    assign in33_2 = {pp1[15],pp1[16],pp1[17],pp1[18],pp1[19],pp1[20],pp1[21],pp1[22],pp1[23],pp1[24],pp1[25],pp1[26],pp1[27],pp1[28],pp1[29],pp1[30],pp3[29],pp5[28],pp7[27],pp9[26],pp11[25],pp13[24],pp15[23],pp17[22],pp19[21],pp21[20],pp23[19],pp25[18],pp27[17],pp29[16],pp31[15],pp33[14],pp35[13],pp37[12],pp39[11],pp41[10],pp43[9],pp45[8],pp47[7],pp49[6],pp51[5],pp53[4],pp55[3],pp57[2],pp59[1],pp61[0],s1[30],s2[30],s2[31],s2[32],s1[34],pp63[4],pp62[6],pp61[8],pp60[10],pp59[12],pp58[14],pp57[16],pp56[18],pp55[20],pp54[22],pp53[24],pp52[26],pp51[28],pp50[30],pp49[32],pp48[34],pp47[36],pp46[38],pp45[40],pp44[42],pp43[44],pp42[46],pp41[48],pp40[50],pp39[52],pp38[54],pp37[56],pp36[58],pp35[60],pp34[62],pp35[62],pp36[62],pp37[62],pp38[62],pp39[62],pp40[62],pp41[62],pp42[62],pp43[62],pp44[62],pp45[62],pp46[62],pp47[62],pp48[62],pp49[62]};
    CLA_96 KS_33(s33, c33, in33_1, in33_2);
    wire[93:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp2[15],pp2[16],pp2[17],pp2[18],pp2[19],pp2[20],pp2[21],pp2[22],pp2[23],pp2[24],pp2[25],pp2[26],pp2[27],pp2[28],pp2[29],pp4[28],pp6[27],pp8[26],pp10[25],pp12[24],pp14[23],pp16[22],pp18[21],pp20[20],pp22[19],pp24[18],pp26[17],pp28[16],pp30[15],pp32[14],pp34[13],pp36[12],pp38[11],pp40[10],pp42[9],pp44[8],pp46[7],pp48[6],pp50[5],pp52[4],pp54[3],pp56[2],pp58[1],pp60[0],s1[29],s2[29],s3[29],s3[30],s3[31],s2[33],s1[35],pp63[5],pp62[7],pp61[9],pp60[11],pp59[13],pp58[15],pp57[17],pp56[19],pp55[21],pp54[23],pp53[25],pp52[27],pp51[29],pp50[31],pp49[33],pp48[35],pp47[37],pp46[39],pp45[41],pp44[43],pp43[45],pp42[47],pp41[49],pp40[51],pp39[53],pp38[55],pp37[57],pp36[59],pp35[61],pp36[61],pp37[61],pp38[61],pp39[61],pp40[61],pp41[61],pp42[61],pp43[61],pp44[61],pp45[61],pp46[61],pp47[61],pp48[61],pp49[61]};
    assign in34_2 = {pp3[14],pp3[15],pp3[16],pp3[17],pp3[18],pp3[19],pp3[20],pp3[21],pp3[22],pp3[23],pp3[24],pp3[25],pp3[26],pp3[27],pp3[28],pp5[27],pp7[26],pp9[25],pp11[24],pp13[23],pp15[22],pp17[21],pp19[20],pp21[19],pp23[18],pp25[17],pp27[16],pp29[15],pp31[14],pp33[13],pp35[12],pp37[11],pp39[10],pp41[9],pp43[8],pp45[7],pp47[6],pp49[5],pp51[4],pp53[3],pp55[2],pp57[1],pp59[0],s1[28],s2[28],s3[28],s4[28],s4[29],s4[30],s3[32],s2[34],s1[36],pp63[6],pp62[8],pp61[10],pp60[12],pp59[14],pp58[16],pp57[18],pp56[20],pp55[22],pp54[24],pp53[26],pp52[28],pp51[30],pp50[32],pp49[34],pp48[36],pp47[38],pp46[40],pp45[42],pp44[44],pp43[46],pp42[48],pp41[50],pp40[52],pp39[54],pp38[56],pp37[58],pp36[60],pp37[60],pp38[60],pp39[60],pp40[60],pp41[60],pp42[60],pp43[60],pp44[60],pp45[60],pp46[60],pp47[60],pp48[60],pp49[60],pp50[60]};
    CLA_94 KS_34(s34, c34, in34_1, in34_2);
    wire[91:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp4[14],pp4[15],pp4[16],pp4[17],pp4[18],pp4[19],pp4[20],pp4[21],pp4[22],pp4[23],pp4[24],pp4[25],pp4[26],pp4[27],pp6[26],pp8[25],pp10[24],pp12[23],pp14[22],pp16[21],pp18[20],pp20[19],pp22[18],pp24[17],pp26[16],pp28[15],pp30[14],pp32[13],pp34[12],pp36[11],pp38[10],pp40[9],pp42[8],pp44[7],pp46[6],pp48[5],pp50[4],pp52[3],pp54[2],pp56[1],pp58[0],s1[27],s2[27],s3[27],s4[27],s5[27],s5[28],s5[29],s4[31],s3[33],s2[35],s1[37],pp63[7],pp62[9],pp61[11],pp60[13],pp59[15],pp58[17],pp57[19],pp56[21],pp55[23],pp54[25],pp53[27],pp52[29],pp51[31],pp50[33],pp49[35],pp48[37],pp47[39],pp46[41],pp45[43],pp44[45],pp43[47],pp42[49],pp41[51],pp40[53],pp39[55],pp38[57],pp37[59],pp38[59],pp39[59],pp40[59],pp41[59],pp42[59],pp43[59],pp44[59],pp45[59],pp46[59],pp47[59],pp48[59],pp49[59],pp50[59]};
    assign in35_2 = {pp5[13],pp5[14],pp5[15],pp5[16],pp5[17],pp5[18],pp5[19],pp5[20],pp5[21],pp5[22],pp5[23],pp5[24],pp5[25],pp5[26],pp7[25],pp9[24],pp11[23],pp13[22],pp15[21],pp17[20],pp19[19],pp21[18],pp23[17],pp25[16],pp27[15],pp29[14],pp31[13],pp33[12],pp35[11],pp37[10],pp39[9],pp41[8],pp43[7],pp45[6],pp47[5],pp49[4],pp51[3],pp53[2],pp55[1],pp57[0],s1[26],s2[26],s3[26],s4[26],s5[26],s6[26],s6[27],s6[28],s5[30],s4[32],s3[34],s2[36],s1[38],pp63[8],pp62[10],pp61[12],pp60[14],pp59[16],pp58[18],pp57[20],pp56[22],pp55[24],pp54[26],pp53[28],pp52[30],pp51[32],pp50[34],pp49[36],pp48[38],pp47[40],pp46[42],pp45[44],pp44[46],pp43[48],pp42[50],pp41[52],pp40[54],pp39[56],pp38[58],pp39[58],pp40[58],pp41[58],pp42[58],pp43[58],pp44[58],pp45[58],pp46[58],pp47[58],pp48[58],pp49[58],pp50[58],pp51[58]};
    CLA_92 KS_35(s35, c35, in35_1, in35_2);
    wire[89:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp6[13],pp6[14],pp6[15],pp6[16],pp6[17],pp6[18],pp6[19],pp6[20],pp6[21],pp6[22],pp6[23],pp6[24],pp6[25],pp8[24],pp10[23],pp12[22],pp14[21],pp16[20],pp18[19],pp20[18],pp22[17],pp24[16],pp26[15],pp28[14],pp30[13],pp32[12],pp34[11],pp36[10],pp38[9],pp40[8],pp42[7],pp44[6],pp46[5],pp48[4],pp50[3],pp52[2],pp54[1],pp56[0],s1[25],s2[25],s3[25],s4[25],s5[25],s6[25],s7[25],s7[26],s7[27],s6[29],s5[31],s4[33],s3[35],s2[37],s1[39],pp63[9],pp62[11],pp61[13],pp60[15],pp59[17],pp58[19],pp57[21],pp56[23],pp55[25],pp54[27],pp53[29],pp52[31],pp51[33],pp50[35],pp49[37],pp48[39],pp47[41],pp46[43],pp45[45],pp44[47],pp43[49],pp42[51],pp41[53],pp40[55],pp39[57],pp40[57],pp41[57],pp42[57],pp43[57],pp44[57],pp45[57],pp46[57],pp47[57],pp48[57],pp49[57],pp50[57],pp51[57]};
    assign in36_2 = {pp7[12],pp7[13],pp7[14],pp7[15],pp7[16],pp7[17],pp7[18],pp7[19],pp7[20],pp7[21],pp7[22],pp7[23],pp7[24],pp9[23],pp11[22],pp13[21],pp15[20],pp17[19],pp19[18],pp21[17],pp23[16],pp25[15],pp27[14],pp29[13],pp31[12],pp33[11],pp35[10],pp37[9],pp39[8],pp41[7],pp43[6],pp45[5],pp47[4],pp49[3],pp51[2],pp53[1],pp55[0],s1[24],s2[24],s3[24],s4[24],s5[24],s6[24],s7[24],s8[24],s8[25],s8[26],s7[28],s6[30],s5[32],s4[34],s3[36],s2[38],s1[40],pp63[10],pp62[12],pp61[14],pp60[16],pp59[18],pp58[20],pp57[22],pp56[24],pp55[26],pp54[28],pp53[30],pp52[32],pp51[34],pp50[36],pp49[38],pp48[40],pp47[42],pp46[44],pp45[46],pp44[48],pp43[50],pp42[52],pp41[54],pp40[56],pp41[56],pp42[56],pp43[56],pp44[56],pp45[56],pp46[56],pp47[56],pp48[56],pp49[56],pp50[56],pp51[56],pp52[56]};
    CLA_90 KS_36(s36, c36, in36_1, in36_2);
    wire[87:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp8[12],pp8[13],pp8[14],pp8[15],pp8[16],pp8[17],pp8[18],pp8[19],pp8[20],pp8[21],pp8[22],pp8[23],pp10[22],pp12[21],pp14[20],pp16[19],pp18[18],pp20[17],pp22[16],pp24[15],pp26[14],pp28[13],pp30[12],pp32[11],pp34[10],pp36[9],pp38[8],pp40[7],pp42[6],pp44[5],pp46[4],pp48[3],pp50[2],pp52[1],pp54[0],s1[23],s2[23],s3[23],s4[23],s5[23],s6[23],s7[23],s8[23],s9[23],s9[24],s9[25],s8[27],s7[29],s6[31],s5[33],s4[35],s3[37],s2[39],s1[41],pp63[11],pp62[13],pp61[15],pp60[17],pp59[19],pp58[21],pp57[23],pp56[25],pp55[27],pp54[29],pp53[31],pp52[33],pp51[35],pp50[37],pp49[39],pp48[41],pp47[43],pp46[45],pp45[47],pp44[49],pp43[51],pp42[53],pp41[55],pp42[55],pp43[55],pp44[55],pp45[55],pp46[55],pp47[55],pp48[55],pp49[55],pp50[55],pp51[55],pp52[55]};
    assign in37_2 = {pp9[11],pp9[12],pp9[13],pp9[14],pp9[15],pp9[16],pp9[17],pp9[18],pp9[19],pp9[20],pp9[21],pp9[22],pp11[21],pp13[20],pp15[19],pp17[18],pp19[17],pp21[16],pp23[15],pp25[14],pp27[13],pp29[12],pp31[11],pp33[10],pp35[9],pp37[8],pp39[7],pp41[6],pp43[5],pp45[4],pp47[3],pp49[2],pp51[1],pp53[0],s1[22],s2[22],s3[22],s4[22],s5[22],s6[22],s7[22],s8[22],s9[22],s10[22],s10[23],s10[24],s9[26],s8[28],s7[30],s6[32],s5[34],s4[36],s3[38],s2[40],s1[42],pp63[12],pp62[14],pp61[16],pp60[18],pp59[20],pp58[22],pp57[24],pp56[26],pp55[28],pp54[30],pp53[32],pp52[34],pp51[36],pp50[38],pp49[40],pp48[42],pp47[44],pp46[46],pp45[48],pp44[50],pp43[52],pp42[54],pp43[54],pp44[54],pp45[54],pp46[54],pp47[54],pp48[54],pp49[54],pp50[54],pp51[54],pp52[54],pp53[54]};
    CLA_88 KS_37(s37, c37, in37_1, in37_2);
    wire[85:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp10[11],pp10[12],pp10[13],pp10[14],pp10[15],pp10[16],pp10[17],pp10[18],pp10[19],pp10[20],pp10[21],pp12[20],pp14[19],pp16[18],pp18[17],pp20[16],pp22[15],pp24[14],pp26[13],pp28[12],pp30[11],pp32[10],pp34[9],pp36[8],pp38[7],pp40[6],pp42[5],pp44[4],pp46[3],pp48[2],pp50[1],pp52[0],s1[21],s2[21],s3[21],s4[21],s5[21],s6[21],s7[21],s8[21],s9[21],s10[21],s11[21],s11[22],s11[23],s10[25],s9[27],s8[29],s7[31],s6[33],s5[35],s4[37],s3[39],s2[41],s1[43],pp63[13],pp62[15],pp61[17],pp60[19],pp59[21],pp58[23],pp57[25],pp56[27],pp55[29],pp54[31],pp53[33],pp52[35],pp51[37],pp50[39],pp49[41],pp48[43],pp47[45],pp46[47],pp45[49],pp44[51],pp43[53],pp44[53],pp45[53],pp46[53],pp47[53],pp48[53],pp49[53],pp50[53],pp51[53],pp52[53],pp53[53]};
    assign in38_2 = {pp11[10],pp11[11],pp11[12],pp11[13],pp11[14],pp11[15],pp11[16],pp11[17],pp11[18],pp11[19],pp11[20],pp13[19],pp15[18],pp17[17],pp19[16],pp21[15],pp23[14],pp25[13],pp27[12],pp29[11],pp31[10],pp33[9],pp35[8],pp37[7],pp39[6],pp41[5],pp43[4],pp45[3],pp47[2],pp49[1],pp51[0],s1[20],s2[20],s3[20],s4[20],s5[20],s6[20],s7[20],s8[20],s9[20],s10[20],s11[20],s12[20],s12[21],s12[22],s11[24],s10[26],s9[28],s8[30],s7[32],s6[34],s5[36],s4[38],s3[40],s2[42],s1[44],pp63[14],pp62[16],pp61[18],pp60[20],pp59[22],pp58[24],pp57[26],pp56[28],pp55[30],pp54[32],pp53[34],pp52[36],pp51[38],pp50[40],pp49[42],pp48[44],pp47[46],pp46[48],pp45[50],pp44[52],pp45[52],pp46[52],pp47[52],pp48[52],pp49[52],pp50[52],pp51[52],pp52[52],pp53[52],pp54[52]};
    CLA_86 KS_38(s38, c38, in38_1, in38_2);
    wire[83:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp12[10],pp12[11],pp12[12],pp12[13],pp12[14],pp12[15],pp12[16],pp12[17],pp12[18],pp12[19],pp14[18],pp16[17],pp18[16],pp20[15],pp22[14],pp24[13],pp26[12],pp28[11],pp30[10],pp32[9],pp34[8],pp36[7],pp38[6],pp40[5],pp42[4],pp44[3],pp46[2],pp48[1],pp50[0],s1[19],s2[19],s3[19],s4[19],s5[19],s6[19],s7[19],s8[19],s9[19],s10[19],s11[19],s12[19],s13[19],s13[20],s13[21],s12[23],s11[25],s10[27],s9[29],s8[31],s7[33],s6[35],s5[37],s4[39],s3[41],s2[43],s1[45],pp63[15],pp62[17],pp61[19],pp60[21],pp59[23],pp58[25],pp57[27],pp56[29],pp55[31],pp54[33],pp53[35],pp52[37],pp51[39],pp50[41],pp49[43],pp48[45],pp47[47],pp46[49],pp45[51],pp46[51],pp47[51],pp48[51],pp49[51],pp50[51],pp51[51],pp52[51],pp53[51],pp54[51]};
    assign in39_2 = {pp13[9],pp13[10],pp13[11],pp13[12],pp13[13],pp13[14],pp13[15],pp13[16],pp13[17],pp13[18],pp15[17],pp17[16],pp19[15],pp21[14],pp23[13],pp25[12],pp27[11],pp29[10],pp31[9],pp33[8],pp35[7],pp37[6],pp39[5],pp41[4],pp43[3],pp45[2],pp47[1],pp49[0],s1[18],s2[18],s3[18],s4[18],s5[18],s6[18],s7[18],s8[18],s9[18],s10[18],s11[18],s12[18],s13[18],s14[18],s14[19],s14[20],s13[22],s12[24],s11[26],s10[28],s9[30],s8[32],s7[34],s6[36],s5[38],s4[40],s3[42],s2[44],s1[46],pp63[16],pp62[18],pp61[20],pp60[22],pp59[24],pp58[26],pp57[28],pp56[30],pp55[32],pp54[34],pp53[36],pp52[38],pp51[40],pp50[42],pp49[44],pp48[46],pp47[48],pp46[50],pp47[50],pp48[50],pp49[50],pp50[50],pp51[50],pp52[50],pp53[50],pp54[50],pp55[50]};
    CLA_84 KS_39(s39, c39, in39_1, in39_2);
    wire[81:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp14[9],pp14[10],pp14[11],pp14[12],pp14[13],pp14[14],pp14[15],pp14[16],pp14[17],pp16[16],pp18[15],pp20[14],pp22[13],pp24[12],pp26[11],pp28[10],pp30[9],pp32[8],pp34[7],pp36[6],pp38[5],pp40[4],pp42[3],pp44[2],pp46[1],pp48[0],s1[17],s2[17],s3[17],s4[17],s5[17],s6[17],s7[17],s8[17],s9[17],s10[17],s11[17],s12[17],s13[17],s14[17],s15[17],s15[18],s15[19],s14[21],s13[23],s12[25],s11[27],s10[29],s9[31],s8[33],s7[35],s6[37],s5[39],s4[41],s3[43],s2[45],s1[47],pp63[17],pp62[19],pp61[21],pp60[23],pp59[25],pp58[27],pp57[29],pp56[31],pp55[33],pp54[35],pp53[37],pp52[39],pp51[41],pp50[43],pp49[45],pp48[47],pp47[49],pp48[49],pp49[49],pp50[49],pp51[49],pp52[49],pp53[49],pp54[49],pp55[49]};
    assign in40_2 = {pp15[8],pp15[9],pp15[10],pp15[11],pp15[12],pp15[13],pp15[14],pp15[15],pp15[16],pp17[15],pp19[14],pp21[13],pp23[12],pp25[11],pp27[10],pp29[9],pp31[8],pp33[7],pp35[6],pp37[5],pp39[4],pp41[3],pp43[2],pp45[1],pp47[0],s1[16],s2[16],s3[16],s4[16],s5[16],s6[16],s7[16],s8[16],s9[16],s10[16],s11[16],s12[16],s13[16],s14[16],s15[16],s16[16],s16[17],s16[18],s15[20],s14[22],s13[24],s12[26],s11[28],s10[30],s9[32],s8[34],s7[36],s6[38],s5[40],s4[42],s3[44],s2[46],s1[48],pp63[18],pp62[20],pp61[22],pp60[24],pp59[26],pp58[28],pp57[30],pp56[32],pp55[34],pp54[36],pp53[38],pp52[40],pp51[42],pp50[44],pp49[46],pp48[48],pp49[48],pp50[48],pp51[48],pp52[48],pp53[48],pp54[48],pp55[48],pp56[48]};
    CLA_82 KS_40(s40, c40, in40_1, in40_2);
    wire[79:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp16[8],pp16[9],pp16[10],pp16[11],pp16[12],pp16[13],pp16[14],pp16[15],pp18[14],pp20[13],pp22[12],pp24[11],pp26[10],pp28[9],pp30[8],pp32[7],pp34[6],pp36[5],pp38[4],pp40[3],pp42[2],pp44[1],pp46[0],s1[15],s2[15],s3[15],s4[15],s5[15],s6[15],s7[15],s8[15],s9[15],s10[15],s11[15],s12[15],s13[15],s14[15],s15[15],s16[15],s17[15],s17[16],s17[17],s16[19],s15[21],s14[23],s13[25],s12[27],s11[29],s10[31],s9[33],s8[35],s7[37],s6[39],s5[41],s4[43],s3[45],s2[47],s1[49],pp63[19],pp62[21],pp61[23],pp60[25],pp59[27],pp58[29],pp57[31],pp56[33],pp55[35],pp54[37],pp53[39],pp52[41],pp51[43],pp50[45],pp49[47],pp50[47],pp51[47],pp52[47],pp53[47],pp54[47],pp55[47],pp56[47]};
    assign in41_2 = {pp17[7],pp17[8],pp17[9],pp17[10],pp17[11],pp17[12],pp17[13],pp17[14],pp19[13],pp21[12],pp23[11],pp25[10],pp27[9],pp29[8],pp31[7],pp33[6],pp35[5],pp37[4],pp39[3],pp41[2],pp43[1],pp45[0],s1[14],s2[14],s3[14],s4[14],s5[14],s6[14],s7[14],s8[14],s9[14],s10[14],s11[14],s12[14],s13[14],s14[14],s15[14],s16[14],s17[14],s18[14],s18[15],s18[16],s17[18],s16[20],s15[22],s14[24],s13[26],s12[28],s11[30],s10[32],s9[34],s8[36],s7[38],s6[40],s5[42],s4[44],s3[46],s2[48],s1[50],pp63[20],pp62[22],pp61[24],pp60[26],pp59[28],pp58[30],pp57[32],pp56[34],pp55[36],pp54[38],pp53[40],pp52[42],pp51[44],pp50[46],pp51[46],pp52[46],pp53[46],pp54[46],pp55[46],pp56[46],pp57[46]};
    CLA_80 KS_41(s41, c41, in41_1, in41_2);
    wire[77:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp18[7],pp18[8],pp18[9],pp18[10],pp18[11],pp18[12],pp18[13],pp20[12],pp22[11],pp24[10],pp26[9],pp28[8],pp30[7],pp32[6],pp34[5],pp36[4],pp38[3],pp40[2],pp42[1],pp44[0],s1[13],s2[13],s3[13],s4[13],s5[13],s6[13],s7[13],s8[13],s9[13],s10[13],s11[13],s12[13],s13[13],s14[13],s15[13],s16[13],s17[13],s18[13],s19[13],s19[14],s19[15],s18[17],s17[19],s16[21],s15[23],s14[25],s13[27],s12[29],s11[31],s10[33],s9[35],s8[37],s7[39],s6[41],s5[43],s4[45],s3[47],s2[49],s1[51],pp63[21],pp62[23],pp61[25],pp60[27],pp59[29],pp58[31],pp57[33],pp56[35],pp55[37],pp54[39],pp53[41],pp52[43],pp51[45],pp52[45],pp53[45],pp54[45],pp55[45],pp56[45],pp57[45]};
    assign in42_2 = {pp19[6],pp19[7],pp19[8],pp19[9],pp19[10],pp19[11],pp19[12],pp21[11],pp23[10],pp25[9],pp27[8],pp29[7],pp31[6],pp33[5],pp35[4],pp37[3],pp39[2],pp41[1],pp43[0],s1[12],s2[12],s3[12],s4[12],s5[12],s6[12],s7[12],s8[12],s9[12],s10[12],s11[12],s12[12],s13[12],s14[12],s15[12],s16[12],s17[12],s18[12],s19[12],s20[12],s20[13],s20[14],s19[16],s18[18],s17[20],s16[22],s15[24],s14[26],s13[28],s12[30],s11[32],s10[34],s9[36],s8[38],s7[40],s6[42],s5[44],s4[46],s3[48],s2[50],s1[52],pp63[22],pp62[24],pp61[26],pp60[28],pp59[30],pp58[32],pp57[34],pp56[36],pp55[38],pp54[40],pp53[42],pp52[44],pp53[44],pp54[44],pp55[44],pp56[44],pp57[44],pp58[44]};
    CLA_78 KS_42(s42, c42, in42_1, in42_2);
    wire[75:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp20[6],pp20[7],pp20[8],pp20[9],pp20[10],pp20[11],pp22[10],pp24[9],pp26[8],pp28[7],pp30[6],pp32[5],pp34[4],pp36[3],pp38[2],pp40[1],pp42[0],s1[11],s2[11],s3[11],s4[11],s5[11],s6[11],s7[11],s8[11],s9[11],s10[11],s11[11],s12[11],s13[11],s14[11],s15[11],s16[11],s17[11],s18[11],s19[11],s20[11],s21[11],s21[12],s21[13],s20[15],s19[17],s18[19],s17[21],s16[23],s15[25],s14[27],s13[29],s12[31],s11[33],s10[35],s9[37],s8[39],s7[41],s6[43],s5[45],s4[47],s3[49],s2[51],s1[53],pp63[23],pp62[25],pp61[27],pp60[29],pp59[31],pp58[33],pp57[35],pp56[37],pp55[39],pp54[41],pp53[43],pp54[43],pp55[43],pp56[43],pp57[43],pp58[43]};
    assign in43_2 = {pp21[5],pp21[6],pp21[7],pp21[8],pp21[9],pp21[10],pp23[9],pp25[8],pp27[7],pp29[6],pp31[5],pp33[4],pp35[3],pp37[2],pp39[1],pp41[0],s1[10],s2[10],s3[10],s4[10],s5[10],s6[10],s7[10],s8[10],s9[10],s10[10],s11[10],s12[10],s13[10],s14[10],s15[10],s16[10],s17[10],s18[10],s19[10],s20[10],s21[10],s22[10],s22[11],s22[12],s21[14],s20[16],s19[18],s18[20],s17[22],s16[24],s15[26],s14[28],s13[30],s12[32],s11[34],s10[36],s9[38],s8[40],s7[42],s6[44],s5[46],s4[48],s3[50],s2[52],s1[54],pp63[24],pp62[26],pp61[28],pp60[30],pp59[32],pp58[34],pp57[36],pp56[38],pp55[40],pp54[42],pp55[42],pp56[42],pp57[42],pp58[42],pp59[42]};
    CLA_76 KS_43(s43, c43, in43_1, in43_2);
    wire[73:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[5],pp22[6],pp22[7],pp22[8],pp22[9],pp24[8],pp26[7],pp28[6],pp30[5],pp32[4],pp34[3],pp36[2],pp38[1],pp40[0],s1[9],s2[9],s3[9],s4[9],s5[9],s6[9],s7[9],s8[9],s9[9],s10[9],s11[9],s12[9],s13[9],s14[9],s15[9],s16[9],s17[9],s18[9],s19[9],s20[9],s21[9],s22[9],s23[9],s23[10],s23[11],s22[13],s21[15],s20[17],s19[19],s18[21],s17[23],s16[25],s15[27],s14[29],s13[31],s12[33],s11[35],s10[37],s9[39],s8[41],s7[43],s6[45],s5[47],s4[49],s3[51],s2[53],s1[55],pp63[25],pp62[27],pp61[29],pp60[31],pp59[33],pp58[35],pp57[37],pp56[39],pp55[41],pp56[41],pp57[41],pp58[41],pp59[41]};
    assign in44_2 = {pp23[4],pp23[5],pp23[6],pp23[7],pp23[8],pp25[7],pp27[6],pp29[5],pp31[4],pp33[3],pp35[2],pp37[1],pp39[0],s1[8],s2[8],s3[8],s4[8],s5[8],s6[8],s7[8],s8[8],s9[8],s10[8],s11[8],s12[8],s13[8],s14[8],s15[8],s16[8],s17[8],s18[8],s19[8],s20[8],s21[8],s22[8],s23[8],s24[8],s24[9],s24[10],s23[12],s22[14],s21[16],s20[18],s19[20],s18[22],s17[24],s16[26],s15[28],s14[30],s13[32],s12[34],s11[36],s10[38],s9[40],s8[42],s7[44],s6[46],s5[48],s4[50],s3[52],s2[54],s1[56],pp63[26],pp62[28],pp61[30],pp60[32],pp59[34],pp58[36],pp57[38],pp56[40],pp57[40],pp58[40],pp59[40],pp60[40]};
    CLA_74 KS_44(s44, c44, in44_1, in44_2);
    wire[71:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[4],pp24[5],pp24[6],pp24[7],pp26[6],pp28[5],pp30[4],pp32[3],pp34[2],pp36[1],pp38[0],s1[7],s2[7],s3[7],s4[7],s5[7],s6[7],s7[7],s8[7],s9[7],s10[7],s11[7],s12[7],s13[7],s14[7],s15[7],s16[7],s17[7],s18[7],s19[7],s20[7],s21[7],s22[7],s23[7],s24[7],s25[7],s25[8],s25[9],s24[11],s23[13],s22[15],s21[17],s20[19],s19[21],s18[23],s17[25],s16[27],s15[29],s14[31],s13[33],s12[35],s11[37],s10[39],s9[41],s8[43],s7[45],s6[47],s5[49],s4[51],s3[53],s2[55],s1[57],pp63[27],pp62[29],pp61[31],pp60[33],pp59[35],pp58[37],pp57[39],pp58[39],pp59[39],pp60[39]};
    assign in45_2 = {pp25[3],pp25[4],pp25[5],pp25[6],pp27[5],pp29[4],pp31[3],pp33[2],pp35[1],pp37[0],s1[6],s2[6],s3[6],s4[6],s5[6],s6[6],s7[6],s8[6],s9[6],s10[6],s11[6],s12[6],s13[6],s14[6],s15[6],s16[6],s17[6],s18[6],s19[6],s20[6],s21[6],s22[6],s23[6],s24[6],s25[6],s26[6],s26[7],s26[8],s25[10],s24[12],s23[14],s22[16],s21[18],s20[20],s19[22],s18[24],s17[26],s16[28],s15[30],s14[32],s13[34],s12[36],s11[38],s10[40],s9[42],s8[44],s7[46],s6[48],s5[50],s4[52],s3[54],s2[56],s1[58],pp63[28],pp62[30],pp61[32],pp60[34],pp59[36],pp58[38],pp59[38],pp60[38],pp61[38]};
    CLA_72 KS_45(s45, c45, in45_1, in45_2);
    wire[69:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp26[3],pp26[4],pp26[5],pp28[4],pp30[3],pp32[2],pp34[1],pp36[0],s1[5],s2[5],s3[5],s4[5],s5[5],s6[5],s7[5],s8[5],s9[5],s10[5],s11[5],s12[5],s13[5],s14[5],s15[5],s16[5],s17[5],s18[5],s19[5],s20[5],s21[5],s22[5],s23[5],s24[5],s25[5],s26[5],s27[5],s27[6],s27[7],s26[9],s25[11],s24[13],s23[15],s22[17],s21[19],s20[21],s19[23],s18[25],s17[27],s16[29],s15[31],s14[33],s13[35],s12[37],s11[39],s10[41],s9[43],s8[45],s7[47],s6[49],s5[51],s4[53],s3[55],s2[57],s1[59],pp63[29],pp62[31],pp61[33],pp60[35],pp59[37],pp60[37],pp61[37]};
    assign in46_2 = {pp27[2],pp27[3],pp27[4],pp29[3],pp31[2],pp33[1],pp35[0],s1[4],s2[4],s3[4],s4[4],s5[4],s6[4],s7[4],s8[4],s9[4],s10[4],s11[4],s12[4],s13[4],s14[4],s15[4],s16[4],s17[4],s18[4],s19[4],s20[4],s21[4],s22[4],s23[4],s24[4],s25[4],s26[4],s27[4],s28[4],s28[5],s28[6],s27[8],s26[10],s25[12],s24[14],s23[16],s22[18],s21[20],s20[22],s19[24],s18[26],s17[28],s16[30],s15[32],s14[34],s13[36],s12[38],s11[40],s10[42],s9[44],s8[46],s7[48],s6[50],s5[52],s4[54],s3[56],s2[58],s1[60],pp63[30],pp62[32],pp61[34],pp60[36],pp61[36],pp62[36]};
    CLA_70 KS_46(s46, c46, in46_1, in46_2);
    wire[67:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp28[2],pp28[3],pp30[2],pp32[1],pp34[0],s1[3],s2[3],s3[3],s4[3],s5[3],s6[3],s7[3],s8[3],s9[3],s10[3],s11[3],s12[3],s13[3],s14[3],s15[3],s16[3],s17[3],s18[3],s19[3],s20[3],s21[3],s22[3],s23[3],s24[3],s25[3],s26[3],s27[3],s28[3],s29[3],s29[4],s29[5],s28[7],s27[9],s26[11],s25[13],s24[15],s23[17],s22[19],s21[21],s20[23],s19[25],s18[27],s17[29],s16[31],s15[33],s14[35],s13[37],s12[39],s11[41],s10[43],s9[45],s8[47],s7[49],s6[51],s5[53],s4[55],s3[57],s2[59],s1[61],pp63[31],pp62[33],pp61[35],pp62[35]};
    assign in47_2 = {pp29[1],pp29[2],pp31[1],pp33[0],s1[2],s2[2],s3[2],s4[2],s5[2],s6[2],s7[2],s8[2],s9[2],s10[2],s11[2],s12[2],s13[2],s14[2],s15[2],s16[2],s17[2],s18[2],s19[2],s20[2],s21[2],s22[2],s23[2],s24[2],s25[2],s26[2],s27[2],s28[2],s29[2],s30[2],s30[3],s30[4],s29[6],s28[8],s27[10],s26[12],s25[14],s24[16],s23[18],s22[20],s21[22],s20[24],s19[26],s18[28],s17[30],s16[32],s15[34],s14[36],s13[38],s12[40],s11[42],s10[44],s9[46],s8[48],s7[50],s6[52],s5[54],s4[56],s3[58],s2[60],s1[62],pp63[32],pp62[34],pp63[34]};
    CLA_68 KS_47(s47, c47, in47_1, in47_2);
    wire[65:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp30[1],pp32[0],s1[1],s2[1],s3[1],s4[1],s5[1],s6[1],s7[1],s8[1],s9[1],s10[1],s11[1],s12[1],s13[1],s14[1],s15[1],s16[1],s17[1],s18[1],s19[1],s20[1],s21[1],s22[1],s23[1],s24[1],s25[1],s26[1],s27[1],s28[1],s29[1],s30[1],s31[1],s31[2],s31[3],s30[5],s29[7],s28[9],s27[11],s26[13],s25[15],s24[17],s23[19],s22[21],s21[23],s20[25],s19[27],s18[29],s17[31],s16[33],s15[35],s14[37],s13[39],s12[41],s11[43],s10[45],s9[47],s8[49],s7[51],s6[53],s5[55],s4[57],s3[59],s2[61],s1[63],pp63[33]};
    assign in48_2 = {pp31[0],s1[0],s2[0],s3[0],s4[0],s5[0],s6[0],s7[0],s8[0],s9[0],s10[0],s11[0],s12[0],s13[0],s14[0],s15[0],s16[0],s17[0],s18[0],s19[0],s20[0],s21[0],s22[0],s23[0],s24[0],s25[0],s26[0],s27[0],s28[0],s29[0],s30[0],s31[0],s32[0],s32[1],c32,c31,c30,c29,c28,c27,c26,c25,c24,c23,c22,c21,c20,c19,c18,c17,c16,c15,c14,c13,c12,c11,c10,c9,c8,c7,c6,c5,c4,c3,c2,c1};
    CLA_66 KS_48(s48, c48, in48_1, in48_2);

    /*Stage 3*/
    wire[111:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp0[8],pp0[9],pp0[10],pp0[11],pp0[12],pp0[13],pp0[14],pp0[15],pp2[14],pp4[13],pp6[12],pp8[11],pp10[10],pp12[9],pp14[8],pp16[7],pp18[6],pp20[5],pp22[4],pp24[3],pp26[2],pp28[1],pp30[0],s33[15],s33[16],s33[17],s33[18],s33[19],s33[20],s33[21],s33[22],s33[23],s33[24],s33[25],s33[26],s33[27],s33[28],s33[29],s33[30],s33[31],s33[32],s33[33],s33[34],s33[35],s33[36],s33[37],s33[38],s33[39],s33[40],s33[41],s33[42],s33[43],s33[44],s33[45],s33[46],s33[47],s33[48],s33[49],s33[50],s33[51],s33[52],s33[53],s33[54],s33[55],s33[56],s33[57],s33[58],s33[59],s33[60],s33[61],s33[62],s33[63],s33[64],s33[65],s33[66],s33[67],s33[68],s33[69],s33[70],s33[71],s33[72],s33[73],s33[74],s33[75],s33[76],s33[77],s33[78],s33[79],s33[80],s33[81],pp63[35],pp62[37],pp61[39],pp60[41],pp59[43],pp58[45],pp57[47],pp56[49],pp55[51],pp54[53],pp53[55],pp52[57],pp51[59],pp50[61],pp49[63],pp50[63],pp51[63],pp52[63],pp53[63],pp54[63],pp55[63],pp56[63]};
    assign in49_2 = {pp1[7],pp1[8],pp1[9],pp1[10],pp1[11],pp1[12],pp1[13],pp1[14],pp3[13],pp5[12],pp7[11],pp9[10],pp11[9],pp13[8],pp15[7],pp17[6],pp19[5],pp21[4],pp23[3],pp25[2],pp27[1],pp29[0],s33[14],s34[14],s34[15],s34[16],s34[17],s34[18],s34[19],s34[20],s34[21],s34[22],s34[23],s34[24],s34[25],s34[26],s34[27],s34[28],s34[29],s34[30],s34[31],s34[32],s34[33],s34[34],s34[35],s34[36],s34[37],s34[38],s34[39],s34[40],s34[41],s34[42],s34[43],s34[44],s34[45],s34[46],s34[47],s34[48],s34[49],s34[50],s34[51],s34[52],s34[53],s34[54],s34[55],s34[56],s34[57],s34[58],s34[59],s34[60],s34[61],s34[62],s34[63],s34[64],s34[65],s34[66],s34[67],s34[68],s34[69],s34[70],s34[71],s34[72],s34[73],s34[74],s34[75],s34[76],s34[77],s34[78],s34[79],s34[80],s33[82],pp63[36],pp62[38],pp61[40],pp60[42],pp59[44],pp58[46],pp57[48],pp56[50],pp55[52],pp54[54],pp53[56],pp52[58],pp51[60],pp50[62],pp51[62],pp52[62],pp53[62],pp54[62],pp55[62],pp56[62],pp57[62]};
    CLA_112 KS_49(s49, c49, in49_1, in49_2);
    wire[109:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp2[7],pp2[8],pp2[9],pp2[10],pp2[11],pp2[12],pp2[13],pp4[12],pp6[11],pp8[10],pp10[9],pp12[8],pp14[7],pp16[6],pp18[5],pp20[4],pp22[3],pp24[2],pp26[1],pp28[0],s33[13],s34[13],s35[13],s35[14],s35[15],s35[16],s35[17],s35[18],s35[19],s35[20],s35[21],s35[22],s35[23],s35[24],s35[25],s35[26],s35[27],s35[28],s35[29],s35[30],s35[31],s35[32],s35[33],s35[34],s35[35],s35[36],s35[37],s35[38],s35[39],s35[40],s35[41],s35[42],s35[43],s35[44],s35[45],s35[46],s35[47],s35[48],s35[49],s35[50],s35[51],s35[52],s35[53],s35[54],s35[55],s35[56],s35[57],s35[58],s35[59],s35[60],s35[61],s35[62],s35[63],s35[64],s35[65],s35[66],s35[67],s35[68],s35[69],s35[70],s35[71],s35[72],s35[73],s35[74],s35[75],s35[76],s35[77],s35[78],s35[79],s34[81],s33[83],pp63[37],pp62[39],pp61[41],pp60[43],pp59[45],pp58[47],pp57[49],pp56[51],pp55[53],pp54[55],pp53[57],pp52[59],pp51[61],pp52[61],pp53[61],pp54[61],pp55[61],pp56[61],pp57[61]};
    assign in50_2 = {pp3[6],pp3[7],pp3[8],pp3[9],pp3[10],pp3[11],pp3[12],pp5[11],pp7[10],pp9[9],pp11[8],pp13[7],pp15[6],pp17[5],pp19[4],pp21[3],pp23[2],pp25[1],pp27[0],s33[12],s34[12],s35[12],s36[12],s36[13],s36[14],s36[15],s36[16],s36[17],s36[18],s36[19],s36[20],s36[21],s36[22],s36[23],s36[24],s36[25],s36[26],s36[27],s36[28],s36[29],s36[30],s36[31],s36[32],s36[33],s36[34],s36[35],s36[36],s36[37],s36[38],s36[39],s36[40],s36[41],s36[42],s36[43],s36[44],s36[45],s36[46],s36[47],s36[48],s36[49],s36[50],s36[51],s36[52],s36[53],s36[54],s36[55],s36[56],s36[57],s36[58],s36[59],s36[60],s36[61],s36[62],s36[63],s36[64],s36[65],s36[66],s36[67],s36[68],s36[69],s36[70],s36[71],s36[72],s36[73],s36[74],s36[75],s36[76],s36[77],s36[78],s35[80],s34[82],s33[84],pp63[38],pp62[40],pp61[42],pp60[44],pp59[46],pp58[48],pp57[50],pp56[52],pp55[54],pp54[56],pp53[58],pp52[60],pp53[60],pp54[60],pp55[60],pp56[60],pp57[60],pp58[60]};
    CLA_110 KS_50(s50, c50, in50_1, in50_2);
    wire[107:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp4[6],pp4[7],pp4[8],pp4[9],pp4[10],pp4[11],pp6[10],pp8[9],pp10[8],pp12[7],pp14[6],pp16[5],pp18[4],pp20[3],pp22[2],pp24[1],pp26[0],s33[11],s34[11],s35[11],s36[11],s37[11],s37[12],s37[13],s37[14],s37[15],s37[16],s37[17],s37[18],s37[19],s37[20],s37[21],s37[22],s37[23],s37[24],s37[25],s37[26],s37[27],s37[28],s37[29],s37[30],s37[31],s37[32],s37[33],s37[34],s37[35],s37[36],s37[37],s37[38],s37[39],s37[40],s37[41],s37[42],s37[43],s37[44],s37[45],s37[46],s37[47],s37[48],s37[49],s37[50],s37[51],s37[52],s37[53],s37[54],s37[55],s37[56],s37[57],s37[58],s37[59],s37[60],s37[61],s37[62],s37[63],s37[64],s37[65],s37[66],s37[67],s37[68],s37[69],s37[70],s37[71],s37[72],s37[73],s37[74],s37[75],s37[76],s37[77],s36[79],s35[81],s34[83],s33[85],pp63[39],pp62[41],pp61[43],pp60[45],pp59[47],pp58[49],pp57[51],pp56[53],pp55[55],pp54[57],pp53[59],pp54[59],pp55[59],pp56[59],pp57[59],pp58[59]};
    assign in51_2 = {pp5[5],pp5[6],pp5[7],pp5[8],pp5[9],pp5[10],pp7[9],pp9[8],pp11[7],pp13[6],pp15[5],pp17[4],pp19[3],pp21[2],pp23[1],pp25[0],s33[10],s34[10],s35[10],s36[10],s37[10],s38[10],s38[11],s38[12],s38[13],s38[14],s38[15],s38[16],s38[17],s38[18],s38[19],s38[20],s38[21],s38[22],s38[23],s38[24],s38[25],s38[26],s38[27],s38[28],s38[29],s38[30],s38[31],s38[32],s38[33],s38[34],s38[35],s38[36],s38[37],s38[38],s38[39],s38[40],s38[41],s38[42],s38[43],s38[44],s38[45],s38[46],s38[47],s38[48],s38[49],s38[50],s38[51],s38[52],s38[53],s38[54],s38[55],s38[56],s38[57],s38[58],s38[59],s38[60],s38[61],s38[62],s38[63],s38[64],s38[65],s38[66],s38[67],s38[68],s38[69],s38[70],s38[71],s38[72],s38[73],s38[74],s38[75],s38[76],s37[78],s36[80],s35[82],s34[84],s33[86],pp63[40],pp62[42],pp61[44],pp60[46],pp59[48],pp58[50],pp57[52],pp56[54],pp55[56],pp54[58],pp55[58],pp56[58],pp57[58],pp58[58],pp59[58]};
    CLA_108 KS_51(s51, c51, in51_1, in51_2);
    wire[105:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp6[5],pp6[6],pp6[7],pp6[8],pp6[9],pp8[8],pp10[7],pp12[6],pp14[5],pp16[4],pp18[3],pp20[2],pp22[1],pp24[0],s33[9],s34[9],s35[9],s36[9],s37[9],s38[9],s39[9],s39[10],s39[11],s39[12],s39[13],s39[14],s39[15],s39[16],s39[17],s39[18],s39[19],s39[20],s39[21],s39[22],s39[23],s39[24],s39[25],s39[26],s39[27],s39[28],s39[29],s39[30],s39[31],s39[32],s39[33],s39[34],s39[35],s39[36],s39[37],s39[38],s39[39],s39[40],s39[41],s39[42],s39[43],s39[44],s39[45],s39[46],s39[47],s39[48],s39[49],s39[50],s39[51],s39[52],s39[53],s39[54],s39[55],s39[56],s39[57],s39[58],s39[59],s39[60],s39[61],s39[62],s39[63],s39[64],s39[65],s39[66],s39[67],s39[68],s39[69],s39[70],s39[71],s39[72],s39[73],s39[74],s39[75],s38[77],s37[79],s36[81],s35[83],s34[85],s33[87],pp63[41],pp62[43],pp61[45],pp60[47],pp59[49],pp58[51],pp57[53],pp56[55],pp55[57],pp56[57],pp57[57],pp58[57],pp59[57]};
    assign in52_2 = {pp7[4],pp7[5],pp7[6],pp7[7],pp7[8],pp9[7],pp11[6],pp13[5],pp15[4],pp17[3],pp19[2],pp21[1],pp23[0],s33[8],s34[8],s35[8],s36[8],s37[8],s38[8],s39[8],s40[8],s40[9],s40[10],s40[11],s40[12],s40[13],s40[14],s40[15],s40[16],s40[17],s40[18],s40[19],s40[20],s40[21],s40[22],s40[23],s40[24],s40[25],s40[26],s40[27],s40[28],s40[29],s40[30],s40[31],s40[32],s40[33],s40[34],s40[35],s40[36],s40[37],s40[38],s40[39],s40[40],s40[41],s40[42],s40[43],s40[44],s40[45],s40[46],s40[47],s40[48],s40[49],s40[50],s40[51],s40[52],s40[53],s40[54],s40[55],s40[56],s40[57],s40[58],s40[59],s40[60],s40[61],s40[62],s40[63],s40[64],s40[65],s40[66],s40[67],s40[68],s40[69],s40[70],s40[71],s40[72],s40[73],s40[74],s39[76],s38[78],s37[80],s36[82],s35[84],s34[86],s33[88],pp63[42],pp62[44],pp61[46],pp60[48],pp59[50],pp58[52],pp57[54],pp56[56],pp57[56],pp58[56],pp59[56],pp60[56]};
    CLA_106 KS_52(s52, c52, in52_1, in52_2);
    wire[103:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp8[4],pp8[5],pp8[6],pp8[7],pp10[6],pp12[5],pp14[4],pp16[3],pp18[2],pp20[1],pp22[0],s33[7],s34[7],s35[7],s36[7],s37[7],s38[7],s39[7],s40[7],s41[7],s41[8],s41[9],s41[10],s41[11],s41[12],s41[13],s41[14],s41[15],s41[16],s41[17],s41[18],s41[19],s41[20],s41[21],s41[22],s41[23],s41[24],s41[25],s41[26],s41[27],s41[28],s41[29],s41[30],s41[31],s41[32],s41[33],s41[34],s41[35],s41[36],s41[37],s41[38],s41[39],s41[40],s41[41],s41[42],s41[43],s41[44],s41[45],s41[46],s41[47],s41[48],s41[49],s41[50],s41[51],s41[52],s41[53],s41[54],s41[55],s41[56],s41[57],s41[58],s41[59],s41[60],s41[61],s41[62],s41[63],s41[64],s41[65],s41[66],s41[67],s41[68],s41[69],s41[70],s41[71],s41[72],s41[73],s40[75],s39[77],s38[79],s37[81],s36[83],s35[85],s34[87],s33[89],pp63[43],pp62[45],pp61[47],pp60[49],pp59[51],pp58[53],pp57[55],pp58[55],pp59[55],pp60[55]};
    assign in53_2 = {pp9[3],pp9[4],pp9[5],pp9[6],pp11[5],pp13[4],pp15[3],pp17[2],pp19[1],pp21[0],s33[6],s34[6],s35[6],s36[6],s37[6],s38[6],s39[6],s40[6],s41[6],s42[6],s42[7],s42[8],s42[9],s42[10],s42[11],s42[12],s42[13],s42[14],s42[15],s42[16],s42[17],s42[18],s42[19],s42[20],s42[21],s42[22],s42[23],s42[24],s42[25],s42[26],s42[27],s42[28],s42[29],s42[30],s42[31],s42[32],s42[33],s42[34],s42[35],s42[36],s42[37],s42[38],s42[39],s42[40],s42[41],s42[42],s42[43],s42[44],s42[45],s42[46],s42[47],s42[48],s42[49],s42[50],s42[51],s42[52],s42[53],s42[54],s42[55],s42[56],s42[57],s42[58],s42[59],s42[60],s42[61],s42[62],s42[63],s42[64],s42[65],s42[66],s42[67],s42[68],s42[69],s42[70],s42[71],s42[72],s41[74],s40[76],s39[78],s38[80],s37[82],s36[84],s35[86],s34[88],s33[90],pp63[44],pp62[46],pp61[48],pp60[50],pp59[52],pp58[54],pp59[54],pp60[54],pp61[54]};
    CLA_104 KS_53(s53, c53, in53_1, in53_2);
    wire[101:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp10[3],pp10[4],pp10[5],pp12[4],pp14[3],pp16[2],pp18[1],pp20[0],s33[5],s34[5],s35[5],s36[5],s37[5],s38[5],s39[5],s40[5],s41[5],s42[5],s43[5],s43[6],s43[7],s43[8],s43[9],s43[10],s43[11],s43[12],s43[13],s43[14],s43[15],s43[16],s43[17],s43[18],s43[19],s43[20],s43[21],s43[22],s43[23],s43[24],s43[25],s43[26],s43[27],s43[28],s43[29],s43[30],s43[31],s43[32],s43[33],s43[34],s43[35],s43[36],s43[37],s43[38],s43[39],s43[40],s43[41],s43[42],s43[43],s43[44],s43[45],s43[46],s43[47],s43[48],s43[49],s43[50],s43[51],s43[52],s43[53],s43[54],s43[55],s43[56],s43[57],s43[58],s43[59],s43[60],s43[61],s43[62],s43[63],s43[64],s43[65],s43[66],s43[67],s43[68],s43[69],s43[70],s43[71],s42[73],s41[75],s40[77],s39[79],s38[81],s37[83],s36[85],s35[87],s34[89],s33[91],pp63[45],pp62[47],pp61[49],pp60[51],pp59[53],pp60[53],pp61[53]};
    assign in54_2 = {pp11[2],pp11[3],pp11[4],pp13[3],pp15[2],pp17[1],pp19[0],s33[4],s34[4],s35[4],s36[4],s37[4],s38[4],s39[4],s40[4],s41[4],s42[4],s43[4],s44[4],s44[5],s44[6],s44[7],s44[8],s44[9],s44[10],s44[11],s44[12],s44[13],s44[14],s44[15],s44[16],s44[17],s44[18],s44[19],s44[20],s44[21],s44[22],s44[23],s44[24],s44[25],s44[26],s44[27],s44[28],s44[29],s44[30],s44[31],s44[32],s44[33],s44[34],s44[35],s44[36],s44[37],s44[38],s44[39],s44[40],s44[41],s44[42],s44[43],s44[44],s44[45],s44[46],s44[47],s44[48],s44[49],s44[50],s44[51],s44[52],s44[53],s44[54],s44[55],s44[56],s44[57],s44[58],s44[59],s44[60],s44[61],s44[62],s44[63],s44[64],s44[65],s44[66],s44[67],s44[68],s44[69],s44[70],s43[72],s42[74],s41[76],s40[78],s39[80],s38[82],s37[84],s36[86],s35[88],s34[90],s33[92],pp63[46],pp62[48],pp61[50],pp60[52],pp61[52],pp62[52]};
    CLA_102 KS_54(s54, c54, in54_1, in54_2);
    wire[99:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp12[2],pp12[3],pp14[2],pp16[1],pp18[0],s33[3],s34[3],s35[3],s36[3],s37[3],s38[3],s39[3],s40[3],s41[3],s42[3],s43[3],s44[3],s45[3],s45[4],s45[5],s45[6],s45[7],s45[8],s45[9],s45[10],s45[11],s45[12],s45[13],s45[14],s45[15],s45[16],s45[17],s45[18],s45[19],s45[20],s45[21],s45[22],s45[23],s45[24],s45[25],s45[26],s45[27],s45[28],s45[29],s45[30],s45[31],s45[32],s45[33],s45[34],s45[35],s45[36],s45[37],s45[38],s45[39],s45[40],s45[41],s45[42],s45[43],s45[44],s45[45],s45[46],s45[47],s45[48],s45[49],s45[50],s45[51],s45[52],s45[53],s45[54],s45[55],s45[56],s45[57],s45[58],s45[59],s45[60],s45[61],s45[62],s45[63],s45[64],s45[65],s45[66],s45[67],s45[68],s45[69],s44[71],s43[73],s42[75],s41[77],s40[79],s39[81],s38[83],s37[85],s36[87],s35[89],s34[91],s33[93],pp63[47],pp62[49],pp61[51],pp62[51]};
    assign in55_2 = {pp13[1],pp13[2],pp15[1],pp17[0],s33[2],s34[2],s35[2],s36[2],s37[2],s38[2],s39[2],s40[2],s41[2],s42[2],s43[2],s44[2],s45[2],s46[2],s46[3],s46[4],s46[5],s46[6],s46[7],s46[8],s46[9],s46[10],s46[11],s46[12],s46[13],s46[14],s46[15],s46[16],s46[17],s46[18],s46[19],s46[20],s46[21],s46[22],s46[23],s46[24],s46[25],s46[26],s46[27],s46[28],s46[29],s46[30],s46[31],s46[32],s46[33],s46[34],s46[35],s46[36],s46[37],s46[38],s46[39],s46[40],s46[41],s46[42],s46[43],s46[44],s46[45],s46[46],s46[47],s46[48],s46[49],s46[50],s46[51],s46[52],s46[53],s46[54],s46[55],s46[56],s46[57],s46[58],s46[59],s46[60],s46[61],s46[62],s46[63],s46[64],s46[65],s46[66],s46[67],s46[68],s45[70],s44[72],s43[74],s42[76],s41[78],s40[80],s39[82],s38[84],s37[86],s36[88],s35[90],s34[92],s33[94],pp63[48],pp62[50],pp63[50]};
    CLA_100 KS_55(s55, c55, in55_1, in55_2);
    wire[97:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp14[1],pp16[0],s33[1],s34[1],s35[1],s36[1],s37[1],s38[1],s39[1],s40[1],s41[1],s42[1],s43[1],s44[1],s45[1],s46[1],s47[1],s47[2],s47[3],s47[4],s47[5],s47[6],s47[7],s47[8],s47[9],s47[10],s47[11],s47[12],s47[13],s47[14],s47[15],s47[16],s47[17],s47[18],s47[19],s47[20],s47[21],s47[22],s47[23],s47[24],s47[25],s47[26],s47[27],s47[28],s47[29],s47[30],s47[31],s47[32],s47[33],s47[34],s47[35],s47[36],s47[37],s47[38],s47[39],s47[40],s47[41],s47[42],s47[43],s47[44],s47[45],s47[46],s47[47],s47[48],s47[49],s47[50],s47[51],s47[52],s47[53],s47[54],s47[55],s47[56],s47[57],s47[58],s47[59],s47[60],s47[61],s47[62],s47[63],s47[64],s47[65],s47[66],s47[67],s46[69],s45[71],s44[73],s43[75],s42[77],s41[79],s40[81],s39[83],s38[85],s37[87],s36[89],s35[91],s34[93],s33[95],pp63[49]};
    assign in56_2 = {pp15[0],s33[0],s34[0],s35[0],s36[0],s37[0],s38[0],s39[0],s40[0],s41[0],s42[0],s43[0],s44[0],s45[0],s46[0],s47[0],s48[0],s48[1],s48[2],s48[3],s48[4],s48[5],s48[6],s48[7],s48[8],s48[9],s48[10],s48[11],s48[12],s48[13],s48[14],s48[15],s48[16],s48[17],s48[18],s48[19],s48[20],s48[21],s48[22],s48[23],s48[24],s48[25],s48[26],s48[27],s48[28],s48[29],s48[30],s48[31],s48[32],s48[33],s48[34],s48[35],s48[36],s48[37],s48[38],s48[39],s48[40],s48[41],s48[42],s48[43],s48[44],s48[45],s48[46],s48[47],s48[48],s48[49],s48[50],s48[51],s48[52],s48[53],s48[54],s48[55],s48[56],s48[57],s48[58],s48[59],s48[60],s48[61],s48[62],s48[63],s48[64],s48[65],c48,c47,c46,c45,c44,c43,c42,c41,c40,c39,c38,c37,c36,c35,c34,c33};
    CLA_98 KS_56(s56, c56, in56_1, in56_2);

    /*Stage 4*/
    wire[119:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp0[4],pp0[5],pp0[6],pp0[7],pp2[6],pp4[5],pp6[4],pp8[3],pp10[2],pp12[1],pp14[0],s49[7],s49[8],s49[9],s49[10],s49[11],s49[12],s49[13],s49[14],s49[15],s49[16],s49[17],s49[18],s49[19],s49[20],s49[21],s49[22],s49[23],s49[24],s49[25],s49[26],s49[27],s49[28],s49[29],s49[30],s49[31],s49[32],s49[33],s49[34],s49[35],s49[36],s49[37],s49[38],s49[39],s49[40],s49[41],s49[42],s49[43],s49[44],s49[45],s49[46],s49[47],s49[48],s49[49],s49[50],s49[51],s49[52],s49[53],s49[54],s49[55],s49[56],s49[57],s49[58],s49[59],s49[60],s49[61],s49[62],s49[63],s49[64],s49[65],s49[66],s49[67],s49[68],s49[69],s49[70],s49[71],s49[72],s49[73],s49[74],s49[75],s49[76],s49[77],s49[78],s49[79],s49[80],s49[81],s49[82],s49[83],s49[84],s49[85],s49[86],s49[87],s49[88],s49[89],s49[90],s49[91],s49[92],s49[93],s49[94],s49[95],s49[96],s49[97],s49[98],s49[99],s49[100],s49[101],s49[102],s49[103],s49[104],s49[105],pp63[51],pp62[53],pp61[55],pp60[57],pp59[59],pp58[61],pp57[63],pp58[63],pp59[63],pp60[63]};
    assign in57_2 = {pp1[3],pp1[4],pp1[5],pp1[6],pp3[5],pp5[4],pp7[3],pp9[2],pp11[1],pp13[0],s49[6],s50[6],s50[7],s50[8],s50[9],s50[10],s50[11],s50[12],s50[13],s50[14],s50[15],s50[16],s50[17],s50[18],s50[19],s50[20],s50[21],s50[22],s50[23],s50[24],s50[25],s50[26],s50[27],s50[28],s50[29],s50[30],s50[31],s50[32],s50[33],s50[34],s50[35],s50[36],s50[37],s50[38],s50[39],s50[40],s50[41],s50[42],s50[43],s50[44],s50[45],s50[46],s50[47],s50[48],s50[49],s50[50],s50[51],s50[52],s50[53],s50[54],s50[55],s50[56],s50[57],s50[58],s50[59],s50[60],s50[61],s50[62],s50[63],s50[64],s50[65],s50[66],s50[67],s50[68],s50[69],s50[70],s50[71],s50[72],s50[73],s50[74],s50[75],s50[76],s50[77],s50[78],s50[79],s50[80],s50[81],s50[82],s50[83],s50[84],s50[85],s50[86],s50[87],s50[88],s50[89],s50[90],s50[91],s50[92],s50[93],s50[94],s50[95],s50[96],s50[97],s50[98],s50[99],s50[100],s50[101],s50[102],s50[103],s50[104],s49[106],pp63[52],pp62[54],pp61[56],pp60[58],pp59[60],pp58[62],pp59[62],pp60[62],pp61[62]};
    CLA_120 KS_57(s57, c57, in57_1, in57_2);
    wire[117:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp2[3],pp2[4],pp2[5],pp4[4],pp6[3],pp8[2],pp10[1],pp12[0],s49[5],s50[5],s51[5],s51[6],s51[7],s51[8],s51[9],s51[10],s51[11],s51[12],s51[13],s51[14],s51[15],s51[16],s51[17],s51[18],s51[19],s51[20],s51[21],s51[22],s51[23],s51[24],s51[25],s51[26],s51[27],s51[28],s51[29],s51[30],s51[31],s51[32],s51[33],s51[34],s51[35],s51[36],s51[37],s51[38],s51[39],s51[40],s51[41],s51[42],s51[43],s51[44],s51[45],s51[46],s51[47],s51[48],s51[49],s51[50],s51[51],s51[52],s51[53],s51[54],s51[55],s51[56],s51[57],s51[58],s51[59],s51[60],s51[61],s51[62],s51[63],s51[64],s51[65],s51[66],s51[67],s51[68],s51[69],s51[70],s51[71],s51[72],s51[73],s51[74],s51[75],s51[76],s51[77],s51[78],s51[79],s51[80],s51[81],s51[82],s51[83],s51[84],s51[85],s51[86],s51[87],s51[88],s51[89],s51[90],s51[91],s51[92],s51[93],s51[94],s51[95],s51[96],s51[97],s51[98],s51[99],s51[100],s51[101],s51[102],s51[103],s50[105],s49[107],pp63[53],pp62[55],pp61[57],pp60[59],pp59[61],pp60[61],pp61[61]};
    assign in58_2 = {pp3[2],pp3[3],pp3[4],pp5[3],pp7[2],pp9[1],pp11[0],s49[4],s50[4],s51[4],s52[4],s52[5],s52[6],s52[7],s52[8],s52[9],s52[10],s52[11],s52[12],s52[13],s52[14],s52[15],s52[16],s52[17],s52[18],s52[19],s52[20],s52[21],s52[22],s52[23],s52[24],s52[25],s52[26],s52[27],s52[28],s52[29],s52[30],s52[31],s52[32],s52[33],s52[34],s52[35],s52[36],s52[37],s52[38],s52[39],s52[40],s52[41],s52[42],s52[43],s52[44],s52[45],s52[46],s52[47],s52[48],s52[49],s52[50],s52[51],s52[52],s52[53],s52[54],s52[55],s52[56],s52[57],s52[58],s52[59],s52[60],s52[61],s52[62],s52[63],s52[64],s52[65],s52[66],s52[67],s52[68],s52[69],s52[70],s52[71],s52[72],s52[73],s52[74],s52[75],s52[76],s52[77],s52[78],s52[79],s52[80],s52[81],s52[82],s52[83],s52[84],s52[85],s52[86],s52[87],s52[88],s52[89],s52[90],s52[91],s52[92],s52[93],s52[94],s52[95],s52[96],s52[97],s52[98],s52[99],s52[100],s52[101],s52[102],s51[104],s50[106],s49[108],pp63[54],pp62[56],pp61[58],pp60[60],pp61[60],pp62[60]};
    CLA_118 KS_58(s58, c58, in58_1, in58_2);
    wire[115:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp4[2],pp4[3],pp6[2],pp8[1],pp10[0],s49[3],s50[3],s51[3],s52[3],s53[3],s53[4],s53[5],s53[6],s53[7],s53[8],s53[9],s53[10],s53[11],s53[12],s53[13],s53[14],s53[15],s53[16],s53[17],s53[18],s53[19],s53[20],s53[21],s53[22],s53[23],s53[24],s53[25],s53[26],s53[27],s53[28],s53[29],s53[30],s53[31],s53[32],s53[33],s53[34],s53[35],s53[36],s53[37],s53[38],s53[39],s53[40],s53[41],s53[42],s53[43],s53[44],s53[45],s53[46],s53[47],s53[48],s53[49],s53[50],s53[51],s53[52],s53[53],s53[54],s53[55],s53[56],s53[57],s53[58],s53[59],s53[60],s53[61],s53[62],s53[63],s53[64],s53[65],s53[66],s53[67],s53[68],s53[69],s53[70],s53[71],s53[72],s53[73],s53[74],s53[75],s53[76],s53[77],s53[78],s53[79],s53[80],s53[81],s53[82],s53[83],s53[84],s53[85],s53[86],s53[87],s53[88],s53[89],s53[90],s53[91],s53[92],s53[93],s53[94],s53[95],s53[96],s53[97],s53[98],s53[99],s53[100],s53[101],s52[103],s51[105],s50[107],s49[109],pp63[55],pp62[57],pp61[59],pp62[59]};
    assign in59_2 = {pp5[1],pp5[2],pp7[1],pp9[0],s49[2],s50[2],s51[2],s52[2],s53[2],s54[2],s54[3],s54[4],s54[5],s54[6],s54[7],s54[8],s54[9],s54[10],s54[11],s54[12],s54[13],s54[14],s54[15],s54[16],s54[17],s54[18],s54[19],s54[20],s54[21],s54[22],s54[23],s54[24],s54[25],s54[26],s54[27],s54[28],s54[29],s54[30],s54[31],s54[32],s54[33],s54[34],s54[35],s54[36],s54[37],s54[38],s54[39],s54[40],s54[41],s54[42],s54[43],s54[44],s54[45],s54[46],s54[47],s54[48],s54[49],s54[50],s54[51],s54[52],s54[53],s54[54],s54[55],s54[56],s54[57],s54[58],s54[59],s54[60],s54[61],s54[62],s54[63],s54[64],s54[65],s54[66],s54[67],s54[68],s54[69],s54[70],s54[71],s54[72],s54[73],s54[74],s54[75],s54[76],s54[77],s54[78],s54[79],s54[80],s54[81],s54[82],s54[83],s54[84],s54[85],s54[86],s54[87],s54[88],s54[89],s54[90],s54[91],s54[92],s54[93],s54[94],s54[95],s54[96],s54[97],s54[98],s54[99],s54[100],s53[102],s52[104],s51[106],s50[108],s49[110],pp63[56],pp62[58],pp63[58]};
    CLA_116 KS_59(s59, c59, in59_1, in59_2);
    wire[113:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp6[1],pp8[0],s49[1],s50[1],s51[1],s52[1],s53[1],s54[1],s55[1],s55[2],s55[3],s55[4],s55[5],s55[6],s55[7],s55[8],s55[9],s55[10],s55[11],s55[12],s55[13],s55[14],s55[15],s55[16],s55[17],s55[18],s55[19],s55[20],s55[21],s55[22],s55[23],s55[24],s55[25],s55[26],s55[27],s55[28],s55[29],s55[30],s55[31],s55[32],s55[33],s55[34],s55[35],s55[36],s55[37],s55[38],s55[39],s55[40],s55[41],s55[42],s55[43],s55[44],s55[45],s55[46],s55[47],s55[48],s55[49],s55[50],s55[51],s55[52],s55[53],s55[54],s55[55],s55[56],s55[57],s55[58],s55[59],s55[60],s55[61],s55[62],s55[63],s55[64],s55[65],s55[66],s55[67],s55[68],s55[69],s55[70],s55[71],s55[72],s55[73],s55[74],s55[75],s55[76],s55[77],s55[78],s55[79],s55[80],s55[81],s55[82],s55[83],s55[84],s55[85],s55[86],s55[87],s55[88],s55[89],s55[90],s55[91],s55[92],s55[93],s55[94],s55[95],s55[96],s55[97],s55[98],s55[99],s54[101],s53[103],s52[105],s51[107],s50[109],s49[111],pp63[57]};
    assign in60_2 = {pp7[0],s49[0],s50[0],s51[0],s52[0],s53[0],s54[0],s55[0],s56[0],s56[1],s56[2],s56[3],s56[4],s56[5],s56[6],s56[7],s56[8],s56[9],s56[10],s56[11],s56[12],s56[13],s56[14],s56[15],s56[16],s56[17],s56[18],s56[19],s56[20],s56[21],s56[22],s56[23],s56[24],s56[25],s56[26],s56[27],s56[28],s56[29],s56[30],s56[31],s56[32],s56[33],s56[34],s56[35],s56[36],s56[37],s56[38],s56[39],s56[40],s56[41],s56[42],s56[43],s56[44],s56[45],s56[46],s56[47],s56[48],s56[49],s56[50],s56[51],s56[52],s56[53],s56[54],s56[55],s56[56],s56[57],s56[58],s56[59],s56[60],s56[61],s56[62],s56[63],s56[64],s56[65],s56[66],s56[67],s56[68],s56[69],s56[70],s56[71],s56[72],s56[73],s56[74],s56[75],s56[76],s56[77],s56[78],s56[79],s56[80],s56[81],s56[82],s56[83],s56[84],s56[85],s56[86],s56[87],s56[88],s56[89],s56[90],s56[91],s56[92],s56[93],s56[94],s56[95],s56[96],s56[97],c56,c55,c54,c53,c52,c51,c50,c49};
    CLA_114 KS_60(s60, c60, in60_1, in60_2);

    /*Stage 5*/
    wire[123:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp0[2],pp0[3],pp2[2],pp4[1],pp6[0],s57[3],s57[4],s57[5],s57[6],s57[7],s57[8],s57[9],s57[10],s57[11],s57[12],s57[13],s57[14],s57[15],s57[16],s57[17],s57[18],s57[19],s57[20],s57[21],s57[22],s57[23],s57[24],s57[25],s57[26],s57[27],s57[28],s57[29],s57[30],s57[31],s57[32],s57[33],s57[34],s57[35],s57[36],s57[37],s57[38],s57[39],s57[40],s57[41],s57[42],s57[43],s57[44],s57[45],s57[46],s57[47],s57[48],s57[49],s57[50],s57[51],s57[52],s57[53],s57[54],s57[55],s57[56],s57[57],s57[58],s57[59],s57[60],s57[61],s57[62],s57[63],s57[64],s57[65],s57[66],s57[67],s57[68],s57[69],s57[70],s57[71],s57[72],s57[73],s57[74],s57[75],s57[76],s57[77],s57[78],s57[79],s57[80],s57[81],s57[82],s57[83],s57[84],s57[85],s57[86],s57[87],s57[88],s57[89],s57[90],s57[91],s57[92],s57[93],s57[94],s57[95],s57[96],s57[97],s57[98],s57[99],s57[100],s57[101],s57[102],s57[103],s57[104],s57[105],s57[106],s57[107],s57[108],s57[109],s57[110],s57[111],s57[112],s57[113],s57[114],s57[115],s57[116],s57[117],pp63[59],pp62[61],pp61[63],pp62[63]};
    assign in61_2 = {pp1[1],pp1[2],pp3[1],pp5[0],s57[2],s58[2],s58[3],s58[4],s58[5],s58[6],s58[7],s58[8],s58[9],s58[10],s58[11],s58[12],s58[13],s58[14],s58[15],s58[16],s58[17],s58[18],s58[19],s58[20],s58[21],s58[22],s58[23],s58[24],s58[25],s58[26],s58[27],s58[28],s58[29],s58[30],s58[31],s58[32],s58[33],s58[34],s58[35],s58[36],s58[37],s58[38],s58[39],s58[40],s58[41],s58[42],s58[43],s58[44],s58[45],s58[46],s58[47],s58[48],s58[49],s58[50],s58[51],s58[52],s58[53],s58[54],s58[55],s58[56],s58[57],s58[58],s58[59],s58[60],s58[61],s58[62],s58[63],s58[64],s58[65],s58[66],s58[67],s58[68],s58[69],s58[70],s58[71],s58[72],s58[73],s58[74],s58[75],s58[76],s58[77],s58[78],s58[79],s58[80],s58[81],s58[82],s58[83],s58[84],s58[85],s58[86],s58[87],s58[88],s58[89],s58[90],s58[91],s58[92],s58[93],s58[94],s58[95],s58[96],s58[97],s58[98],s58[99],s58[100],s58[101],s58[102],s58[103],s58[104],s58[105],s58[106],s58[107],s58[108],s58[109],s58[110],s58[111],s58[112],s58[113],s58[114],s58[115],s58[116],s57[118],pp63[60],pp62[62],pp63[62]};
    CLA_124 KS_61(s61, c61, in61_1, in61_2);
    wire[121:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp2[1],pp4[0],s57[1],s58[1],s59[1],s59[2],s59[3],s59[4],s59[5],s59[6],s59[7],s59[8],s59[9],s59[10],s59[11],s59[12],s59[13],s59[14],s59[15],s59[16],s59[17],s59[18],s59[19],s59[20],s59[21],s59[22],s59[23],s59[24],s59[25],s59[26],s59[27],s59[28],s59[29],s59[30],s59[31],s59[32],s59[33],s59[34],s59[35],s59[36],s59[37],s59[38],s59[39],s59[40],s59[41],s59[42],s59[43],s59[44],s59[45],s59[46],s59[47],s59[48],s59[49],s59[50],s59[51],s59[52],s59[53],s59[54],s59[55],s59[56],s59[57],s59[58],s59[59],s59[60],s59[61],s59[62],s59[63],s59[64],s59[65],s59[66],s59[67],s59[68],s59[69],s59[70],s59[71],s59[72],s59[73],s59[74],s59[75],s59[76],s59[77],s59[78],s59[79],s59[80],s59[81],s59[82],s59[83],s59[84],s59[85],s59[86],s59[87],s59[88],s59[89],s59[90],s59[91],s59[92],s59[93],s59[94],s59[95],s59[96],s59[97],s59[98],s59[99],s59[100],s59[101],s59[102],s59[103],s59[104],s59[105],s59[106],s59[107],s59[108],s59[109],s59[110],s59[111],s59[112],s59[113],s59[114],s59[115],s58[117],s57[119],pp63[61]};
    assign in62_2 = {pp3[0],s57[0],s58[0],s59[0],s60[0],s60[1],s60[2],s60[3],s60[4],s60[5],s60[6],s60[7],s60[8],s60[9],s60[10],s60[11],s60[12],s60[13],s60[14],s60[15],s60[16],s60[17],s60[18],s60[19],s60[20],s60[21],s60[22],s60[23],s60[24],s60[25],s60[26],s60[27],s60[28],s60[29],s60[30],s60[31],s60[32],s60[33],s60[34],s60[35],s60[36],s60[37],s60[38],s60[39],s60[40],s60[41],s60[42],s60[43],s60[44],s60[45],s60[46],s60[47],s60[48],s60[49],s60[50],s60[51],s60[52],s60[53],s60[54],s60[55],s60[56],s60[57],s60[58],s60[59],s60[60],s60[61],s60[62],s60[63],s60[64],s60[65],s60[66],s60[67],s60[68],s60[69],s60[70],s60[71],s60[72],s60[73],s60[74],s60[75],s60[76],s60[77],s60[78],s60[79],s60[80],s60[81],s60[82],s60[83],s60[84],s60[85],s60[86],s60[87],s60[88],s60[89],s60[90],s60[91],s60[92],s60[93],s60[94],s60[95],s60[96],s60[97],s60[98],s60[99],s60[100],s60[101],s60[102],s60[103],s60[104],s60[105],s60[106],s60[107],s60[108],s60[109],s60[110],s60[111],s60[112],s60[113],c60,c59,c58,c57};
    CLA_122 KS_62(s62, c62, in62_1, in62_2);


    /*Final Stage 5*/
    wire[125:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],s61[1],s61[2],s61[3],s61[4],s61[5],s61[6],s61[7],s61[8],s61[9],s61[10],s61[11],s61[12],s61[13],s61[14],s61[15],s61[16],s61[17],s61[18],s61[19],s61[20],s61[21],s61[22],s61[23],s61[24],s61[25],s61[26],s61[27],s61[28],s61[29],s61[30],s61[31],s61[32],s61[33],s61[34],s61[35],s61[36],s61[37],s61[38],s61[39],s61[40],s61[41],s61[42],s61[43],s61[44],s61[45],s61[46],s61[47],s61[48],s61[49],s61[50],s61[51],s61[52],s61[53],s61[54],s61[55],s61[56],s61[57],s61[58],s61[59],s61[60],s61[61],s61[62],s61[63],s61[64],s61[65],s61[66],s61[67],s61[68],s61[69],s61[70],s61[71],s61[72],s61[73],s61[74],s61[75],s61[76],s61[77],s61[78],s61[79],s61[80],s61[81],s61[82],s61[83],s61[84],s61[85],s61[86],s61[87],s61[88],s61[89],s61[90],s61[91],s61[92],s61[93],s61[94],s61[95],s61[96],s61[97],s61[98],s61[99],s61[100],s61[101],s61[102],s61[103],s61[104],s61[105],s61[106],s61[107],s61[108],s61[109],s61[110],s61[111],s61[112],s61[113],s61[114],s61[115],s61[116],s61[117],s61[118],s61[119],s61[120],s61[121],s61[122],s61[123],pp63[63]};
    assign in_2 = {pp1[0],s61[0],s62[0],s62[1],s62[2],s62[3],s62[4],s62[5],s62[6],s62[7],s62[8],s62[9],s62[10],s62[11],s62[12],s62[13],s62[14],s62[15],s62[16],s62[17],s62[18],s62[19],s62[20],s62[21],s62[22],s62[23],s62[24],s62[25],s62[26],s62[27],s62[28],s62[29],s62[30],s62[31],s62[32],s62[33],s62[34],s62[35],s62[36],s62[37],s62[38],s62[39],s62[40],s62[41],s62[42],s62[43],s62[44],s62[45],s62[46],s62[47],s62[48],s62[49],s62[50],s62[51],s62[52],s62[53],s62[54],s62[55],s62[56],s62[57],s62[58],s62[59],s62[60],s62[61],s62[62],s62[63],s62[64],s62[65],s62[66],s62[67],s62[68],s62[69],s62[70],s62[71],s62[72],s62[73],s62[74],s62[75],s62[76],s62[77],s62[78],s62[79],s62[80],s62[81],s62[82],s62[83],s62[84],s62[85],s62[86],s62[87],s62[88],s62[89],s62[90],s62[91],s62[92],s62[93],s62[94],s62[95],s62[96],s62[97],s62[98],s62[99],s62[100],s62[101],s62[102],s62[103],s62[104],s62[105],s62[106],s62[107],s62[108],s62[109],s62[110],s62[111],s62[112],s62[113],s62[114],s62[115],s62[116],s62[117],s62[118],s62[119],s62[120],s62[121],c62,c61};
    CLA_126(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = c;
endmodule

module CLA_128(output [127:0] sum, output cout, input [127:0] in1, input [127:0] in2);

    wire[127:0] G;
    wire[127:0] C;
    wire[127:0] P;

    assign G[0] = in1[127] & in2[127];
    assign P[0] = in1[127] ^ in2[127];
    assign G[1] = in1[126] & in2[126];
    assign P[1] = in1[126] ^ in2[126];
    assign G[2] = in1[125] & in2[125];
    assign P[2] = in1[125] ^ in2[125];
    assign G[3] = in1[124] & in2[124];
    assign P[3] = in1[124] ^ in2[124];
    assign G[4] = in1[123] & in2[123];
    assign P[4] = in1[123] ^ in2[123];
    assign G[5] = in1[122] & in2[122];
    assign P[5] = in1[122] ^ in2[122];
    assign G[6] = in1[121] & in2[121];
    assign P[6] = in1[121] ^ in2[121];
    assign G[7] = in1[120] & in2[120];
    assign P[7] = in1[120] ^ in2[120];
    assign G[8] = in1[119] & in2[119];
    assign P[8] = in1[119] ^ in2[119];
    assign G[9] = in1[118] & in2[118];
    assign P[9] = in1[118] ^ in2[118];
    assign G[10] = in1[117] & in2[117];
    assign P[10] = in1[117] ^ in2[117];
    assign G[11] = in1[116] & in2[116];
    assign P[11] = in1[116] ^ in2[116];
    assign G[12] = in1[115] & in2[115];
    assign P[12] = in1[115] ^ in2[115];
    assign G[13] = in1[114] & in2[114];
    assign P[13] = in1[114] ^ in2[114];
    assign G[14] = in1[113] & in2[113];
    assign P[14] = in1[113] ^ in2[113];
    assign G[15] = in1[112] & in2[112];
    assign P[15] = in1[112] ^ in2[112];
    assign G[16] = in1[111] & in2[111];
    assign P[16] = in1[111] ^ in2[111];
    assign G[17] = in1[110] & in2[110];
    assign P[17] = in1[110] ^ in2[110];
    assign G[18] = in1[109] & in2[109];
    assign P[18] = in1[109] ^ in2[109];
    assign G[19] = in1[108] & in2[108];
    assign P[19] = in1[108] ^ in2[108];
    assign G[20] = in1[107] & in2[107];
    assign P[20] = in1[107] ^ in2[107];
    assign G[21] = in1[106] & in2[106];
    assign P[21] = in1[106] ^ in2[106];
    assign G[22] = in1[105] & in2[105];
    assign P[22] = in1[105] ^ in2[105];
    assign G[23] = in1[104] & in2[104];
    assign P[23] = in1[104] ^ in2[104];
    assign G[24] = in1[103] & in2[103];
    assign P[24] = in1[103] ^ in2[103];
    assign G[25] = in1[102] & in2[102];
    assign P[25] = in1[102] ^ in2[102];
    assign G[26] = in1[101] & in2[101];
    assign P[26] = in1[101] ^ in2[101];
    assign G[27] = in1[100] & in2[100];
    assign P[27] = in1[100] ^ in2[100];
    assign G[28] = in1[99] & in2[99];
    assign P[28] = in1[99] ^ in2[99];
    assign G[29] = in1[98] & in2[98];
    assign P[29] = in1[98] ^ in2[98];
    assign G[30] = in1[97] & in2[97];
    assign P[30] = in1[97] ^ in2[97];
    assign G[31] = in1[96] & in2[96];
    assign P[31] = in1[96] ^ in2[96];
    assign G[32] = in1[95] & in2[95];
    assign P[32] = in1[95] ^ in2[95];
    assign G[33] = in1[94] & in2[94];
    assign P[33] = in1[94] ^ in2[94];
    assign G[34] = in1[93] & in2[93];
    assign P[34] = in1[93] ^ in2[93];
    assign G[35] = in1[92] & in2[92];
    assign P[35] = in1[92] ^ in2[92];
    assign G[36] = in1[91] & in2[91];
    assign P[36] = in1[91] ^ in2[91];
    assign G[37] = in1[90] & in2[90];
    assign P[37] = in1[90] ^ in2[90];
    assign G[38] = in1[89] & in2[89];
    assign P[38] = in1[89] ^ in2[89];
    assign G[39] = in1[88] & in2[88];
    assign P[39] = in1[88] ^ in2[88];
    assign G[40] = in1[87] & in2[87];
    assign P[40] = in1[87] ^ in2[87];
    assign G[41] = in1[86] & in2[86];
    assign P[41] = in1[86] ^ in2[86];
    assign G[42] = in1[85] & in2[85];
    assign P[42] = in1[85] ^ in2[85];
    assign G[43] = in1[84] & in2[84];
    assign P[43] = in1[84] ^ in2[84];
    assign G[44] = in1[83] & in2[83];
    assign P[44] = in1[83] ^ in2[83];
    assign G[45] = in1[82] & in2[82];
    assign P[45] = in1[82] ^ in2[82];
    assign G[46] = in1[81] & in2[81];
    assign P[46] = in1[81] ^ in2[81];
    assign G[47] = in1[80] & in2[80];
    assign P[47] = in1[80] ^ in2[80];
    assign G[48] = in1[79] & in2[79];
    assign P[48] = in1[79] ^ in2[79];
    assign G[49] = in1[78] & in2[78];
    assign P[49] = in1[78] ^ in2[78];
    assign G[50] = in1[77] & in2[77];
    assign P[50] = in1[77] ^ in2[77];
    assign G[51] = in1[76] & in2[76];
    assign P[51] = in1[76] ^ in2[76];
    assign G[52] = in1[75] & in2[75];
    assign P[52] = in1[75] ^ in2[75];
    assign G[53] = in1[74] & in2[74];
    assign P[53] = in1[74] ^ in2[74];
    assign G[54] = in1[73] & in2[73];
    assign P[54] = in1[73] ^ in2[73];
    assign G[55] = in1[72] & in2[72];
    assign P[55] = in1[72] ^ in2[72];
    assign G[56] = in1[71] & in2[71];
    assign P[56] = in1[71] ^ in2[71];
    assign G[57] = in1[70] & in2[70];
    assign P[57] = in1[70] ^ in2[70];
    assign G[58] = in1[69] & in2[69];
    assign P[58] = in1[69] ^ in2[69];
    assign G[59] = in1[68] & in2[68];
    assign P[59] = in1[68] ^ in2[68];
    assign G[60] = in1[67] & in2[67];
    assign P[60] = in1[67] ^ in2[67];
    assign G[61] = in1[66] & in2[66];
    assign P[61] = in1[66] ^ in2[66];
    assign G[62] = in1[65] & in2[65];
    assign P[62] = in1[65] ^ in2[65];
    assign G[63] = in1[64] & in2[64];
    assign P[63] = in1[64] ^ in2[64];
    assign G[64] = in1[63] & in2[63];
    assign P[64] = in1[63] ^ in2[63];
    assign G[65] = in1[62] & in2[62];
    assign P[65] = in1[62] ^ in2[62];
    assign G[66] = in1[61] & in2[61];
    assign P[66] = in1[61] ^ in2[61];
    assign G[67] = in1[60] & in2[60];
    assign P[67] = in1[60] ^ in2[60];
    assign G[68] = in1[59] & in2[59];
    assign P[68] = in1[59] ^ in2[59];
    assign G[69] = in1[58] & in2[58];
    assign P[69] = in1[58] ^ in2[58];
    assign G[70] = in1[57] & in2[57];
    assign P[70] = in1[57] ^ in2[57];
    assign G[71] = in1[56] & in2[56];
    assign P[71] = in1[56] ^ in2[56];
    assign G[72] = in1[55] & in2[55];
    assign P[72] = in1[55] ^ in2[55];
    assign G[73] = in1[54] & in2[54];
    assign P[73] = in1[54] ^ in2[54];
    assign G[74] = in1[53] & in2[53];
    assign P[74] = in1[53] ^ in2[53];
    assign G[75] = in1[52] & in2[52];
    assign P[75] = in1[52] ^ in2[52];
    assign G[76] = in1[51] & in2[51];
    assign P[76] = in1[51] ^ in2[51];
    assign G[77] = in1[50] & in2[50];
    assign P[77] = in1[50] ^ in2[50];
    assign G[78] = in1[49] & in2[49];
    assign P[78] = in1[49] ^ in2[49];
    assign G[79] = in1[48] & in2[48];
    assign P[79] = in1[48] ^ in2[48];
    assign G[80] = in1[47] & in2[47];
    assign P[80] = in1[47] ^ in2[47];
    assign G[81] = in1[46] & in2[46];
    assign P[81] = in1[46] ^ in2[46];
    assign G[82] = in1[45] & in2[45];
    assign P[82] = in1[45] ^ in2[45];
    assign G[83] = in1[44] & in2[44];
    assign P[83] = in1[44] ^ in2[44];
    assign G[84] = in1[43] & in2[43];
    assign P[84] = in1[43] ^ in2[43];
    assign G[85] = in1[42] & in2[42];
    assign P[85] = in1[42] ^ in2[42];
    assign G[86] = in1[41] & in2[41];
    assign P[86] = in1[41] ^ in2[41];
    assign G[87] = in1[40] & in2[40];
    assign P[87] = in1[40] ^ in2[40];
    assign G[88] = in1[39] & in2[39];
    assign P[88] = in1[39] ^ in2[39];
    assign G[89] = in1[38] & in2[38];
    assign P[89] = in1[38] ^ in2[38];
    assign G[90] = in1[37] & in2[37];
    assign P[90] = in1[37] ^ in2[37];
    assign G[91] = in1[36] & in2[36];
    assign P[91] = in1[36] ^ in2[36];
    assign G[92] = in1[35] & in2[35];
    assign P[92] = in1[35] ^ in2[35];
    assign G[93] = in1[34] & in2[34];
    assign P[93] = in1[34] ^ in2[34];
    assign G[94] = in1[33] & in2[33];
    assign P[94] = in1[33] ^ in2[33];
    assign G[95] = in1[32] & in2[32];
    assign P[95] = in1[32] ^ in2[32];
    assign G[96] = in1[31] & in2[31];
    assign P[96] = in1[31] ^ in2[31];
    assign G[97] = in1[30] & in2[30];
    assign P[97] = in1[30] ^ in2[30];
    assign G[98] = in1[29] & in2[29];
    assign P[98] = in1[29] ^ in2[29];
    assign G[99] = in1[28] & in2[28];
    assign P[99] = in1[28] ^ in2[28];
    assign G[100] = in1[27] & in2[27];
    assign P[100] = in1[27] ^ in2[27];
    assign G[101] = in1[26] & in2[26];
    assign P[101] = in1[26] ^ in2[26];
    assign G[102] = in1[25] & in2[25];
    assign P[102] = in1[25] ^ in2[25];
    assign G[103] = in1[24] & in2[24];
    assign P[103] = in1[24] ^ in2[24];
    assign G[104] = in1[23] & in2[23];
    assign P[104] = in1[23] ^ in2[23];
    assign G[105] = in1[22] & in2[22];
    assign P[105] = in1[22] ^ in2[22];
    assign G[106] = in1[21] & in2[21];
    assign P[106] = in1[21] ^ in2[21];
    assign G[107] = in1[20] & in2[20];
    assign P[107] = in1[20] ^ in2[20];
    assign G[108] = in1[19] & in2[19];
    assign P[108] = in1[19] ^ in2[19];
    assign G[109] = in1[18] & in2[18];
    assign P[109] = in1[18] ^ in2[18];
    assign G[110] = in1[17] & in2[17];
    assign P[110] = in1[17] ^ in2[17];
    assign G[111] = in1[16] & in2[16];
    assign P[111] = in1[16] ^ in2[16];
    assign G[112] = in1[15] & in2[15];
    assign P[112] = in1[15] ^ in2[15];
    assign G[113] = in1[14] & in2[14];
    assign P[113] = in1[14] ^ in2[14];
    assign G[114] = in1[13] & in2[13];
    assign P[114] = in1[13] ^ in2[13];
    assign G[115] = in1[12] & in2[12];
    assign P[115] = in1[12] ^ in2[12];
    assign G[116] = in1[11] & in2[11];
    assign P[116] = in1[11] ^ in2[11];
    assign G[117] = in1[10] & in2[10];
    assign P[117] = in1[10] ^ in2[10];
    assign G[118] = in1[9] & in2[9];
    assign P[118] = in1[9] ^ in2[9];
    assign G[119] = in1[8] & in2[8];
    assign P[119] = in1[8] ^ in2[8];
    assign G[120] = in1[7] & in2[7];
    assign P[120] = in1[7] ^ in2[7];
    assign G[121] = in1[6] & in2[6];
    assign P[121] = in1[6] ^ in2[6];
    assign G[122] = in1[5] & in2[5];
    assign P[122] = in1[5] ^ in2[5];
    assign G[123] = in1[4] & in2[4];
    assign P[123] = in1[4] ^ in2[4];
    assign G[124] = in1[3] & in2[3];
    assign P[124] = in1[3] ^ in2[3];
    assign G[125] = in1[2] & in2[2];
    assign P[125] = in1[2] ^ in2[2];
    assign G[126] = in1[1] & in2[1];
    assign P[126] = in1[1] ^ in2[1];
    assign G[127] = in1[0] & in2[0];
    assign P[127] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign cout = G[127] | (P[127] & C[127]);
    assign sum = P ^ C;
endmodule

module CLA_127(output [126:0] sum, output cout, input [126:0] in1, input [126:0] in2);

    wire[126:0] G;
    wire[126:0] C;
    wire[126:0] P;

    assign G[0] = in1[126] & in2[126];
    assign P[0] = in1[126] ^ in2[126];
    assign G[1] = in1[125] & in2[125];
    assign P[1] = in1[125] ^ in2[125];
    assign G[2] = in1[124] & in2[124];
    assign P[2] = in1[124] ^ in2[124];
    assign G[3] = in1[123] & in2[123];
    assign P[3] = in1[123] ^ in2[123];
    assign G[4] = in1[122] & in2[122];
    assign P[4] = in1[122] ^ in2[122];
    assign G[5] = in1[121] & in2[121];
    assign P[5] = in1[121] ^ in2[121];
    assign G[6] = in1[120] & in2[120];
    assign P[6] = in1[120] ^ in2[120];
    assign G[7] = in1[119] & in2[119];
    assign P[7] = in1[119] ^ in2[119];
    assign G[8] = in1[118] & in2[118];
    assign P[8] = in1[118] ^ in2[118];
    assign G[9] = in1[117] & in2[117];
    assign P[9] = in1[117] ^ in2[117];
    assign G[10] = in1[116] & in2[116];
    assign P[10] = in1[116] ^ in2[116];
    assign G[11] = in1[115] & in2[115];
    assign P[11] = in1[115] ^ in2[115];
    assign G[12] = in1[114] & in2[114];
    assign P[12] = in1[114] ^ in2[114];
    assign G[13] = in1[113] & in2[113];
    assign P[13] = in1[113] ^ in2[113];
    assign G[14] = in1[112] & in2[112];
    assign P[14] = in1[112] ^ in2[112];
    assign G[15] = in1[111] & in2[111];
    assign P[15] = in1[111] ^ in2[111];
    assign G[16] = in1[110] & in2[110];
    assign P[16] = in1[110] ^ in2[110];
    assign G[17] = in1[109] & in2[109];
    assign P[17] = in1[109] ^ in2[109];
    assign G[18] = in1[108] & in2[108];
    assign P[18] = in1[108] ^ in2[108];
    assign G[19] = in1[107] & in2[107];
    assign P[19] = in1[107] ^ in2[107];
    assign G[20] = in1[106] & in2[106];
    assign P[20] = in1[106] ^ in2[106];
    assign G[21] = in1[105] & in2[105];
    assign P[21] = in1[105] ^ in2[105];
    assign G[22] = in1[104] & in2[104];
    assign P[22] = in1[104] ^ in2[104];
    assign G[23] = in1[103] & in2[103];
    assign P[23] = in1[103] ^ in2[103];
    assign G[24] = in1[102] & in2[102];
    assign P[24] = in1[102] ^ in2[102];
    assign G[25] = in1[101] & in2[101];
    assign P[25] = in1[101] ^ in2[101];
    assign G[26] = in1[100] & in2[100];
    assign P[26] = in1[100] ^ in2[100];
    assign G[27] = in1[99] & in2[99];
    assign P[27] = in1[99] ^ in2[99];
    assign G[28] = in1[98] & in2[98];
    assign P[28] = in1[98] ^ in2[98];
    assign G[29] = in1[97] & in2[97];
    assign P[29] = in1[97] ^ in2[97];
    assign G[30] = in1[96] & in2[96];
    assign P[30] = in1[96] ^ in2[96];
    assign G[31] = in1[95] & in2[95];
    assign P[31] = in1[95] ^ in2[95];
    assign G[32] = in1[94] & in2[94];
    assign P[32] = in1[94] ^ in2[94];
    assign G[33] = in1[93] & in2[93];
    assign P[33] = in1[93] ^ in2[93];
    assign G[34] = in1[92] & in2[92];
    assign P[34] = in1[92] ^ in2[92];
    assign G[35] = in1[91] & in2[91];
    assign P[35] = in1[91] ^ in2[91];
    assign G[36] = in1[90] & in2[90];
    assign P[36] = in1[90] ^ in2[90];
    assign G[37] = in1[89] & in2[89];
    assign P[37] = in1[89] ^ in2[89];
    assign G[38] = in1[88] & in2[88];
    assign P[38] = in1[88] ^ in2[88];
    assign G[39] = in1[87] & in2[87];
    assign P[39] = in1[87] ^ in2[87];
    assign G[40] = in1[86] & in2[86];
    assign P[40] = in1[86] ^ in2[86];
    assign G[41] = in1[85] & in2[85];
    assign P[41] = in1[85] ^ in2[85];
    assign G[42] = in1[84] & in2[84];
    assign P[42] = in1[84] ^ in2[84];
    assign G[43] = in1[83] & in2[83];
    assign P[43] = in1[83] ^ in2[83];
    assign G[44] = in1[82] & in2[82];
    assign P[44] = in1[82] ^ in2[82];
    assign G[45] = in1[81] & in2[81];
    assign P[45] = in1[81] ^ in2[81];
    assign G[46] = in1[80] & in2[80];
    assign P[46] = in1[80] ^ in2[80];
    assign G[47] = in1[79] & in2[79];
    assign P[47] = in1[79] ^ in2[79];
    assign G[48] = in1[78] & in2[78];
    assign P[48] = in1[78] ^ in2[78];
    assign G[49] = in1[77] & in2[77];
    assign P[49] = in1[77] ^ in2[77];
    assign G[50] = in1[76] & in2[76];
    assign P[50] = in1[76] ^ in2[76];
    assign G[51] = in1[75] & in2[75];
    assign P[51] = in1[75] ^ in2[75];
    assign G[52] = in1[74] & in2[74];
    assign P[52] = in1[74] ^ in2[74];
    assign G[53] = in1[73] & in2[73];
    assign P[53] = in1[73] ^ in2[73];
    assign G[54] = in1[72] & in2[72];
    assign P[54] = in1[72] ^ in2[72];
    assign G[55] = in1[71] & in2[71];
    assign P[55] = in1[71] ^ in2[71];
    assign G[56] = in1[70] & in2[70];
    assign P[56] = in1[70] ^ in2[70];
    assign G[57] = in1[69] & in2[69];
    assign P[57] = in1[69] ^ in2[69];
    assign G[58] = in1[68] & in2[68];
    assign P[58] = in1[68] ^ in2[68];
    assign G[59] = in1[67] & in2[67];
    assign P[59] = in1[67] ^ in2[67];
    assign G[60] = in1[66] & in2[66];
    assign P[60] = in1[66] ^ in2[66];
    assign G[61] = in1[65] & in2[65];
    assign P[61] = in1[65] ^ in2[65];
    assign G[62] = in1[64] & in2[64];
    assign P[62] = in1[64] ^ in2[64];
    assign G[63] = in1[63] & in2[63];
    assign P[63] = in1[63] ^ in2[63];
    assign G[64] = in1[62] & in2[62];
    assign P[64] = in1[62] ^ in2[62];
    assign G[65] = in1[61] & in2[61];
    assign P[65] = in1[61] ^ in2[61];
    assign G[66] = in1[60] & in2[60];
    assign P[66] = in1[60] ^ in2[60];
    assign G[67] = in1[59] & in2[59];
    assign P[67] = in1[59] ^ in2[59];
    assign G[68] = in1[58] & in2[58];
    assign P[68] = in1[58] ^ in2[58];
    assign G[69] = in1[57] & in2[57];
    assign P[69] = in1[57] ^ in2[57];
    assign G[70] = in1[56] & in2[56];
    assign P[70] = in1[56] ^ in2[56];
    assign G[71] = in1[55] & in2[55];
    assign P[71] = in1[55] ^ in2[55];
    assign G[72] = in1[54] & in2[54];
    assign P[72] = in1[54] ^ in2[54];
    assign G[73] = in1[53] & in2[53];
    assign P[73] = in1[53] ^ in2[53];
    assign G[74] = in1[52] & in2[52];
    assign P[74] = in1[52] ^ in2[52];
    assign G[75] = in1[51] & in2[51];
    assign P[75] = in1[51] ^ in2[51];
    assign G[76] = in1[50] & in2[50];
    assign P[76] = in1[50] ^ in2[50];
    assign G[77] = in1[49] & in2[49];
    assign P[77] = in1[49] ^ in2[49];
    assign G[78] = in1[48] & in2[48];
    assign P[78] = in1[48] ^ in2[48];
    assign G[79] = in1[47] & in2[47];
    assign P[79] = in1[47] ^ in2[47];
    assign G[80] = in1[46] & in2[46];
    assign P[80] = in1[46] ^ in2[46];
    assign G[81] = in1[45] & in2[45];
    assign P[81] = in1[45] ^ in2[45];
    assign G[82] = in1[44] & in2[44];
    assign P[82] = in1[44] ^ in2[44];
    assign G[83] = in1[43] & in2[43];
    assign P[83] = in1[43] ^ in2[43];
    assign G[84] = in1[42] & in2[42];
    assign P[84] = in1[42] ^ in2[42];
    assign G[85] = in1[41] & in2[41];
    assign P[85] = in1[41] ^ in2[41];
    assign G[86] = in1[40] & in2[40];
    assign P[86] = in1[40] ^ in2[40];
    assign G[87] = in1[39] & in2[39];
    assign P[87] = in1[39] ^ in2[39];
    assign G[88] = in1[38] & in2[38];
    assign P[88] = in1[38] ^ in2[38];
    assign G[89] = in1[37] & in2[37];
    assign P[89] = in1[37] ^ in2[37];
    assign G[90] = in1[36] & in2[36];
    assign P[90] = in1[36] ^ in2[36];
    assign G[91] = in1[35] & in2[35];
    assign P[91] = in1[35] ^ in2[35];
    assign G[92] = in1[34] & in2[34];
    assign P[92] = in1[34] ^ in2[34];
    assign G[93] = in1[33] & in2[33];
    assign P[93] = in1[33] ^ in2[33];
    assign G[94] = in1[32] & in2[32];
    assign P[94] = in1[32] ^ in2[32];
    assign G[95] = in1[31] & in2[31];
    assign P[95] = in1[31] ^ in2[31];
    assign G[96] = in1[30] & in2[30];
    assign P[96] = in1[30] ^ in2[30];
    assign G[97] = in1[29] & in2[29];
    assign P[97] = in1[29] ^ in2[29];
    assign G[98] = in1[28] & in2[28];
    assign P[98] = in1[28] ^ in2[28];
    assign G[99] = in1[27] & in2[27];
    assign P[99] = in1[27] ^ in2[27];
    assign G[100] = in1[26] & in2[26];
    assign P[100] = in1[26] ^ in2[26];
    assign G[101] = in1[25] & in2[25];
    assign P[101] = in1[25] ^ in2[25];
    assign G[102] = in1[24] & in2[24];
    assign P[102] = in1[24] ^ in2[24];
    assign G[103] = in1[23] & in2[23];
    assign P[103] = in1[23] ^ in2[23];
    assign G[104] = in1[22] & in2[22];
    assign P[104] = in1[22] ^ in2[22];
    assign G[105] = in1[21] & in2[21];
    assign P[105] = in1[21] ^ in2[21];
    assign G[106] = in1[20] & in2[20];
    assign P[106] = in1[20] ^ in2[20];
    assign G[107] = in1[19] & in2[19];
    assign P[107] = in1[19] ^ in2[19];
    assign G[108] = in1[18] & in2[18];
    assign P[108] = in1[18] ^ in2[18];
    assign G[109] = in1[17] & in2[17];
    assign P[109] = in1[17] ^ in2[17];
    assign G[110] = in1[16] & in2[16];
    assign P[110] = in1[16] ^ in2[16];
    assign G[111] = in1[15] & in2[15];
    assign P[111] = in1[15] ^ in2[15];
    assign G[112] = in1[14] & in2[14];
    assign P[112] = in1[14] ^ in2[14];
    assign G[113] = in1[13] & in2[13];
    assign P[113] = in1[13] ^ in2[13];
    assign G[114] = in1[12] & in2[12];
    assign P[114] = in1[12] ^ in2[12];
    assign G[115] = in1[11] & in2[11];
    assign P[115] = in1[11] ^ in2[11];
    assign G[116] = in1[10] & in2[10];
    assign P[116] = in1[10] ^ in2[10];
    assign G[117] = in1[9] & in2[9];
    assign P[117] = in1[9] ^ in2[9];
    assign G[118] = in1[8] & in2[8];
    assign P[118] = in1[8] ^ in2[8];
    assign G[119] = in1[7] & in2[7];
    assign P[119] = in1[7] ^ in2[7];
    assign G[120] = in1[6] & in2[6];
    assign P[120] = in1[6] ^ in2[6];
    assign G[121] = in1[5] & in2[5];
    assign P[121] = in1[5] ^ in2[5];
    assign G[122] = in1[4] & in2[4];
    assign P[122] = in1[4] ^ in2[4];
    assign G[123] = in1[3] & in2[3];
    assign P[123] = in1[3] ^ in2[3];
    assign G[124] = in1[2] & in2[2];
    assign P[124] = in1[2] ^ in2[2];
    assign G[125] = in1[1] & in2[1];
    assign P[125] = in1[1] ^ in2[1];
    assign G[126] = in1[0] & in2[0];
    assign P[126] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign cout = G[126] | (P[126] & C[126]);
    assign sum = P ^ C;
endmodule

module CLA_126(output [125:0] sum, output cout, input [125:0] in1, input [125:0] in2);

    wire[125:0] G;
    wire[125:0] C;
    wire[125:0] P;

    assign G[0] = in1[125] & in2[125];
    assign P[0] = in1[125] ^ in2[125];
    assign G[1] = in1[124] & in2[124];
    assign P[1] = in1[124] ^ in2[124];
    assign G[2] = in1[123] & in2[123];
    assign P[2] = in1[123] ^ in2[123];
    assign G[3] = in1[122] & in2[122];
    assign P[3] = in1[122] ^ in2[122];
    assign G[4] = in1[121] & in2[121];
    assign P[4] = in1[121] ^ in2[121];
    assign G[5] = in1[120] & in2[120];
    assign P[5] = in1[120] ^ in2[120];
    assign G[6] = in1[119] & in2[119];
    assign P[6] = in1[119] ^ in2[119];
    assign G[7] = in1[118] & in2[118];
    assign P[7] = in1[118] ^ in2[118];
    assign G[8] = in1[117] & in2[117];
    assign P[8] = in1[117] ^ in2[117];
    assign G[9] = in1[116] & in2[116];
    assign P[9] = in1[116] ^ in2[116];
    assign G[10] = in1[115] & in2[115];
    assign P[10] = in1[115] ^ in2[115];
    assign G[11] = in1[114] & in2[114];
    assign P[11] = in1[114] ^ in2[114];
    assign G[12] = in1[113] & in2[113];
    assign P[12] = in1[113] ^ in2[113];
    assign G[13] = in1[112] & in2[112];
    assign P[13] = in1[112] ^ in2[112];
    assign G[14] = in1[111] & in2[111];
    assign P[14] = in1[111] ^ in2[111];
    assign G[15] = in1[110] & in2[110];
    assign P[15] = in1[110] ^ in2[110];
    assign G[16] = in1[109] & in2[109];
    assign P[16] = in1[109] ^ in2[109];
    assign G[17] = in1[108] & in2[108];
    assign P[17] = in1[108] ^ in2[108];
    assign G[18] = in1[107] & in2[107];
    assign P[18] = in1[107] ^ in2[107];
    assign G[19] = in1[106] & in2[106];
    assign P[19] = in1[106] ^ in2[106];
    assign G[20] = in1[105] & in2[105];
    assign P[20] = in1[105] ^ in2[105];
    assign G[21] = in1[104] & in2[104];
    assign P[21] = in1[104] ^ in2[104];
    assign G[22] = in1[103] & in2[103];
    assign P[22] = in1[103] ^ in2[103];
    assign G[23] = in1[102] & in2[102];
    assign P[23] = in1[102] ^ in2[102];
    assign G[24] = in1[101] & in2[101];
    assign P[24] = in1[101] ^ in2[101];
    assign G[25] = in1[100] & in2[100];
    assign P[25] = in1[100] ^ in2[100];
    assign G[26] = in1[99] & in2[99];
    assign P[26] = in1[99] ^ in2[99];
    assign G[27] = in1[98] & in2[98];
    assign P[27] = in1[98] ^ in2[98];
    assign G[28] = in1[97] & in2[97];
    assign P[28] = in1[97] ^ in2[97];
    assign G[29] = in1[96] & in2[96];
    assign P[29] = in1[96] ^ in2[96];
    assign G[30] = in1[95] & in2[95];
    assign P[30] = in1[95] ^ in2[95];
    assign G[31] = in1[94] & in2[94];
    assign P[31] = in1[94] ^ in2[94];
    assign G[32] = in1[93] & in2[93];
    assign P[32] = in1[93] ^ in2[93];
    assign G[33] = in1[92] & in2[92];
    assign P[33] = in1[92] ^ in2[92];
    assign G[34] = in1[91] & in2[91];
    assign P[34] = in1[91] ^ in2[91];
    assign G[35] = in1[90] & in2[90];
    assign P[35] = in1[90] ^ in2[90];
    assign G[36] = in1[89] & in2[89];
    assign P[36] = in1[89] ^ in2[89];
    assign G[37] = in1[88] & in2[88];
    assign P[37] = in1[88] ^ in2[88];
    assign G[38] = in1[87] & in2[87];
    assign P[38] = in1[87] ^ in2[87];
    assign G[39] = in1[86] & in2[86];
    assign P[39] = in1[86] ^ in2[86];
    assign G[40] = in1[85] & in2[85];
    assign P[40] = in1[85] ^ in2[85];
    assign G[41] = in1[84] & in2[84];
    assign P[41] = in1[84] ^ in2[84];
    assign G[42] = in1[83] & in2[83];
    assign P[42] = in1[83] ^ in2[83];
    assign G[43] = in1[82] & in2[82];
    assign P[43] = in1[82] ^ in2[82];
    assign G[44] = in1[81] & in2[81];
    assign P[44] = in1[81] ^ in2[81];
    assign G[45] = in1[80] & in2[80];
    assign P[45] = in1[80] ^ in2[80];
    assign G[46] = in1[79] & in2[79];
    assign P[46] = in1[79] ^ in2[79];
    assign G[47] = in1[78] & in2[78];
    assign P[47] = in1[78] ^ in2[78];
    assign G[48] = in1[77] & in2[77];
    assign P[48] = in1[77] ^ in2[77];
    assign G[49] = in1[76] & in2[76];
    assign P[49] = in1[76] ^ in2[76];
    assign G[50] = in1[75] & in2[75];
    assign P[50] = in1[75] ^ in2[75];
    assign G[51] = in1[74] & in2[74];
    assign P[51] = in1[74] ^ in2[74];
    assign G[52] = in1[73] & in2[73];
    assign P[52] = in1[73] ^ in2[73];
    assign G[53] = in1[72] & in2[72];
    assign P[53] = in1[72] ^ in2[72];
    assign G[54] = in1[71] & in2[71];
    assign P[54] = in1[71] ^ in2[71];
    assign G[55] = in1[70] & in2[70];
    assign P[55] = in1[70] ^ in2[70];
    assign G[56] = in1[69] & in2[69];
    assign P[56] = in1[69] ^ in2[69];
    assign G[57] = in1[68] & in2[68];
    assign P[57] = in1[68] ^ in2[68];
    assign G[58] = in1[67] & in2[67];
    assign P[58] = in1[67] ^ in2[67];
    assign G[59] = in1[66] & in2[66];
    assign P[59] = in1[66] ^ in2[66];
    assign G[60] = in1[65] & in2[65];
    assign P[60] = in1[65] ^ in2[65];
    assign G[61] = in1[64] & in2[64];
    assign P[61] = in1[64] ^ in2[64];
    assign G[62] = in1[63] & in2[63];
    assign P[62] = in1[63] ^ in2[63];
    assign G[63] = in1[62] & in2[62];
    assign P[63] = in1[62] ^ in2[62];
    assign G[64] = in1[61] & in2[61];
    assign P[64] = in1[61] ^ in2[61];
    assign G[65] = in1[60] & in2[60];
    assign P[65] = in1[60] ^ in2[60];
    assign G[66] = in1[59] & in2[59];
    assign P[66] = in1[59] ^ in2[59];
    assign G[67] = in1[58] & in2[58];
    assign P[67] = in1[58] ^ in2[58];
    assign G[68] = in1[57] & in2[57];
    assign P[68] = in1[57] ^ in2[57];
    assign G[69] = in1[56] & in2[56];
    assign P[69] = in1[56] ^ in2[56];
    assign G[70] = in1[55] & in2[55];
    assign P[70] = in1[55] ^ in2[55];
    assign G[71] = in1[54] & in2[54];
    assign P[71] = in1[54] ^ in2[54];
    assign G[72] = in1[53] & in2[53];
    assign P[72] = in1[53] ^ in2[53];
    assign G[73] = in1[52] & in2[52];
    assign P[73] = in1[52] ^ in2[52];
    assign G[74] = in1[51] & in2[51];
    assign P[74] = in1[51] ^ in2[51];
    assign G[75] = in1[50] & in2[50];
    assign P[75] = in1[50] ^ in2[50];
    assign G[76] = in1[49] & in2[49];
    assign P[76] = in1[49] ^ in2[49];
    assign G[77] = in1[48] & in2[48];
    assign P[77] = in1[48] ^ in2[48];
    assign G[78] = in1[47] & in2[47];
    assign P[78] = in1[47] ^ in2[47];
    assign G[79] = in1[46] & in2[46];
    assign P[79] = in1[46] ^ in2[46];
    assign G[80] = in1[45] & in2[45];
    assign P[80] = in1[45] ^ in2[45];
    assign G[81] = in1[44] & in2[44];
    assign P[81] = in1[44] ^ in2[44];
    assign G[82] = in1[43] & in2[43];
    assign P[82] = in1[43] ^ in2[43];
    assign G[83] = in1[42] & in2[42];
    assign P[83] = in1[42] ^ in2[42];
    assign G[84] = in1[41] & in2[41];
    assign P[84] = in1[41] ^ in2[41];
    assign G[85] = in1[40] & in2[40];
    assign P[85] = in1[40] ^ in2[40];
    assign G[86] = in1[39] & in2[39];
    assign P[86] = in1[39] ^ in2[39];
    assign G[87] = in1[38] & in2[38];
    assign P[87] = in1[38] ^ in2[38];
    assign G[88] = in1[37] & in2[37];
    assign P[88] = in1[37] ^ in2[37];
    assign G[89] = in1[36] & in2[36];
    assign P[89] = in1[36] ^ in2[36];
    assign G[90] = in1[35] & in2[35];
    assign P[90] = in1[35] ^ in2[35];
    assign G[91] = in1[34] & in2[34];
    assign P[91] = in1[34] ^ in2[34];
    assign G[92] = in1[33] & in2[33];
    assign P[92] = in1[33] ^ in2[33];
    assign G[93] = in1[32] & in2[32];
    assign P[93] = in1[32] ^ in2[32];
    assign G[94] = in1[31] & in2[31];
    assign P[94] = in1[31] ^ in2[31];
    assign G[95] = in1[30] & in2[30];
    assign P[95] = in1[30] ^ in2[30];
    assign G[96] = in1[29] & in2[29];
    assign P[96] = in1[29] ^ in2[29];
    assign G[97] = in1[28] & in2[28];
    assign P[97] = in1[28] ^ in2[28];
    assign G[98] = in1[27] & in2[27];
    assign P[98] = in1[27] ^ in2[27];
    assign G[99] = in1[26] & in2[26];
    assign P[99] = in1[26] ^ in2[26];
    assign G[100] = in1[25] & in2[25];
    assign P[100] = in1[25] ^ in2[25];
    assign G[101] = in1[24] & in2[24];
    assign P[101] = in1[24] ^ in2[24];
    assign G[102] = in1[23] & in2[23];
    assign P[102] = in1[23] ^ in2[23];
    assign G[103] = in1[22] & in2[22];
    assign P[103] = in1[22] ^ in2[22];
    assign G[104] = in1[21] & in2[21];
    assign P[104] = in1[21] ^ in2[21];
    assign G[105] = in1[20] & in2[20];
    assign P[105] = in1[20] ^ in2[20];
    assign G[106] = in1[19] & in2[19];
    assign P[106] = in1[19] ^ in2[19];
    assign G[107] = in1[18] & in2[18];
    assign P[107] = in1[18] ^ in2[18];
    assign G[108] = in1[17] & in2[17];
    assign P[108] = in1[17] ^ in2[17];
    assign G[109] = in1[16] & in2[16];
    assign P[109] = in1[16] ^ in2[16];
    assign G[110] = in1[15] & in2[15];
    assign P[110] = in1[15] ^ in2[15];
    assign G[111] = in1[14] & in2[14];
    assign P[111] = in1[14] ^ in2[14];
    assign G[112] = in1[13] & in2[13];
    assign P[112] = in1[13] ^ in2[13];
    assign G[113] = in1[12] & in2[12];
    assign P[113] = in1[12] ^ in2[12];
    assign G[114] = in1[11] & in2[11];
    assign P[114] = in1[11] ^ in2[11];
    assign G[115] = in1[10] & in2[10];
    assign P[115] = in1[10] ^ in2[10];
    assign G[116] = in1[9] & in2[9];
    assign P[116] = in1[9] ^ in2[9];
    assign G[117] = in1[8] & in2[8];
    assign P[117] = in1[8] ^ in2[8];
    assign G[118] = in1[7] & in2[7];
    assign P[118] = in1[7] ^ in2[7];
    assign G[119] = in1[6] & in2[6];
    assign P[119] = in1[6] ^ in2[6];
    assign G[120] = in1[5] & in2[5];
    assign P[120] = in1[5] ^ in2[5];
    assign G[121] = in1[4] & in2[4];
    assign P[121] = in1[4] ^ in2[4];
    assign G[122] = in1[3] & in2[3];
    assign P[122] = in1[3] ^ in2[3];
    assign G[123] = in1[2] & in2[2];
    assign P[123] = in1[2] ^ in2[2];
    assign G[124] = in1[1] & in2[1];
    assign P[124] = in1[1] ^ in2[1];
    assign G[125] = in1[0] & in2[0];
    assign P[125] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign cout = G[125] | (P[125] & C[125]);
    assign sum = P ^ C;
endmodule

module CLA_125(output [124:0] sum, output cout, input [124:0] in1, input [124:0] in2);

    wire[124:0] G;
    wire[124:0] C;
    wire[124:0] P;

    assign G[0] = in1[124] & in2[124];
    assign P[0] = in1[124] ^ in2[124];
    assign G[1] = in1[123] & in2[123];
    assign P[1] = in1[123] ^ in2[123];
    assign G[2] = in1[122] & in2[122];
    assign P[2] = in1[122] ^ in2[122];
    assign G[3] = in1[121] & in2[121];
    assign P[3] = in1[121] ^ in2[121];
    assign G[4] = in1[120] & in2[120];
    assign P[4] = in1[120] ^ in2[120];
    assign G[5] = in1[119] & in2[119];
    assign P[5] = in1[119] ^ in2[119];
    assign G[6] = in1[118] & in2[118];
    assign P[6] = in1[118] ^ in2[118];
    assign G[7] = in1[117] & in2[117];
    assign P[7] = in1[117] ^ in2[117];
    assign G[8] = in1[116] & in2[116];
    assign P[8] = in1[116] ^ in2[116];
    assign G[9] = in1[115] & in2[115];
    assign P[9] = in1[115] ^ in2[115];
    assign G[10] = in1[114] & in2[114];
    assign P[10] = in1[114] ^ in2[114];
    assign G[11] = in1[113] & in2[113];
    assign P[11] = in1[113] ^ in2[113];
    assign G[12] = in1[112] & in2[112];
    assign P[12] = in1[112] ^ in2[112];
    assign G[13] = in1[111] & in2[111];
    assign P[13] = in1[111] ^ in2[111];
    assign G[14] = in1[110] & in2[110];
    assign P[14] = in1[110] ^ in2[110];
    assign G[15] = in1[109] & in2[109];
    assign P[15] = in1[109] ^ in2[109];
    assign G[16] = in1[108] & in2[108];
    assign P[16] = in1[108] ^ in2[108];
    assign G[17] = in1[107] & in2[107];
    assign P[17] = in1[107] ^ in2[107];
    assign G[18] = in1[106] & in2[106];
    assign P[18] = in1[106] ^ in2[106];
    assign G[19] = in1[105] & in2[105];
    assign P[19] = in1[105] ^ in2[105];
    assign G[20] = in1[104] & in2[104];
    assign P[20] = in1[104] ^ in2[104];
    assign G[21] = in1[103] & in2[103];
    assign P[21] = in1[103] ^ in2[103];
    assign G[22] = in1[102] & in2[102];
    assign P[22] = in1[102] ^ in2[102];
    assign G[23] = in1[101] & in2[101];
    assign P[23] = in1[101] ^ in2[101];
    assign G[24] = in1[100] & in2[100];
    assign P[24] = in1[100] ^ in2[100];
    assign G[25] = in1[99] & in2[99];
    assign P[25] = in1[99] ^ in2[99];
    assign G[26] = in1[98] & in2[98];
    assign P[26] = in1[98] ^ in2[98];
    assign G[27] = in1[97] & in2[97];
    assign P[27] = in1[97] ^ in2[97];
    assign G[28] = in1[96] & in2[96];
    assign P[28] = in1[96] ^ in2[96];
    assign G[29] = in1[95] & in2[95];
    assign P[29] = in1[95] ^ in2[95];
    assign G[30] = in1[94] & in2[94];
    assign P[30] = in1[94] ^ in2[94];
    assign G[31] = in1[93] & in2[93];
    assign P[31] = in1[93] ^ in2[93];
    assign G[32] = in1[92] & in2[92];
    assign P[32] = in1[92] ^ in2[92];
    assign G[33] = in1[91] & in2[91];
    assign P[33] = in1[91] ^ in2[91];
    assign G[34] = in1[90] & in2[90];
    assign P[34] = in1[90] ^ in2[90];
    assign G[35] = in1[89] & in2[89];
    assign P[35] = in1[89] ^ in2[89];
    assign G[36] = in1[88] & in2[88];
    assign P[36] = in1[88] ^ in2[88];
    assign G[37] = in1[87] & in2[87];
    assign P[37] = in1[87] ^ in2[87];
    assign G[38] = in1[86] & in2[86];
    assign P[38] = in1[86] ^ in2[86];
    assign G[39] = in1[85] & in2[85];
    assign P[39] = in1[85] ^ in2[85];
    assign G[40] = in1[84] & in2[84];
    assign P[40] = in1[84] ^ in2[84];
    assign G[41] = in1[83] & in2[83];
    assign P[41] = in1[83] ^ in2[83];
    assign G[42] = in1[82] & in2[82];
    assign P[42] = in1[82] ^ in2[82];
    assign G[43] = in1[81] & in2[81];
    assign P[43] = in1[81] ^ in2[81];
    assign G[44] = in1[80] & in2[80];
    assign P[44] = in1[80] ^ in2[80];
    assign G[45] = in1[79] & in2[79];
    assign P[45] = in1[79] ^ in2[79];
    assign G[46] = in1[78] & in2[78];
    assign P[46] = in1[78] ^ in2[78];
    assign G[47] = in1[77] & in2[77];
    assign P[47] = in1[77] ^ in2[77];
    assign G[48] = in1[76] & in2[76];
    assign P[48] = in1[76] ^ in2[76];
    assign G[49] = in1[75] & in2[75];
    assign P[49] = in1[75] ^ in2[75];
    assign G[50] = in1[74] & in2[74];
    assign P[50] = in1[74] ^ in2[74];
    assign G[51] = in1[73] & in2[73];
    assign P[51] = in1[73] ^ in2[73];
    assign G[52] = in1[72] & in2[72];
    assign P[52] = in1[72] ^ in2[72];
    assign G[53] = in1[71] & in2[71];
    assign P[53] = in1[71] ^ in2[71];
    assign G[54] = in1[70] & in2[70];
    assign P[54] = in1[70] ^ in2[70];
    assign G[55] = in1[69] & in2[69];
    assign P[55] = in1[69] ^ in2[69];
    assign G[56] = in1[68] & in2[68];
    assign P[56] = in1[68] ^ in2[68];
    assign G[57] = in1[67] & in2[67];
    assign P[57] = in1[67] ^ in2[67];
    assign G[58] = in1[66] & in2[66];
    assign P[58] = in1[66] ^ in2[66];
    assign G[59] = in1[65] & in2[65];
    assign P[59] = in1[65] ^ in2[65];
    assign G[60] = in1[64] & in2[64];
    assign P[60] = in1[64] ^ in2[64];
    assign G[61] = in1[63] & in2[63];
    assign P[61] = in1[63] ^ in2[63];
    assign G[62] = in1[62] & in2[62];
    assign P[62] = in1[62] ^ in2[62];
    assign G[63] = in1[61] & in2[61];
    assign P[63] = in1[61] ^ in2[61];
    assign G[64] = in1[60] & in2[60];
    assign P[64] = in1[60] ^ in2[60];
    assign G[65] = in1[59] & in2[59];
    assign P[65] = in1[59] ^ in2[59];
    assign G[66] = in1[58] & in2[58];
    assign P[66] = in1[58] ^ in2[58];
    assign G[67] = in1[57] & in2[57];
    assign P[67] = in1[57] ^ in2[57];
    assign G[68] = in1[56] & in2[56];
    assign P[68] = in1[56] ^ in2[56];
    assign G[69] = in1[55] & in2[55];
    assign P[69] = in1[55] ^ in2[55];
    assign G[70] = in1[54] & in2[54];
    assign P[70] = in1[54] ^ in2[54];
    assign G[71] = in1[53] & in2[53];
    assign P[71] = in1[53] ^ in2[53];
    assign G[72] = in1[52] & in2[52];
    assign P[72] = in1[52] ^ in2[52];
    assign G[73] = in1[51] & in2[51];
    assign P[73] = in1[51] ^ in2[51];
    assign G[74] = in1[50] & in2[50];
    assign P[74] = in1[50] ^ in2[50];
    assign G[75] = in1[49] & in2[49];
    assign P[75] = in1[49] ^ in2[49];
    assign G[76] = in1[48] & in2[48];
    assign P[76] = in1[48] ^ in2[48];
    assign G[77] = in1[47] & in2[47];
    assign P[77] = in1[47] ^ in2[47];
    assign G[78] = in1[46] & in2[46];
    assign P[78] = in1[46] ^ in2[46];
    assign G[79] = in1[45] & in2[45];
    assign P[79] = in1[45] ^ in2[45];
    assign G[80] = in1[44] & in2[44];
    assign P[80] = in1[44] ^ in2[44];
    assign G[81] = in1[43] & in2[43];
    assign P[81] = in1[43] ^ in2[43];
    assign G[82] = in1[42] & in2[42];
    assign P[82] = in1[42] ^ in2[42];
    assign G[83] = in1[41] & in2[41];
    assign P[83] = in1[41] ^ in2[41];
    assign G[84] = in1[40] & in2[40];
    assign P[84] = in1[40] ^ in2[40];
    assign G[85] = in1[39] & in2[39];
    assign P[85] = in1[39] ^ in2[39];
    assign G[86] = in1[38] & in2[38];
    assign P[86] = in1[38] ^ in2[38];
    assign G[87] = in1[37] & in2[37];
    assign P[87] = in1[37] ^ in2[37];
    assign G[88] = in1[36] & in2[36];
    assign P[88] = in1[36] ^ in2[36];
    assign G[89] = in1[35] & in2[35];
    assign P[89] = in1[35] ^ in2[35];
    assign G[90] = in1[34] & in2[34];
    assign P[90] = in1[34] ^ in2[34];
    assign G[91] = in1[33] & in2[33];
    assign P[91] = in1[33] ^ in2[33];
    assign G[92] = in1[32] & in2[32];
    assign P[92] = in1[32] ^ in2[32];
    assign G[93] = in1[31] & in2[31];
    assign P[93] = in1[31] ^ in2[31];
    assign G[94] = in1[30] & in2[30];
    assign P[94] = in1[30] ^ in2[30];
    assign G[95] = in1[29] & in2[29];
    assign P[95] = in1[29] ^ in2[29];
    assign G[96] = in1[28] & in2[28];
    assign P[96] = in1[28] ^ in2[28];
    assign G[97] = in1[27] & in2[27];
    assign P[97] = in1[27] ^ in2[27];
    assign G[98] = in1[26] & in2[26];
    assign P[98] = in1[26] ^ in2[26];
    assign G[99] = in1[25] & in2[25];
    assign P[99] = in1[25] ^ in2[25];
    assign G[100] = in1[24] & in2[24];
    assign P[100] = in1[24] ^ in2[24];
    assign G[101] = in1[23] & in2[23];
    assign P[101] = in1[23] ^ in2[23];
    assign G[102] = in1[22] & in2[22];
    assign P[102] = in1[22] ^ in2[22];
    assign G[103] = in1[21] & in2[21];
    assign P[103] = in1[21] ^ in2[21];
    assign G[104] = in1[20] & in2[20];
    assign P[104] = in1[20] ^ in2[20];
    assign G[105] = in1[19] & in2[19];
    assign P[105] = in1[19] ^ in2[19];
    assign G[106] = in1[18] & in2[18];
    assign P[106] = in1[18] ^ in2[18];
    assign G[107] = in1[17] & in2[17];
    assign P[107] = in1[17] ^ in2[17];
    assign G[108] = in1[16] & in2[16];
    assign P[108] = in1[16] ^ in2[16];
    assign G[109] = in1[15] & in2[15];
    assign P[109] = in1[15] ^ in2[15];
    assign G[110] = in1[14] & in2[14];
    assign P[110] = in1[14] ^ in2[14];
    assign G[111] = in1[13] & in2[13];
    assign P[111] = in1[13] ^ in2[13];
    assign G[112] = in1[12] & in2[12];
    assign P[112] = in1[12] ^ in2[12];
    assign G[113] = in1[11] & in2[11];
    assign P[113] = in1[11] ^ in2[11];
    assign G[114] = in1[10] & in2[10];
    assign P[114] = in1[10] ^ in2[10];
    assign G[115] = in1[9] & in2[9];
    assign P[115] = in1[9] ^ in2[9];
    assign G[116] = in1[8] & in2[8];
    assign P[116] = in1[8] ^ in2[8];
    assign G[117] = in1[7] & in2[7];
    assign P[117] = in1[7] ^ in2[7];
    assign G[118] = in1[6] & in2[6];
    assign P[118] = in1[6] ^ in2[6];
    assign G[119] = in1[5] & in2[5];
    assign P[119] = in1[5] ^ in2[5];
    assign G[120] = in1[4] & in2[4];
    assign P[120] = in1[4] ^ in2[4];
    assign G[121] = in1[3] & in2[3];
    assign P[121] = in1[3] ^ in2[3];
    assign G[122] = in1[2] & in2[2];
    assign P[122] = in1[2] ^ in2[2];
    assign G[123] = in1[1] & in2[1];
    assign P[123] = in1[1] ^ in2[1];
    assign G[124] = in1[0] & in2[0];
    assign P[124] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign cout = G[124] | (P[124] & C[124]);
    assign sum = P ^ C;
endmodule

module CLA_124(output [123:0] sum, output cout, input [123:0] in1, input [123:0] in2);

    wire[123:0] G;
    wire[123:0] C;
    wire[123:0] P;

    assign G[0] = in1[123] & in2[123];
    assign P[0] = in1[123] ^ in2[123];
    assign G[1] = in1[122] & in2[122];
    assign P[1] = in1[122] ^ in2[122];
    assign G[2] = in1[121] & in2[121];
    assign P[2] = in1[121] ^ in2[121];
    assign G[3] = in1[120] & in2[120];
    assign P[3] = in1[120] ^ in2[120];
    assign G[4] = in1[119] & in2[119];
    assign P[4] = in1[119] ^ in2[119];
    assign G[5] = in1[118] & in2[118];
    assign P[5] = in1[118] ^ in2[118];
    assign G[6] = in1[117] & in2[117];
    assign P[6] = in1[117] ^ in2[117];
    assign G[7] = in1[116] & in2[116];
    assign P[7] = in1[116] ^ in2[116];
    assign G[8] = in1[115] & in2[115];
    assign P[8] = in1[115] ^ in2[115];
    assign G[9] = in1[114] & in2[114];
    assign P[9] = in1[114] ^ in2[114];
    assign G[10] = in1[113] & in2[113];
    assign P[10] = in1[113] ^ in2[113];
    assign G[11] = in1[112] & in2[112];
    assign P[11] = in1[112] ^ in2[112];
    assign G[12] = in1[111] & in2[111];
    assign P[12] = in1[111] ^ in2[111];
    assign G[13] = in1[110] & in2[110];
    assign P[13] = in1[110] ^ in2[110];
    assign G[14] = in1[109] & in2[109];
    assign P[14] = in1[109] ^ in2[109];
    assign G[15] = in1[108] & in2[108];
    assign P[15] = in1[108] ^ in2[108];
    assign G[16] = in1[107] & in2[107];
    assign P[16] = in1[107] ^ in2[107];
    assign G[17] = in1[106] & in2[106];
    assign P[17] = in1[106] ^ in2[106];
    assign G[18] = in1[105] & in2[105];
    assign P[18] = in1[105] ^ in2[105];
    assign G[19] = in1[104] & in2[104];
    assign P[19] = in1[104] ^ in2[104];
    assign G[20] = in1[103] & in2[103];
    assign P[20] = in1[103] ^ in2[103];
    assign G[21] = in1[102] & in2[102];
    assign P[21] = in1[102] ^ in2[102];
    assign G[22] = in1[101] & in2[101];
    assign P[22] = in1[101] ^ in2[101];
    assign G[23] = in1[100] & in2[100];
    assign P[23] = in1[100] ^ in2[100];
    assign G[24] = in1[99] & in2[99];
    assign P[24] = in1[99] ^ in2[99];
    assign G[25] = in1[98] & in2[98];
    assign P[25] = in1[98] ^ in2[98];
    assign G[26] = in1[97] & in2[97];
    assign P[26] = in1[97] ^ in2[97];
    assign G[27] = in1[96] & in2[96];
    assign P[27] = in1[96] ^ in2[96];
    assign G[28] = in1[95] & in2[95];
    assign P[28] = in1[95] ^ in2[95];
    assign G[29] = in1[94] & in2[94];
    assign P[29] = in1[94] ^ in2[94];
    assign G[30] = in1[93] & in2[93];
    assign P[30] = in1[93] ^ in2[93];
    assign G[31] = in1[92] & in2[92];
    assign P[31] = in1[92] ^ in2[92];
    assign G[32] = in1[91] & in2[91];
    assign P[32] = in1[91] ^ in2[91];
    assign G[33] = in1[90] & in2[90];
    assign P[33] = in1[90] ^ in2[90];
    assign G[34] = in1[89] & in2[89];
    assign P[34] = in1[89] ^ in2[89];
    assign G[35] = in1[88] & in2[88];
    assign P[35] = in1[88] ^ in2[88];
    assign G[36] = in1[87] & in2[87];
    assign P[36] = in1[87] ^ in2[87];
    assign G[37] = in1[86] & in2[86];
    assign P[37] = in1[86] ^ in2[86];
    assign G[38] = in1[85] & in2[85];
    assign P[38] = in1[85] ^ in2[85];
    assign G[39] = in1[84] & in2[84];
    assign P[39] = in1[84] ^ in2[84];
    assign G[40] = in1[83] & in2[83];
    assign P[40] = in1[83] ^ in2[83];
    assign G[41] = in1[82] & in2[82];
    assign P[41] = in1[82] ^ in2[82];
    assign G[42] = in1[81] & in2[81];
    assign P[42] = in1[81] ^ in2[81];
    assign G[43] = in1[80] & in2[80];
    assign P[43] = in1[80] ^ in2[80];
    assign G[44] = in1[79] & in2[79];
    assign P[44] = in1[79] ^ in2[79];
    assign G[45] = in1[78] & in2[78];
    assign P[45] = in1[78] ^ in2[78];
    assign G[46] = in1[77] & in2[77];
    assign P[46] = in1[77] ^ in2[77];
    assign G[47] = in1[76] & in2[76];
    assign P[47] = in1[76] ^ in2[76];
    assign G[48] = in1[75] & in2[75];
    assign P[48] = in1[75] ^ in2[75];
    assign G[49] = in1[74] & in2[74];
    assign P[49] = in1[74] ^ in2[74];
    assign G[50] = in1[73] & in2[73];
    assign P[50] = in1[73] ^ in2[73];
    assign G[51] = in1[72] & in2[72];
    assign P[51] = in1[72] ^ in2[72];
    assign G[52] = in1[71] & in2[71];
    assign P[52] = in1[71] ^ in2[71];
    assign G[53] = in1[70] & in2[70];
    assign P[53] = in1[70] ^ in2[70];
    assign G[54] = in1[69] & in2[69];
    assign P[54] = in1[69] ^ in2[69];
    assign G[55] = in1[68] & in2[68];
    assign P[55] = in1[68] ^ in2[68];
    assign G[56] = in1[67] & in2[67];
    assign P[56] = in1[67] ^ in2[67];
    assign G[57] = in1[66] & in2[66];
    assign P[57] = in1[66] ^ in2[66];
    assign G[58] = in1[65] & in2[65];
    assign P[58] = in1[65] ^ in2[65];
    assign G[59] = in1[64] & in2[64];
    assign P[59] = in1[64] ^ in2[64];
    assign G[60] = in1[63] & in2[63];
    assign P[60] = in1[63] ^ in2[63];
    assign G[61] = in1[62] & in2[62];
    assign P[61] = in1[62] ^ in2[62];
    assign G[62] = in1[61] & in2[61];
    assign P[62] = in1[61] ^ in2[61];
    assign G[63] = in1[60] & in2[60];
    assign P[63] = in1[60] ^ in2[60];
    assign G[64] = in1[59] & in2[59];
    assign P[64] = in1[59] ^ in2[59];
    assign G[65] = in1[58] & in2[58];
    assign P[65] = in1[58] ^ in2[58];
    assign G[66] = in1[57] & in2[57];
    assign P[66] = in1[57] ^ in2[57];
    assign G[67] = in1[56] & in2[56];
    assign P[67] = in1[56] ^ in2[56];
    assign G[68] = in1[55] & in2[55];
    assign P[68] = in1[55] ^ in2[55];
    assign G[69] = in1[54] & in2[54];
    assign P[69] = in1[54] ^ in2[54];
    assign G[70] = in1[53] & in2[53];
    assign P[70] = in1[53] ^ in2[53];
    assign G[71] = in1[52] & in2[52];
    assign P[71] = in1[52] ^ in2[52];
    assign G[72] = in1[51] & in2[51];
    assign P[72] = in1[51] ^ in2[51];
    assign G[73] = in1[50] & in2[50];
    assign P[73] = in1[50] ^ in2[50];
    assign G[74] = in1[49] & in2[49];
    assign P[74] = in1[49] ^ in2[49];
    assign G[75] = in1[48] & in2[48];
    assign P[75] = in1[48] ^ in2[48];
    assign G[76] = in1[47] & in2[47];
    assign P[76] = in1[47] ^ in2[47];
    assign G[77] = in1[46] & in2[46];
    assign P[77] = in1[46] ^ in2[46];
    assign G[78] = in1[45] & in2[45];
    assign P[78] = in1[45] ^ in2[45];
    assign G[79] = in1[44] & in2[44];
    assign P[79] = in1[44] ^ in2[44];
    assign G[80] = in1[43] & in2[43];
    assign P[80] = in1[43] ^ in2[43];
    assign G[81] = in1[42] & in2[42];
    assign P[81] = in1[42] ^ in2[42];
    assign G[82] = in1[41] & in2[41];
    assign P[82] = in1[41] ^ in2[41];
    assign G[83] = in1[40] & in2[40];
    assign P[83] = in1[40] ^ in2[40];
    assign G[84] = in1[39] & in2[39];
    assign P[84] = in1[39] ^ in2[39];
    assign G[85] = in1[38] & in2[38];
    assign P[85] = in1[38] ^ in2[38];
    assign G[86] = in1[37] & in2[37];
    assign P[86] = in1[37] ^ in2[37];
    assign G[87] = in1[36] & in2[36];
    assign P[87] = in1[36] ^ in2[36];
    assign G[88] = in1[35] & in2[35];
    assign P[88] = in1[35] ^ in2[35];
    assign G[89] = in1[34] & in2[34];
    assign P[89] = in1[34] ^ in2[34];
    assign G[90] = in1[33] & in2[33];
    assign P[90] = in1[33] ^ in2[33];
    assign G[91] = in1[32] & in2[32];
    assign P[91] = in1[32] ^ in2[32];
    assign G[92] = in1[31] & in2[31];
    assign P[92] = in1[31] ^ in2[31];
    assign G[93] = in1[30] & in2[30];
    assign P[93] = in1[30] ^ in2[30];
    assign G[94] = in1[29] & in2[29];
    assign P[94] = in1[29] ^ in2[29];
    assign G[95] = in1[28] & in2[28];
    assign P[95] = in1[28] ^ in2[28];
    assign G[96] = in1[27] & in2[27];
    assign P[96] = in1[27] ^ in2[27];
    assign G[97] = in1[26] & in2[26];
    assign P[97] = in1[26] ^ in2[26];
    assign G[98] = in1[25] & in2[25];
    assign P[98] = in1[25] ^ in2[25];
    assign G[99] = in1[24] & in2[24];
    assign P[99] = in1[24] ^ in2[24];
    assign G[100] = in1[23] & in2[23];
    assign P[100] = in1[23] ^ in2[23];
    assign G[101] = in1[22] & in2[22];
    assign P[101] = in1[22] ^ in2[22];
    assign G[102] = in1[21] & in2[21];
    assign P[102] = in1[21] ^ in2[21];
    assign G[103] = in1[20] & in2[20];
    assign P[103] = in1[20] ^ in2[20];
    assign G[104] = in1[19] & in2[19];
    assign P[104] = in1[19] ^ in2[19];
    assign G[105] = in1[18] & in2[18];
    assign P[105] = in1[18] ^ in2[18];
    assign G[106] = in1[17] & in2[17];
    assign P[106] = in1[17] ^ in2[17];
    assign G[107] = in1[16] & in2[16];
    assign P[107] = in1[16] ^ in2[16];
    assign G[108] = in1[15] & in2[15];
    assign P[108] = in1[15] ^ in2[15];
    assign G[109] = in1[14] & in2[14];
    assign P[109] = in1[14] ^ in2[14];
    assign G[110] = in1[13] & in2[13];
    assign P[110] = in1[13] ^ in2[13];
    assign G[111] = in1[12] & in2[12];
    assign P[111] = in1[12] ^ in2[12];
    assign G[112] = in1[11] & in2[11];
    assign P[112] = in1[11] ^ in2[11];
    assign G[113] = in1[10] & in2[10];
    assign P[113] = in1[10] ^ in2[10];
    assign G[114] = in1[9] & in2[9];
    assign P[114] = in1[9] ^ in2[9];
    assign G[115] = in1[8] & in2[8];
    assign P[115] = in1[8] ^ in2[8];
    assign G[116] = in1[7] & in2[7];
    assign P[116] = in1[7] ^ in2[7];
    assign G[117] = in1[6] & in2[6];
    assign P[117] = in1[6] ^ in2[6];
    assign G[118] = in1[5] & in2[5];
    assign P[118] = in1[5] ^ in2[5];
    assign G[119] = in1[4] & in2[4];
    assign P[119] = in1[4] ^ in2[4];
    assign G[120] = in1[3] & in2[3];
    assign P[120] = in1[3] ^ in2[3];
    assign G[121] = in1[2] & in2[2];
    assign P[121] = in1[2] ^ in2[2];
    assign G[122] = in1[1] & in2[1];
    assign P[122] = in1[1] ^ in2[1];
    assign G[123] = in1[0] & in2[0];
    assign P[123] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign cout = G[123] | (P[123] & C[123]);
    assign sum = P ^ C;
endmodule

module CLA_123(output [122:0] sum, output cout, input [122:0] in1, input [122:0] in2);

    wire[122:0] G;
    wire[122:0] C;
    wire[122:0] P;

    assign G[0] = in1[122] & in2[122];
    assign P[0] = in1[122] ^ in2[122];
    assign G[1] = in1[121] & in2[121];
    assign P[1] = in1[121] ^ in2[121];
    assign G[2] = in1[120] & in2[120];
    assign P[2] = in1[120] ^ in2[120];
    assign G[3] = in1[119] & in2[119];
    assign P[3] = in1[119] ^ in2[119];
    assign G[4] = in1[118] & in2[118];
    assign P[4] = in1[118] ^ in2[118];
    assign G[5] = in1[117] & in2[117];
    assign P[5] = in1[117] ^ in2[117];
    assign G[6] = in1[116] & in2[116];
    assign P[6] = in1[116] ^ in2[116];
    assign G[7] = in1[115] & in2[115];
    assign P[7] = in1[115] ^ in2[115];
    assign G[8] = in1[114] & in2[114];
    assign P[8] = in1[114] ^ in2[114];
    assign G[9] = in1[113] & in2[113];
    assign P[9] = in1[113] ^ in2[113];
    assign G[10] = in1[112] & in2[112];
    assign P[10] = in1[112] ^ in2[112];
    assign G[11] = in1[111] & in2[111];
    assign P[11] = in1[111] ^ in2[111];
    assign G[12] = in1[110] & in2[110];
    assign P[12] = in1[110] ^ in2[110];
    assign G[13] = in1[109] & in2[109];
    assign P[13] = in1[109] ^ in2[109];
    assign G[14] = in1[108] & in2[108];
    assign P[14] = in1[108] ^ in2[108];
    assign G[15] = in1[107] & in2[107];
    assign P[15] = in1[107] ^ in2[107];
    assign G[16] = in1[106] & in2[106];
    assign P[16] = in1[106] ^ in2[106];
    assign G[17] = in1[105] & in2[105];
    assign P[17] = in1[105] ^ in2[105];
    assign G[18] = in1[104] & in2[104];
    assign P[18] = in1[104] ^ in2[104];
    assign G[19] = in1[103] & in2[103];
    assign P[19] = in1[103] ^ in2[103];
    assign G[20] = in1[102] & in2[102];
    assign P[20] = in1[102] ^ in2[102];
    assign G[21] = in1[101] & in2[101];
    assign P[21] = in1[101] ^ in2[101];
    assign G[22] = in1[100] & in2[100];
    assign P[22] = in1[100] ^ in2[100];
    assign G[23] = in1[99] & in2[99];
    assign P[23] = in1[99] ^ in2[99];
    assign G[24] = in1[98] & in2[98];
    assign P[24] = in1[98] ^ in2[98];
    assign G[25] = in1[97] & in2[97];
    assign P[25] = in1[97] ^ in2[97];
    assign G[26] = in1[96] & in2[96];
    assign P[26] = in1[96] ^ in2[96];
    assign G[27] = in1[95] & in2[95];
    assign P[27] = in1[95] ^ in2[95];
    assign G[28] = in1[94] & in2[94];
    assign P[28] = in1[94] ^ in2[94];
    assign G[29] = in1[93] & in2[93];
    assign P[29] = in1[93] ^ in2[93];
    assign G[30] = in1[92] & in2[92];
    assign P[30] = in1[92] ^ in2[92];
    assign G[31] = in1[91] & in2[91];
    assign P[31] = in1[91] ^ in2[91];
    assign G[32] = in1[90] & in2[90];
    assign P[32] = in1[90] ^ in2[90];
    assign G[33] = in1[89] & in2[89];
    assign P[33] = in1[89] ^ in2[89];
    assign G[34] = in1[88] & in2[88];
    assign P[34] = in1[88] ^ in2[88];
    assign G[35] = in1[87] & in2[87];
    assign P[35] = in1[87] ^ in2[87];
    assign G[36] = in1[86] & in2[86];
    assign P[36] = in1[86] ^ in2[86];
    assign G[37] = in1[85] & in2[85];
    assign P[37] = in1[85] ^ in2[85];
    assign G[38] = in1[84] & in2[84];
    assign P[38] = in1[84] ^ in2[84];
    assign G[39] = in1[83] & in2[83];
    assign P[39] = in1[83] ^ in2[83];
    assign G[40] = in1[82] & in2[82];
    assign P[40] = in1[82] ^ in2[82];
    assign G[41] = in1[81] & in2[81];
    assign P[41] = in1[81] ^ in2[81];
    assign G[42] = in1[80] & in2[80];
    assign P[42] = in1[80] ^ in2[80];
    assign G[43] = in1[79] & in2[79];
    assign P[43] = in1[79] ^ in2[79];
    assign G[44] = in1[78] & in2[78];
    assign P[44] = in1[78] ^ in2[78];
    assign G[45] = in1[77] & in2[77];
    assign P[45] = in1[77] ^ in2[77];
    assign G[46] = in1[76] & in2[76];
    assign P[46] = in1[76] ^ in2[76];
    assign G[47] = in1[75] & in2[75];
    assign P[47] = in1[75] ^ in2[75];
    assign G[48] = in1[74] & in2[74];
    assign P[48] = in1[74] ^ in2[74];
    assign G[49] = in1[73] & in2[73];
    assign P[49] = in1[73] ^ in2[73];
    assign G[50] = in1[72] & in2[72];
    assign P[50] = in1[72] ^ in2[72];
    assign G[51] = in1[71] & in2[71];
    assign P[51] = in1[71] ^ in2[71];
    assign G[52] = in1[70] & in2[70];
    assign P[52] = in1[70] ^ in2[70];
    assign G[53] = in1[69] & in2[69];
    assign P[53] = in1[69] ^ in2[69];
    assign G[54] = in1[68] & in2[68];
    assign P[54] = in1[68] ^ in2[68];
    assign G[55] = in1[67] & in2[67];
    assign P[55] = in1[67] ^ in2[67];
    assign G[56] = in1[66] & in2[66];
    assign P[56] = in1[66] ^ in2[66];
    assign G[57] = in1[65] & in2[65];
    assign P[57] = in1[65] ^ in2[65];
    assign G[58] = in1[64] & in2[64];
    assign P[58] = in1[64] ^ in2[64];
    assign G[59] = in1[63] & in2[63];
    assign P[59] = in1[63] ^ in2[63];
    assign G[60] = in1[62] & in2[62];
    assign P[60] = in1[62] ^ in2[62];
    assign G[61] = in1[61] & in2[61];
    assign P[61] = in1[61] ^ in2[61];
    assign G[62] = in1[60] & in2[60];
    assign P[62] = in1[60] ^ in2[60];
    assign G[63] = in1[59] & in2[59];
    assign P[63] = in1[59] ^ in2[59];
    assign G[64] = in1[58] & in2[58];
    assign P[64] = in1[58] ^ in2[58];
    assign G[65] = in1[57] & in2[57];
    assign P[65] = in1[57] ^ in2[57];
    assign G[66] = in1[56] & in2[56];
    assign P[66] = in1[56] ^ in2[56];
    assign G[67] = in1[55] & in2[55];
    assign P[67] = in1[55] ^ in2[55];
    assign G[68] = in1[54] & in2[54];
    assign P[68] = in1[54] ^ in2[54];
    assign G[69] = in1[53] & in2[53];
    assign P[69] = in1[53] ^ in2[53];
    assign G[70] = in1[52] & in2[52];
    assign P[70] = in1[52] ^ in2[52];
    assign G[71] = in1[51] & in2[51];
    assign P[71] = in1[51] ^ in2[51];
    assign G[72] = in1[50] & in2[50];
    assign P[72] = in1[50] ^ in2[50];
    assign G[73] = in1[49] & in2[49];
    assign P[73] = in1[49] ^ in2[49];
    assign G[74] = in1[48] & in2[48];
    assign P[74] = in1[48] ^ in2[48];
    assign G[75] = in1[47] & in2[47];
    assign P[75] = in1[47] ^ in2[47];
    assign G[76] = in1[46] & in2[46];
    assign P[76] = in1[46] ^ in2[46];
    assign G[77] = in1[45] & in2[45];
    assign P[77] = in1[45] ^ in2[45];
    assign G[78] = in1[44] & in2[44];
    assign P[78] = in1[44] ^ in2[44];
    assign G[79] = in1[43] & in2[43];
    assign P[79] = in1[43] ^ in2[43];
    assign G[80] = in1[42] & in2[42];
    assign P[80] = in1[42] ^ in2[42];
    assign G[81] = in1[41] & in2[41];
    assign P[81] = in1[41] ^ in2[41];
    assign G[82] = in1[40] & in2[40];
    assign P[82] = in1[40] ^ in2[40];
    assign G[83] = in1[39] & in2[39];
    assign P[83] = in1[39] ^ in2[39];
    assign G[84] = in1[38] & in2[38];
    assign P[84] = in1[38] ^ in2[38];
    assign G[85] = in1[37] & in2[37];
    assign P[85] = in1[37] ^ in2[37];
    assign G[86] = in1[36] & in2[36];
    assign P[86] = in1[36] ^ in2[36];
    assign G[87] = in1[35] & in2[35];
    assign P[87] = in1[35] ^ in2[35];
    assign G[88] = in1[34] & in2[34];
    assign P[88] = in1[34] ^ in2[34];
    assign G[89] = in1[33] & in2[33];
    assign P[89] = in1[33] ^ in2[33];
    assign G[90] = in1[32] & in2[32];
    assign P[90] = in1[32] ^ in2[32];
    assign G[91] = in1[31] & in2[31];
    assign P[91] = in1[31] ^ in2[31];
    assign G[92] = in1[30] & in2[30];
    assign P[92] = in1[30] ^ in2[30];
    assign G[93] = in1[29] & in2[29];
    assign P[93] = in1[29] ^ in2[29];
    assign G[94] = in1[28] & in2[28];
    assign P[94] = in1[28] ^ in2[28];
    assign G[95] = in1[27] & in2[27];
    assign P[95] = in1[27] ^ in2[27];
    assign G[96] = in1[26] & in2[26];
    assign P[96] = in1[26] ^ in2[26];
    assign G[97] = in1[25] & in2[25];
    assign P[97] = in1[25] ^ in2[25];
    assign G[98] = in1[24] & in2[24];
    assign P[98] = in1[24] ^ in2[24];
    assign G[99] = in1[23] & in2[23];
    assign P[99] = in1[23] ^ in2[23];
    assign G[100] = in1[22] & in2[22];
    assign P[100] = in1[22] ^ in2[22];
    assign G[101] = in1[21] & in2[21];
    assign P[101] = in1[21] ^ in2[21];
    assign G[102] = in1[20] & in2[20];
    assign P[102] = in1[20] ^ in2[20];
    assign G[103] = in1[19] & in2[19];
    assign P[103] = in1[19] ^ in2[19];
    assign G[104] = in1[18] & in2[18];
    assign P[104] = in1[18] ^ in2[18];
    assign G[105] = in1[17] & in2[17];
    assign P[105] = in1[17] ^ in2[17];
    assign G[106] = in1[16] & in2[16];
    assign P[106] = in1[16] ^ in2[16];
    assign G[107] = in1[15] & in2[15];
    assign P[107] = in1[15] ^ in2[15];
    assign G[108] = in1[14] & in2[14];
    assign P[108] = in1[14] ^ in2[14];
    assign G[109] = in1[13] & in2[13];
    assign P[109] = in1[13] ^ in2[13];
    assign G[110] = in1[12] & in2[12];
    assign P[110] = in1[12] ^ in2[12];
    assign G[111] = in1[11] & in2[11];
    assign P[111] = in1[11] ^ in2[11];
    assign G[112] = in1[10] & in2[10];
    assign P[112] = in1[10] ^ in2[10];
    assign G[113] = in1[9] & in2[9];
    assign P[113] = in1[9] ^ in2[9];
    assign G[114] = in1[8] & in2[8];
    assign P[114] = in1[8] ^ in2[8];
    assign G[115] = in1[7] & in2[7];
    assign P[115] = in1[7] ^ in2[7];
    assign G[116] = in1[6] & in2[6];
    assign P[116] = in1[6] ^ in2[6];
    assign G[117] = in1[5] & in2[5];
    assign P[117] = in1[5] ^ in2[5];
    assign G[118] = in1[4] & in2[4];
    assign P[118] = in1[4] ^ in2[4];
    assign G[119] = in1[3] & in2[3];
    assign P[119] = in1[3] ^ in2[3];
    assign G[120] = in1[2] & in2[2];
    assign P[120] = in1[2] ^ in2[2];
    assign G[121] = in1[1] & in2[1];
    assign P[121] = in1[1] ^ in2[1];
    assign G[122] = in1[0] & in2[0];
    assign P[122] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign cout = G[122] | (P[122] & C[122]);
    assign sum = P ^ C;
endmodule

module CLA_122(output [121:0] sum, output cout, input [121:0] in1, input [121:0] in2);

    wire[121:0] G;
    wire[121:0] C;
    wire[121:0] P;

    assign G[0] = in1[121] & in2[121];
    assign P[0] = in1[121] ^ in2[121];
    assign G[1] = in1[120] & in2[120];
    assign P[1] = in1[120] ^ in2[120];
    assign G[2] = in1[119] & in2[119];
    assign P[2] = in1[119] ^ in2[119];
    assign G[3] = in1[118] & in2[118];
    assign P[3] = in1[118] ^ in2[118];
    assign G[4] = in1[117] & in2[117];
    assign P[4] = in1[117] ^ in2[117];
    assign G[5] = in1[116] & in2[116];
    assign P[5] = in1[116] ^ in2[116];
    assign G[6] = in1[115] & in2[115];
    assign P[6] = in1[115] ^ in2[115];
    assign G[7] = in1[114] & in2[114];
    assign P[7] = in1[114] ^ in2[114];
    assign G[8] = in1[113] & in2[113];
    assign P[8] = in1[113] ^ in2[113];
    assign G[9] = in1[112] & in2[112];
    assign P[9] = in1[112] ^ in2[112];
    assign G[10] = in1[111] & in2[111];
    assign P[10] = in1[111] ^ in2[111];
    assign G[11] = in1[110] & in2[110];
    assign P[11] = in1[110] ^ in2[110];
    assign G[12] = in1[109] & in2[109];
    assign P[12] = in1[109] ^ in2[109];
    assign G[13] = in1[108] & in2[108];
    assign P[13] = in1[108] ^ in2[108];
    assign G[14] = in1[107] & in2[107];
    assign P[14] = in1[107] ^ in2[107];
    assign G[15] = in1[106] & in2[106];
    assign P[15] = in1[106] ^ in2[106];
    assign G[16] = in1[105] & in2[105];
    assign P[16] = in1[105] ^ in2[105];
    assign G[17] = in1[104] & in2[104];
    assign P[17] = in1[104] ^ in2[104];
    assign G[18] = in1[103] & in2[103];
    assign P[18] = in1[103] ^ in2[103];
    assign G[19] = in1[102] & in2[102];
    assign P[19] = in1[102] ^ in2[102];
    assign G[20] = in1[101] & in2[101];
    assign P[20] = in1[101] ^ in2[101];
    assign G[21] = in1[100] & in2[100];
    assign P[21] = in1[100] ^ in2[100];
    assign G[22] = in1[99] & in2[99];
    assign P[22] = in1[99] ^ in2[99];
    assign G[23] = in1[98] & in2[98];
    assign P[23] = in1[98] ^ in2[98];
    assign G[24] = in1[97] & in2[97];
    assign P[24] = in1[97] ^ in2[97];
    assign G[25] = in1[96] & in2[96];
    assign P[25] = in1[96] ^ in2[96];
    assign G[26] = in1[95] & in2[95];
    assign P[26] = in1[95] ^ in2[95];
    assign G[27] = in1[94] & in2[94];
    assign P[27] = in1[94] ^ in2[94];
    assign G[28] = in1[93] & in2[93];
    assign P[28] = in1[93] ^ in2[93];
    assign G[29] = in1[92] & in2[92];
    assign P[29] = in1[92] ^ in2[92];
    assign G[30] = in1[91] & in2[91];
    assign P[30] = in1[91] ^ in2[91];
    assign G[31] = in1[90] & in2[90];
    assign P[31] = in1[90] ^ in2[90];
    assign G[32] = in1[89] & in2[89];
    assign P[32] = in1[89] ^ in2[89];
    assign G[33] = in1[88] & in2[88];
    assign P[33] = in1[88] ^ in2[88];
    assign G[34] = in1[87] & in2[87];
    assign P[34] = in1[87] ^ in2[87];
    assign G[35] = in1[86] & in2[86];
    assign P[35] = in1[86] ^ in2[86];
    assign G[36] = in1[85] & in2[85];
    assign P[36] = in1[85] ^ in2[85];
    assign G[37] = in1[84] & in2[84];
    assign P[37] = in1[84] ^ in2[84];
    assign G[38] = in1[83] & in2[83];
    assign P[38] = in1[83] ^ in2[83];
    assign G[39] = in1[82] & in2[82];
    assign P[39] = in1[82] ^ in2[82];
    assign G[40] = in1[81] & in2[81];
    assign P[40] = in1[81] ^ in2[81];
    assign G[41] = in1[80] & in2[80];
    assign P[41] = in1[80] ^ in2[80];
    assign G[42] = in1[79] & in2[79];
    assign P[42] = in1[79] ^ in2[79];
    assign G[43] = in1[78] & in2[78];
    assign P[43] = in1[78] ^ in2[78];
    assign G[44] = in1[77] & in2[77];
    assign P[44] = in1[77] ^ in2[77];
    assign G[45] = in1[76] & in2[76];
    assign P[45] = in1[76] ^ in2[76];
    assign G[46] = in1[75] & in2[75];
    assign P[46] = in1[75] ^ in2[75];
    assign G[47] = in1[74] & in2[74];
    assign P[47] = in1[74] ^ in2[74];
    assign G[48] = in1[73] & in2[73];
    assign P[48] = in1[73] ^ in2[73];
    assign G[49] = in1[72] & in2[72];
    assign P[49] = in1[72] ^ in2[72];
    assign G[50] = in1[71] & in2[71];
    assign P[50] = in1[71] ^ in2[71];
    assign G[51] = in1[70] & in2[70];
    assign P[51] = in1[70] ^ in2[70];
    assign G[52] = in1[69] & in2[69];
    assign P[52] = in1[69] ^ in2[69];
    assign G[53] = in1[68] & in2[68];
    assign P[53] = in1[68] ^ in2[68];
    assign G[54] = in1[67] & in2[67];
    assign P[54] = in1[67] ^ in2[67];
    assign G[55] = in1[66] & in2[66];
    assign P[55] = in1[66] ^ in2[66];
    assign G[56] = in1[65] & in2[65];
    assign P[56] = in1[65] ^ in2[65];
    assign G[57] = in1[64] & in2[64];
    assign P[57] = in1[64] ^ in2[64];
    assign G[58] = in1[63] & in2[63];
    assign P[58] = in1[63] ^ in2[63];
    assign G[59] = in1[62] & in2[62];
    assign P[59] = in1[62] ^ in2[62];
    assign G[60] = in1[61] & in2[61];
    assign P[60] = in1[61] ^ in2[61];
    assign G[61] = in1[60] & in2[60];
    assign P[61] = in1[60] ^ in2[60];
    assign G[62] = in1[59] & in2[59];
    assign P[62] = in1[59] ^ in2[59];
    assign G[63] = in1[58] & in2[58];
    assign P[63] = in1[58] ^ in2[58];
    assign G[64] = in1[57] & in2[57];
    assign P[64] = in1[57] ^ in2[57];
    assign G[65] = in1[56] & in2[56];
    assign P[65] = in1[56] ^ in2[56];
    assign G[66] = in1[55] & in2[55];
    assign P[66] = in1[55] ^ in2[55];
    assign G[67] = in1[54] & in2[54];
    assign P[67] = in1[54] ^ in2[54];
    assign G[68] = in1[53] & in2[53];
    assign P[68] = in1[53] ^ in2[53];
    assign G[69] = in1[52] & in2[52];
    assign P[69] = in1[52] ^ in2[52];
    assign G[70] = in1[51] & in2[51];
    assign P[70] = in1[51] ^ in2[51];
    assign G[71] = in1[50] & in2[50];
    assign P[71] = in1[50] ^ in2[50];
    assign G[72] = in1[49] & in2[49];
    assign P[72] = in1[49] ^ in2[49];
    assign G[73] = in1[48] & in2[48];
    assign P[73] = in1[48] ^ in2[48];
    assign G[74] = in1[47] & in2[47];
    assign P[74] = in1[47] ^ in2[47];
    assign G[75] = in1[46] & in2[46];
    assign P[75] = in1[46] ^ in2[46];
    assign G[76] = in1[45] & in2[45];
    assign P[76] = in1[45] ^ in2[45];
    assign G[77] = in1[44] & in2[44];
    assign P[77] = in1[44] ^ in2[44];
    assign G[78] = in1[43] & in2[43];
    assign P[78] = in1[43] ^ in2[43];
    assign G[79] = in1[42] & in2[42];
    assign P[79] = in1[42] ^ in2[42];
    assign G[80] = in1[41] & in2[41];
    assign P[80] = in1[41] ^ in2[41];
    assign G[81] = in1[40] & in2[40];
    assign P[81] = in1[40] ^ in2[40];
    assign G[82] = in1[39] & in2[39];
    assign P[82] = in1[39] ^ in2[39];
    assign G[83] = in1[38] & in2[38];
    assign P[83] = in1[38] ^ in2[38];
    assign G[84] = in1[37] & in2[37];
    assign P[84] = in1[37] ^ in2[37];
    assign G[85] = in1[36] & in2[36];
    assign P[85] = in1[36] ^ in2[36];
    assign G[86] = in1[35] & in2[35];
    assign P[86] = in1[35] ^ in2[35];
    assign G[87] = in1[34] & in2[34];
    assign P[87] = in1[34] ^ in2[34];
    assign G[88] = in1[33] & in2[33];
    assign P[88] = in1[33] ^ in2[33];
    assign G[89] = in1[32] & in2[32];
    assign P[89] = in1[32] ^ in2[32];
    assign G[90] = in1[31] & in2[31];
    assign P[90] = in1[31] ^ in2[31];
    assign G[91] = in1[30] & in2[30];
    assign P[91] = in1[30] ^ in2[30];
    assign G[92] = in1[29] & in2[29];
    assign P[92] = in1[29] ^ in2[29];
    assign G[93] = in1[28] & in2[28];
    assign P[93] = in1[28] ^ in2[28];
    assign G[94] = in1[27] & in2[27];
    assign P[94] = in1[27] ^ in2[27];
    assign G[95] = in1[26] & in2[26];
    assign P[95] = in1[26] ^ in2[26];
    assign G[96] = in1[25] & in2[25];
    assign P[96] = in1[25] ^ in2[25];
    assign G[97] = in1[24] & in2[24];
    assign P[97] = in1[24] ^ in2[24];
    assign G[98] = in1[23] & in2[23];
    assign P[98] = in1[23] ^ in2[23];
    assign G[99] = in1[22] & in2[22];
    assign P[99] = in1[22] ^ in2[22];
    assign G[100] = in1[21] & in2[21];
    assign P[100] = in1[21] ^ in2[21];
    assign G[101] = in1[20] & in2[20];
    assign P[101] = in1[20] ^ in2[20];
    assign G[102] = in1[19] & in2[19];
    assign P[102] = in1[19] ^ in2[19];
    assign G[103] = in1[18] & in2[18];
    assign P[103] = in1[18] ^ in2[18];
    assign G[104] = in1[17] & in2[17];
    assign P[104] = in1[17] ^ in2[17];
    assign G[105] = in1[16] & in2[16];
    assign P[105] = in1[16] ^ in2[16];
    assign G[106] = in1[15] & in2[15];
    assign P[106] = in1[15] ^ in2[15];
    assign G[107] = in1[14] & in2[14];
    assign P[107] = in1[14] ^ in2[14];
    assign G[108] = in1[13] & in2[13];
    assign P[108] = in1[13] ^ in2[13];
    assign G[109] = in1[12] & in2[12];
    assign P[109] = in1[12] ^ in2[12];
    assign G[110] = in1[11] & in2[11];
    assign P[110] = in1[11] ^ in2[11];
    assign G[111] = in1[10] & in2[10];
    assign P[111] = in1[10] ^ in2[10];
    assign G[112] = in1[9] & in2[9];
    assign P[112] = in1[9] ^ in2[9];
    assign G[113] = in1[8] & in2[8];
    assign P[113] = in1[8] ^ in2[8];
    assign G[114] = in1[7] & in2[7];
    assign P[114] = in1[7] ^ in2[7];
    assign G[115] = in1[6] & in2[6];
    assign P[115] = in1[6] ^ in2[6];
    assign G[116] = in1[5] & in2[5];
    assign P[116] = in1[5] ^ in2[5];
    assign G[117] = in1[4] & in2[4];
    assign P[117] = in1[4] ^ in2[4];
    assign G[118] = in1[3] & in2[3];
    assign P[118] = in1[3] ^ in2[3];
    assign G[119] = in1[2] & in2[2];
    assign P[119] = in1[2] ^ in2[2];
    assign G[120] = in1[1] & in2[1];
    assign P[120] = in1[1] ^ in2[1];
    assign G[121] = in1[0] & in2[0];
    assign P[121] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign cout = G[121] | (P[121] & C[121]);
    assign sum = P ^ C;
endmodule

module CLA_121(output [120:0] sum, output cout, input [120:0] in1, input [120:0] in2);

    wire[120:0] G;
    wire[120:0] C;
    wire[120:0] P;

    assign G[0] = in1[120] & in2[120];
    assign P[0] = in1[120] ^ in2[120];
    assign G[1] = in1[119] & in2[119];
    assign P[1] = in1[119] ^ in2[119];
    assign G[2] = in1[118] & in2[118];
    assign P[2] = in1[118] ^ in2[118];
    assign G[3] = in1[117] & in2[117];
    assign P[3] = in1[117] ^ in2[117];
    assign G[4] = in1[116] & in2[116];
    assign P[4] = in1[116] ^ in2[116];
    assign G[5] = in1[115] & in2[115];
    assign P[5] = in1[115] ^ in2[115];
    assign G[6] = in1[114] & in2[114];
    assign P[6] = in1[114] ^ in2[114];
    assign G[7] = in1[113] & in2[113];
    assign P[7] = in1[113] ^ in2[113];
    assign G[8] = in1[112] & in2[112];
    assign P[8] = in1[112] ^ in2[112];
    assign G[9] = in1[111] & in2[111];
    assign P[9] = in1[111] ^ in2[111];
    assign G[10] = in1[110] & in2[110];
    assign P[10] = in1[110] ^ in2[110];
    assign G[11] = in1[109] & in2[109];
    assign P[11] = in1[109] ^ in2[109];
    assign G[12] = in1[108] & in2[108];
    assign P[12] = in1[108] ^ in2[108];
    assign G[13] = in1[107] & in2[107];
    assign P[13] = in1[107] ^ in2[107];
    assign G[14] = in1[106] & in2[106];
    assign P[14] = in1[106] ^ in2[106];
    assign G[15] = in1[105] & in2[105];
    assign P[15] = in1[105] ^ in2[105];
    assign G[16] = in1[104] & in2[104];
    assign P[16] = in1[104] ^ in2[104];
    assign G[17] = in1[103] & in2[103];
    assign P[17] = in1[103] ^ in2[103];
    assign G[18] = in1[102] & in2[102];
    assign P[18] = in1[102] ^ in2[102];
    assign G[19] = in1[101] & in2[101];
    assign P[19] = in1[101] ^ in2[101];
    assign G[20] = in1[100] & in2[100];
    assign P[20] = in1[100] ^ in2[100];
    assign G[21] = in1[99] & in2[99];
    assign P[21] = in1[99] ^ in2[99];
    assign G[22] = in1[98] & in2[98];
    assign P[22] = in1[98] ^ in2[98];
    assign G[23] = in1[97] & in2[97];
    assign P[23] = in1[97] ^ in2[97];
    assign G[24] = in1[96] & in2[96];
    assign P[24] = in1[96] ^ in2[96];
    assign G[25] = in1[95] & in2[95];
    assign P[25] = in1[95] ^ in2[95];
    assign G[26] = in1[94] & in2[94];
    assign P[26] = in1[94] ^ in2[94];
    assign G[27] = in1[93] & in2[93];
    assign P[27] = in1[93] ^ in2[93];
    assign G[28] = in1[92] & in2[92];
    assign P[28] = in1[92] ^ in2[92];
    assign G[29] = in1[91] & in2[91];
    assign P[29] = in1[91] ^ in2[91];
    assign G[30] = in1[90] & in2[90];
    assign P[30] = in1[90] ^ in2[90];
    assign G[31] = in1[89] & in2[89];
    assign P[31] = in1[89] ^ in2[89];
    assign G[32] = in1[88] & in2[88];
    assign P[32] = in1[88] ^ in2[88];
    assign G[33] = in1[87] & in2[87];
    assign P[33] = in1[87] ^ in2[87];
    assign G[34] = in1[86] & in2[86];
    assign P[34] = in1[86] ^ in2[86];
    assign G[35] = in1[85] & in2[85];
    assign P[35] = in1[85] ^ in2[85];
    assign G[36] = in1[84] & in2[84];
    assign P[36] = in1[84] ^ in2[84];
    assign G[37] = in1[83] & in2[83];
    assign P[37] = in1[83] ^ in2[83];
    assign G[38] = in1[82] & in2[82];
    assign P[38] = in1[82] ^ in2[82];
    assign G[39] = in1[81] & in2[81];
    assign P[39] = in1[81] ^ in2[81];
    assign G[40] = in1[80] & in2[80];
    assign P[40] = in1[80] ^ in2[80];
    assign G[41] = in1[79] & in2[79];
    assign P[41] = in1[79] ^ in2[79];
    assign G[42] = in1[78] & in2[78];
    assign P[42] = in1[78] ^ in2[78];
    assign G[43] = in1[77] & in2[77];
    assign P[43] = in1[77] ^ in2[77];
    assign G[44] = in1[76] & in2[76];
    assign P[44] = in1[76] ^ in2[76];
    assign G[45] = in1[75] & in2[75];
    assign P[45] = in1[75] ^ in2[75];
    assign G[46] = in1[74] & in2[74];
    assign P[46] = in1[74] ^ in2[74];
    assign G[47] = in1[73] & in2[73];
    assign P[47] = in1[73] ^ in2[73];
    assign G[48] = in1[72] & in2[72];
    assign P[48] = in1[72] ^ in2[72];
    assign G[49] = in1[71] & in2[71];
    assign P[49] = in1[71] ^ in2[71];
    assign G[50] = in1[70] & in2[70];
    assign P[50] = in1[70] ^ in2[70];
    assign G[51] = in1[69] & in2[69];
    assign P[51] = in1[69] ^ in2[69];
    assign G[52] = in1[68] & in2[68];
    assign P[52] = in1[68] ^ in2[68];
    assign G[53] = in1[67] & in2[67];
    assign P[53] = in1[67] ^ in2[67];
    assign G[54] = in1[66] & in2[66];
    assign P[54] = in1[66] ^ in2[66];
    assign G[55] = in1[65] & in2[65];
    assign P[55] = in1[65] ^ in2[65];
    assign G[56] = in1[64] & in2[64];
    assign P[56] = in1[64] ^ in2[64];
    assign G[57] = in1[63] & in2[63];
    assign P[57] = in1[63] ^ in2[63];
    assign G[58] = in1[62] & in2[62];
    assign P[58] = in1[62] ^ in2[62];
    assign G[59] = in1[61] & in2[61];
    assign P[59] = in1[61] ^ in2[61];
    assign G[60] = in1[60] & in2[60];
    assign P[60] = in1[60] ^ in2[60];
    assign G[61] = in1[59] & in2[59];
    assign P[61] = in1[59] ^ in2[59];
    assign G[62] = in1[58] & in2[58];
    assign P[62] = in1[58] ^ in2[58];
    assign G[63] = in1[57] & in2[57];
    assign P[63] = in1[57] ^ in2[57];
    assign G[64] = in1[56] & in2[56];
    assign P[64] = in1[56] ^ in2[56];
    assign G[65] = in1[55] & in2[55];
    assign P[65] = in1[55] ^ in2[55];
    assign G[66] = in1[54] & in2[54];
    assign P[66] = in1[54] ^ in2[54];
    assign G[67] = in1[53] & in2[53];
    assign P[67] = in1[53] ^ in2[53];
    assign G[68] = in1[52] & in2[52];
    assign P[68] = in1[52] ^ in2[52];
    assign G[69] = in1[51] & in2[51];
    assign P[69] = in1[51] ^ in2[51];
    assign G[70] = in1[50] & in2[50];
    assign P[70] = in1[50] ^ in2[50];
    assign G[71] = in1[49] & in2[49];
    assign P[71] = in1[49] ^ in2[49];
    assign G[72] = in1[48] & in2[48];
    assign P[72] = in1[48] ^ in2[48];
    assign G[73] = in1[47] & in2[47];
    assign P[73] = in1[47] ^ in2[47];
    assign G[74] = in1[46] & in2[46];
    assign P[74] = in1[46] ^ in2[46];
    assign G[75] = in1[45] & in2[45];
    assign P[75] = in1[45] ^ in2[45];
    assign G[76] = in1[44] & in2[44];
    assign P[76] = in1[44] ^ in2[44];
    assign G[77] = in1[43] & in2[43];
    assign P[77] = in1[43] ^ in2[43];
    assign G[78] = in1[42] & in2[42];
    assign P[78] = in1[42] ^ in2[42];
    assign G[79] = in1[41] & in2[41];
    assign P[79] = in1[41] ^ in2[41];
    assign G[80] = in1[40] & in2[40];
    assign P[80] = in1[40] ^ in2[40];
    assign G[81] = in1[39] & in2[39];
    assign P[81] = in1[39] ^ in2[39];
    assign G[82] = in1[38] & in2[38];
    assign P[82] = in1[38] ^ in2[38];
    assign G[83] = in1[37] & in2[37];
    assign P[83] = in1[37] ^ in2[37];
    assign G[84] = in1[36] & in2[36];
    assign P[84] = in1[36] ^ in2[36];
    assign G[85] = in1[35] & in2[35];
    assign P[85] = in1[35] ^ in2[35];
    assign G[86] = in1[34] & in2[34];
    assign P[86] = in1[34] ^ in2[34];
    assign G[87] = in1[33] & in2[33];
    assign P[87] = in1[33] ^ in2[33];
    assign G[88] = in1[32] & in2[32];
    assign P[88] = in1[32] ^ in2[32];
    assign G[89] = in1[31] & in2[31];
    assign P[89] = in1[31] ^ in2[31];
    assign G[90] = in1[30] & in2[30];
    assign P[90] = in1[30] ^ in2[30];
    assign G[91] = in1[29] & in2[29];
    assign P[91] = in1[29] ^ in2[29];
    assign G[92] = in1[28] & in2[28];
    assign P[92] = in1[28] ^ in2[28];
    assign G[93] = in1[27] & in2[27];
    assign P[93] = in1[27] ^ in2[27];
    assign G[94] = in1[26] & in2[26];
    assign P[94] = in1[26] ^ in2[26];
    assign G[95] = in1[25] & in2[25];
    assign P[95] = in1[25] ^ in2[25];
    assign G[96] = in1[24] & in2[24];
    assign P[96] = in1[24] ^ in2[24];
    assign G[97] = in1[23] & in2[23];
    assign P[97] = in1[23] ^ in2[23];
    assign G[98] = in1[22] & in2[22];
    assign P[98] = in1[22] ^ in2[22];
    assign G[99] = in1[21] & in2[21];
    assign P[99] = in1[21] ^ in2[21];
    assign G[100] = in1[20] & in2[20];
    assign P[100] = in1[20] ^ in2[20];
    assign G[101] = in1[19] & in2[19];
    assign P[101] = in1[19] ^ in2[19];
    assign G[102] = in1[18] & in2[18];
    assign P[102] = in1[18] ^ in2[18];
    assign G[103] = in1[17] & in2[17];
    assign P[103] = in1[17] ^ in2[17];
    assign G[104] = in1[16] & in2[16];
    assign P[104] = in1[16] ^ in2[16];
    assign G[105] = in1[15] & in2[15];
    assign P[105] = in1[15] ^ in2[15];
    assign G[106] = in1[14] & in2[14];
    assign P[106] = in1[14] ^ in2[14];
    assign G[107] = in1[13] & in2[13];
    assign P[107] = in1[13] ^ in2[13];
    assign G[108] = in1[12] & in2[12];
    assign P[108] = in1[12] ^ in2[12];
    assign G[109] = in1[11] & in2[11];
    assign P[109] = in1[11] ^ in2[11];
    assign G[110] = in1[10] & in2[10];
    assign P[110] = in1[10] ^ in2[10];
    assign G[111] = in1[9] & in2[9];
    assign P[111] = in1[9] ^ in2[9];
    assign G[112] = in1[8] & in2[8];
    assign P[112] = in1[8] ^ in2[8];
    assign G[113] = in1[7] & in2[7];
    assign P[113] = in1[7] ^ in2[7];
    assign G[114] = in1[6] & in2[6];
    assign P[114] = in1[6] ^ in2[6];
    assign G[115] = in1[5] & in2[5];
    assign P[115] = in1[5] ^ in2[5];
    assign G[116] = in1[4] & in2[4];
    assign P[116] = in1[4] ^ in2[4];
    assign G[117] = in1[3] & in2[3];
    assign P[117] = in1[3] ^ in2[3];
    assign G[118] = in1[2] & in2[2];
    assign P[118] = in1[2] ^ in2[2];
    assign G[119] = in1[1] & in2[1];
    assign P[119] = in1[1] ^ in2[1];
    assign G[120] = in1[0] & in2[0];
    assign P[120] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign cout = G[120] | (P[120] & C[120]);
    assign sum = P ^ C;
endmodule

module CLA_120(output [119:0] sum, output cout, input [119:0] in1, input [119:0] in2);

    wire[119:0] G;
    wire[119:0] C;
    wire[119:0] P;

    assign G[0] = in1[119] & in2[119];
    assign P[0] = in1[119] ^ in2[119];
    assign G[1] = in1[118] & in2[118];
    assign P[1] = in1[118] ^ in2[118];
    assign G[2] = in1[117] & in2[117];
    assign P[2] = in1[117] ^ in2[117];
    assign G[3] = in1[116] & in2[116];
    assign P[3] = in1[116] ^ in2[116];
    assign G[4] = in1[115] & in2[115];
    assign P[4] = in1[115] ^ in2[115];
    assign G[5] = in1[114] & in2[114];
    assign P[5] = in1[114] ^ in2[114];
    assign G[6] = in1[113] & in2[113];
    assign P[6] = in1[113] ^ in2[113];
    assign G[7] = in1[112] & in2[112];
    assign P[7] = in1[112] ^ in2[112];
    assign G[8] = in1[111] & in2[111];
    assign P[8] = in1[111] ^ in2[111];
    assign G[9] = in1[110] & in2[110];
    assign P[9] = in1[110] ^ in2[110];
    assign G[10] = in1[109] & in2[109];
    assign P[10] = in1[109] ^ in2[109];
    assign G[11] = in1[108] & in2[108];
    assign P[11] = in1[108] ^ in2[108];
    assign G[12] = in1[107] & in2[107];
    assign P[12] = in1[107] ^ in2[107];
    assign G[13] = in1[106] & in2[106];
    assign P[13] = in1[106] ^ in2[106];
    assign G[14] = in1[105] & in2[105];
    assign P[14] = in1[105] ^ in2[105];
    assign G[15] = in1[104] & in2[104];
    assign P[15] = in1[104] ^ in2[104];
    assign G[16] = in1[103] & in2[103];
    assign P[16] = in1[103] ^ in2[103];
    assign G[17] = in1[102] & in2[102];
    assign P[17] = in1[102] ^ in2[102];
    assign G[18] = in1[101] & in2[101];
    assign P[18] = in1[101] ^ in2[101];
    assign G[19] = in1[100] & in2[100];
    assign P[19] = in1[100] ^ in2[100];
    assign G[20] = in1[99] & in2[99];
    assign P[20] = in1[99] ^ in2[99];
    assign G[21] = in1[98] & in2[98];
    assign P[21] = in1[98] ^ in2[98];
    assign G[22] = in1[97] & in2[97];
    assign P[22] = in1[97] ^ in2[97];
    assign G[23] = in1[96] & in2[96];
    assign P[23] = in1[96] ^ in2[96];
    assign G[24] = in1[95] & in2[95];
    assign P[24] = in1[95] ^ in2[95];
    assign G[25] = in1[94] & in2[94];
    assign P[25] = in1[94] ^ in2[94];
    assign G[26] = in1[93] & in2[93];
    assign P[26] = in1[93] ^ in2[93];
    assign G[27] = in1[92] & in2[92];
    assign P[27] = in1[92] ^ in2[92];
    assign G[28] = in1[91] & in2[91];
    assign P[28] = in1[91] ^ in2[91];
    assign G[29] = in1[90] & in2[90];
    assign P[29] = in1[90] ^ in2[90];
    assign G[30] = in1[89] & in2[89];
    assign P[30] = in1[89] ^ in2[89];
    assign G[31] = in1[88] & in2[88];
    assign P[31] = in1[88] ^ in2[88];
    assign G[32] = in1[87] & in2[87];
    assign P[32] = in1[87] ^ in2[87];
    assign G[33] = in1[86] & in2[86];
    assign P[33] = in1[86] ^ in2[86];
    assign G[34] = in1[85] & in2[85];
    assign P[34] = in1[85] ^ in2[85];
    assign G[35] = in1[84] & in2[84];
    assign P[35] = in1[84] ^ in2[84];
    assign G[36] = in1[83] & in2[83];
    assign P[36] = in1[83] ^ in2[83];
    assign G[37] = in1[82] & in2[82];
    assign P[37] = in1[82] ^ in2[82];
    assign G[38] = in1[81] & in2[81];
    assign P[38] = in1[81] ^ in2[81];
    assign G[39] = in1[80] & in2[80];
    assign P[39] = in1[80] ^ in2[80];
    assign G[40] = in1[79] & in2[79];
    assign P[40] = in1[79] ^ in2[79];
    assign G[41] = in1[78] & in2[78];
    assign P[41] = in1[78] ^ in2[78];
    assign G[42] = in1[77] & in2[77];
    assign P[42] = in1[77] ^ in2[77];
    assign G[43] = in1[76] & in2[76];
    assign P[43] = in1[76] ^ in2[76];
    assign G[44] = in1[75] & in2[75];
    assign P[44] = in1[75] ^ in2[75];
    assign G[45] = in1[74] & in2[74];
    assign P[45] = in1[74] ^ in2[74];
    assign G[46] = in1[73] & in2[73];
    assign P[46] = in1[73] ^ in2[73];
    assign G[47] = in1[72] & in2[72];
    assign P[47] = in1[72] ^ in2[72];
    assign G[48] = in1[71] & in2[71];
    assign P[48] = in1[71] ^ in2[71];
    assign G[49] = in1[70] & in2[70];
    assign P[49] = in1[70] ^ in2[70];
    assign G[50] = in1[69] & in2[69];
    assign P[50] = in1[69] ^ in2[69];
    assign G[51] = in1[68] & in2[68];
    assign P[51] = in1[68] ^ in2[68];
    assign G[52] = in1[67] & in2[67];
    assign P[52] = in1[67] ^ in2[67];
    assign G[53] = in1[66] & in2[66];
    assign P[53] = in1[66] ^ in2[66];
    assign G[54] = in1[65] & in2[65];
    assign P[54] = in1[65] ^ in2[65];
    assign G[55] = in1[64] & in2[64];
    assign P[55] = in1[64] ^ in2[64];
    assign G[56] = in1[63] & in2[63];
    assign P[56] = in1[63] ^ in2[63];
    assign G[57] = in1[62] & in2[62];
    assign P[57] = in1[62] ^ in2[62];
    assign G[58] = in1[61] & in2[61];
    assign P[58] = in1[61] ^ in2[61];
    assign G[59] = in1[60] & in2[60];
    assign P[59] = in1[60] ^ in2[60];
    assign G[60] = in1[59] & in2[59];
    assign P[60] = in1[59] ^ in2[59];
    assign G[61] = in1[58] & in2[58];
    assign P[61] = in1[58] ^ in2[58];
    assign G[62] = in1[57] & in2[57];
    assign P[62] = in1[57] ^ in2[57];
    assign G[63] = in1[56] & in2[56];
    assign P[63] = in1[56] ^ in2[56];
    assign G[64] = in1[55] & in2[55];
    assign P[64] = in1[55] ^ in2[55];
    assign G[65] = in1[54] & in2[54];
    assign P[65] = in1[54] ^ in2[54];
    assign G[66] = in1[53] & in2[53];
    assign P[66] = in1[53] ^ in2[53];
    assign G[67] = in1[52] & in2[52];
    assign P[67] = in1[52] ^ in2[52];
    assign G[68] = in1[51] & in2[51];
    assign P[68] = in1[51] ^ in2[51];
    assign G[69] = in1[50] & in2[50];
    assign P[69] = in1[50] ^ in2[50];
    assign G[70] = in1[49] & in2[49];
    assign P[70] = in1[49] ^ in2[49];
    assign G[71] = in1[48] & in2[48];
    assign P[71] = in1[48] ^ in2[48];
    assign G[72] = in1[47] & in2[47];
    assign P[72] = in1[47] ^ in2[47];
    assign G[73] = in1[46] & in2[46];
    assign P[73] = in1[46] ^ in2[46];
    assign G[74] = in1[45] & in2[45];
    assign P[74] = in1[45] ^ in2[45];
    assign G[75] = in1[44] & in2[44];
    assign P[75] = in1[44] ^ in2[44];
    assign G[76] = in1[43] & in2[43];
    assign P[76] = in1[43] ^ in2[43];
    assign G[77] = in1[42] & in2[42];
    assign P[77] = in1[42] ^ in2[42];
    assign G[78] = in1[41] & in2[41];
    assign P[78] = in1[41] ^ in2[41];
    assign G[79] = in1[40] & in2[40];
    assign P[79] = in1[40] ^ in2[40];
    assign G[80] = in1[39] & in2[39];
    assign P[80] = in1[39] ^ in2[39];
    assign G[81] = in1[38] & in2[38];
    assign P[81] = in1[38] ^ in2[38];
    assign G[82] = in1[37] & in2[37];
    assign P[82] = in1[37] ^ in2[37];
    assign G[83] = in1[36] & in2[36];
    assign P[83] = in1[36] ^ in2[36];
    assign G[84] = in1[35] & in2[35];
    assign P[84] = in1[35] ^ in2[35];
    assign G[85] = in1[34] & in2[34];
    assign P[85] = in1[34] ^ in2[34];
    assign G[86] = in1[33] & in2[33];
    assign P[86] = in1[33] ^ in2[33];
    assign G[87] = in1[32] & in2[32];
    assign P[87] = in1[32] ^ in2[32];
    assign G[88] = in1[31] & in2[31];
    assign P[88] = in1[31] ^ in2[31];
    assign G[89] = in1[30] & in2[30];
    assign P[89] = in1[30] ^ in2[30];
    assign G[90] = in1[29] & in2[29];
    assign P[90] = in1[29] ^ in2[29];
    assign G[91] = in1[28] & in2[28];
    assign P[91] = in1[28] ^ in2[28];
    assign G[92] = in1[27] & in2[27];
    assign P[92] = in1[27] ^ in2[27];
    assign G[93] = in1[26] & in2[26];
    assign P[93] = in1[26] ^ in2[26];
    assign G[94] = in1[25] & in2[25];
    assign P[94] = in1[25] ^ in2[25];
    assign G[95] = in1[24] & in2[24];
    assign P[95] = in1[24] ^ in2[24];
    assign G[96] = in1[23] & in2[23];
    assign P[96] = in1[23] ^ in2[23];
    assign G[97] = in1[22] & in2[22];
    assign P[97] = in1[22] ^ in2[22];
    assign G[98] = in1[21] & in2[21];
    assign P[98] = in1[21] ^ in2[21];
    assign G[99] = in1[20] & in2[20];
    assign P[99] = in1[20] ^ in2[20];
    assign G[100] = in1[19] & in2[19];
    assign P[100] = in1[19] ^ in2[19];
    assign G[101] = in1[18] & in2[18];
    assign P[101] = in1[18] ^ in2[18];
    assign G[102] = in1[17] & in2[17];
    assign P[102] = in1[17] ^ in2[17];
    assign G[103] = in1[16] & in2[16];
    assign P[103] = in1[16] ^ in2[16];
    assign G[104] = in1[15] & in2[15];
    assign P[104] = in1[15] ^ in2[15];
    assign G[105] = in1[14] & in2[14];
    assign P[105] = in1[14] ^ in2[14];
    assign G[106] = in1[13] & in2[13];
    assign P[106] = in1[13] ^ in2[13];
    assign G[107] = in1[12] & in2[12];
    assign P[107] = in1[12] ^ in2[12];
    assign G[108] = in1[11] & in2[11];
    assign P[108] = in1[11] ^ in2[11];
    assign G[109] = in1[10] & in2[10];
    assign P[109] = in1[10] ^ in2[10];
    assign G[110] = in1[9] & in2[9];
    assign P[110] = in1[9] ^ in2[9];
    assign G[111] = in1[8] & in2[8];
    assign P[111] = in1[8] ^ in2[8];
    assign G[112] = in1[7] & in2[7];
    assign P[112] = in1[7] ^ in2[7];
    assign G[113] = in1[6] & in2[6];
    assign P[113] = in1[6] ^ in2[6];
    assign G[114] = in1[5] & in2[5];
    assign P[114] = in1[5] ^ in2[5];
    assign G[115] = in1[4] & in2[4];
    assign P[115] = in1[4] ^ in2[4];
    assign G[116] = in1[3] & in2[3];
    assign P[116] = in1[3] ^ in2[3];
    assign G[117] = in1[2] & in2[2];
    assign P[117] = in1[2] ^ in2[2];
    assign G[118] = in1[1] & in2[1];
    assign P[118] = in1[1] ^ in2[1];
    assign G[119] = in1[0] & in2[0];
    assign P[119] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign cout = G[119] | (P[119] & C[119]);
    assign sum = P ^ C;
endmodule

module CLA_119(output [118:0] sum, output cout, input [118:0] in1, input [118:0] in2);

    wire[118:0] G;
    wire[118:0] C;
    wire[118:0] P;

    assign G[0] = in1[118] & in2[118];
    assign P[0] = in1[118] ^ in2[118];
    assign G[1] = in1[117] & in2[117];
    assign P[1] = in1[117] ^ in2[117];
    assign G[2] = in1[116] & in2[116];
    assign P[2] = in1[116] ^ in2[116];
    assign G[3] = in1[115] & in2[115];
    assign P[3] = in1[115] ^ in2[115];
    assign G[4] = in1[114] & in2[114];
    assign P[4] = in1[114] ^ in2[114];
    assign G[5] = in1[113] & in2[113];
    assign P[5] = in1[113] ^ in2[113];
    assign G[6] = in1[112] & in2[112];
    assign P[6] = in1[112] ^ in2[112];
    assign G[7] = in1[111] & in2[111];
    assign P[7] = in1[111] ^ in2[111];
    assign G[8] = in1[110] & in2[110];
    assign P[8] = in1[110] ^ in2[110];
    assign G[9] = in1[109] & in2[109];
    assign P[9] = in1[109] ^ in2[109];
    assign G[10] = in1[108] & in2[108];
    assign P[10] = in1[108] ^ in2[108];
    assign G[11] = in1[107] & in2[107];
    assign P[11] = in1[107] ^ in2[107];
    assign G[12] = in1[106] & in2[106];
    assign P[12] = in1[106] ^ in2[106];
    assign G[13] = in1[105] & in2[105];
    assign P[13] = in1[105] ^ in2[105];
    assign G[14] = in1[104] & in2[104];
    assign P[14] = in1[104] ^ in2[104];
    assign G[15] = in1[103] & in2[103];
    assign P[15] = in1[103] ^ in2[103];
    assign G[16] = in1[102] & in2[102];
    assign P[16] = in1[102] ^ in2[102];
    assign G[17] = in1[101] & in2[101];
    assign P[17] = in1[101] ^ in2[101];
    assign G[18] = in1[100] & in2[100];
    assign P[18] = in1[100] ^ in2[100];
    assign G[19] = in1[99] & in2[99];
    assign P[19] = in1[99] ^ in2[99];
    assign G[20] = in1[98] & in2[98];
    assign P[20] = in1[98] ^ in2[98];
    assign G[21] = in1[97] & in2[97];
    assign P[21] = in1[97] ^ in2[97];
    assign G[22] = in1[96] & in2[96];
    assign P[22] = in1[96] ^ in2[96];
    assign G[23] = in1[95] & in2[95];
    assign P[23] = in1[95] ^ in2[95];
    assign G[24] = in1[94] & in2[94];
    assign P[24] = in1[94] ^ in2[94];
    assign G[25] = in1[93] & in2[93];
    assign P[25] = in1[93] ^ in2[93];
    assign G[26] = in1[92] & in2[92];
    assign P[26] = in1[92] ^ in2[92];
    assign G[27] = in1[91] & in2[91];
    assign P[27] = in1[91] ^ in2[91];
    assign G[28] = in1[90] & in2[90];
    assign P[28] = in1[90] ^ in2[90];
    assign G[29] = in1[89] & in2[89];
    assign P[29] = in1[89] ^ in2[89];
    assign G[30] = in1[88] & in2[88];
    assign P[30] = in1[88] ^ in2[88];
    assign G[31] = in1[87] & in2[87];
    assign P[31] = in1[87] ^ in2[87];
    assign G[32] = in1[86] & in2[86];
    assign P[32] = in1[86] ^ in2[86];
    assign G[33] = in1[85] & in2[85];
    assign P[33] = in1[85] ^ in2[85];
    assign G[34] = in1[84] & in2[84];
    assign P[34] = in1[84] ^ in2[84];
    assign G[35] = in1[83] & in2[83];
    assign P[35] = in1[83] ^ in2[83];
    assign G[36] = in1[82] & in2[82];
    assign P[36] = in1[82] ^ in2[82];
    assign G[37] = in1[81] & in2[81];
    assign P[37] = in1[81] ^ in2[81];
    assign G[38] = in1[80] & in2[80];
    assign P[38] = in1[80] ^ in2[80];
    assign G[39] = in1[79] & in2[79];
    assign P[39] = in1[79] ^ in2[79];
    assign G[40] = in1[78] & in2[78];
    assign P[40] = in1[78] ^ in2[78];
    assign G[41] = in1[77] & in2[77];
    assign P[41] = in1[77] ^ in2[77];
    assign G[42] = in1[76] & in2[76];
    assign P[42] = in1[76] ^ in2[76];
    assign G[43] = in1[75] & in2[75];
    assign P[43] = in1[75] ^ in2[75];
    assign G[44] = in1[74] & in2[74];
    assign P[44] = in1[74] ^ in2[74];
    assign G[45] = in1[73] & in2[73];
    assign P[45] = in1[73] ^ in2[73];
    assign G[46] = in1[72] & in2[72];
    assign P[46] = in1[72] ^ in2[72];
    assign G[47] = in1[71] & in2[71];
    assign P[47] = in1[71] ^ in2[71];
    assign G[48] = in1[70] & in2[70];
    assign P[48] = in1[70] ^ in2[70];
    assign G[49] = in1[69] & in2[69];
    assign P[49] = in1[69] ^ in2[69];
    assign G[50] = in1[68] & in2[68];
    assign P[50] = in1[68] ^ in2[68];
    assign G[51] = in1[67] & in2[67];
    assign P[51] = in1[67] ^ in2[67];
    assign G[52] = in1[66] & in2[66];
    assign P[52] = in1[66] ^ in2[66];
    assign G[53] = in1[65] & in2[65];
    assign P[53] = in1[65] ^ in2[65];
    assign G[54] = in1[64] & in2[64];
    assign P[54] = in1[64] ^ in2[64];
    assign G[55] = in1[63] & in2[63];
    assign P[55] = in1[63] ^ in2[63];
    assign G[56] = in1[62] & in2[62];
    assign P[56] = in1[62] ^ in2[62];
    assign G[57] = in1[61] & in2[61];
    assign P[57] = in1[61] ^ in2[61];
    assign G[58] = in1[60] & in2[60];
    assign P[58] = in1[60] ^ in2[60];
    assign G[59] = in1[59] & in2[59];
    assign P[59] = in1[59] ^ in2[59];
    assign G[60] = in1[58] & in2[58];
    assign P[60] = in1[58] ^ in2[58];
    assign G[61] = in1[57] & in2[57];
    assign P[61] = in1[57] ^ in2[57];
    assign G[62] = in1[56] & in2[56];
    assign P[62] = in1[56] ^ in2[56];
    assign G[63] = in1[55] & in2[55];
    assign P[63] = in1[55] ^ in2[55];
    assign G[64] = in1[54] & in2[54];
    assign P[64] = in1[54] ^ in2[54];
    assign G[65] = in1[53] & in2[53];
    assign P[65] = in1[53] ^ in2[53];
    assign G[66] = in1[52] & in2[52];
    assign P[66] = in1[52] ^ in2[52];
    assign G[67] = in1[51] & in2[51];
    assign P[67] = in1[51] ^ in2[51];
    assign G[68] = in1[50] & in2[50];
    assign P[68] = in1[50] ^ in2[50];
    assign G[69] = in1[49] & in2[49];
    assign P[69] = in1[49] ^ in2[49];
    assign G[70] = in1[48] & in2[48];
    assign P[70] = in1[48] ^ in2[48];
    assign G[71] = in1[47] & in2[47];
    assign P[71] = in1[47] ^ in2[47];
    assign G[72] = in1[46] & in2[46];
    assign P[72] = in1[46] ^ in2[46];
    assign G[73] = in1[45] & in2[45];
    assign P[73] = in1[45] ^ in2[45];
    assign G[74] = in1[44] & in2[44];
    assign P[74] = in1[44] ^ in2[44];
    assign G[75] = in1[43] & in2[43];
    assign P[75] = in1[43] ^ in2[43];
    assign G[76] = in1[42] & in2[42];
    assign P[76] = in1[42] ^ in2[42];
    assign G[77] = in1[41] & in2[41];
    assign P[77] = in1[41] ^ in2[41];
    assign G[78] = in1[40] & in2[40];
    assign P[78] = in1[40] ^ in2[40];
    assign G[79] = in1[39] & in2[39];
    assign P[79] = in1[39] ^ in2[39];
    assign G[80] = in1[38] & in2[38];
    assign P[80] = in1[38] ^ in2[38];
    assign G[81] = in1[37] & in2[37];
    assign P[81] = in1[37] ^ in2[37];
    assign G[82] = in1[36] & in2[36];
    assign P[82] = in1[36] ^ in2[36];
    assign G[83] = in1[35] & in2[35];
    assign P[83] = in1[35] ^ in2[35];
    assign G[84] = in1[34] & in2[34];
    assign P[84] = in1[34] ^ in2[34];
    assign G[85] = in1[33] & in2[33];
    assign P[85] = in1[33] ^ in2[33];
    assign G[86] = in1[32] & in2[32];
    assign P[86] = in1[32] ^ in2[32];
    assign G[87] = in1[31] & in2[31];
    assign P[87] = in1[31] ^ in2[31];
    assign G[88] = in1[30] & in2[30];
    assign P[88] = in1[30] ^ in2[30];
    assign G[89] = in1[29] & in2[29];
    assign P[89] = in1[29] ^ in2[29];
    assign G[90] = in1[28] & in2[28];
    assign P[90] = in1[28] ^ in2[28];
    assign G[91] = in1[27] & in2[27];
    assign P[91] = in1[27] ^ in2[27];
    assign G[92] = in1[26] & in2[26];
    assign P[92] = in1[26] ^ in2[26];
    assign G[93] = in1[25] & in2[25];
    assign P[93] = in1[25] ^ in2[25];
    assign G[94] = in1[24] & in2[24];
    assign P[94] = in1[24] ^ in2[24];
    assign G[95] = in1[23] & in2[23];
    assign P[95] = in1[23] ^ in2[23];
    assign G[96] = in1[22] & in2[22];
    assign P[96] = in1[22] ^ in2[22];
    assign G[97] = in1[21] & in2[21];
    assign P[97] = in1[21] ^ in2[21];
    assign G[98] = in1[20] & in2[20];
    assign P[98] = in1[20] ^ in2[20];
    assign G[99] = in1[19] & in2[19];
    assign P[99] = in1[19] ^ in2[19];
    assign G[100] = in1[18] & in2[18];
    assign P[100] = in1[18] ^ in2[18];
    assign G[101] = in1[17] & in2[17];
    assign P[101] = in1[17] ^ in2[17];
    assign G[102] = in1[16] & in2[16];
    assign P[102] = in1[16] ^ in2[16];
    assign G[103] = in1[15] & in2[15];
    assign P[103] = in1[15] ^ in2[15];
    assign G[104] = in1[14] & in2[14];
    assign P[104] = in1[14] ^ in2[14];
    assign G[105] = in1[13] & in2[13];
    assign P[105] = in1[13] ^ in2[13];
    assign G[106] = in1[12] & in2[12];
    assign P[106] = in1[12] ^ in2[12];
    assign G[107] = in1[11] & in2[11];
    assign P[107] = in1[11] ^ in2[11];
    assign G[108] = in1[10] & in2[10];
    assign P[108] = in1[10] ^ in2[10];
    assign G[109] = in1[9] & in2[9];
    assign P[109] = in1[9] ^ in2[9];
    assign G[110] = in1[8] & in2[8];
    assign P[110] = in1[8] ^ in2[8];
    assign G[111] = in1[7] & in2[7];
    assign P[111] = in1[7] ^ in2[7];
    assign G[112] = in1[6] & in2[6];
    assign P[112] = in1[6] ^ in2[6];
    assign G[113] = in1[5] & in2[5];
    assign P[113] = in1[5] ^ in2[5];
    assign G[114] = in1[4] & in2[4];
    assign P[114] = in1[4] ^ in2[4];
    assign G[115] = in1[3] & in2[3];
    assign P[115] = in1[3] ^ in2[3];
    assign G[116] = in1[2] & in2[2];
    assign P[116] = in1[2] ^ in2[2];
    assign G[117] = in1[1] & in2[1];
    assign P[117] = in1[1] ^ in2[1];
    assign G[118] = in1[0] & in2[0];
    assign P[118] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign cout = G[118] | (P[118] & C[118]);
    assign sum = P ^ C;
endmodule

module CLA_118(output [117:0] sum, output cout, input [117:0] in1, input [117:0] in2);

    wire[117:0] G;
    wire[117:0] C;
    wire[117:0] P;

    assign G[0] = in1[117] & in2[117];
    assign P[0] = in1[117] ^ in2[117];
    assign G[1] = in1[116] & in2[116];
    assign P[1] = in1[116] ^ in2[116];
    assign G[2] = in1[115] & in2[115];
    assign P[2] = in1[115] ^ in2[115];
    assign G[3] = in1[114] & in2[114];
    assign P[3] = in1[114] ^ in2[114];
    assign G[4] = in1[113] & in2[113];
    assign P[4] = in1[113] ^ in2[113];
    assign G[5] = in1[112] & in2[112];
    assign P[5] = in1[112] ^ in2[112];
    assign G[6] = in1[111] & in2[111];
    assign P[6] = in1[111] ^ in2[111];
    assign G[7] = in1[110] & in2[110];
    assign P[7] = in1[110] ^ in2[110];
    assign G[8] = in1[109] & in2[109];
    assign P[8] = in1[109] ^ in2[109];
    assign G[9] = in1[108] & in2[108];
    assign P[9] = in1[108] ^ in2[108];
    assign G[10] = in1[107] & in2[107];
    assign P[10] = in1[107] ^ in2[107];
    assign G[11] = in1[106] & in2[106];
    assign P[11] = in1[106] ^ in2[106];
    assign G[12] = in1[105] & in2[105];
    assign P[12] = in1[105] ^ in2[105];
    assign G[13] = in1[104] & in2[104];
    assign P[13] = in1[104] ^ in2[104];
    assign G[14] = in1[103] & in2[103];
    assign P[14] = in1[103] ^ in2[103];
    assign G[15] = in1[102] & in2[102];
    assign P[15] = in1[102] ^ in2[102];
    assign G[16] = in1[101] & in2[101];
    assign P[16] = in1[101] ^ in2[101];
    assign G[17] = in1[100] & in2[100];
    assign P[17] = in1[100] ^ in2[100];
    assign G[18] = in1[99] & in2[99];
    assign P[18] = in1[99] ^ in2[99];
    assign G[19] = in1[98] & in2[98];
    assign P[19] = in1[98] ^ in2[98];
    assign G[20] = in1[97] & in2[97];
    assign P[20] = in1[97] ^ in2[97];
    assign G[21] = in1[96] & in2[96];
    assign P[21] = in1[96] ^ in2[96];
    assign G[22] = in1[95] & in2[95];
    assign P[22] = in1[95] ^ in2[95];
    assign G[23] = in1[94] & in2[94];
    assign P[23] = in1[94] ^ in2[94];
    assign G[24] = in1[93] & in2[93];
    assign P[24] = in1[93] ^ in2[93];
    assign G[25] = in1[92] & in2[92];
    assign P[25] = in1[92] ^ in2[92];
    assign G[26] = in1[91] & in2[91];
    assign P[26] = in1[91] ^ in2[91];
    assign G[27] = in1[90] & in2[90];
    assign P[27] = in1[90] ^ in2[90];
    assign G[28] = in1[89] & in2[89];
    assign P[28] = in1[89] ^ in2[89];
    assign G[29] = in1[88] & in2[88];
    assign P[29] = in1[88] ^ in2[88];
    assign G[30] = in1[87] & in2[87];
    assign P[30] = in1[87] ^ in2[87];
    assign G[31] = in1[86] & in2[86];
    assign P[31] = in1[86] ^ in2[86];
    assign G[32] = in1[85] & in2[85];
    assign P[32] = in1[85] ^ in2[85];
    assign G[33] = in1[84] & in2[84];
    assign P[33] = in1[84] ^ in2[84];
    assign G[34] = in1[83] & in2[83];
    assign P[34] = in1[83] ^ in2[83];
    assign G[35] = in1[82] & in2[82];
    assign P[35] = in1[82] ^ in2[82];
    assign G[36] = in1[81] & in2[81];
    assign P[36] = in1[81] ^ in2[81];
    assign G[37] = in1[80] & in2[80];
    assign P[37] = in1[80] ^ in2[80];
    assign G[38] = in1[79] & in2[79];
    assign P[38] = in1[79] ^ in2[79];
    assign G[39] = in1[78] & in2[78];
    assign P[39] = in1[78] ^ in2[78];
    assign G[40] = in1[77] & in2[77];
    assign P[40] = in1[77] ^ in2[77];
    assign G[41] = in1[76] & in2[76];
    assign P[41] = in1[76] ^ in2[76];
    assign G[42] = in1[75] & in2[75];
    assign P[42] = in1[75] ^ in2[75];
    assign G[43] = in1[74] & in2[74];
    assign P[43] = in1[74] ^ in2[74];
    assign G[44] = in1[73] & in2[73];
    assign P[44] = in1[73] ^ in2[73];
    assign G[45] = in1[72] & in2[72];
    assign P[45] = in1[72] ^ in2[72];
    assign G[46] = in1[71] & in2[71];
    assign P[46] = in1[71] ^ in2[71];
    assign G[47] = in1[70] & in2[70];
    assign P[47] = in1[70] ^ in2[70];
    assign G[48] = in1[69] & in2[69];
    assign P[48] = in1[69] ^ in2[69];
    assign G[49] = in1[68] & in2[68];
    assign P[49] = in1[68] ^ in2[68];
    assign G[50] = in1[67] & in2[67];
    assign P[50] = in1[67] ^ in2[67];
    assign G[51] = in1[66] & in2[66];
    assign P[51] = in1[66] ^ in2[66];
    assign G[52] = in1[65] & in2[65];
    assign P[52] = in1[65] ^ in2[65];
    assign G[53] = in1[64] & in2[64];
    assign P[53] = in1[64] ^ in2[64];
    assign G[54] = in1[63] & in2[63];
    assign P[54] = in1[63] ^ in2[63];
    assign G[55] = in1[62] & in2[62];
    assign P[55] = in1[62] ^ in2[62];
    assign G[56] = in1[61] & in2[61];
    assign P[56] = in1[61] ^ in2[61];
    assign G[57] = in1[60] & in2[60];
    assign P[57] = in1[60] ^ in2[60];
    assign G[58] = in1[59] & in2[59];
    assign P[58] = in1[59] ^ in2[59];
    assign G[59] = in1[58] & in2[58];
    assign P[59] = in1[58] ^ in2[58];
    assign G[60] = in1[57] & in2[57];
    assign P[60] = in1[57] ^ in2[57];
    assign G[61] = in1[56] & in2[56];
    assign P[61] = in1[56] ^ in2[56];
    assign G[62] = in1[55] & in2[55];
    assign P[62] = in1[55] ^ in2[55];
    assign G[63] = in1[54] & in2[54];
    assign P[63] = in1[54] ^ in2[54];
    assign G[64] = in1[53] & in2[53];
    assign P[64] = in1[53] ^ in2[53];
    assign G[65] = in1[52] & in2[52];
    assign P[65] = in1[52] ^ in2[52];
    assign G[66] = in1[51] & in2[51];
    assign P[66] = in1[51] ^ in2[51];
    assign G[67] = in1[50] & in2[50];
    assign P[67] = in1[50] ^ in2[50];
    assign G[68] = in1[49] & in2[49];
    assign P[68] = in1[49] ^ in2[49];
    assign G[69] = in1[48] & in2[48];
    assign P[69] = in1[48] ^ in2[48];
    assign G[70] = in1[47] & in2[47];
    assign P[70] = in1[47] ^ in2[47];
    assign G[71] = in1[46] & in2[46];
    assign P[71] = in1[46] ^ in2[46];
    assign G[72] = in1[45] & in2[45];
    assign P[72] = in1[45] ^ in2[45];
    assign G[73] = in1[44] & in2[44];
    assign P[73] = in1[44] ^ in2[44];
    assign G[74] = in1[43] & in2[43];
    assign P[74] = in1[43] ^ in2[43];
    assign G[75] = in1[42] & in2[42];
    assign P[75] = in1[42] ^ in2[42];
    assign G[76] = in1[41] & in2[41];
    assign P[76] = in1[41] ^ in2[41];
    assign G[77] = in1[40] & in2[40];
    assign P[77] = in1[40] ^ in2[40];
    assign G[78] = in1[39] & in2[39];
    assign P[78] = in1[39] ^ in2[39];
    assign G[79] = in1[38] & in2[38];
    assign P[79] = in1[38] ^ in2[38];
    assign G[80] = in1[37] & in2[37];
    assign P[80] = in1[37] ^ in2[37];
    assign G[81] = in1[36] & in2[36];
    assign P[81] = in1[36] ^ in2[36];
    assign G[82] = in1[35] & in2[35];
    assign P[82] = in1[35] ^ in2[35];
    assign G[83] = in1[34] & in2[34];
    assign P[83] = in1[34] ^ in2[34];
    assign G[84] = in1[33] & in2[33];
    assign P[84] = in1[33] ^ in2[33];
    assign G[85] = in1[32] & in2[32];
    assign P[85] = in1[32] ^ in2[32];
    assign G[86] = in1[31] & in2[31];
    assign P[86] = in1[31] ^ in2[31];
    assign G[87] = in1[30] & in2[30];
    assign P[87] = in1[30] ^ in2[30];
    assign G[88] = in1[29] & in2[29];
    assign P[88] = in1[29] ^ in2[29];
    assign G[89] = in1[28] & in2[28];
    assign P[89] = in1[28] ^ in2[28];
    assign G[90] = in1[27] & in2[27];
    assign P[90] = in1[27] ^ in2[27];
    assign G[91] = in1[26] & in2[26];
    assign P[91] = in1[26] ^ in2[26];
    assign G[92] = in1[25] & in2[25];
    assign P[92] = in1[25] ^ in2[25];
    assign G[93] = in1[24] & in2[24];
    assign P[93] = in1[24] ^ in2[24];
    assign G[94] = in1[23] & in2[23];
    assign P[94] = in1[23] ^ in2[23];
    assign G[95] = in1[22] & in2[22];
    assign P[95] = in1[22] ^ in2[22];
    assign G[96] = in1[21] & in2[21];
    assign P[96] = in1[21] ^ in2[21];
    assign G[97] = in1[20] & in2[20];
    assign P[97] = in1[20] ^ in2[20];
    assign G[98] = in1[19] & in2[19];
    assign P[98] = in1[19] ^ in2[19];
    assign G[99] = in1[18] & in2[18];
    assign P[99] = in1[18] ^ in2[18];
    assign G[100] = in1[17] & in2[17];
    assign P[100] = in1[17] ^ in2[17];
    assign G[101] = in1[16] & in2[16];
    assign P[101] = in1[16] ^ in2[16];
    assign G[102] = in1[15] & in2[15];
    assign P[102] = in1[15] ^ in2[15];
    assign G[103] = in1[14] & in2[14];
    assign P[103] = in1[14] ^ in2[14];
    assign G[104] = in1[13] & in2[13];
    assign P[104] = in1[13] ^ in2[13];
    assign G[105] = in1[12] & in2[12];
    assign P[105] = in1[12] ^ in2[12];
    assign G[106] = in1[11] & in2[11];
    assign P[106] = in1[11] ^ in2[11];
    assign G[107] = in1[10] & in2[10];
    assign P[107] = in1[10] ^ in2[10];
    assign G[108] = in1[9] & in2[9];
    assign P[108] = in1[9] ^ in2[9];
    assign G[109] = in1[8] & in2[8];
    assign P[109] = in1[8] ^ in2[8];
    assign G[110] = in1[7] & in2[7];
    assign P[110] = in1[7] ^ in2[7];
    assign G[111] = in1[6] & in2[6];
    assign P[111] = in1[6] ^ in2[6];
    assign G[112] = in1[5] & in2[5];
    assign P[112] = in1[5] ^ in2[5];
    assign G[113] = in1[4] & in2[4];
    assign P[113] = in1[4] ^ in2[4];
    assign G[114] = in1[3] & in2[3];
    assign P[114] = in1[3] ^ in2[3];
    assign G[115] = in1[2] & in2[2];
    assign P[115] = in1[2] ^ in2[2];
    assign G[116] = in1[1] & in2[1];
    assign P[116] = in1[1] ^ in2[1];
    assign G[117] = in1[0] & in2[0];
    assign P[117] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign cout = G[117] | (P[117] & C[117]);
    assign sum = P ^ C;
endmodule

module CLA_117(output [116:0] sum, output cout, input [116:0] in1, input [116:0] in2);

    wire[116:0] G;
    wire[116:0] C;
    wire[116:0] P;

    assign G[0] = in1[116] & in2[116];
    assign P[0] = in1[116] ^ in2[116];
    assign G[1] = in1[115] & in2[115];
    assign P[1] = in1[115] ^ in2[115];
    assign G[2] = in1[114] & in2[114];
    assign P[2] = in1[114] ^ in2[114];
    assign G[3] = in1[113] & in2[113];
    assign P[3] = in1[113] ^ in2[113];
    assign G[4] = in1[112] & in2[112];
    assign P[4] = in1[112] ^ in2[112];
    assign G[5] = in1[111] & in2[111];
    assign P[5] = in1[111] ^ in2[111];
    assign G[6] = in1[110] & in2[110];
    assign P[6] = in1[110] ^ in2[110];
    assign G[7] = in1[109] & in2[109];
    assign P[7] = in1[109] ^ in2[109];
    assign G[8] = in1[108] & in2[108];
    assign P[8] = in1[108] ^ in2[108];
    assign G[9] = in1[107] & in2[107];
    assign P[9] = in1[107] ^ in2[107];
    assign G[10] = in1[106] & in2[106];
    assign P[10] = in1[106] ^ in2[106];
    assign G[11] = in1[105] & in2[105];
    assign P[11] = in1[105] ^ in2[105];
    assign G[12] = in1[104] & in2[104];
    assign P[12] = in1[104] ^ in2[104];
    assign G[13] = in1[103] & in2[103];
    assign P[13] = in1[103] ^ in2[103];
    assign G[14] = in1[102] & in2[102];
    assign P[14] = in1[102] ^ in2[102];
    assign G[15] = in1[101] & in2[101];
    assign P[15] = in1[101] ^ in2[101];
    assign G[16] = in1[100] & in2[100];
    assign P[16] = in1[100] ^ in2[100];
    assign G[17] = in1[99] & in2[99];
    assign P[17] = in1[99] ^ in2[99];
    assign G[18] = in1[98] & in2[98];
    assign P[18] = in1[98] ^ in2[98];
    assign G[19] = in1[97] & in2[97];
    assign P[19] = in1[97] ^ in2[97];
    assign G[20] = in1[96] & in2[96];
    assign P[20] = in1[96] ^ in2[96];
    assign G[21] = in1[95] & in2[95];
    assign P[21] = in1[95] ^ in2[95];
    assign G[22] = in1[94] & in2[94];
    assign P[22] = in1[94] ^ in2[94];
    assign G[23] = in1[93] & in2[93];
    assign P[23] = in1[93] ^ in2[93];
    assign G[24] = in1[92] & in2[92];
    assign P[24] = in1[92] ^ in2[92];
    assign G[25] = in1[91] & in2[91];
    assign P[25] = in1[91] ^ in2[91];
    assign G[26] = in1[90] & in2[90];
    assign P[26] = in1[90] ^ in2[90];
    assign G[27] = in1[89] & in2[89];
    assign P[27] = in1[89] ^ in2[89];
    assign G[28] = in1[88] & in2[88];
    assign P[28] = in1[88] ^ in2[88];
    assign G[29] = in1[87] & in2[87];
    assign P[29] = in1[87] ^ in2[87];
    assign G[30] = in1[86] & in2[86];
    assign P[30] = in1[86] ^ in2[86];
    assign G[31] = in1[85] & in2[85];
    assign P[31] = in1[85] ^ in2[85];
    assign G[32] = in1[84] & in2[84];
    assign P[32] = in1[84] ^ in2[84];
    assign G[33] = in1[83] & in2[83];
    assign P[33] = in1[83] ^ in2[83];
    assign G[34] = in1[82] & in2[82];
    assign P[34] = in1[82] ^ in2[82];
    assign G[35] = in1[81] & in2[81];
    assign P[35] = in1[81] ^ in2[81];
    assign G[36] = in1[80] & in2[80];
    assign P[36] = in1[80] ^ in2[80];
    assign G[37] = in1[79] & in2[79];
    assign P[37] = in1[79] ^ in2[79];
    assign G[38] = in1[78] & in2[78];
    assign P[38] = in1[78] ^ in2[78];
    assign G[39] = in1[77] & in2[77];
    assign P[39] = in1[77] ^ in2[77];
    assign G[40] = in1[76] & in2[76];
    assign P[40] = in1[76] ^ in2[76];
    assign G[41] = in1[75] & in2[75];
    assign P[41] = in1[75] ^ in2[75];
    assign G[42] = in1[74] & in2[74];
    assign P[42] = in1[74] ^ in2[74];
    assign G[43] = in1[73] & in2[73];
    assign P[43] = in1[73] ^ in2[73];
    assign G[44] = in1[72] & in2[72];
    assign P[44] = in1[72] ^ in2[72];
    assign G[45] = in1[71] & in2[71];
    assign P[45] = in1[71] ^ in2[71];
    assign G[46] = in1[70] & in2[70];
    assign P[46] = in1[70] ^ in2[70];
    assign G[47] = in1[69] & in2[69];
    assign P[47] = in1[69] ^ in2[69];
    assign G[48] = in1[68] & in2[68];
    assign P[48] = in1[68] ^ in2[68];
    assign G[49] = in1[67] & in2[67];
    assign P[49] = in1[67] ^ in2[67];
    assign G[50] = in1[66] & in2[66];
    assign P[50] = in1[66] ^ in2[66];
    assign G[51] = in1[65] & in2[65];
    assign P[51] = in1[65] ^ in2[65];
    assign G[52] = in1[64] & in2[64];
    assign P[52] = in1[64] ^ in2[64];
    assign G[53] = in1[63] & in2[63];
    assign P[53] = in1[63] ^ in2[63];
    assign G[54] = in1[62] & in2[62];
    assign P[54] = in1[62] ^ in2[62];
    assign G[55] = in1[61] & in2[61];
    assign P[55] = in1[61] ^ in2[61];
    assign G[56] = in1[60] & in2[60];
    assign P[56] = in1[60] ^ in2[60];
    assign G[57] = in1[59] & in2[59];
    assign P[57] = in1[59] ^ in2[59];
    assign G[58] = in1[58] & in2[58];
    assign P[58] = in1[58] ^ in2[58];
    assign G[59] = in1[57] & in2[57];
    assign P[59] = in1[57] ^ in2[57];
    assign G[60] = in1[56] & in2[56];
    assign P[60] = in1[56] ^ in2[56];
    assign G[61] = in1[55] & in2[55];
    assign P[61] = in1[55] ^ in2[55];
    assign G[62] = in1[54] & in2[54];
    assign P[62] = in1[54] ^ in2[54];
    assign G[63] = in1[53] & in2[53];
    assign P[63] = in1[53] ^ in2[53];
    assign G[64] = in1[52] & in2[52];
    assign P[64] = in1[52] ^ in2[52];
    assign G[65] = in1[51] & in2[51];
    assign P[65] = in1[51] ^ in2[51];
    assign G[66] = in1[50] & in2[50];
    assign P[66] = in1[50] ^ in2[50];
    assign G[67] = in1[49] & in2[49];
    assign P[67] = in1[49] ^ in2[49];
    assign G[68] = in1[48] & in2[48];
    assign P[68] = in1[48] ^ in2[48];
    assign G[69] = in1[47] & in2[47];
    assign P[69] = in1[47] ^ in2[47];
    assign G[70] = in1[46] & in2[46];
    assign P[70] = in1[46] ^ in2[46];
    assign G[71] = in1[45] & in2[45];
    assign P[71] = in1[45] ^ in2[45];
    assign G[72] = in1[44] & in2[44];
    assign P[72] = in1[44] ^ in2[44];
    assign G[73] = in1[43] & in2[43];
    assign P[73] = in1[43] ^ in2[43];
    assign G[74] = in1[42] & in2[42];
    assign P[74] = in1[42] ^ in2[42];
    assign G[75] = in1[41] & in2[41];
    assign P[75] = in1[41] ^ in2[41];
    assign G[76] = in1[40] & in2[40];
    assign P[76] = in1[40] ^ in2[40];
    assign G[77] = in1[39] & in2[39];
    assign P[77] = in1[39] ^ in2[39];
    assign G[78] = in1[38] & in2[38];
    assign P[78] = in1[38] ^ in2[38];
    assign G[79] = in1[37] & in2[37];
    assign P[79] = in1[37] ^ in2[37];
    assign G[80] = in1[36] & in2[36];
    assign P[80] = in1[36] ^ in2[36];
    assign G[81] = in1[35] & in2[35];
    assign P[81] = in1[35] ^ in2[35];
    assign G[82] = in1[34] & in2[34];
    assign P[82] = in1[34] ^ in2[34];
    assign G[83] = in1[33] & in2[33];
    assign P[83] = in1[33] ^ in2[33];
    assign G[84] = in1[32] & in2[32];
    assign P[84] = in1[32] ^ in2[32];
    assign G[85] = in1[31] & in2[31];
    assign P[85] = in1[31] ^ in2[31];
    assign G[86] = in1[30] & in2[30];
    assign P[86] = in1[30] ^ in2[30];
    assign G[87] = in1[29] & in2[29];
    assign P[87] = in1[29] ^ in2[29];
    assign G[88] = in1[28] & in2[28];
    assign P[88] = in1[28] ^ in2[28];
    assign G[89] = in1[27] & in2[27];
    assign P[89] = in1[27] ^ in2[27];
    assign G[90] = in1[26] & in2[26];
    assign P[90] = in1[26] ^ in2[26];
    assign G[91] = in1[25] & in2[25];
    assign P[91] = in1[25] ^ in2[25];
    assign G[92] = in1[24] & in2[24];
    assign P[92] = in1[24] ^ in2[24];
    assign G[93] = in1[23] & in2[23];
    assign P[93] = in1[23] ^ in2[23];
    assign G[94] = in1[22] & in2[22];
    assign P[94] = in1[22] ^ in2[22];
    assign G[95] = in1[21] & in2[21];
    assign P[95] = in1[21] ^ in2[21];
    assign G[96] = in1[20] & in2[20];
    assign P[96] = in1[20] ^ in2[20];
    assign G[97] = in1[19] & in2[19];
    assign P[97] = in1[19] ^ in2[19];
    assign G[98] = in1[18] & in2[18];
    assign P[98] = in1[18] ^ in2[18];
    assign G[99] = in1[17] & in2[17];
    assign P[99] = in1[17] ^ in2[17];
    assign G[100] = in1[16] & in2[16];
    assign P[100] = in1[16] ^ in2[16];
    assign G[101] = in1[15] & in2[15];
    assign P[101] = in1[15] ^ in2[15];
    assign G[102] = in1[14] & in2[14];
    assign P[102] = in1[14] ^ in2[14];
    assign G[103] = in1[13] & in2[13];
    assign P[103] = in1[13] ^ in2[13];
    assign G[104] = in1[12] & in2[12];
    assign P[104] = in1[12] ^ in2[12];
    assign G[105] = in1[11] & in2[11];
    assign P[105] = in1[11] ^ in2[11];
    assign G[106] = in1[10] & in2[10];
    assign P[106] = in1[10] ^ in2[10];
    assign G[107] = in1[9] & in2[9];
    assign P[107] = in1[9] ^ in2[9];
    assign G[108] = in1[8] & in2[8];
    assign P[108] = in1[8] ^ in2[8];
    assign G[109] = in1[7] & in2[7];
    assign P[109] = in1[7] ^ in2[7];
    assign G[110] = in1[6] & in2[6];
    assign P[110] = in1[6] ^ in2[6];
    assign G[111] = in1[5] & in2[5];
    assign P[111] = in1[5] ^ in2[5];
    assign G[112] = in1[4] & in2[4];
    assign P[112] = in1[4] ^ in2[4];
    assign G[113] = in1[3] & in2[3];
    assign P[113] = in1[3] ^ in2[3];
    assign G[114] = in1[2] & in2[2];
    assign P[114] = in1[2] ^ in2[2];
    assign G[115] = in1[1] & in2[1];
    assign P[115] = in1[1] ^ in2[1];
    assign G[116] = in1[0] & in2[0];
    assign P[116] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign cout = G[116] | (P[116] & C[116]);
    assign sum = P ^ C;
endmodule

module CLA_116(output [115:0] sum, output cout, input [115:0] in1, input [115:0] in2);

    wire[115:0] G;
    wire[115:0] C;
    wire[115:0] P;

    assign G[0] = in1[115] & in2[115];
    assign P[0] = in1[115] ^ in2[115];
    assign G[1] = in1[114] & in2[114];
    assign P[1] = in1[114] ^ in2[114];
    assign G[2] = in1[113] & in2[113];
    assign P[2] = in1[113] ^ in2[113];
    assign G[3] = in1[112] & in2[112];
    assign P[3] = in1[112] ^ in2[112];
    assign G[4] = in1[111] & in2[111];
    assign P[4] = in1[111] ^ in2[111];
    assign G[5] = in1[110] & in2[110];
    assign P[5] = in1[110] ^ in2[110];
    assign G[6] = in1[109] & in2[109];
    assign P[6] = in1[109] ^ in2[109];
    assign G[7] = in1[108] & in2[108];
    assign P[7] = in1[108] ^ in2[108];
    assign G[8] = in1[107] & in2[107];
    assign P[8] = in1[107] ^ in2[107];
    assign G[9] = in1[106] & in2[106];
    assign P[9] = in1[106] ^ in2[106];
    assign G[10] = in1[105] & in2[105];
    assign P[10] = in1[105] ^ in2[105];
    assign G[11] = in1[104] & in2[104];
    assign P[11] = in1[104] ^ in2[104];
    assign G[12] = in1[103] & in2[103];
    assign P[12] = in1[103] ^ in2[103];
    assign G[13] = in1[102] & in2[102];
    assign P[13] = in1[102] ^ in2[102];
    assign G[14] = in1[101] & in2[101];
    assign P[14] = in1[101] ^ in2[101];
    assign G[15] = in1[100] & in2[100];
    assign P[15] = in1[100] ^ in2[100];
    assign G[16] = in1[99] & in2[99];
    assign P[16] = in1[99] ^ in2[99];
    assign G[17] = in1[98] & in2[98];
    assign P[17] = in1[98] ^ in2[98];
    assign G[18] = in1[97] & in2[97];
    assign P[18] = in1[97] ^ in2[97];
    assign G[19] = in1[96] & in2[96];
    assign P[19] = in1[96] ^ in2[96];
    assign G[20] = in1[95] & in2[95];
    assign P[20] = in1[95] ^ in2[95];
    assign G[21] = in1[94] & in2[94];
    assign P[21] = in1[94] ^ in2[94];
    assign G[22] = in1[93] & in2[93];
    assign P[22] = in1[93] ^ in2[93];
    assign G[23] = in1[92] & in2[92];
    assign P[23] = in1[92] ^ in2[92];
    assign G[24] = in1[91] & in2[91];
    assign P[24] = in1[91] ^ in2[91];
    assign G[25] = in1[90] & in2[90];
    assign P[25] = in1[90] ^ in2[90];
    assign G[26] = in1[89] & in2[89];
    assign P[26] = in1[89] ^ in2[89];
    assign G[27] = in1[88] & in2[88];
    assign P[27] = in1[88] ^ in2[88];
    assign G[28] = in1[87] & in2[87];
    assign P[28] = in1[87] ^ in2[87];
    assign G[29] = in1[86] & in2[86];
    assign P[29] = in1[86] ^ in2[86];
    assign G[30] = in1[85] & in2[85];
    assign P[30] = in1[85] ^ in2[85];
    assign G[31] = in1[84] & in2[84];
    assign P[31] = in1[84] ^ in2[84];
    assign G[32] = in1[83] & in2[83];
    assign P[32] = in1[83] ^ in2[83];
    assign G[33] = in1[82] & in2[82];
    assign P[33] = in1[82] ^ in2[82];
    assign G[34] = in1[81] & in2[81];
    assign P[34] = in1[81] ^ in2[81];
    assign G[35] = in1[80] & in2[80];
    assign P[35] = in1[80] ^ in2[80];
    assign G[36] = in1[79] & in2[79];
    assign P[36] = in1[79] ^ in2[79];
    assign G[37] = in1[78] & in2[78];
    assign P[37] = in1[78] ^ in2[78];
    assign G[38] = in1[77] & in2[77];
    assign P[38] = in1[77] ^ in2[77];
    assign G[39] = in1[76] & in2[76];
    assign P[39] = in1[76] ^ in2[76];
    assign G[40] = in1[75] & in2[75];
    assign P[40] = in1[75] ^ in2[75];
    assign G[41] = in1[74] & in2[74];
    assign P[41] = in1[74] ^ in2[74];
    assign G[42] = in1[73] & in2[73];
    assign P[42] = in1[73] ^ in2[73];
    assign G[43] = in1[72] & in2[72];
    assign P[43] = in1[72] ^ in2[72];
    assign G[44] = in1[71] & in2[71];
    assign P[44] = in1[71] ^ in2[71];
    assign G[45] = in1[70] & in2[70];
    assign P[45] = in1[70] ^ in2[70];
    assign G[46] = in1[69] & in2[69];
    assign P[46] = in1[69] ^ in2[69];
    assign G[47] = in1[68] & in2[68];
    assign P[47] = in1[68] ^ in2[68];
    assign G[48] = in1[67] & in2[67];
    assign P[48] = in1[67] ^ in2[67];
    assign G[49] = in1[66] & in2[66];
    assign P[49] = in1[66] ^ in2[66];
    assign G[50] = in1[65] & in2[65];
    assign P[50] = in1[65] ^ in2[65];
    assign G[51] = in1[64] & in2[64];
    assign P[51] = in1[64] ^ in2[64];
    assign G[52] = in1[63] & in2[63];
    assign P[52] = in1[63] ^ in2[63];
    assign G[53] = in1[62] & in2[62];
    assign P[53] = in1[62] ^ in2[62];
    assign G[54] = in1[61] & in2[61];
    assign P[54] = in1[61] ^ in2[61];
    assign G[55] = in1[60] & in2[60];
    assign P[55] = in1[60] ^ in2[60];
    assign G[56] = in1[59] & in2[59];
    assign P[56] = in1[59] ^ in2[59];
    assign G[57] = in1[58] & in2[58];
    assign P[57] = in1[58] ^ in2[58];
    assign G[58] = in1[57] & in2[57];
    assign P[58] = in1[57] ^ in2[57];
    assign G[59] = in1[56] & in2[56];
    assign P[59] = in1[56] ^ in2[56];
    assign G[60] = in1[55] & in2[55];
    assign P[60] = in1[55] ^ in2[55];
    assign G[61] = in1[54] & in2[54];
    assign P[61] = in1[54] ^ in2[54];
    assign G[62] = in1[53] & in2[53];
    assign P[62] = in1[53] ^ in2[53];
    assign G[63] = in1[52] & in2[52];
    assign P[63] = in1[52] ^ in2[52];
    assign G[64] = in1[51] & in2[51];
    assign P[64] = in1[51] ^ in2[51];
    assign G[65] = in1[50] & in2[50];
    assign P[65] = in1[50] ^ in2[50];
    assign G[66] = in1[49] & in2[49];
    assign P[66] = in1[49] ^ in2[49];
    assign G[67] = in1[48] & in2[48];
    assign P[67] = in1[48] ^ in2[48];
    assign G[68] = in1[47] & in2[47];
    assign P[68] = in1[47] ^ in2[47];
    assign G[69] = in1[46] & in2[46];
    assign P[69] = in1[46] ^ in2[46];
    assign G[70] = in1[45] & in2[45];
    assign P[70] = in1[45] ^ in2[45];
    assign G[71] = in1[44] & in2[44];
    assign P[71] = in1[44] ^ in2[44];
    assign G[72] = in1[43] & in2[43];
    assign P[72] = in1[43] ^ in2[43];
    assign G[73] = in1[42] & in2[42];
    assign P[73] = in1[42] ^ in2[42];
    assign G[74] = in1[41] & in2[41];
    assign P[74] = in1[41] ^ in2[41];
    assign G[75] = in1[40] & in2[40];
    assign P[75] = in1[40] ^ in2[40];
    assign G[76] = in1[39] & in2[39];
    assign P[76] = in1[39] ^ in2[39];
    assign G[77] = in1[38] & in2[38];
    assign P[77] = in1[38] ^ in2[38];
    assign G[78] = in1[37] & in2[37];
    assign P[78] = in1[37] ^ in2[37];
    assign G[79] = in1[36] & in2[36];
    assign P[79] = in1[36] ^ in2[36];
    assign G[80] = in1[35] & in2[35];
    assign P[80] = in1[35] ^ in2[35];
    assign G[81] = in1[34] & in2[34];
    assign P[81] = in1[34] ^ in2[34];
    assign G[82] = in1[33] & in2[33];
    assign P[82] = in1[33] ^ in2[33];
    assign G[83] = in1[32] & in2[32];
    assign P[83] = in1[32] ^ in2[32];
    assign G[84] = in1[31] & in2[31];
    assign P[84] = in1[31] ^ in2[31];
    assign G[85] = in1[30] & in2[30];
    assign P[85] = in1[30] ^ in2[30];
    assign G[86] = in1[29] & in2[29];
    assign P[86] = in1[29] ^ in2[29];
    assign G[87] = in1[28] & in2[28];
    assign P[87] = in1[28] ^ in2[28];
    assign G[88] = in1[27] & in2[27];
    assign P[88] = in1[27] ^ in2[27];
    assign G[89] = in1[26] & in2[26];
    assign P[89] = in1[26] ^ in2[26];
    assign G[90] = in1[25] & in2[25];
    assign P[90] = in1[25] ^ in2[25];
    assign G[91] = in1[24] & in2[24];
    assign P[91] = in1[24] ^ in2[24];
    assign G[92] = in1[23] & in2[23];
    assign P[92] = in1[23] ^ in2[23];
    assign G[93] = in1[22] & in2[22];
    assign P[93] = in1[22] ^ in2[22];
    assign G[94] = in1[21] & in2[21];
    assign P[94] = in1[21] ^ in2[21];
    assign G[95] = in1[20] & in2[20];
    assign P[95] = in1[20] ^ in2[20];
    assign G[96] = in1[19] & in2[19];
    assign P[96] = in1[19] ^ in2[19];
    assign G[97] = in1[18] & in2[18];
    assign P[97] = in1[18] ^ in2[18];
    assign G[98] = in1[17] & in2[17];
    assign P[98] = in1[17] ^ in2[17];
    assign G[99] = in1[16] & in2[16];
    assign P[99] = in1[16] ^ in2[16];
    assign G[100] = in1[15] & in2[15];
    assign P[100] = in1[15] ^ in2[15];
    assign G[101] = in1[14] & in2[14];
    assign P[101] = in1[14] ^ in2[14];
    assign G[102] = in1[13] & in2[13];
    assign P[102] = in1[13] ^ in2[13];
    assign G[103] = in1[12] & in2[12];
    assign P[103] = in1[12] ^ in2[12];
    assign G[104] = in1[11] & in2[11];
    assign P[104] = in1[11] ^ in2[11];
    assign G[105] = in1[10] & in2[10];
    assign P[105] = in1[10] ^ in2[10];
    assign G[106] = in1[9] & in2[9];
    assign P[106] = in1[9] ^ in2[9];
    assign G[107] = in1[8] & in2[8];
    assign P[107] = in1[8] ^ in2[8];
    assign G[108] = in1[7] & in2[7];
    assign P[108] = in1[7] ^ in2[7];
    assign G[109] = in1[6] & in2[6];
    assign P[109] = in1[6] ^ in2[6];
    assign G[110] = in1[5] & in2[5];
    assign P[110] = in1[5] ^ in2[5];
    assign G[111] = in1[4] & in2[4];
    assign P[111] = in1[4] ^ in2[4];
    assign G[112] = in1[3] & in2[3];
    assign P[112] = in1[3] ^ in2[3];
    assign G[113] = in1[2] & in2[2];
    assign P[113] = in1[2] ^ in2[2];
    assign G[114] = in1[1] & in2[1];
    assign P[114] = in1[1] ^ in2[1];
    assign G[115] = in1[0] & in2[0];
    assign P[115] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign cout = G[115] | (P[115] & C[115]);
    assign sum = P ^ C;
endmodule

module CLA_115(output [114:0] sum, output cout, input [114:0] in1, input [114:0] in2);

    wire[114:0] G;
    wire[114:0] C;
    wire[114:0] P;

    assign G[0] = in1[114] & in2[114];
    assign P[0] = in1[114] ^ in2[114];
    assign G[1] = in1[113] & in2[113];
    assign P[1] = in1[113] ^ in2[113];
    assign G[2] = in1[112] & in2[112];
    assign P[2] = in1[112] ^ in2[112];
    assign G[3] = in1[111] & in2[111];
    assign P[3] = in1[111] ^ in2[111];
    assign G[4] = in1[110] & in2[110];
    assign P[4] = in1[110] ^ in2[110];
    assign G[5] = in1[109] & in2[109];
    assign P[5] = in1[109] ^ in2[109];
    assign G[6] = in1[108] & in2[108];
    assign P[6] = in1[108] ^ in2[108];
    assign G[7] = in1[107] & in2[107];
    assign P[7] = in1[107] ^ in2[107];
    assign G[8] = in1[106] & in2[106];
    assign P[8] = in1[106] ^ in2[106];
    assign G[9] = in1[105] & in2[105];
    assign P[9] = in1[105] ^ in2[105];
    assign G[10] = in1[104] & in2[104];
    assign P[10] = in1[104] ^ in2[104];
    assign G[11] = in1[103] & in2[103];
    assign P[11] = in1[103] ^ in2[103];
    assign G[12] = in1[102] & in2[102];
    assign P[12] = in1[102] ^ in2[102];
    assign G[13] = in1[101] & in2[101];
    assign P[13] = in1[101] ^ in2[101];
    assign G[14] = in1[100] & in2[100];
    assign P[14] = in1[100] ^ in2[100];
    assign G[15] = in1[99] & in2[99];
    assign P[15] = in1[99] ^ in2[99];
    assign G[16] = in1[98] & in2[98];
    assign P[16] = in1[98] ^ in2[98];
    assign G[17] = in1[97] & in2[97];
    assign P[17] = in1[97] ^ in2[97];
    assign G[18] = in1[96] & in2[96];
    assign P[18] = in1[96] ^ in2[96];
    assign G[19] = in1[95] & in2[95];
    assign P[19] = in1[95] ^ in2[95];
    assign G[20] = in1[94] & in2[94];
    assign P[20] = in1[94] ^ in2[94];
    assign G[21] = in1[93] & in2[93];
    assign P[21] = in1[93] ^ in2[93];
    assign G[22] = in1[92] & in2[92];
    assign P[22] = in1[92] ^ in2[92];
    assign G[23] = in1[91] & in2[91];
    assign P[23] = in1[91] ^ in2[91];
    assign G[24] = in1[90] & in2[90];
    assign P[24] = in1[90] ^ in2[90];
    assign G[25] = in1[89] & in2[89];
    assign P[25] = in1[89] ^ in2[89];
    assign G[26] = in1[88] & in2[88];
    assign P[26] = in1[88] ^ in2[88];
    assign G[27] = in1[87] & in2[87];
    assign P[27] = in1[87] ^ in2[87];
    assign G[28] = in1[86] & in2[86];
    assign P[28] = in1[86] ^ in2[86];
    assign G[29] = in1[85] & in2[85];
    assign P[29] = in1[85] ^ in2[85];
    assign G[30] = in1[84] & in2[84];
    assign P[30] = in1[84] ^ in2[84];
    assign G[31] = in1[83] & in2[83];
    assign P[31] = in1[83] ^ in2[83];
    assign G[32] = in1[82] & in2[82];
    assign P[32] = in1[82] ^ in2[82];
    assign G[33] = in1[81] & in2[81];
    assign P[33] = in1[81] ^ in2[81];
    assign G[34] = in1[80] & in2[80];
    assign P[34] = in1[80] ^ in2[80];
    assign G[35] = in1[79] & in2[79];
    assign P[35] = in1[79] ^ in2[79];
    assign G[36] = in1[78] & in2[78];
    assign P[36] = in1[78] ^ in2[78];
    assign G[37] = in1[77] & in2[77];
    assign P[37] = in1[77] ^ in2[77];
    assign G[38] = in1[76] & in2[76];
    assign P[38] = in1[76] ^ in2[76];
    assign G[39] = in1[75] & in2[75];
    assign P[39] = in1[75] ^ in2[75];
    assign G[40] = in1[74] & in2[74];
    assign P[40] = in1[74] ^ in2[74];
    assign G[41] = in1[73] & in2[73];
    assign P[41] = in1[73] ^ in2[73];
    assign G[42] = in1[72] & in2[72];
    assign P[42] = in1[72] ^ in2[72];
    assign G[43] = in1[71] & in2[71];
    assign P[43] = in1[71] ^ in2[71];
    assign G[44] = in1[70] & in2[70];
    assign P[44] = in1[70] ^ in2[70];
    assign G[45] = in1[69] & in2[69];
    assign P[45] = in1[69] ^ in2[69];
    assign G[46] = in1[68] & in2[68];
    assign P[46] = in1[68] ^ in2[68];
    assign G[47] = in1[67] & in2[67];
    assign P[47] = in1[67] ^ in2[67];
    assign G[48] = in1[66] & in2[66];
    assign P[48] = in1[66] ^ in2[66];
    assign G[49] = in1[65] & in2[65];
    assign P[49] = in1[65] ^ in2[65];
    assign G[50] = in1[64] & in2[64];
    assign P[50] = in1[64] ^ in2[64];
    assign G[51] = in1[63] & in2[63];
    assign P[51] = in1[63] ^ in2[63];
    assign G[52] = in1[62] & in2[62];
    assign P[52] = in1[62] ^ in2[62];
    assign G[53] = in1[61] & in2[61];
    assign P[53] = in1[61] ^ in2[61];
    assign G[54] = in1[60] & in2[60];
    assign P[54] = in1[60] ^ in2[60];
    assign G[55] = in1[59] & in2[59];
    assign P[55] = in1[59] ^ in2[59];
    assign G[56] = in1[58] & in2[58];
    assign P[56] = in1[58] ^ in2[58];
    assign G[57] = in1[57] & in2[57];
    assign P[57] = in1[57] ^ in2[57];
    assign G[58] = in1[56] & in2[56];
    assign P[58] = in1[56] ^ in2[56];
    assign G[59] = in1[55] & in2[55];
    assign P[59] = in1[55] ^ in2[55];
    assign G[60] = in1[54] & in2[54];
    assign P[60] = in1[54] ^ in2[54];
    assign G[61] = in1[53] & in2[53];
    assign P[61] = in1[53] ^ in2[53];
    assign G[62] = in1[52] & in2[52];
    assign P[62] = in1[52] ^ in2[52];
    assign G[63] = in1[51] & in2[51];
    assign P[63] = in1[51] ^ in2[51];
    assign G[64] = in1[50] & in2[50];
    assign P[64] = in1[50] ^ in2[50];
    assign G[65] = in1[49] & in2[49];
    assign P[65] = in1[49] ^ in2[49];
    assign G[66] = in1[48] & in2[48];
    assign P[66] = in1[48] ^ in2[48];
    assign G[67] = in1[47] & in2[47];
    assign P[67] = in1[47] ^ in2[47];
    assign G[68] = in1[46] & in2[46];
    assign P[68] = in1[46] ^ in2[46];
    assign G[69] = in1[45] & in2[45];
    assign P[69] = in1[45] ^ in2[45];
    assign G[70] = in1[44] & in2[44];
    assign P[70] = in1[44] ^ in2[44];
    assign G[71] = in1[43] & in2[43];
    assign P[71] = in1[43] ^ in2[43];
    assign G[72] = in1[42] & in2[42];
    assign P[72] = in1[42] ^ in2[42];
    assign G[73] = in1[41] & in2[41];
    assign P[73] = in1[41] ^ in2[41];
    assign G[74] = in1[40] & in2[40];
    assign P[74] = in1[40] ^ in2[40];
    assign G[75] = in1[39] & in2[39];
    assign P[75] = in1[39] ^ in2[39];
    assign G[76] = in1[38] & in2[38];
    assign P[76] = in1[38] ^ in2[38];
    assign G[77] = in1[37] & in2[37];
    assign P[77] = in1[37] ^ in2[37];
    assign G[78] = in1[36] & in2[36];
    assign P[78] = in1[36] ^ in2[36];
    assign G[79] = in1[35] & in2[35];
    assign P[79] = in1[35] ^ in2[35];
    assign G[80] = in1[34] & in2[34];
    assign P[80] = in1[34] ^ in2[34];
    assign G[81] = in1[33] & in2[33];
    assign P[81] = in1[33] ^ in2[33];
    assign G[82] = in1[32] & in2[32];
    assign P[82] = in1[32] ^ in2[32];
    assign G[83] = in1[31] & in2[31];
    assign P[83] = in1[31] ^ in2[31];
    assign G[84] = in1[30] & in2[30];
    assign P[84] = in1[30] ^ in2[30];
    assign G[85] = in1[29] & in2[29];
    assign P[85] = in1[29] ^ in2[29];
    assign G[86] = in1[28] & in2[28];
    assign P[86] = in1[28] ^ in2[28];
    assign G[87] = in1[27] & in2[27];
    assign P[87] = in1[27] ^ in2[27];
    assign G[88] = in1[26] & in2[26];
    assign P[88] = in1[26] ^ in2[26];
    assign G[89] = in1[25] & in2[25];
    assign P[89] = in1[25] ^ in2[25];
    assign G[90] = in1[24] & in2[24];
    assign P[90] = in1[24] ^ in2[24];
    assign G[91] = in1[23] & in2[23];
    assign P[91] = in1[23] ^ in2[23];
    assign G[92] = in1[22] & in2[22];
    assign P[92] = in1[22] ^ in2[22];
    assign G[93] = in1[21] & in2[21];
    assign P[93] = in1[21] ^ in2[21];
    assign G[94] = in1[20] & in2[20];
    assign P[94] = in1[20] ^ in2[20];
    assign G[95] = in1[19] & in2[19];
    assign P[95] = in1[19] ^ in2[19];
    assign G[96] = in1[18] & in2[18];
    assign P[96] = in1[18] ^ in2[18];
    assign G[97] = in1[17] & in2[17];
    assign P[97] = in1[17] ^ in2[17];
    assign G[98] = in1[16] & in2[16];
    assign P[98] = in1[16] ^ in2[16];
    assign G[99] = in1[15] & in2[15];
    assign P[99] = in1[15] ^ in2[15];
    assign G[100] = in1[14] & in2[14];
    assign P[100] = in1[14] ^ in2[14];
    assign G[101] = in1[13] & in2[13];
    assign P[101] = in1[13] ^ in2[13];
    assign G[102] = in1[12] & in2[12];
    assign P[102] = in1[12] ^ in2[12];
    assign G[103] = in1[11] & in2[11];
    assign P[103] = in1[11] ^ in2[11];
    assign G[104] = in1[10] & in2[10];
    assign P[104] = in1[10] ^ in2[10];
    assign G[105] = in1[9] & in2[9];
    assign P[105] = in1[9] ^ in2[9];
    assign G[106] = in1[8] & in2[8];
    assign P[106] = in1[8] ^ in2[8];
    assign G[107] = in1[7] & in2[7];
    assign P[107] = in1[7] ^ in2[7];
    assign G[108] = in1[6] & in2[6];
    assign P[108] = in1[6] ^ in2[6];
    assign G[109] = in1[5] & in2[5];
    assign P[109] = in1[5] ^ in2[5];
    assign G[110] = in1[4] & in2[4];
    assign P[110] = in1[4] ^ in2[4];
    assign G[111] = in1[3] & in2[3];
    assign P[111] = in1[3] ^ in2[3];
    assign G[112] = in1[2] & in2[2];
    assign P[112] = in1[2] ^ in2[2];
    assign G[113] = in1[1] & in2[1];
    assign P[113] = in1[1] ^ in2[1];
    assign G[114] = in1[0] & in2[0];
    assign P[114] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign cout = G[114] | (P[114] & C[114]);
    assign sum = P ^ C;
endmodule

module CLA_114(output [113:0] sum, output cout, input [113:0] in1, input [113:0] in2);

    wire[113:0] G;
    wire[113:0] C;
    wire[113:0] P;

    assign G[0] = in1[113] & in2[113];
    assign P[0] = in1[113] ^ in2[113];
    assign G[1] = in1[112] & in2[112];
    assign P[1] = in1[112] ^ in2[112];
    assign G[2] = in1[111] & in2[111];
    assign P[2] = in1[111] ^ in2[111];
    assign G[3] = in1[110] & in2[110];
    assign P[3] = in1[110] ^ in2[110];
    assign G[4] = in1[109] & in2[109];
    assign P[4] = in1[109] ^ in2[109];
    assign G[5] = in1[108] & in2[108];
    assign P[5] = in1[108] ^ in2[108];
    assign G[6] = in1[107] & in2[107];
    assign P[6] = in1[107] ^ in2[107];
    assign G[7] = in1[106] & in2[106];
    assign P[7] = in1[106] ^ in2[106];
    assign G[8] = in1[105] & in2[105];
    assign P[8] = in1[105] ^ in2[105];
    assign G[9] = in1[104] & in2[104];
    assign P[9] = in1[104] ^ in2[104];
    assign G[10] = in1[103] & in2[103];
    assign P[10] = in1[103] ^ in2[103];
    assign G[11] = in1[102] & in2[102];
    assign P[11] = in1[102] ^ in2[102];
    assign G[12] = in1[101] & in2[101];
    assign P[12] = in1[101] ^ in2[101];
    assign G[13] = in1[100] & in2[100];
    assign P[13] = in1[100] ^ in2[100];
    assign G[14] = in1[99] & in2[99];
    assign P[14] = in1[99] ^ in2[99];
    assign G[15] = in1[98] & in2[98];
    assign P[15] = in1[98] ^ in2[98];
    assign G[16] = in1[97] & in2[97];
    assign P[16] = in1[97] ^ in2[97];
    assign G[17] = in1[96] & in2[96];
    assign P[17] = in1[96] ^ in2[96];
    assign G[18] = in1[95] & in2[95];
    assign P[18] = in1[95] ^ in2[95];
    assign G[19] = in1[94] & in2[94];
    assign P[19] = in1[94] ^ in2[94];
    assign G[20] = in1[93] & in2[93];
    assign P[20] = in1[93] ^ in2[93];
    assign G[21] = in1[92] & in2[92];
    assign P[21] = in1[92] ^ in2[92];
    assign G[22] = in1[91] & in2[91];
    assign P[22] = in1[91] ^ in2[91];
    assign G[23] = in1[90] & in2[90];
    assign P[23] = in1[90] ^ in2[90];
    assign G[24] = in1[89] & in2[89];
    assign P[24] = in1[89] ^ in2[89];
    assign G[25] = in1[88] & in2[88];
    assign P[25] = in1[88] ^ in2[88];
    assign G[26] = in1[87] & in2[87];
    assign P[26] = in1[87] ^ in2[87];
    assign G[27] = in1[86] & in2[86];
    assign P[27] = in1[86] ^ in2[86];
    assign G[28] = in1[85] & in2[85];
    assign P[28] = in1[85] ^ in2[85];
    assign G[29] = in1[84] & in2[84];
    assign P[29] = in1[84] ^ in2[84];
    assign G[30] = in1[83] & in2[83];
    assign P[30] = in1[83] ^ in2[83];
    assign G[31] = in1[82] & in2[82];
    assign P[31] = in1[82] ^ in2[82];
    assign G[32] = in1[81] & in2[81];
    assign P[32] = in1[81] ^ in2[81];
    assign G[33] = in1[80] & in2[80];
    assign P[33] = in1[80] ^ in2[80];
    assign G[34] = in1[79] & in2[79];
    assign P[34] = in1[79] ^ in2[79];
    assign G[35] = in1[78] & in2[78];
    assign P[35] = in1[78] ^ in2[78];
    assign G[36] = in1[77] & in2[77];
    assign P[36] = in1[77] ^ in2[77];
    assign G[37] = in1[76] & in2[76];
    assign P[37] = in1[76] ^ in2[76];
    assign G[38] = in1[75] & in2[75];
    assign P[38] = in1[75] ^ in2[75];
    assign G[39] = in1[74] & in2[74];
    assign P[39] = in1[74] ^ in2[74];
    assign G[40] = in1[73] & in2[73];
    assign P[40] = in1[73] ^ in2[73];
    assign G[41] = in1[72] & in2[72];
    assign P[41] = in1[72] ^ in2[72];
    assign G[42] = in1[71] & in2[71];
    assign P[42] = in1[71] ^ in2[71];
    assign G[43] = in1[70] & in2[70];
    assign P[43] = in1[70] ^ in2[70];
    assign G[44] = in1[69] & in2[69];
    assign P[44] = in1[69] ^ in2[69];
    assign G[45] = in1[68] & in2[68];
    assign P[45] = in1[68] ^ in2[68];
    assign G[46] = in1[67] & in2[67];
    assign P[46] = in1[67] ^ in2[67];
    assign G[47] = in1[66] & in2[66];
    assign P[47] = in1[66] ^ in2[66];
    assign G[48] = in1[65] & in2[65];
    assign P[48] = in1[65] ^ in2[65];
    assign G[49] = in1[64] & in2[64];
    assign P[49] = in1[64] ^ in2[64];
    assign G[50] = in1[63] & in2[63];
    assign P[50] = in1[63] ^ in2[63];
    assign G[51] = in1[62] & in2[62];
    assign P[51] = in1[62] ^ in2[62];
    assign G[52] = in1[61] & in2[61];
    assign P[52] = in1[61] ^ in2[61];
    assign G[53] = in1[60] & in2[60];
    assign P[53] = in1[60] ^ in2[60];
    assign G[54] = in1[59] & in2[59];
    assign P[54] = in1[59] ^ in2[59];
    assign G[55] = in1[58] & in2[58];
    assign P[55] = in1[58] ^ in2[58];
    assign G[56] = in1[57] & in2[57];
    assign P[56] = in1[57] ^ in2[57];
    assign G[57] = in1[56] & in2[56];
    assign P[57] = in1[56] ^ in2[56];
    assign G[58] = in1[55] & in2[55];
    assign P[58] = in1[55] ^ in2[55];
    assign G[59] = in1[54] & in2[54];
    assign P[59] = in1[54] ^ in2[54];
    assign G[60] = in1[53] & in2[53];
    assign P[60] = in1[53] ^ in2[53];
    assign G[61] = in1[52] & in2[52];
    assign P[61] = in1[52] ^ in2[52];
    assign G[62] = in1[51] & in2[51];
    assign P[62] = in1[51] ^ in2[51];
    assign G[63] = in1[50] & in2[50];
    assign P[63] = in1[50] ^ in2[50];
    assign G[64] = in1[49] & in2[49];
    assign P[64] = in1[49] ^ in2[49];
    assign G[65] = in1[48] & in2[48];
    assign P[65] = in1[48] ^ in2[48];
    assign G[66] = in1[47] & in2[47];
    assign P[66] = in1[47] ^ in2[47];
    assign G[67] = in1[46] & in2[46];
    assign P[67] = in1[46] ^ in2[46];
    assign G[68] = in1[45] & in2[45];
    assign P[68] = in1[45] ^ in2[45];
    assign G[69] = in1[44] & in2[44];
    assign P[69] = in1[44] ^ in2[44];
    assign G[70] = in1[43] & in2[43];
    assign P[70] = in1[43] ^ in2[43];
    assign G[71] = in1[42] & in2[42];
    assign P[71] = in1[42] ^ in2[42];
    assign G[72] = in1[41] & in2[41];
    assign P[72] = in1[41] ^ in2[41];
    assign G[73] = in1[40] & in2[40];
    assign P[73] = in1[40] ^ in2[40];
    assign G[74] = in1[39] & in2[39];
    assign P[74] = in1[39] ^ in2[39];
    assign G[75] = in1[38] & in2[38];
    assign P[75] = in1[38] ^ in2[38];
    assign G[76] = in1[37] & in2[37];
    assign P[76] = in1[37] ^ in2[37];
    assign G[77] = in1[36] & in2[36];
    assign P[77] = in1[36] ^ in2[36];
    assign G[78] = in1[35] & in2[35];
    assign P[78] = in1[35] ^ in2[35];
    assign G[79] = in1[34] & in2[34];
    assign P[79] = in1[34] ^ in2[34];
    assign G[80] = in1[33] & in2[33];
    assign P[80] = in1[33] ^ in2[33];
    assign G[81] = in1[32] & in2[32];
    assign P[81] = in1[32] ^ in2[32];
    assign G[82] = in1[31] & in2[31];
    assign P[82] = in1[31] ^ in2[31];
    assign G[83] = in1[30] & in2[30];
    assign P[83] = in1[30] ^ in2[30];
    assign G[84] = in1[29] & in2[29];
    assign P[84] = in1[29] ^ in2[29];
    assign G[85] = in1[28] & in2[28];
    assign P[85] = in1[28] ^ in2[28];
    assign G[86] = in1[27] & in2[27];
    assign P[86] = in1[27] ^ in2[27];
    assign G[87] = in1[26] & in2[26];
    assign P[87] = in1[26] ^ in2[26];
    assign G[88] = in1[25] & in2[25];
    assign P[88] = in1[25] ^ in2[25];
    assign G[89] = in1[24] & in2[24];
    assign P[89] = in1[24] ^ in2[24];
    assign G[90] = in1[23] & in2[23];
    assign P[90] = in1[23] ^ in2[23];
    assign G[91] = in1[22] & in2[22];
    assign P[91] = in1[22] ^ in2[22];
    assign G[92] = in1[21] & in2[21];
    assign P[92] = in1[21] ^ in2[21];
    assign G[93] = in1[20] & in2[20];
    assign P[93] = in1[20] ^ in2[20];
    assign G[94] = in1[19] & in2[19];
    assign P[94] = in1[19] ^ in2[19];
    assign G[95] = in1[18] & in2[18];
    assign P[95] = in1[18] ^ in2[18];
    assign G[96] = in1[17] & in2[17];
    assign P[96] = in1[17] ^ in2[17];
    assign G[97] = in1[16] & in2[16];
    assign P[97] = in1[16] ^ in2[16];
    assign G[98] = in1[15] & in2[15];
    assign P[98] = in1[15] ^ in2[15];
    assign G[99] = in1[14] & in2[14];
    assign P[99] = in1[14] ^ in2[14];
    assign G[100] = in1[13] & in2[13];
    assign P[100] = in1[13] ^ in2[13];
    assign G[101] = in1[12] & in2[12];
    assign P[101] = in1[12] ^ in2[12];
    assign G[102] = in1[11] & in2[11];
    assign P[102] = in1[11] ^ in2[11];
    assign G[103] = in1[10] & in2[10];
    assign P[103] = in1[10] ^ in2[10];
    assign G[104] = in1[9] & in2[9];
    assign P[104] = in1[9] ^ in2[9];
    assign G[105] = in1[8] & in2[8];
    assign P[105] = in1[8] ^ in2[8];
    assign G[106] = in1[7] & in2[7];
    assign P[106] = in1[7] ^ in2[7];
    assign G[107] = in1[6] & in2[6];
    assign P[107] = in1[6] ^ in2[6];
    assign G[108] = in1[5] & in2[5];
    assign P[108] = in1[5] ^ in2[5];
    assign G[109] = in1[4] & in2[4];
    assign P[109] = in1[4] ^ in2[4];
    assign G[110] = in1[3] & in2[3];
    assign P[110] = in1[3] ^ in2[3];
    assign G[111] = in1[2] & in2[2];
    assign P[111] = in1[2] ^ in2[2];
    assign G[112] = in1[1] & in2[1];
    assign P[112] = in1[1] ^ in2[1];
    assign G[113] = in1[0] & in2[0];
    assign P[113] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign cout = G[113] | (P[113] & C[113]);
    assign sum = P ^ C;
endmodule

module CLA_113(output [112:0] sum, output cout, input [112:0] in1, input [112:0] in2);

    wire[112:0] G;
    wire[112:0] C;
    wire[112:0] P;

    assign G[0] = in1[112] & in2[112];
    assign P[0] = in1[112] ^ in2[112];
    assign G[1] = in1[111] & in2[111];
    assign P[1] = in1[111] ^ in2[111];
    assign G[2] = in1[110] & in2[110];
    assign P[2] = in1[110] ^ in2[110];
    assign G[3] = in1[109] & in2[109];
    assign P[3] = in1[109] ^ in2[109];
    assign G[4] = in1[108] & in2[108];
    assign P[4] = in1[108] ^ in2[108];
    assign G[5] = in1[107] & in2[107];
    assign P[5] = in1[107] ^ in2[107];
    assign G[6] = in1[106] & in2[106];
    assign P[6] = in1[106] ^ in2[106];
    assign G[7] = in1[105] & in2[105];
    assign P[7] = in1[105] ^ in2[105];
    assign G[8] = in1[104] & in2[104];
    assign P[8] = in1[104] ^ in2[104];
    assign G[9] = in1[103] & in2[103];
    assign P[9] = in1[103] ^ in2[103];
    assign G[10] = in1[102] & in2[102];
    assign P[10] = in1[102] ^ in2[102];
    assign G[11] = in1[101] & in2[101];
    assign P[11] = in1[101] ^ in2[101];
    assign G[12] = in1[100] & in2[100];
    assign P[12] = in1[100] ^ in2[100];
    assign G[13] = in1[99] & in2[99];
    assign P[13] = in1[99] ^ in2[99];
    assign G[14] = in1[98] & in2[98];
    assign P[14] = in1[98] ^ in2[98];
    assign G[15] = in1[97] & in2[97];
    assign P[15] = in1[97] ^ in2[97];
    assign G[16] = in1[96] & in2[96];
    assign P[16] = in1[96] ^ in2[96];
    assign G[17] = in1[95] & in2[95];
    assign P[17] = in1[95] ^ in2[95];
    assign G[18] = in1[94] & in2[94];
    assign P[18] = in1[94] ^ in2[94];
    assign G[19] = in1[93] & in2[93];
    assign P[19] = in1[93] ^ in2[93];
    assign G[20] = in1[92] & in2[92];
    assign P[20] = in1[92] ^ in2[92];
    assign G[21] = in1[91] & in2[91];
    assign P[21] = in1[91] ^ in2[91];
    assign G[22] = in1[90] & in2[90];
    assign P[22] = in1[90] ^ in2[90];
    assign G[23] = in1[89] & in2[89];
    assign P[23] = in1[89] ^ in2[89];
    assign G[24] = in1[88] & in2[88];
    assign P[24] = in1[88] ^ in2[88];
    assign G[25] = in1[87] & in2[87];
    assign P[25] = in1[87] ^ in2[87];
    assign G[26] = in1[86] & in2[86];
    assign P[26] = in1[86] ^ in2[86];
    assign G[27] = in1[85] & in2[85];
    assign P[27] = in1[85] ^ in2[85];
    assign G[28] = in1[84] & in2[84];
    assign P[28] = in1[84] ^ in2[84];
    assign G[29] = in1[83] & in2[83];
    assign P[29] = in1[83] ^ in2[83];
    assign G[30] = in1[82] & in2[82];
    assign P[30] = in1[82] ^ in2[82];
    assign G[31] = in1[81] & in2[81];
    assign P[31] = in1[81] ^ in2[81];
    assign G[32] = in1[80] & in2[80];
    assign P[32] = in1[80] ^ in2[80];
    assign G[33] = in1[79] & in2[79];
    assign P[33] = in1[79] ^ in2[79];
    assign G[34] = in1[78] & in2[78];
    assign P[34] = in1[78] ^ in2[78];
    assign G[35] = in1[77] & in2[77];
    assign P[35] = in1[77] ^ in2[77];
    assign G[36] = in1[76] & in2[76];
    assign P[36] = in1[76] ^ in2[76];
    assign G[37] = in1[75] & in2[75];
    assign P[37] = in1[75] ^ in2[75];
    assign G[38] = in1[74] & in2[74];
    assign P[38] = in1[74] ^ in2[74];
    assign G[39] = in1[73] & in2[73];
    assign P[39] = in1[73] ^ in2[73];
    assign G[40] = in1[72] & in2[72];
    assign P[40] = in1[72] ^ in2[72];
    assign G[41] = in1[71] & in2[71];
    assign P[41] = in1[71] ^ in2[71];
    assign G[42] = in1[70] & in2[70];
    assign P[42] = in1[70] ^ in2[70];
    assign G[43] = in1[69] & in2[69];
    assign P[43] = in1[69] ^ in2[69];
    assign G[44] = in1[68] & in2[68];
    assign P[44] = in1[68] ^ in2[68];
    assign G[45] = in1[67] & in2[67];
    assign P[45] = in1[67] ^ in2[67];
    assign G[46] = in1[66] & in2[66];
    assign P[46] = in1[66] ^ in2[66];
    assign G[47] = in1[65] & in2[65];
    assign P[47] = in1[65] ^ in2[65];
    assign G[48] = in1[64] & in2[64];
    assign P[48] = in1[64] ^ in2[64];
    assign G[49] = in1[63] & in2[63];
    assign P[49] = in1[63] ^ in2[63];
    assign G[50] = in1[62] & in2[62];
    assign P[50] = in1[62] ^ in2[62];
    assign G[51] = in1[61] & in2[61];
    assign P[51] = in1[61] ^ in2[61];
    assign G[52] = in1[60] & in2[60];
    assign P[52] = in1[60] ^ in2[60];
    assign G[53] = in1[59] & in2[59];
    assign P[53] = in1[59] ^ in2[59];
    assign G[54] = in1[58] & in2[58];
    assign P[54] = in1[58] ^ in2[58];
    assign G[55] = in1[57] & in2[57];
    assign P[55] = in1[57] ^ in2[57];
    assign G[56] = in1[56] & in2[56];
    assign P[56] = in1[56] ^ in2[56];
    assign G[57] = in1[55] & in2[55];
    assign P[57] = in1[55] ^ in2[55];
    assign G[58] = in1[54] & in2[54];
    assign P[58] = in1[54] ^ in2[54];
    assign G[59] = in1[53] & in2[53];
    assign P[59] = in1[53] ^ in2[53];
    assign G[60] = in1[52] & in2[52];
    assign P[60] = in1[52] ^ in2[52];
    assign G[61] = in1[51] & in2[51];
    assign P[61] = in1[51] ^ in2[51];
    assign G[62] = in1[50] & in2[50];
    assign P[62] = in1[50] ^ in2[50];
    assign G[63] = in1[49] & in2[49];
    assign P[63] = in1[49] ^ in2[49];
    assign G[64] = in1[48] & in2[48];
    assign P[64] = in1[48] ^ in2[48];
    assign G[65] = in1[47] & in2[47];
    assign P[65] = in1[47] ^ in2[47];
    assign G[66] = in1[46] & in2[46];
    assign P[66] = in1[46] ^ in2[46];
    assign G[67] = in1[45] & in2[45];
    assign P[67] = in1[45] ^ in2[45];
    assign G[68] = in1[44] & in2[44];
    assign P[68] = in1[44] ^ in2[44];
    assign G[69] = in1[43] & in2[43];
    assign P[69] = in1[43] ^ in2[43];
    assign G[70] = in1[42] & in2[42];
    assign P[70] = in1[42] ^ in2[42];
    assign G[71] = in1[41] & in2[41];
    assign P[71] = in1[41] ^ in2[41];
    assign G[72] = in1[40] & in2[40];
    assign P[72] = in1[40] ^ in2[40];
    assign G[73] = in1[39] & in2[39];
    assign P[73] = in1[39] ^ in2[39];
    assign G[74] = in1[38] & in2[38];
    assign P[74] = in1[38] ^ in2[38];
    assign G[75] = in1[37] & in2[37];
    assign P[75] = in1[37] ^ in2[37];
    assign G[76] = in1[36] & in2[36];
    assign P[76] = in1[36] ^ in2[36];
    assign G[77] = in1[35] & in2[35];
    assign P[77] = in1[35] ^ in2[35];
    assign G[78] = in1[34] & in2[34];
    assign P[78] = in1[34] ^ in2[34];
    assign G[79] = in1[33] & in2[33];
    assign P[79] = in1[33] ^ in2[33];
    assign G[80] = in1[32] & in2[32];
    assign P[80] = in1[32] ^ in2[32];
    assign G[81] = in1[31] & in2[31];
    assign P[81] = in1[31] ^ in2[31];
    assign G[82] = in1[30] & in2[30];
    assign P[82] = in1[30] ^ in2[30];
    assign G[83] = in1[29] & in2[29];
    assign P[83] = in1[29] ^ in2[29];
    assign G[84] = in1[28] & in2[28];
    assign P[84] = in1[28] ^ in2[28];
    assign G[85] = in1[27] & in2[27];
    assign P[85] = in1[27] ^ in2[27];
    assign G[86] = in1[26] & in2[26];
    assign P[86] = in1[26] ^ in2[26];
    assign G[87] = in1[25] & in2[25];
    assign P[87] = in1[25] ^ in2[25];
    assign G[88] = in1[24] & in2[24];
    assign P[88] = in1[24] ^ in2[24];
    assign G[89] = in1[23] & in2[23];
    assign P[89] = in1[23] ^ in2[23];
    assign G[90] = in1[22] & in2[22];
    assign P[90] = in1[22] ^ in2[22];
    assign G[91] = in1[21] & in2[21];
    assign P[91] = in1[21] ^ in2[21];
    assign G[92] = in1[20] & in2[20];
    assign P[92] = in1[20] ^ in2[20];
    assign G[93] = in1[19] & in2[19];
    assign P[93] = in1[19] ^ in2[19];
    assign G[94] = in1[18] & in2[18];
    assign P[94] = in1[18] ^ in2[18];
    assign G[95] = in1[17] & in2[17];
    assign P[95] = in1[17] ^ in2[17];
    assign G[96] = in1[16] & in2[16];
    assign P[96] = in1[16] ^ in2[16];
    assign G[97] = in1[15] & in2[15];
    assign P[97] = in1[15] ^ in2[15];
    assign G[98] = in1[14] & in2[14];
    assign P[98] = in1[14] ^ in2[14];
    assign G[99] = in1[13] & in2[13];
    assign P[99] = in1[13] ^ in2[13];
    assign G[100] = in1[12] & in2[12];
    assign P[100] = in1[12] ^ in2[12];
    assign G[101] = in1[11] & in2[11];
    assign P[101] = in1[11] ^ in2[11];
    assign G[102] = in1[10] & in2[10];
    assign P[102] = in1[10] ^ in2[10];
    assign G[103] = in1[9] & in2[9];
    assign P[103] = in1[9] ^ in2[9];
    assign G[104] = in1[8] & in2[8];
    assign P[104] = in1[8] ^ in2[8];
    assign G[105] = in1[7] & in2[7];
    assign P[105] = in1[7] ^ in2[7];
    assign G[106] = in1[6] & in2[6];
    assign P[106] = in1[6] ^ in2[6];
    assign G[107] = in1[5] & in2[5];
    assign P[107] = in1[5] ^ in2[5];
    assign G[108] = in1[4] & in2[4];
    assign P[108] = in1[4] ^ in2[4];
    assign G[109] = in1[3] & in2[3];
    assign P[109] = in1[3] ^ in2[3];
    assign G[110] = in1[2] & in2[2];
    assign P[110] = in1[2] ^ in2[2];
    assign G[111] = in1[1] & in2[1];
    assign P[111] = in1[1] ^ in2[1];
    assign G[112] = in1[0] & in2[0];
    assign P[112] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign cout = G[112] | (P[112] & C[112]);
    assign sum = P ^ C;
endmodule

module CLA_112(output [111:0] sum, output cout, input [111:0] in1, input [111:0] in2);

    wire[111:0] G;
    wire[111:0] C;
    wire[111:0] P;

    assign G[0] = in1[111] & in2[111];
    assign P[0] = in1[111] ^ in2[111];
    assign G[1] = in1[110] & in2[110];
    assign P[1] = in1[110] ^ in2[110];
    assign G[2] = in1[109] & in2[109];
    assign P[2] = in1[109] ^ in2[109];
    assign G[3] = in1[108] & in2[108];
    assign P[3] = in1[108] ^ in2[108];
    assign G[4] = in1[107] & in2[107];
    assign P[4] = in1[107] ^ in2[107];
    assign G[5] = in1[106] & in2[106];
    assign P[5] = in1[106] ^ in2[106];
    assign G[6] = in1[105] & in2[105];
    assign P[6] = in1[105] ^ in2[105];
    assign G[7] = in1[104] & in2[104];
    assign P[7] = in1[104] ^ in2[104];
    assign G[8] = in1[103] & in2[103];
    assign P[8] = in1[103] ^ in2[103];
    assign G[9] = in1[102] & in2[102];
    assign P[9] = in1[102] ^ in2[102];
    assign G[10] = in1[101] & in2[101];
    assign P[10] = in1[101] ^ in2[101];
    assign G[11] = in1[100] & in2[100];
    assign P[11] = in1[100] ^ in2[100];
    assign G[12] = in1[99] & in2[99];
    assign P[12] = in1[99] ^ in2[99];
    assign G[13] = in1[98] & in2[98];
    assign P[13] = in1[98] ^ in2[98];
    assign G[14] = in1[97] & in2[97];
    assign P[14] = in1[97] ^ in2[97];
    assign G[15] = in1[96] & in2[96];
    assign P[15] = in1[96] ^ in2[96];
    assign G[16] = in1[95] & in2[95];
    assign P[16] = in1[95] ^ in2[95];
    assign G[17] = in1[94] & in2[94];
    assign P[17] = in1[94] ^ in2[94];
    assign G[18] = in1[93] & in2[93];
    assign P[18] = in1[93] ^ in2[93];
    assign G[19] = in1[92] & in2[92];
    assign P[19] = in1[92] ^ in2[92];
    assign G[20] = in1[91] & in2[91];
    assign P[20] = in1[91] ^ in2[91];
    assign G[21] = in1[90] & in2[90];
    assign P[21] = in1[90] ^ in2[90];
    assign G[22] = in1[89] & in2[89];
    assign P[22] = in1[89] ^ in2[89];
    assign G[23] = in1[88] & in2[88];
    assign P[23] = in1[88] ^ in2[88];
    assign G[24] = in1[87] & in2[87];
    assign P[24] = in1[87] ^ in2[87];
    assign G[25] = in1[86] & in2[86];
    assign P[25] = in1[86] ^ in2[86];
    assign G[26] = in1[85] & in2[85];
    assign P[26] = in1[85] ^ in2[85];
    assign G[27] = in1[84] & in2[84];
    assign P[27] = in1[84] ^ in2[84];
    assign G[28] = in1[83] & in2[83];
    assign P[28] = in1[83] ^ in2[83];
    assign G[29] = in1[82] & in2[82];
    assign P[29] = in1[82] ^ in2[82];
    assign G[30] = in1[81] & in2[81];
    assign P[30] = in1[81] ^ in2[81];
    assign G[31] = in1[80] & in2[80];
    assign P[31] = in1[80] ^ in2[80];
    assign G[32] = in1[79] & in2[79];
    assign P[32] = in1[79] ^ in2[79];
    assign G[33] = in1[78] & in2[78];
    assign P[33] = in1[78] ^ in2[78];
    assign G[34] = in1[77] & in2[77];
    assign P[34] = in1[77] ^ in2[77];
    assign G[35] = in1[76] & in2[76];
    assign P[35] = in1[76] ^ in2[76];
    assign G[36] = in1[75] & in2[75];
    assign P[36] = in1[75] ^ in2[75];
    assign G[37] = in1[74] & in2[74];
    assign P[37] = in1[74] ^ in2[74];
    assign G[38] = in1[73] & in2[73];
    assign P[38] = in1[73] ^ in2[73];
    assign G[39] = in1[72] & in2[72];
    assign P[39] = in1[72] ^ in2[72];
    assign G[40] = in1[71] & in2[71];
    assign P[40] = in1[71] ^ in2[71];
    assign G[41] = in1[70] & in2[70];
    assign P[41] = in1[70] ^ in2[70];
    assign G[42] = in1[69] & in2[69];
    assign P[42] = in1[69] ^ in2[69];
    assign G[43] = in1[68] & in2[68];
    assign P[43] = in1[68] ^ in2[68];
    assign G[44] = in1[67] & in2[67];
    assign P[44] = in1[67] ^ in2[67];
    assign G[45] = in1[66] & in2[66];
    assign P[45] = in1[66] ^ in2[66];
    assign G[46] = in1[65] & in2[65];
    assign P[46] = in1[65] ^ in2[65];
    assign G[47] = in1[64] & in2[64];
    assign P[47] = in1[64] ^ in2[64];
    assign G[48] = in1[63] & in2[63];
    assign P[48] = in1[63] ^ in2[63];
    assign G[49] = in1[62] & in2[62];
    assign P[49] = in1[62] ^ in2[62];
    assign G[50] = in1[61] & in2[61];
    assign P[50] = in1[61] ^ in2[61];
    assign G[51] = in1[60] & in2[60];
    assign P[51] = in1[60] ^ in2[60];
    assign G[52] = in1[59] & in2[59];
    assign P[52] = in1[59] ^ in2[59];
    assign G[53] = in1[58] & in2[58];
    assign P[53] = in1[58] ^ in2[58];
    assign G[54] = in1[57] & in2[57];
    assign P[54] = in1[57] ^ in2[57];
    assign G[55] = in1[56] & in2[56];
    assign P[55] = in1[56] ^ in2[56];
    assign G[56] = in1[55] & in2[55];
    assign P[56] = in1[55] ^ in2[55];
    assign G[57] = in1[54] & in2[54];
    assign P[57] = in1[54] ^ in2[54];
    assign G[58] = in1[53] & in2[53];
    assign P[58] = in1[53] ^ in2[53];
    assign G[59] = in1[52] & in2[52];
    assign P[59] = in1[52] ^ in2[52];
    assign G[60] = in1[51] & in2[51];
    assign P[60] = in1[51] ^ in2[51];
    assign G[61] = in1[50] & in2[50];
    assign P[61] = in1[50] ^ in2[50];
    assign G[62] = in1[49] & in2[49];
    assign P[62] = in1[49] ^ in2[49];
    assign G[63] = in1[48] & in2[48];
    assign P[63] = in1[48] ^ in2[48];
    assign G[64] = in1[47] & in2[47];
    assign P[64] = in1[47] ^ in2[47];
    assign G[65] = in1[46] & in2[46];
    assign P[65] = in1[46] ^ in2[46];
    assign G[66] = in1[45] & in2[45];
    assign P[66] = in1[45] ^ in2[45];
    assign G[67] = in1[44] & in2[44];
    assign P[67] = in1[44] ^ in2[44];
    assign G[68] = in1[43] & in2[43];
    assign P[68] = in1[43] ^ in2[43];
    assign G[69] = in1[42] & in2[42];
    assign P[69] = in1[42] ^ in2[42];
    assign G[70] = in1[41] & in2[41];
    assign P[70] = in1[41] ^ in2[41];
    assign G[71] = in1[40] & in2[40];
    assign P[71] = in1[40] ^ in2[40];
    assign G[72] = in1[39] & in2[39];
    assign P[72] = in1[39] ^ in2[39];
    assign G[73] = in1[38] & in2[38];
    assign P[73] = in1[38] ^ in2[38];
    assign G[74] = in1[37] & in2[37];
    assign P[74] = in1[37] ^ in2[37];
    assign G[75] = in1[36] & in2[36];
    assign P[75] = in1[36] ^ in2[36];
    assign G[76] = in1[35] & in2[35];
    assign P[76] = in1[35] ^ in2[35];
    assign G[77] = in1[34] & in2[34];
    assign P[77] = in1[34] ^ in2[34];
    assign G[78] = in1[33] & in2[33];
    assign P[78] = in1[33] ^ in2[33];
    assign G[79] = in1[32] & in2[32];
    assign P[79] = in1[32] ^ in2[32];
    assign G[80] = in1[31] & in2[31];
    assign P[80] = in1[31] ^ in2[31];
    assign G[81] = in1[30] & in2[30];
    assign P[81] = in1[30] ^ in2[30];
    assign G[82] = in1[29] & in2[29];
    assign P[82] = in1[29] ^ in2[29];
    assign G[83] = in1[28] & in2[28];
    assign P[83] = in1[28] ^ in2[28];
    assign G[84] = in1[27] & in2[27];
    assign P[84] = in1[27] ^ in2[27];
    assign G[85] = in1[26] & in2[26];
    assign P[85] = in1[26] ^ in2[26];
    assign G[86] = in1[25] & in2[25];
    assign P[86] = in1[25] ^ in2[25];
    assign G[87] = in1[24] & in2[24];
    assign P[87] = in1[24] ^ in2[24];
    assign G[88] = in1[23] & in2[23];
    assign P[88] = in1[23] ^ in2[23];
    assign G[89] = in1[22] & in2[22];
    assign P[89] = in1[22] ^ in2[22];
    assign G[90] = in1[21] & in2[21];
    assign P[90] = in1[21] ^ in2[21];
    assign G[91] = in1[20] & in2[20];
    assign P[91] = in1[20] ^ in2[20];
    assign G[92] = in1[19] & in2[19];
    assign P[92] = in1[19] ^ in2[19];
    assign G[93] = in1[18] & in2[18];
    assign P[93] = in1[18] ^ in2[18];
    assign G[94] = in1[17] & in2[17];
    assign P[94] = in1[17] ^ in2[17];
    assign G[95] = in1[16] & in2[16];
    assign P[95] = in1[16] ^ in2[16];
    assign G[96] = in1[15] & in2[15];
    assign P[96] = in1[15] ^ in2[15];
    assign G[97] = in1[14] & in2[14];
    assign P[97] = in1[14] ^ in2[14];
    assign G[98] = in1[13] & in2[13];
    assign P[98] = in1[13] ^ in2[13];
    assign G[99] = in1[12] & in2[12];
    assign P[99] = in1[12] ^ in2[12];
    assign G[100] = in1[11] & in2[11];
    assign P[100] = in1[11] ^ in2[11];
    assign G[101] = in1[10] & in2[10];
    assign P[101] = in1[10] ^ in2[10];
    assign G[102] = in1[9] & in2[9];
    assign P[102] = in1[9] ^ in2[9];
    assign G[103] = in1[8] & in2[8];
    assign P[103] = in1[8] ^ in2[8];
    assign G[104] = in1[7] & in2[7];
    assign P[104] = in1[7] ^ in2[7];
    assign G[105] = in1[6] & in2[6];
    assign P[105] = in1[6] ^ in2[6];
    assign G[106] = in1[5] & in2[5];
    assign P[106] = in1[5] ^ in2[5];
    assign G[107] = in1[4] & in2[4];
    assign P[107] = in1[4] ^ in2[4];
    assign G[108] = in1[3] & in2[3];
    assign P[108] = in1[3] ^ in2[3];
    assign G[109] = in1[2] & in2[2];
    assign P[109] = in1[2] ^ in2[2];
    assign G[110] = in1[1] & in2[1];
    assign P[110] = in1[1] ^ in2[1];
    assign G[111] = in1[0] & in2[0];
    assign P[111] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign cout = G[111] | (P[111] & C[111]);
    assign sum = P ^ C;
endmodule

module CLA_111(output [110:0] sum, output cout, input [110:0] in1, input [110:0] in2);

    wire[110:0] G;
    wire[110:0] C;
    wire[110:0] P;

    assign G[0] = in1[110] & in2[110];
    assign P[0] = in1[110] ^ in2[110];
    assign G[1] = in1[109] & in2[109];
    assign P[1] = in1[109] ^ in2[109];
    assign G[2] = in1[108] & in2[108];
    assign P[2] = in1[108] ^ in2[108];
    assign G[3] = in1[107] & in2[107];
    assign P[3] = in1[107] ^ in2[107];
    assign G[4] = in1[106] & in2[106];
    assign P[4] = in1[106] ^ in2[106];
    assign G[5] = in1[105] & in2[105];
    assign P[5] = in1[105] ^ in2[105];
    assign G[6] = in1[104] & in2[104];
    assign P[6] = in1[104] ^ in2[104];
    assign G[7] = in1[103] & in2[103];
    assign P[7] = in1[103] ^ in2[103];
    assign G[8] = in1[102] & in2[102];
    assign P[8] = in1[102] ^ in2[102];
    assign G[9] = in1[101] & in2[101];
    assign P[9] = in1[101] ^ in2[101];
    assign G[10] = in1[100] & in2[100];
    assign P[10] = in1[100] ^ in2[100];
    assign G[11] = in1[99] & in2[99];
    assign P[11] = in1[99] ^ in2[99];
    assign G[12] = in1[98] & in2[98];
    assign P[12] = in1[98] ^ in2[98];
    assign G[13] = in1[97] & in2[97];
    assign P[13] = in1[97] ^ in2[97];
    assign G[14] = in1[96] & in2[96];
    assign P[14] = in1[96] ^ in2[96];
    assign G[15] = in1[95] & in2[95];
    assign P[15] = in1[95] ^ in2[95];
    assign G[16] = in1[94] & in2[94];
    assign P[16] = in1[94] ^ in2[94];
    assign G[17] = in1[93] & in2[93];
    assign P[17] = in1[93] ^ in2[93];
    assign G[18] = in1[92] & in2[92];
    assign P[18] = in1[92] ^ in2[92];
    assign G[19] = in1[91] & in2[91];
    assign P[19] = in1[91] ^ in2[91];
    assign G[20] = in1[90] & in2[90];
    assign P[20] = in1[90] ^ in2[90];
    assign G[21] = in1[89] & in2[89];
    assign P[21] = in1[89] ^ in2[89];
    assign G[22] = in1[88] & in2[88];
    assign P[22] = in1[88] ^ in2[88];
    assign G[23] = in1[87] & in2[87];
    assign P[23] = in1[87] ^ in2[87];
    assign G[24] = in1[86] & in2[86];
    assign P[24] = in1[86] ^ in2[86];
    assign G[25] = in1[85] & in2[85];
    assign P[25] = in1[85] ^ in2[85];
    assign G[26] = in1[84] & in2[84];
    assign P[26] = in1[84] ^ in2[84];
    assign G[27] = in1[83] & in2[83];
    assign P[27] = in1[83] ^ in2[83];
    assign G[28] = in1[82] & in2[82];
    assign P[28] = in1[82] ^ in2[82];
    assign G[29] = in1[81] & in2[81];
    assign P[29] = in1[81] ^ in2[81];
    assign G[30] = in1[80] & in2[80];
    assign P[30] = in1[80] ^ in2[80];
    assign G[31] = in1[79] & in2[79];
    assign P[31] = in1[79] ^ in2[79];
    assign G[32] = in1[78] & in2[78];
    assign P[32] = in1[78] ^ in2[78];
    assign G[33] = in1[77] & in2[77];
    assign P[33] = in1[77] ^ in2[77];
    assign G[34] = in1[76] & in2[76];
    assign P[34] = in1[76] ^ in2[76];
    assign G[35] = in1[75] & in2[75];
    assign P[35] = in1[75] ^ in2[75];
    assign G[36] = in1[74] & in2[74];
    assign P[36] = in1[74] ^ in2[74];
    assign G[37] = in1[73] & in2[73];
    assign P[37] = in1[73] ^ in2[73];
    assign G[38] = in1[72] & in2[72];
    assign P[38] = in1[72] ^ in2[72];
    assign G[39] = in1[71] & in2[71];
    assign P[39] = in1[71] ^ in2[71];
    assign G[40] = in1[70] & in2[70];
    assign P[40] = in1[70] ^ in2[70];
    assign G[41] = in1[69] & in2[69];
    assign P[41] = in1[69] ^ in2[69];
    assign G[42] = in1[68] & in2[68];
    assign P[42] = in1[68] ^ in2[68];
    assign G[43] = in1[67] & in2[67];
    assign P[43] = in1[67] ^ in2[67];
    assign G[44] = in1[66] & in2[66];
    assign P[44] = in1[66] ^ in2[66];
    assign G[45] = in1[65] & in2[65];
    assign P[45] = in1[65] ^ in2[65];
    assign G[46] = in1[64] & in2[64];
    assign P[46] = in1[64] ^ in2[64];
    assign G[47] = in1[63] & in2[63];
    assign P[47] = in1[63] ^ in2[63];
    assign G[48] = in1[62] & in2[62];
    assign P[48] = in1[62] ^ in2[62];
    assign G[49] = in1[61] & in2[61];
    assign P[49] = in1[61] ^ in2[61];
    assign G[50] = in1[60] & in2[60];
    assign P[50] = in1[60] ^ in2[60];
    assign G[51] = in1[59] & in2[59];
    assign P[51] = in1[59] ^ in2[59];
    assign G[52] = in1[58] & in2[58];
    assign P[52] = in1[58] ^ in2[58];
    assign G[53] = in1[57] & in2[57];
    assign P[53] = in1[57] ^ in2[57];
    assign G[54] = in1[56] & in2[56];
    assign P[54] = in1[56] ^ in2[56];
    assign G[55] = in1[55] & in2[55];
    assign P[55] = in1[55] ^ in2[55];
    assign G[56] = in1[54] & in2[54];
    assign P[56] = in1[54] ^ in2[54];
    assign G[57] = in1[53] & in2[53];
    assign P[57] = in1[53] ^ in2[53];
    assign G[58] = in1[52] & in2[52];
    assign P[58] = in1[52] ^ in2[52];
    assign G[59] = in1[51] & in2[51];
    assign P[59] = in1[51] ^ in2[51];
    assign G[60] = in1[50] & in2[50];
    assign P[60] = in1[50] ^ in2[50];
    assign G[61] = in1[49] & in2[49];
    assign P[61] = in1[49] ^ in2[49];
    assign G[62] = in1[48] & in2[48];
    assign P[62] = in1[48] ^ in2[48];
    assign G[63] = in1[47] & in2[47];
    assign P[63] = in1[47] ^ in2[47];
    assign G[64] = in1[46] & in2[46];
    assign P[64] = in1[46] ^ in2[46];
    assign G[65] = in1[45] & in2[45];
    assign P[65] = in1[45] ^ in2[45];
    assign G[66] = in1[44] & in2[44];
    assign P[66] = in1[44] ^ in2[44];
    assign G[67] = in1[43] & in2[43];
    assign P[67] = in1[43] ^ in2[43];
    assign G[68] = in1[42] & in2[42];
    assign P[68] = in1[42] ^ in2[42];
    assign G[69] = in1[41] & in2[41];
    assign P[69] = in1[41] ^ in2[41];
    assign G[70] = in1[40] & in2[40];
    assign P[70] = in1[40] ^ in2[40];
    assign G[71] = in1[39] & in2[39];
    assign P[71] = in1[39] ^ in2[39];
    assign G[72] = in1[38] & in2[38];
    assign P[72] = in1[38] ^ in2[38];
    assign G[73] = in1[37] & in2[37];
    assign P[73] = in1[37] ^ in2[37];
    assign G[74] = in1[36] & in2[36];
    assign P[74] = in1[36] ^ in2[36];
    assign G[75] = in1[35] & in2[35];
    assign P[75] = in1[35] ^ in2[35];
    assign G[76] = in1[34] & in2[34];
    assign P[76] = in1[34] ^ in2[34];
    assign G[77] = in1[33] & in2[33];
    assign P[77] = in1[33] ^ in2[33];
    assign G[78] = in1[32] & in2[32];
    assign P[78] = in1[32] ^ in2[32];
    assign G[79] = in1[31] & in2[31];
    assign P[79] = in1[31] ^ in2[31];
    assign G[80] = in1[30] & in2[30];
    assign P[80] = in1[30] ^ in2[30];
    assign G[81] = in1[29] & in2[29];
    assign P[81] = in1[29] ^ in2[29];
    assign G[82] = in1[28] & in2[28];
    assign P[82] = in1[28] ^ in2[28];
    assign G[83] = in1[27] & in2[27];
    assign P[83] = in1[27] ^ in2[27];
    assign G[84] = in1[26] & in2[26];
    assign P[84] = in1[26] ^ in2[26];
    assign G[85] = in1[25] & in2[25];
    assign P[85] = in1[25] ^ in2[25];
    assign G[86] = in1[24] & in2[24];
    assign P[86] = in1[24] ^ in2[24];
    assign G[87] = in1[23] & in2[23];
    assign P[87] = in1[23] ^ in2[23];
    assign G[88] = in1[22] & in2[22];
    assign P[88] = in1[22] ^ in2[22];
    assign G[89] = in1[21] & in2[21];
    assign P[89] = in1[21] ^ in2[21];
    assign G[90] = in1[20] & in2[20];
    assign P[90] = in1[20] ^ in2[20];
    assign G[91] = in1[19] & in2[19];
    assign P[91] = in1[19] ^ in2[19];
    assign G[92] = in1[18] & in2[18];
    assign P[92] = in1[18] ^ in2[18];
    assign G[93] = in1[17] & in2[17];
    assign P[93] = in1[17] ^ in2[17];
    assign G[94] = in1[16] & in2[16];
    assign P[94] = in1[16] ^ in2[16];
    assign G[95] = in1[15] & in2[15];
    assign P[95] = in1[15] ^ in2[15];
    assign G[96] = in1[14] & in2[14];
    assign P[96] = in1[14] ^ in2[14];
    assign G[97] = in1[13] & in2[13];
    assign P[97] = in1[13] ^ in2[13];
    assign G[98] = in1[12] & in2[12];
    assign P[98] = in1[12] ^ in2[12];
    assign G[99] = in1[11] & in2[11];
    assign P[99] = in1[11] ^ in2[11];
    assign G[100] = in1[10] & in2[10];
    assign P[100] = in1[10] ^ in2[10];
    assign G[101] = in1[9] & in2[9];
    assign P[101] = in1[9] ^ in2[9];
    assign G[102] = in1[8] & in2[8];
    assign P[102] = in1[8] ^ in2[8];
    assign G[103] = in1[7] & in2[7];
    assign P[103] = in1[7] ^ in2[7];
    assign G[104] = in1[6] & in2[6];
    assign P[104] = in1[6] ^ in2[6];
    assign G[105] = in1[5] & in2[5];
    assign P[105] = in1[5] ^ in2[5];
    assign G[106] = in1[4] & in2[4];
    assign P[106] = in1[4] ^ in2[4];
    assign G[107] = in1[3] & in2[3];
    assign P[107] = in1[3] ^ in2[3];
    assign G[108] = in1[2] & in2[2];
    assign P[108] = in1[2] ^ in2[2];
    assign G[109] = in1[1] & in2[1];
    assign P[109] = in1[1] ^ in2[1];
    assign G[110] = in1[0] & in2[0];
    assign P[110] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign cout = G[110] | (P[110] & C[110]);
    assign sum = P ^ C;
endmodule

module CLA_110(output [109:0] sum, output cout, input [109:0] in1, input [109:0] in2);

    wire[109:0] G;
    wire[109:0] C;
    wire[109:0] P;

    assign G[0] = in1[109] & in2[109];
    assign P[0] = in1[109] ^ in2[109];
    assign G[1] = in1[108] & in2[108];
    assign P[1] = in1[108] ^ in2[108];
    assign G[2] = in1[107] & in2[107];
    assign P[2] = in1[107] ^ in2[107];
    assign G[3] = in1[106] & in2[106];
    assign P[3] = in1[106] ^ in2[106];
    assign G[4] = in1[105] & in2[105];
    assign P[4] = in1[105] ^ in2[105];
    assign G[5] = in1[104] & in2[104];
    assign P[5] = in1[104] ^ in2[104];
    assign G[6] = in1[103] & in2[103];
    assign P[6] = in1[103] ^ in2[103];
    assign G[7] = in1[102] & in2[102];
    assign P[7] = in1[102] ^ in2[102];
    assign G[8] = in1[101] & in2[101];
    assign P[8] = in1[101] ^ in2[101];
    assign G[9] = in1[100] & in2[100];
    assign P[9] = in1[100] ^ in2[100];
    assign G[10] = in1[99] & in2[99];
    assign P[10] = in1[99] ^ in2[99];
    assign G[11] = in1[98] & in2[98];
    assign P[11] = in1[98] ^ in2[98];
    assign G[12] = in1[97] & in2[97];
    assign P[12] = in1[97] ^ in2[97];
    assign G[13] = in1[96] & in2[96];
    assign P[13] = in1[96] ^ in2[96];
    assign G[14] = in1[95] & in2[95];
    assign P[14] = in1[95] ^ in2[95];
    assign G[15] = in1[94] & in2[94];
    assign P[15] = in1[94] ^ in2[94];
    assign G[16] = in1[93] & in2[93];
    assign P[16] = in1[93] ^ in2[93];
    assign G[17] = in1[92] & in2[92];
    assign P[17] = in1[92] ^ in2[92];
    assign G[18] = in1[91] & in2[91];
    assign P[18] = in1[91] ^ in2[91];
    assign G[19] = in1[90] & in2[90];
    assign P[19] = in1[90] ^ in2[90];
    assign G[20] = in1[89] & in2[89];
    assign P[20] = in1[89] ^ in2[89];
    assign G[21] = in1[88] & in2[88];
    assign P[21] = in1[88] ^ in2[88];
    assign G[22] = in1[87] & in2[87];
    assign P[22] = in1[87] ^ in2[87];
    assign G[23] = in1[86] & in2[86];
    assign P[23] = in1[86] ^ in2[86];
    assign G[24] = in1[85] & in2[85];
    assign P[24] = in1[85] ^ in2[85];
    assign G[25] = in1[84] & in2[84];
    assign P[25] = in1[84] ^ in2[84];
    assign G[26] = in1[83] & in2[83];
    assign P[26] = in1[83] ^ in2[83];
    assign G[27] = in1[82] & in2[82];
    assign P[27] = in1[82] ^ in2[82];
    assign G[28] = in1[81] & in2[81];
    assign P[28] = in1[81] ^ in2[81];
    assign G[29] = in1[80] & in2[80];
    assign P[29] = in1[80] ^ in2[80];
    assign G[30] = in1[79] & in2[79];
    assign P[30] = in1[79] ^ in2[79];
    assign G[31] = in1[78] & in2[78];
    assign P[31] = in1[78] ^ in2[78];
    assign G[32] = in1[77] & in2[77];
    assign P[32] = in1[77] ^ in2[77];
    assign G[33] = in1[76] & in2[76];
    assign P[33] = in1[76] ^ in2[76];
    assign G[34] = in1[75] & in2[75];
    assign P[34] = in1[75] ^ in2[75];
    assign G[35] = in1[74] & in2[74];
    assign P[35] = in1[74] ^ in2[74];
    assign G[36] = in1[73] & in2[73];
    assign P[36] = in1[73] ^ in2[73];
    assign G[37] = in1[72] & in2[72];
    assign P[37] = in1[72] ^ in2[72];
    assign G[38] = in1[71] & in2[71];
    assign P[38] = in1[71] ^ in2[71];
    assign G[39] = in1[70] & in2[70];
    assign P[39] = in1[70] ^ in2[70];
    assign G[40] = in1[69] & in2[69];
    assign P[40] = in1[69] ^ in2[69];
    assign G[41] = in1[68] & in2[68];
    assign P[41] = in1[68] ^ in2[68];
    assign G[42] = in1[67] & in2[67];
    assign P[42] = in1[67] ^ in2[67];
    assign G[43] = in1[66] & in2[66];
    assign P[43] = in1[66] ^ in2[66];
    assign G[44] = in1[65] & in2[65];
    assign P[44] = in1[65] ^ in2[65];
    assign G[45] = in1[64] & in2[64];
    assign P[45] = in1[64] ^ in2[64];
    assign G[46] = in1[63] & in2[63];
    assign P[46] = in1[63] ^ in2[63];
    assign G[47] = in1[62] & in2[62];
    assign P[47] = in1[62] ^ in2[62];
    assign G[48] = in1[61] & in2[61];
    assign P[48] = in1[61] ^ in2[61];
    assign G[49] = in1[60] & in2[60];
    assign P[49] = in1[60] ^ in2[60];
    assign G[50] = in1[59] & in2[59];
    assign P[50] = in1[59] ^ in2[59];
    assign G[51] = in1[58] & in2[58];
    assign P[51] = in1[58] ^ in2[58];
    assign G[52] = in1[57] & in2[57];
    assign P[52] = in1[57] ^ in2[57];
    assign G[53] = in1[56] & in2[56];
    assign P[53] = in1[56] ^ in2[56];
    assign G[54] = in1[55] & in2[55];
    assign P[54] = in1[55] ^ in2[55];
    assign G[55] = in1[54] & in2[54];
    assign P[55] = in1[54] ^ in2[54];
    assign G[56] = in1[53] & in2[53];
    assign P[56] = in1[53] ^ in2[53];
    assign G[57] = in1[52] & in2[52];
    assign P[57] = in1[52] ^ in2[52];
    assign G[58] = in1[51] & in2[51];
    assign P[58] = in1[51] ^ in2[51];
    assign G[59] = in1[50] & in2[50];
    assign P[59] = in1[50] ^ in2[50];
    assign G[60] = in1[49] & in2[49];
    assign P[60] = in1[49] ^ in2[49];
    assign G[61] = in1[48] & in2[48];
    assign P[61] = in1[48] ^ in2[48];
    assign G[62] = in1[47] & in2[47];
    assign P[62] = in1[47] ^ in2[47];
    assign G[63] = in1[46] & in2[46];
    assign P[63] = in1[46] ^ in2[46];
    assign G[64] = in1[45] & in2[45];
    assign P[64] = in1[45] ^ in2[45];
    assign G[65] = in1[44] & in2[44];
    assign P[65] = in1[44] ^ in2[44];
    assign G[66] = in1[43] & in2[43];
    assign P[66] = in1[43] ^ in2[43];
    assign G[67] = in1[42] & in2[42];
    assign P[67] = in1[42] ^ in2[42];
    assign G[68] = in1[41] & in2[41];
    assign P[68] = in1[41] ^ in2[41];
    assign G[69] = in1[40] & in2[40];
    assign P[69] = in1[40] ^ in2[40];
    assign G[70] = in1[39] & in2[39];
    assign P[70] = in1[39] ^ in2[39];
    assign G[71] = in1[38] & in2[38];
    assign P[71] = in1[38] ^ in2[38];
    assign G[72] = in1[37] & in2[37];
    assign P[72] = in1[37] ^ in2[37];
    assign G[73] = in1[36] & in2[36];
    assign P[73] = in1[36] ^ in2[36];
    assign G[74] = in1[35] & in2[35];
    assign P[74] = in1[35] ^ in2[35];
    assign G[75] = in1[34] & in2[34];
    assign P[75] = in1[34] ^ in2[34];
    assign G[76] = in1[33] & in2[33];
    assign P[76] = in1[33] ^ in2[33];
    assign G[77] = in1[32] & in2[32];
    assign P[77] = in1[32] ^ in2[32];
    assign G[78] = in1[31] & in2[31];
    assign P[78] = in1[31] ^ in2[31];
    assign G[79] = in1[30] & in2[30];
    assign P[79] = in1[30] ^ in2[30];
    assign G[80] = in1[29] & in2[29];
    assign P[80] = in1[29] ^ in2[29];
    assign G[81] = in1[28] & in2[28];
    assign P[81] = in1[28] ^ in2[28];
    assign G[82] = in1[27] & in2[27];
    assign P[82] = in1[27] ^ in2[27];
    assign G[83] = in1[26] & in2[26];
    assign P[83] = in1[26] ^ in2[26];
    assign G[84] = in1[25] & in2[25];
    assign P[84] = in1[25] ^ in2[25];
    assign G[85] = in1[24] & in2[24];
    assign P[85] = in1[24] ^ in2[24];
    assign G[86] = in1[23] & in2[23];
    assign P[86] = in1[23] ^ in2[23];
    assign G[87] = in1[22] & in2[22];
    assign P[87] = in1[22] ^ in2[22];
    assign G[88] = in1[21] & in2[21];
    assign P[88] = in1[21] ^ in2[21];
    assign G[89] = in1[20] & in2[20];
    assign P[89] = in1[20] ^ in2[20];
    assign G[90] = in1[19] & in2[19];
    assign P[90] = in1[19] ^ in2[19];
    assign G[91] = in1[18] & in2[18];
    assign P[91] = in1[18] ^ in2[18];
    assign G[92] = in1[17] & in2[17];
    assign P[92] = in1[17] ^ in2[17];
    assign G[93] = in1[16] & in2[16];
    assign P[93] = in1[16] ^ in2[16];
    assign G[94] = in1[15] & in2[15];
    assign P[94] = in1[15] ^ in2[15];
    assign G[95] = in1[14] & in2[14];
    assign P[95] = in1[14] ^ in2[14];
    assign G[96] = in1[13] & in2[13];
    assign P[96] = in1[13] ^ in2[13];
    assign G[97] = in1[12] & in2[12];
    assign P[97] = in1[12] ^ in2[12];
    assign G[98] = in1[11] & in2[11];
    assign P[98] = in1[11] ^ in2[11];
    assign G[99] = in1[10] & in2[10];
    assign P[99] = in1[10] ^ in2[10];
    assign G[100] = in1[9] & in2[9];
    assign P[100] = in1[9] ^ in2[9];
    assign G[101] = in1[8] & in2[8];
    assign P[101] = in1[8] ^ in2[8];
    assign G[102] = in1[7] & in2[7];
    assign P[102] = in1[7] ^ in2[7];
    assign G[103] = in1[6] & in2[6];
    assign P[103] = in1[6] ^ in2[6];
    assign G[104] = in1[5] & in2[5];
    assign P[104] = in1[5] ^ in2[5];
    assign G[105] = in1[4] & in2[4];
    assign P[105] = in1[4] ^ in2[4];
    assign G[106] = in1[3] & in2[3];
    assign P[106] = in1[3] ^ in2[3];
    assign G[107] = in1[2] & in2[2];
    assign P[107] = in1[2] ^ in2[2];
    assign G[108] = in1[1] & in2[1];
    assign P[108] = in1[1] ^ in2[1];
    assign G[109] = in1[0] & in2[0];
    assign P[109] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign cout = G[109] | (P[109] & C[109]);
    assign sum = P ^ C;
endmodule

module CLA_109(output [108:0] sum, output cout, input [108:0] in1, input [108:0] in2);

    wire[108:0] G;
    wire[108:0] C;
    wire[108:0] P;

    assign G[0] = in1[108] & in2[108];
    assign P[0] = in1[108] ^ in2[108];
    assign G[1] = in1[107] & in2[107];
    assign P[1] = in1[107] ^ in2[107];
    assign G[2] = in1[106] & in2[106];
    assign P[2] = in1[106] ^ in2[106];
    assign G[3] = in1[105] & in2[105];
    assign P[3] = in1[105] ^ in2[105];
    assign G[4] = in1[104] & in2[104];
    assign P[4] = in1[104] ^ in2[104];
    assign G[5] = in1[103] & in2[103];
    assign P[5] = in1[103] ^ in2[103];
    assign G[6] = in1[102] & in2[102];
    assign P[6] = in1[102] ^ in2[102];
    assign G[7] = in1[101] & in2[101];
    assign P[7] = in1[101] ^ in2[101];
    assign G[8] = in1[100] & in2[100];
    assign P[8] = in1[100] ^ in2[100];
    assign G[9] = in1[99] & in2[99];
    assign P[9] = in1[99] ^ in2[99];
    assign G[10] = in1[98] & in2[98];
    assign P[10] = in1[98] ^ in2[98];
    assign G[11] = in1[97] & in2[97];
    assign P[11] = in1[97] ^ in2[97];
    assign G[12] = in1[96] & in2[96];
    assign P[12] = in1[96] ^ in2[96];
    assign G[13] = in1[95] & in2[95];
    assign P[13] = in1[95] ^ in2[95];
    assign G[14] = in1[94] & in2[94];
    assign P[14] = in1[94] ^ in2[94];
    assign G[15] = in1[93] & in2[93];
    assign P[15] = in1[93] ^ in2[93];
    assign G[16] = in1[92] & in2[92];
    assign P[16] = in1[92] ^ in2[92];
    assign G[17] = in1[91] & in2[91];
    assign P[17] = in1[91] ^ in2[91];
    assign G[18] = in1[90] & in2[90];
    assign P[18] = in1[90] ^ in2[90];
    assign G[19] = in1[89] & in2[89];
    assign P[19] = in1[89] ^ in2[89];
    assign G[20] = in1[88] & in2[88];
    assign P[20] = in1[88] ^ in2[88];
    assign G[21] = in1[87] & in2[87];
    assign P[21] = in1[87] ^ in2[87];
    assign G[22] = in1[86] & in2[86];
    assign P[22] = in1[86] ^ in2[86];
    assign G[23] = in1[85] & in2[85];
    assign P[23] = in1[85] ^ in2[85];
    assign G[24] = in1[84] & in2[84];
    assign P[24] = in1[84] ^ in2[84];
    assign G[25] = in1[83] & in2[83];
    assign P[25] = in1[83] ^ in2[83];
    assign G[26] = in1[82] & in2[82];
    assign P[26] = in1[82] ^ in2[82];
    assign G[27] = in1[81] & in2[81];
    assign P[27] = in1[81] ^ in2[81];
    assign G[28] = in1[80] & in2[80];
    assign P[28] = in1[80] ^ in2[80];
    assign G[29] = in1[79] & in2[79];
    assign P[29] = in1[79] ^ in2[79];
    assign G[30] = in1[78] & in2[78];
    assign P[30] = in1[78] ^ in2[78];
    assign G[31] = in1[77] & in2[77];
    assign P[31] = in1[77] ^ in2[77];
    assign G[32] = in1[76] & in2[76];
    assign P[32] = in1[76] ^ in2[76];
    assign G[33] = in1[75] & in2[75];
    assign P[33] = in1[75] ^ in2[75];
    assign G[34] = in1[74] & in2[74];
    assign P[34] = in1[74] ^ in2[74];
    assign G[35] = in1[73] & in2[73];
    assign P[35] = in1[73] ^ in2[73];
    assign G[36] = in1[72] & in2[72];
    assign P[36] = in1[72] ^ in2[72];
    assign G[37] = in1[71] & in2[71];
    assign P[37] = in1[71] ^ in2[71];
    assign G[38] = in1[70] & in2[70];
    assign P[38] = in1[70] ^ in2[70];
    assign G[39] = in1[69] & in2[69];
    assign P[39] = in1[69] ^ in2[69];
    assign G[40] = in1[68] & in2[68];
    assign P[40] = in1[68] ^ in2[68];
    assign G[41] = in1[67] & in2[67];
    assign P[41] = in1[67] ^ in2[67];
    assign G[42] = in1[66] & in2[66];
    assign P[42] = in1[66] ^ in2[66];
    assign G[43] = in1[65] & in2[65];
    assign P[43] = in1[65] ^ in2[65];
    assign G[44] = in1[64] & in2[64];
    assign P[44] = in1[64] ^ in2[64];
    assign G[45] = in1[63] & in2[63];
    assign P[45] = in1[63] ^ in2[63];
    assign G[46] = in1[62] & in2[62];
    assign P[46] = in1[62] ^ in2[62];
    assign G[47] = in1[61] & in2[61];
    assign P[47] = in1[61] ^ in2[61];
    assign G[48] = in1[60] & in2[60];
    assign P[48] = in1[60] ^ in2[60];
    assign G[49] = in1[59] & in2[59];
    assign P[49] = in1[59] ^ in2[59];
    assign G[50] = in1[58] & in2[58];
    assign P[50] = in1[58] ^ in2[58];
    assign G[51] = in1[57] & in2[57];
    assign P[51] = in1[57] ^ in2[57];
    assign G[52] = in1[56] & in2[56];
    assign P[52] = in1[56] ^ in2[56];
    assign G[53] = in1[55] & in2[55];
    assign P[53] = in1[55] ^ in2[55];
    assign G[54] = in1[54] & in2[54];
    assign P[54] = in1[54] ^ in2[54];
    assign G[55] = in1[53] & in2[53];
    assign P[55] = in1[53] ^ in2[53];
    assign G[56] = in1[52] & in2[52];
    assign P[56] = in1[52] ^ in2[52];
    assign G[57] = in1[51] & in2[51];
    assign P[57] = in1[51] ^ in2[51];
    assign G[58] = in1[50] & in2[50];
    assign P[58] = in1[50] ^ in2[50];
    assign G[59] = in1[49] & in2[49];
    assign P[59] = in1[49] ^ in2[49];
    assign G[60] = in1[48] & in2[48];
    assign P[60] = in1[48] ^ in2[48];
    assign G[61] = in1[47] & in2[47];
    assign P[61] = in1[47] ^ in2[47];
    assign G[62] = in1[46] & in2[46];
    assign P[62] = in1[46] ^ in2[46];
    assign G[63] = in1[45] & in2[45];
    assign P[63] = in1[45] ^ in2[45];
    assign G[64] = in1[44] & in2[44];
    assign P[64] = in1[44] ^ in2[44];
    assign G[65] = in1[43] & in2[43];
    assign P[65] = in1[43] ^ in2[43];
    assign G[66] = in1[42] & in2[42];
    assign P[66] = in1[42] ^ in2[42];
    assign G[67] = in1[41] & in2[41];
    assign P[67] = in1[41] ^ in2[41];
    assign G[68] = in1[40] & in2[40];
    assign P[68] = in1[40] ^ in2[40];
    assign G[69] = in1[39] & in2[39];
    assign P[69] = in1[39] ^ in2[39];
    assign G[70] = in1[38] & in2[38];
    assign P[70] = in1[38] ^ in2[38];
    assign G[71] = in1[37] & in2[37];
    assign P[71] = in1[37] ^ in2[37];
    assign G[72] = in1[36] & in2[36];
    assign P[72] = in1[36] ^ in2[36];
    assign G[73] = in1[35] & in2[35];
    assign P[73] = in1[35] ^ in2[35];
    assign G[74] = in1[34] & in2[34];
    assign P[74] = in1[34] ^ in2[34];
    assign G[75] = in1[33] & in2[33];
    assign P[75] = in1[33] ^ in2[33];
    assign G[76] = in1[32] & in2[32];
    assign P[76] = in1[32] ^ in2[32];
    assign G[77] = in1[31] & in2[31];
    assign P[77] = in1[31] ^ in2[31];
    assign G[78] = in1[30] & in2[30];
    assign P[78] = in1[30] ^ in2[30];
    assign G[79] = in1[29] & in2[29];
    assign P[79] = in1[29] ^ in2[29];
    assign G[80] = in1[28] & in2[28];
    assign P[80] = in1[28] ^ in2[28];
    assign G[81] = in1[27] & in2[27];
    assign P[81] = in1[27] ^ in2[27];
    assign G[82] = in1[26] & in2[26];
    assign P[82] = in1[26] ^ in2[26];
    assign G[83] = in1[25] & in2[25];
    assign P[83] = in1[25] ^ in2[25];
    assign G[84] = in1[24] & in2[24];
    assign P[84] = in1[24] ^ in2[24];
    assign G[85] = in1[23] & in2[23];
    assign P[85] = in1[23] ^ in2[23];
    assign G[86] = in1[22] & in2[22];
    assign P[86] = in1[22] ^ in2[22];
    assign G[87] = in1[21] & in2[21];
    assign P[87] = in1[21] ^ in2[21];
    assign G[88] = in1[20] & in2[20];
    assign P[88] = in1[20] ^ in2[20];
    assign G[89] = in1[19] & in2[19];
    assign P[89] = in1[19] ^ in2[19];
    assign G[90] = in1[18] & in2[18];
    assign P[90] = in1[18] ^ in2[18];
    assign G[91] = in1[17] & in2[17];
    assign P[91] = in1[17] ^ in2[17];
    assign G[92] = in1[16] & in2[16];
    assign P[92] = in1[16] ^ in2[16];
    assign G[93] = in1[15] & in2[15];
    assign P[93] = in1[15] ^ in2[15];
    assign G[94] = in1[14] & in2[14];
    assign P[94] = in1[14] ^ in2[14];
    assign G[95] = in1[13] & in2[13];
    assign P[95] = in1[13] ^ in2[13];
    assign G[96] = in1[12] & in2[12];
    assign P[96] = in1[12] ^ in2[12];
    assign G[97] = in1[11] & in2[11];
    assign P[97] = in1[11] ^ in2[11];
    assign G[98] = in1[10] & in2[10];
    assign P[98] = in1[10] ^ in2[10];
    assign G[99] = in1[9] & in2[9];
    assign P[99] = in1[9] ^ in2[9];
    assign G[100] = in1[8] & in2[8];
    assign P[100] = in1[8] ^ in2[8];
    assign G[101] = in1[7] & in2[7];
    assign P[101] = in1[7] ^ in2[7];
    assign G[102] = in1[6] & in2[6];
    assign P[102] = in1[6] ^ in2[6];
    assign G[103] = in1[5] & in2[5];
    assign P[103] = in1[5] ^ in2[5];
    assign G[104] = in1[4] & in2[4];
    assign P[104] = in1[4] ^ in2[4];
    assign G[105] = in1[3] & in2[3];
    assign P[105] = in1[3] ^ in2[3];
    assign G[106] = in1[2] & in2[2];
    assign P[106] = in1[2] ^ in2[2];
    assign G[107] = in1[1] & in2[1];
    assign P[107] = in1[1] ^ in2[1];
    assign G[108] = in1[0] & in2[0];
    assign P[108] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign cout = G[108] | (P[108] & C[108]);
    assign sum = P ^ C;
endmodule

module CLA_108(output [107:0] sum, output cout, input [107:0] in1, input [107:0] in2);

    wire[107:0] G;
    wire[107:0] C;
    wire[107:0] P;

    assign G[0] = in1[107] & in2[107];
    assign P[0] = in1[107] ^ in2[107];
    assign G[1] = in1[106] & in2[106];
    assign P[1] = in1[106] ^ in2[106];
    assign G[2] = in1[105] & in2[105];
    assign P[2] = in1[105] ^ in2[105];
    assign G[3] = in1[104] & in2[104];
    assign P[3] = in1[104] ^ in2[104];
    assign G[4] = in1[103] & in2[103];
    assign P[4] = in1[103] ^ in2[103];
    assign G[5] = in1[102] & in2[102];
    assign P[5] = in1[102] ^ in2[102];
    assign G[6] = in1[101] & in2[101];
    assign P[6] = in1[101] ^ in2[101];
    assign G[7] = in1[100] & in2[100];
    assign P[7] = in1[100] ^ in2[100];
    assign G[8] = in1[99] & in2[99];
    assign P[8] = in1[99] ^ in2[99];
    assign G[9] = in1[98] & in2[98];
    assign P[9] = in1[98] ^ in2[98];
    assign G[10] = in1[97] & in2[97];
    assign P[10] = in1[97] ^ in2[97];
    assign G[11] = in1[96] & in2[96];
    assign P[11] = in1[96] ^ in2[96];
    assign G[12] = in1[95] & in2[95];
    assign P[12] = in1[95] ^ in2[95];
    assign G[13] = in1[94] & in2[94];
    assign P[13] = in1[94] ^ in2[94];
    assign G[14] = in1[93] & in2[93];
    assign P[14] = in1[93] ^ in2[93];
    assign G[15] = in1[92] & in2[92];
    assign P[15] = in1[92] ^ in2[92];
    assign G[16] = in1[91] & in2[91];
    assign P[16] = in1[91] ^ in2[91];
    assign G[17] = in1[90] & in2[90];
    assign P[17] = in1[90] ^ in2[90];
    assign G[18] = in1[89] & in2[89];
    assign P[18] = in1[89] ^ in2[89];
    assign G[19] = in1[88] & in2[88];
    assign P[19] = in1[88] ^ in2[88];
    assign G[20] = in1[87] & in2[87];
    assign P[20] = in1[87] ^ in2[87];
    assign G[21] = in1[86] & in2[86];
    assign P[21] = in1[86] ^ in2[86];
    assign G[22] = in1[85] & in2[85];
    assign P[22] = in1[85] ^ in2[85];
    assign G[23] = in1[84] & in2[84];
    assign P[23] = in1[84] ^ in2[84];
    assign G[24] = in1[83] & in2[83];
    assign P[24] = in1[83] ^ in2[83];
    assign G[25] = in1[82] & in2[82];
    assign P[25] = in1[82] ^ in2[82];
    assign G[26] = in1[81] & in2[81];
    assign P[26] = in1[81] ^ in2[81];
    assign G[27] = in1[80] & in2[80];
    assign P[27] = in1[80] ^ in2[80];
    assign G[28] = in1[79] & in2[79];
    assign P[28] = in1[79] ^ in2[79];
    assign G[29] = in1[78] & in2[78];
    assign P[29] = in1[78] ^ in2[78];
    assign G[30] = in1[77] & in2[77];
    assign P[30] = in1[77] ^ in2[77];
    assign G[31] = in1[76] & in2[76];
    assign P[31] = in1[76] ^ in2[76];
    assign G[32] = in1[75] & in2[75];
    assign P[32] = in1[75] ^ in2[75];
    assign G[33] = in1[74] & in2[74];
    assign P[33] = in1[74] ^ in2[74];
    assign G[34] = in1[73] & in2[73];
    assign P[34] = in1[73] ^ in2[73];
    assign G[35] = in1[72] & in2[72];
    assign P[35] = in1[72] ^ in2[72];
    assign G[36] = in1[71] & in2[71];
    assign P[36] = in1[71] ^ in2[71];
    assign G[37] = in1[70] & in2[70];
    assign P[37] = in1[70] ^ in2[70];
    assign G[38] = in1[69] & in2[69];
    assign P[38] = in1[69] ^ in2[69];
    assign G[39] = in1[68] & in2[68];
    assign P[39] = in1[68] ^ in2[68];
    assign G[40] = in1[67] & in2[67];
    assign P[40] = in1[67] ^ in2[67];
    assign G[41] = in1[66] & in2[66];
    assign P[41] = in1[66] ^ in2[66];
    assign G[42] = in1[65] & in2[65];
    assign P[42] = in1[65] ^ in2[65];
    assign G[43] = in1[64] & in2[64];
    assign P[43] = in1[64] ^ in2[64];
    assign G[44] = in1[63] & in2[63];
    assign P[44] = in1[63] ^ in2[63];
    assign G[45] = in1[62] & in2[62];
    assign P[45] = in1[62] ^ in2[62];
    assign G[46] = in1[61] & in2[61];
    assign P[46] = in1[61] ^ in2[61];
    assign G[47] = in1[60] & in2[60];
    assign P[47] = in1[60] ^ in2[60];
    assign G[48] = in1[59] & in2[59];
    assign P[48] = in1[59] ^ in2[59];
    assign G[49] = in1[58] & in2[58];
    assign P[49] = in1[58] ^ in2[58];
    assign G[50] = in1[57] & in2[57];
    assign P[50] = in1[57] ^ in2[57];
    assign G[51] = in1[56] & in2[56];
    assign P[51] = in1[56] ^ in2[56];
    assign G[52] = in1[55] & in2[55];
    assign P[52] = in1[55] ^ in2[55];
    assign G[53] = in1[54] & in2[54];
    assign P[53] = in1[54] ^ in2[54];
    assign G[54] = in1[53] & in2[53];
    assign P[54] = in1[53] ^ in2[53];
    assign G[55] = in1[52] & in2[52];
    assign P[55] = in1[52] ^ in2[52];
    assign G[56] = in1[51] & in2[51];
    assign P[56] = in1[51] ^ in2[51];
    assign G[57] = in1[50] & in2[50];
    assign P[57] = in1[50] ^ in2[50];
    assign G[58] = in1[49] & in2[49];
    assign P[58] = in1[49] ^ in2[49];
    assign G[59] = in1[48] & in2[48];
    assign P[59] = in1[48] ^ in2[48];
    assign G[60] = in1[47] & in2[47];
    assign P[60] = in1[47] ^ in2[47];
    assign G[61] = in1[46] & in2[46];
    assign P[61] = in1[46] ^ in2[46];
    assign G[62] = in1[45] & in2[45];
    assign P[62] = in1[45] ^ in2[45];
    assign G[63] = in1[44] & in2[44];
    assign P[63] = in1[44] ^ in2[44];
    assign G[64] = in1[43] & in2[43];
    assign P[64] = in1[43] ^ in2[43];
    assign G[65] = in1[42] & in2[42];
    assign P[65] = in1[42] ^ in2[42];
    assign G[66] = in1[41] & in2[41];
    assign P[66] = in1[41] ^ in2[41];
    assign G[67] = in1[40] & in2[40];
    assign P[67] = in1[40] ^ in2[40];
    assign G[68] = in1[39] & in2[39];
    assign P[68] = in1[39] ^ in2[39];
    assign G[69] = in1[38] & in2[38];
    assign P[69] = in1[38] ^ in2[38];
    assign G[70] = in1[37] & in2[37];
    assign P[70] = in1[37] ^ in2[37];
    assign G[71] = in1[36] & in2[36];
    assign P[71] = in1[36] ^ in2[36];
    assign G[72] = in1[35] & in2[35];
    assign P[72] = in1[35] ^ in2[35];
    assign G[73] = in1[34] & in2[34];
    assign P[73] = in1[34] ^ in2[34];
    assign G[74] = in1[33] & in2[33];
    assign P[74] = in1[33] ^ in2[33];
    assign G[75] = in1[32] & in2[32];
    assign P[75] = in1[32] ^ in2[32];
    assign G[76] = in1[31] & in2[31];
    assign P[76] = in1[31] ^ in2[31];
    assign G[77] = in1[30] & in2[30];
    assign P[77] = in1[30] ^ in2[30];
    assign G[78] = in1[29] & in2[29];
    assign P[78] = in1[29] ^ in2[29];
    assign G[79] = in1[28] & in2[28];
    assign P[79] = in1[28] ^ in2[28];
    assign G[80] = in1[27] & in2[27];
    assign P[80] = in1[27] ^ in2[27];
    assign G[81] = in1[26] & in2[26];
    assign P[81] = in1[26] ^ in2[26];
    assign G[82] = in1[25] & in2[25];
    assign P[82] = in1[25] ^ in2[25];
    assign G[83] = in1[24] & in2[24];
    assign P[83] = in1[24] ^ in2[24];
    assign G[84] = in1[23] & in2[23];
    assign P[84] = in1[23] ^ in2[23];
    assign G[85] = in1[22] & in2[22];
    assign P[85] = in1[22] ^ in2[22];
    assign G[86] = in1[21] & in2[21];
    assign P[86] = in1[21] ^ in2[21];
    assign G[87] = in1[20] & in2[20];
    assign P[87] = in1[20] ^ in2[20];
    assign G[88] = in1[19] & in2[19];
    assign P[88] = in1[19] ^ in2[19];
    assign G[89] = in1[18] & in2[18];
    assign P[89] = in1[18] ^ in2[18];
    assign G[90] = in1[17] & in2[17];
    assign P[90] = in1[17] ^ in2[17];
    assign G[91] = in1[16] & in2[16];
    assign P[91] = in1[16] ^ in2[16];
    assign G[92] = in1[15] & in2[15];
    assign P[92] = in1[15] ^ in2[15];
    assign G[93] = in1[14] & in2[14];
    assign P[93] = in1[14] ^ in2[14];
    assign G[94] = in1[13] & in2[13];
    assign P[94] = in1[13] ^ in2[13];
    assign G[95] = in1[12] & in2[12];
    assign P[95] = in1[12] ^ in2[12];
    assign G[96] = in1[11] & in2[11];
    assign P[96] = in1[11] ^ in2[11];
    assign G[97] = in1[10] & in2[10];
    assign P[97] = in1[10] ^ in2[10];
    assign G[98] = in1[9] & in2[9];
    assign P[98] = in1[9] ^ in2[9];
    assign G[99] = in1[8] & in2[8];
    assign P[99] = in1[8] ^ in2[8];
    assign G[100] = in1[7] & in2[7];
    assign P[100] = in1[7] ^ in2[7];
    assign G[101] = in1[6] & in2[6];
    assign P[101] = in1[6] ^ in2[6];
    assign G[102] = in1[5] & in2[5];
    assign P[102] = in1[5] ^ in2[5];
    assign G[103] = in1[4] & in2[4];
    assign P[103] = in1[4] ^ in2[4];
    assign G[104] = in1[3] & in2[3];
    assign P[104] = in1[3] ^ in2[3];
    assign G[105] = in1[2] & in2[2];
    assign P[105] = in1[2] ^ in2[2];
    assign G[106] = in1[1] & in2[1];
    assign P[106] = in1[1] ^ in2[1];
    assign G[107] = in1[0] & in2[0];
    assign P[107] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign cout = G[107] | (P[107] & C[107]);
    assign sum = P ^ C;
endmodule

module CLA_107(output [106:0] sum, output cout, input [106:0] in1, input [106:0] in2);

    wire[106:0] G;
    wire[106:0] C;
    wire[106:0] P;

    assign G[0] = in1[106] & in2[106];
    assign P[0] = in1[106] ^ in2[106];
    assign G[1] = in1[105] & in2[105];
    assign P[1] = in1[105] ^ in2[105];
    assign G[2] = in1[104] & in2[104];
    assign P[2] = in1[104] ^ in2[104];
    assign G[3] = in1[103] & in2[103];
    assign P[3] = in1[103] ^ in2[103];
    assign G[4] = in1[102] & in2[102];
    assign P[4] = in1[102] ^ in2[102];
    assign G[5] = in1[101] & in2[101];
    assign P[5] = in1[101] ^ in2[101];
    assign G[6] = in1[100] & in2[100];
    assign P[6] = in1[100] ^ in2[100];
    assign G[7] = in1[99] & in2[99];
    assign P[7] = in1[99] ^ in2[99];
    assign G[8] = in1[98] & in2[98];
    assign P[8] = in1[98] ^ in2[98];
    assign G[9] = in1[97] & in2[97];
    assign P[9] = in1[97] ^ in2[97];
    assign G[10] = in1[96] & in2[96];
    assign P[10] = in1[96] ^ in2[96];
    assign G[11] = in1[95] & in2[95];
    assign P[11] = in1[95] ^ in2[95];
    assign G[12] = in1[94] & in2[94];
    assign P[12] = in1[94] ^ in2[94];
    assign G[13] = in1[93] & in2[93];
    assign P[13] = in1[93] ^ in2[93];
    assign G[14] = in1[92] & in2[92];
    assign P[14] = in1[92] ^ in2[92];
    assign G[15] = in1[91] & in2[91];
    assign P[15] = in1[91] ^ in2[91];
    assign G[16] = in1[90] & in2[90];
    assign P[16] = in1[90] ^ in2[90];
    assign G[17] = in1[89] & in2[89];
    assign P[17] = in1[89] ^ in2[89];
    assign G[18] = in1[88] & in2[88];
    assign P[18] = in1[88] ^ in2[88];
    assign G[19] = in1[87] & in2[87];
    assign P[19] = in1[87] ^ in2[87];
    assign G[20] = in1[86] & in2[86];
    assign P[20] = in1[86] ^ in2[86];
    assign G[21] = in1[85] & in2[85];
    assign P[21] = in1[85] ^ in2[85];
    assign G[22] = in1[84] & in2[84];
    assign P[22] = in1[84] ^ in2[84];
    assign G[23] = in1[83] & in2[83];
    assign P[23] = in1[83] ^ in2[83];
    assign G[24] = in1[82] & in2[82];
    assign P[24] = in1[82] ^ in2[82];
    assign G[25] = in1[81] & in2[81];
    assign P[25] = in1[81] ^ in2[81];
    assign G[26] = in1[80] & in2[80];
    assign P[26] = in1[80] ^ in2[80];
    assign G[27] = in1[79] & in2[79];
    assign P[27] = in1[79] ^ in2[79];
    assign G[28] = in1[78] & in2[78];
    assign P[28] = in1[78] ^ in2[78];
    assign G[29] = in1[77] & in2[77];
    assign P[29] = in1[77] ^ in2[77];
    assign G[30] = in1[76] & in2[76];
    assign P[30] = in1[76] ^ in2[76];
    assign G[31] = in1[75] & in2[75];
    assign P[31] = in1[75] ^ in2[75];
    assign G[32] = in1[74] & in2[74];
    assign P[32] = in1[74] ^ in2[74];
    assign G[33] = in1[73] & in2[73];
    assign P[33] = in1[73] ^ in2[73];
    assign G[34] = in1[72] & in2[72];
    assign P[34] = in1[72] ^ in2[72];
    assign G[35] = in1[71] & in2[71];
    assign P[35] = in1[71] ^ in2[71];
    assign G[36] = in1[70] & in2[70];
    assign P[36] = in1[70] ^ in2[70];
    assign G[37] = in1[69] & in2[69];
    assign P[37] = in1[69] ^ in2[69];
    assign G[38] = in1[68] & in2[68];
    assign P[38] = in1[68] ^ in2[68];
    assign G[39] = in1[67] & in2[67];
    assign P[39] = in1[67] ^ in2[67];
    assign G[40] = in1[66] & in2[66];
    assign P[40] = in1[66] ^ in2[66];
    assign G[41] = in1[65] & in2[65];
    assign P[41] = in1[65] ^ in2[65];
    assign G[42] = in1[64] & in2[64];
    assign P[42] = in1[64] ^ in2[64];
    assign G[43] = in1[63] & in2[63];
    assign P[43] = in1[63] ^ in2[63];
    assign G[44] = in1[62] & in2[62];
    assign P[44] = in1[62] ^ in2[62];
    assign G[45] = in1[61] & in2[61];
    assign P[45] = in1[61] ^ in2[61];
    assign G[46] = in1[60] & in2[60];
    assign P[46] = in1[60] ^ in2[60];
    assign G[47] = in1[59] & in2[59];
    assign P[47] = in1[59] ^ in2[59];
    assign G[48] = in1[58] & in2[58];
    assign P[48] = in1[58] ^ in2[58];
    assign G[49] = in1[57] & in2[57];
    assign P[49] = in1[57] ^ in2[57];
    assign G[50] = in1[56] & in2[56];
    assign P[50] = in1[56] ^ in2[56];
    assign G[51] = in1[55] & in2[55];
    assign P[51] = in1[55] ^ in2[55];
    assign G[52] = in1[54] & in2[54];
    assign P[52] = in1[54] ^ in2[54];
    assign G[53] = in1[53] & in2[53];
    assign P[53] = in1[53] ^ in2[53];
    assign G[54] = in1[52] & in2[52];
    assign P[54] = in1[52] ^ in2[52];
    assign G[55] = in1[51] & in2[51];
    assign P[55] = in1[51] ^ in2[51];
    assign G[56] = in1[50] & in2[50];
    assign P[56] = in1[50] ^ in2[50];
    assign G[57] = in1[49] & in2[49];
    assign P[57] = in1[49] ^ in2[49];
    assign G[58] = in1[48] & in2[48];
    assign P[58] = in1[48] ^ in2[48];
    assign G[59] = in1[47] & in2[47];
    assign P[59] = in1[47] ^ in2[47];
    assign G[60] = in1[46] & in2[46];
    assign P[60] = in1[46] ^ in2[46];
    assign G[61] = in1[45] & in2[45];
    assign P[61] = in1[45] ^ in2[45];
    assign G[62] = in1[44] & in2[44];
    assign P[62] = in1[44] ^ in2[44];
    assign G[63] = in1[43] & in2[43];
    assign P[63] = in1[43] ^ in2[43];
    assign G[64] = in1[42] & in2[42];
    assign P[64] = in1[42] ^ in2[42];
    assign G[65] = in1[41] & in2[41];
    assign P[65] = in1[41] ^ in2[41];
    assign G[66] = in1[40] & in2[40];
    assign P[66] = in1[40] ^ in2[40];
    assign G[67] = in1[39] & in2[39];
    assign P[67] = in1[39] ^ in2[39];
    assign G[68] = in1[38] & in2[38];
    assign P[68] = in1[38] ^ in2[38];
    assign G[69] = in1[37] & in2[37];
    assign P[69] = in1[37] ^ in2[37];
    assign G[70] = in1[36] & in2[36];
    assign P[70] = in1[36] ^ in2[36];
    assign G[71] = in1[35] & in2[35];
    assign P[71] = in1[35] ^ in2[35];
    assign G[72] = in1[34] & in2[34];
    assign P[72] = in1[34] ^ in2[34];
    assign G[73] = in1[33] & in2[33];
    assign P[73] = in1[33] ^ in2[33];
    assign G[74] = in1[32] & in2[32];
    assign P[74] = in1[32] ^ in2[32];
    assign G[75] = in1[31] & in2[31];
    assign P[75] = in1[31] ^ in2[31];
    assign G[76] = in1[30] & in2[30];
    assign P[76] = in1[30] ^ in2[30];
    assign G[77] = in1[29] & in2[29];
    assign P[77] = in1[29] ^ in2[29];
    assign G[78] = in1[28] & in2[28];
    assign P[78] = in1[28] ^ in2[28];
    assign G[79] = in1[27] & in2[27];
    assign P[79] = in1[27] ^ in2[27];
    assign G[80] = in1[26] & in2[26];
    assign P[80] = in1[26] ^ in2[26];
    assign G[81] = in1[25] & in2[25];
    assign P[81] = in1[25] ^ in2[25];
    assign G[82] = in1[24] & in2[24];
    assign P[82] = in1[24] ^ in2[24];
    assign G[83] = in1[23] & in2[23];
    assign P[83] = in1[23] ^ in2[23];
    assign G[84] = in1[22] & in2[22];
    assign P[84] = in1[22] ^ in2[22];
    assign G[85] = in1[21] & in2[21];
    assign P[85] = in1[21] ^ in2[21];
    assign G[86] = in1[20] & in2[20];
    assign P[86] = in1[20] ^ in2[20];
    assign G[87] = in1[19] & in2[19];
    assign P[87] = in1[19] ^ in2[19];
    assign G[88] = in1[18] & in2[18];
    assign P[88] = in1[18] ^ in2[18];
    assign G[89] = in1[17] & in2[17];
    assign P[89] = in1[17] ^ in2[17];
    assign G[90] = in1[16] & in2[16];
    assign P[90] = in1[16] ^ in2[16];
    assign G[91] = in1[15] & in2[15];
    assign P[91] = in1[15] ^ in2[15];
    assign G[92] = in1[14] & in2[14];
    assign P[92] = in1[14] ^ in2[14];
    assign G[93] = in1[13] & in2[13];
    assign P[93] = in1[13] ^ in2[13];
    assign G[94] = in1[12] & in2[12];
    assign P[94] = in1[12] ^ in2[12];
    assign G[95] = in1[11] & in2[11];
    assign P[95] = in1[11] ^ in2[11];
    assign G[96] = in1[10] & in2[10];
    assign P[96] = in1[10] ^ in2[10];
    assign G[97] = in1[9] & in2[9];
    assign P[97] = in1[9] ^ in2[9];
    assign G[98] = in1[8] & in2[8];
    assign P[98] = in1[8] ^ in2[8];
    assign G[99] = in1[7] & in2[7];
    assign P[99] = in1[7] ^ in2[7];
    assign G[100] = in1[6] & in2[6];
    assign P[100] = in1[6] ^ in2[6];
    assign G[101] = in1[5] & in2[5];
    assign P[101] = in1[5] ^ in2[5];
    assign G[102] = in1[4] & in2[4];
    assign P[102] = in1[4] ^ in2[4];
    assign G[103] = in1[3] & in2[3];
    assign P[103] = in1[3] ^ in2[3];
    assign G[104] = in1[2] & in2[2];
    assign P[104] = in1[2] ^ in2[2];
    assign G[105] = in1[1] & in2[1];
    assign P[105] = in1[1] ^ in2[1];
    assign G[106] = in1[0] & in2[0];
    assign P[106] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign cout = G[106] | (P[106] & C[106]);
    assign sum = P ^ C;
endmodule

module CLA_106(output [105:0] sum, output cout, input [105:0] in1, input [105:0] in2);

    wire[105:0] G;
    wire[105:0] C;
    wire[105:0] P;

    assign G[0] = in1[105] & in2[105];
    assign P[0] = in1[105] ^ in2[105];
    assign G[1] = in1[104] & in2[104];
    assign P[1] = in1[104] ^ in2[104];
    assign G[2] = in1[103] & in2[103];
    assign P[2] = in1[103] ^ in2[103];
    assign G[3] = in1[102] & in2[102];
    assign P[3] = in1[102] ^ in2[102];
    assign G[4] = in1[101] & in2[101];
    assign P[4] = in1[101] ^ in2[101];
    assign G[5] = in1[100] & in2[100];
    assign P[5] = in1[100] ^ in2[100];
    assign G[6] = in1[99] & in2[99];
    assign P[6] = in1[99] ^ in2[99];
    assign G[7] = in1[98] & in2[98];
    assign P[7] = in1[98] ^ in2[98];
    assign G[8] = in1[97] & in2[97];
    assign P[8] = in1[97] ^ in2[97];
    assign G[9] = in1[96] & in2[96];
    assign P[9] = in1[96] ^ in2[96];
    assign G[10] = in1[95] & in2[95];
    assign P[10] = in1[95] ^ in2[95];
    assign G[11] = in1[94] & in2[94];
    assign P[11] = in1[94] ^ in2[94];
    assign G[12] = in1[93] & in2[93];
    assign P[12] = in1[93] ^ in2[93];
    assign G[13] = in1[92] & in2[92];
    assign P[13] = in1[92] ^ in2[92];
    assign G[14] = in1[91] & in2[91];
    assign P[14] = in1[91] ^ in2[91];
    assign G[15] = in1[90] & in2[90];
    assign P[15] = in1[90] ^ in2[90];
    assign G[16] = in1[89] & in2[89];
    assign P[16] = in1[89] ^ in2[89];
    assign G[17] = in1[88] & in2[88];
    assign P[17] = in1[88] ^ in2[88];
    assign G[18] = in1[87] & in2[87];
    assign P[18] = in1[87] ^ in2[87];
    assign G[19] = in1[86] & in2[86];
    assign P[19] = in1[86] ^ in2[86];
    assign G[20] = in1[85] & in2[85];
    assign P[20] = in1[85] ^ in2[85];
    assign G[21] = in1[84] & in2[84];
    assign P[21] = in1[84] ^ in2[84];
    assign G[22] = in1[83] & in2[83];
    assign P[22] = in1[83] ^ in2[83];
    assign G[23] = in1[82] & in2[82];
    assign P[23] = in1[82] ^ in2[82];
    assign G[24] = in1[81] & in2[81];
    assign P[24] = in1[81] ^ in2[81];
    assign G[25] = in1[80] & in2[80];
    assign P[25] = in1[80] ^ in2[80];
    assign G[26] = in1[79] & in2[79];
    assign P[26] = in1[79] ^ in2[79];
    assign G[27] = in1[78] & in2[78];
    assign P[27] = in1[78] ^ in2[78];
    assign G[28] = in1[77] & in2[77];
    assign P[28] = in1[77] ^ in2[77];
    assign G[29] = in1[76] & in2[76];
    assign P[29] = in1[76] ^ in2[76];
    assign G[30] = in1[75] & in2[75];
    assign P[30] = in1[75] ^ in2[75];
    assign G[31] = in1[74] & in2[74];
    assign P[31] = in1[74] ^ in2[74];
    assign G[32] = in1[73] & in2[73];
    assign P[32] = in1[73] ^ in2[73];
    assign G[33] = in1[72] & in2[72];
    assign P[33] = in1[72] ^ in2[72];
    assign G[34] = in1[71] & in2[71];
    assign P[34] = in1[71] ^ in2[71];
    assign G[35] = in1[70] & in2[70];
    assign P[35] = in1[70] ^ in2[70];
    assign G[36] = in1[69] & in2[69];
    assign P[36] = in1[69] ^ in2[69];
    assign G[37] = in1[68] & in2[68];
    assign P[37] = in1[68] ^ in2[68];
    assign G[38] = in1[67] & in2[67];
    assign P[38] = in1[67] ^ in2[67];
    assign G[39] = in1[66] & in2[66];
    assign P[39] = in1[66] ^ in2[66];
    assign G[40] = in1[65] & in2[65];
    assign P[40] = in1[65] ^ in2[65];
    assign G[41] = in1[64] & in2[64];
    assign P[41] = in1[64] ^ in2[64];
    assign G[42] = in1[63] & in2[63];
    assign P[42] = in1[63] ^ in2[63];
    assign G[43] = in1[62] & in2[62];
    assign P[43] = in1[62] ^ in2[62];
    assign G[44] = in1[61] & in2[61];
    assign P[44] = in1[61] ^ in2[61];
    assign G[45] = in1[60] & in2[60];
    assign P[45] = in1[60] ^ in2[60];
    assign G[46] = in1[59] & in2[59];
    assign P[46] = in1[59] ^ in2[59];
    assign G[47] = in1[58] & in2[58];
    assign P[47] = in1[58] ^ in2[58];
    assign G[48] = in1[57] & in2[57];
    assign P[48] = in1[57] ^ in2[57];
    assign G[49] = in1[56] & in2[56];
    assign P[49] = in1[56] ^ in2[56];
    assign G[50] = in1[55] & in2[55];
    assign P[50] = in1[55] ^ in2[55];
    assign G[51] = in1[54] & in2[54];
    assign P[51] = in1[54] ^ in2[54];
    assign G[52] = in1[53] & in2[53];
    assign P[52] = in1[53] ^ in2[53];
    assign G[53] = in1[52] & in2[52];
    assign P[53] = in1[52] ^ in2[52];
    assign G[54] = in1[51] & in2[51];
    assign P[54] = in1[51] ^ in2[51];
    assign G[55] = in1[50] & in2[50];
    assign P[55] = in1[50] ^ in2[50];
    assign G[56] = in1[49] & in2[49];
    assign P[56] = in1[49] ^ in2[49];
    assign G[57] = in1[48] & in2[48];
    assign P[57] = in1[48] ^ in2[48];
    assign G[58] = in1[47] & in2[47];
    assign P[58] = in1[47] ^ in2[47];
    assign G[59] = in1[46] & in2[46];
    assign P[59] = in1[46] ^ in2[46];
    assign G[60] = in1[45] & in2[45];
    assign P[60] = in1[45] ^ in2[45];
    assign G[61] = in1[44] & in2[44];
    assign P[61] = in1[44] ^ in2[44];
    assign G[62] = in1[43] & in2[43];
    assign P[62] = in1[43] ^ in2[43];
    assign G[63] = in1[42] & in2[42];
    assign P[63] = in1[42] ^ in2[42];
    assign G[64] = in1[41] & in2[41];
    assign P[64] = in1[41] ^ in2[41];
    assign G[65] = in1[40] & in2[40];
    assign P[65] = in1[40] ^ in2[40];
    assign G[66] = in1[39] & in2[39];
    assign P[66] = in1[39] ^ in2[39];
    assign G[67] = in1[38] & in2[38];
    assign P[67] = in1[38] ^ in2[38];
    assign G[68] = in1[37] & in2[37];
    assign P[68] = in1[37] ^ in2[37];
    assign G[69] = in1[36] & in2[36];
    assign P[69] = in1[36] ^ in2[36];
    assign G[70] = in1[35] & in2[35];
    assign P[70] = in1[35] ^ in2[35];
    assign G[71] = in1[34] & in2[34];
    assign P[71] = in1[34] ^ in2[34];
    assign G[72] = in1[33] & in2[33];
    assign P[72] = in1[33] ^ in2[33];
    assign G[73] = in1[32] & in2[32];
    assign P[73] = in1[32] ^ in2[32];
    assign G[74] = in1[31] & in2[31];
    assign P[74] = in1[31] ^ in2[31];
    assign G[75] = in1[30] & in2[30];
    assign P[75] = in1[30] ^ in2[30];
    assign G[76] = in1[29] & in2[29];
    assign P[76] = in1[29] ^ in2[29];
    assign G[77] = in1[28] & in2[28];
    assign P[77] = in1[28] ^ in2[28];
    assign G[78] = in1[27] & in2[27];
    assign P[78] = in1[27] ^ in2[27];
    assign G[79] = in1[26] & in2[26];
    assign P[79] = in1[26] ^ in2[26];
    assign G[80] = in1[25] & in2[25];
    assign P[80] = in1[25] ^ in2[25];
    assign G[81] = in1[24] & in2[24];
    assign P[81] = in1[24] ^ in2[24];
    assign G[82] = in1[23] & in2[23];
    assign P[82] = in1[23] ^ in2[23];
    assign G[83] = in1[22] & in2[22];
    assign P[83] = in1[22] ^ in2[22];
    assign G[84] = in1[21] & in2[21];
    assign P[84] = in1[21] ^ in2[21];
    assign G[85] = in1[20] & in2[20];
    assign P[85] = in1[20] ^ in2[20];
    assign G[86] = in1[19] & in2[19];
    assign P[86] = in1[19] ^ in2[19];
    assign G[87] = in1[18] & in2[18];
    assign P[87] = in1[18] ^ in2[18];
    assign G[88] = in1[17] & in2[17];
    assign P[88] = in1[17] ^ in2[17];
    assign G[89] = in1[16] & in2[16];
    assign P[89] = in1[16] ^ in2[16];
    assign G[90] = in1[15] & in2[15];
    assign P[90] = in1[15] ^ in2[15];
    assign G[91] = in1[14] & in2[14];
    assign P[91] = in1[14] ^ in2[14];
    assign G[92] = in1[13] & in2[13];
    assign P[92] = in1[13] ^ in2[13];
    assign G[93] = in1[12] & in2[12];
    assign P[93] = in1[12] ^ in2[12];
    assign G[94] = in1[11] & in2[11];
    assign P[94] = in1[11] ^ in2[11];
    assign G[95] = in1[10] & in2[10];
    assign P[95] = in1[10] ^ in2[10];
    assign G[96] = in1[9] & in2[9];
    assign P[96] = in1[9] ^ in2[9];
    assign G[97] = in1[8] & in2[8];
    assign P[97] = in1[8] ^ in2[8];
    assign G[98] = in1[7] & in2[7];
    assign P[98] = in1[7] ^ in2[7];
    assign G[99] = in1[6] & in2[6];
    assign P[99] = in1[6] ^ in2[6];
    assign G[100] = in1[5] & in2[5];
    assign P[100] = in1[5] ^ in2[5];
    assign G[101] = in1[4] & in2[4];
    assign P[101] = in1[4] ^ in2[4];
    assign G[102] = in1[3] & in2[3];
    assign P[102] = in1[3] ^ in2[3];
    assign G[103] = in1[2] & in2[2];
    assign P[103] = in1[2] ^ in2[2];
    assign G[104] = in1[1] & in2[1];
    assign P[104] = in1[1] ^ in2[1];
    assign G[105] = in1[0] & in2[0];
    assign P[105] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign cout = G[105] | (P[105] & C[105]);
    assign sum = P ^ C;
endmodule

module CLA_105(output [104:0] sum, output cout, input [104:0] in1, input [104:0] in2);

    wire[104:0] G;
    wire[104:0] C;
    wire[104:0] P;

    assign G[0] = in1[104] & in2[104];
    assign P[0] = in1[104] ^ in2[104];
    assign G[1] = in1[103] & in2[103];
    assign P[1] = in1[103] ^ in2[103];
    assign G[2] = in1[102] & in2[102];
    assign P[2] = in1[102] ^ in2[102];
    assign G[3] = in1[101] & in2[101];
    assign P[3] = in1[101] ^ in2[101];
    assign G[4] = in1[100] & in2[100];
    assign P[4] = in1[100] ^ in2[100];
    assign G[5] = in1[99] & in2[99];
    assign P[5] = in1[99] ^ in2[99];
    assign G[6] = in1[98] & in2[98];
    assign P[6] = in1[98] ^ in2[98];
    assign G[7] = in1[97] & in2[97];
    assign P[7] = in1[97] ^ in2[97];
    assign G[8] = in1[96] & in2[96];
    assign P[8] = in1[96] ^ in2[96];
    assign G[9] = in1[95] & in2[95];
    assign P[9] = in1[95] ^ in2[95];
    assign G[10] = in1[94] & in2[94];
    assign P[10] = in1[94] ^ in2[94];
    assign G[11] = in1[93] & in2[93];
    assign P[11] = in1[93] ^ in2[93];
    assign G[12] = in1[92] & in2[92];
    assign P[12] = in1[92] ^ in2[92];
    assign G[13] = in1[91] & in2[91];
    assign P[13] = in1[91] ^ in2[91];
    assign G[14] = in1[90] & in2[90];
    assign P[14] = in1[90] ^ in2[90];
    assign G[15] = in1[89] & in2[89];
    assign P[15] = in1[89] ^ in2[89];
    assign G[16] = in1[88] & in2[88];
    assign P[16] = in1[88] ^ in2[88];
    assign G[17] = in1[87] & in2[87];
    assign P[17] = in1[87] ^ in2[87];
    assign G[18] = in1[86] & in2[86];
    assign P[18] = in1[86] ^ in2[86];
    assign G[19] = in1[85] & in2[85];
    assign P[19] = in1[85] ^ in2[85];
    assign G[20] = in1[84] & in2[84];
    assign P[20] = in1[84] ^ in2[84];
    assign G[21] = in1[83] & in2[83];
    assign P[21] = in1[83] ^ in2[83];
    assign G[22] = in1[82] & in2[82];
    assign P[22] = in1[82] ^ in2[82];
    assign G[23] = in1[81] & in2[81];
    assign P[23] = in1[81] ^ in2[81];
    assign G[24] = in1[80] & in2[80];
    assign P[24] = in1[80] ^ in2[80];
    assign G[25] = in1[79] & in2[79];
    assign P[25] = in1[79] ^ in2[79];
    assign G[26] = in1[78] & in2[78];
    assign P[26] = in1[78] ^ in2[78];
    assign G[27] = in1[77] & in2[77];
    assign P[27] = in1[77] ^ in2[77];
    assign G[28] = in1[76] & in2[76];
    assign P[28] = in1[76] ^ in2[76];
    assign G[29] = in1[75] & in2[75];
    assign P[29] = in1[75] ^ in2[75];
    assign G[30] = in1[74] & in2[74];
    assign P[30] = in1[74] ^ in2[74];
    assign G[31] = in1[73] & in2[73];
    assign P[31] = in1[73] ^ in2[73];
    assign G[32] = in1[72] & in2[72];
    assign P[32] = in1[72] ^ in2[72];
    assign G[33] = in1[71] & in2[71];
    assign P[33] = in1[71] ^ in2[71];
    assign G[34] = in1[70] & in2[70];
    assign P[34] = in1[70] ^ in2[70];
    assign G[35] = in1[69] & in2[69];
    assign P[35] = in1[69] ^ in2[69];
    assign G[36] = in1[68] & in2[68];
    assign P[36] = in1[68] ^ in2[68];
    assign G[37] = in1[67] & in2[67];
    assign P[37] = in1[67] ^ in2[67];
    assign G[38] = in1[66] & in2[66];
    assign P[38] = in1[66] ^ in2[66];
    assign G[39] = in1[65] & in2[65];
    assign P[39] = in1[65] ^ in2[65];
    assign G[40] = in1[64] & in2[64];
    assign P[40] = in1[64] ^ in2[64];
    assign G[41] = in1[63] & in2[63];
    assign P[41] = in1[63] ^ in2[63];
    assign G[42] = in1[62] & in2[62];
    assign P[42] = in1[62] ^ in2[62];
    assign G[43] = in1[61] & in2[61];
    assign P[43] = in1[61] ^ in2[61];
    assign G[44] = in1[60] & in2[60];
    assign P[44] = in1[60] ^ in2[60];
    assign G[45] = in1[59] & in2[59];
    assign P[45] = in1[59] ^ in2[59];
    assign G[46] = in1[58] & in2[58];
    assign P[46] = in1[58] ^ in2[58];
    assign G[47] = in1[57] & in2[57];
    assign P[47] = in1[57] ^ in2[57];
    assign G[48] = in1[56] & in2[56];
    assign P[48] = in1[56] ^ in2[56];
    assign G[49] = in1[55] & in2[55];
    assign P[49] = in1[55] ^ in2[55];
    assign G[50] = in1[54] & in2[54];
    assign P[50] = in1[54] ^ in2[54];
    assign G[51] = in1[53] & in2[53];
    assign P[51] = in1[53] ^ in2[53];
    assign G[52] = in1[52] & in2[52];
    assign P[52] = in1[52] ^ in2[52];
    assign G[53] = in1[51] & in2[51];
    assign P[53] = in1[51] ^ in2[51];
    assign G[54] = in1[50] & in2[50];
    assign P[54] = in1[50] ^ in2[50];
    assign G[55] = in1[49] & in2[49];
    assign P[55] = in1[49] ^ in2[49];
    assign G[56] = in1[48] & in2[48];
    assign P[56] = in1[48] ^ in2[48];
    assign G[57] = in1[47] & in2[47];
    assign P[57] = in1[47] ^ in2[47];
    assign G[58] = in1[46] & in2[46];
    assign P[58] = in1[46] ^ in2[46];
    assign G[59] = in1[45] & in2[45];
    assign P[59] = in1[45] ^ in2[45];
    assign G[60] = in1[44] & in2[44];
    assign P[60] = in1[44] ^ in2[44];
    assign G[61] = in1[43] & in2[43];
    assign P[61] = in1[43] ^ in2[43];
    assign G[62] = in1[42] & in2[42];
    assign P[62] = in1[42] ^ in2[42];
    assign G[63] = in1[41] & in2[41];
    assign P[63] = in1[41] ^ in2[41];
    assign G[64] = in1[40] & in2[40];
    assign P[64] = in1[40] ^ in2[40];
    assign G[65] = in1[39] & in2[39];
    assign P[65] = in1[39] ^ in2[39];
    assign G[66] = in1[38] & in2[38];
    assign P[66] = in1[38] ^ in2[38];
    assign G[67] = in1[37] & in2[37];
    assign P[67] = in1[37] ^ in2[37];
    assign G[68] = in1[36] & in2[36];
    assign P[68] = in1[36] ^ in2[36];
    assign G[69] = in1[35] & in2[35];
    assign P[69] = in1[35] ^ in2[35];
    assign G[70] = in1[34] & in2[34];
    assign P[70] = in1[34] ^ in2[34];
    assign G[71] = in1[33] & in2[33];
    assign P[71] = in1[33] ^ in2[33];
    assign G[72] = in1[32] & in2[32];
    assign P[72] = in1[32] ^ in2[32];
    assign G[73] = in1[31] & in2[31];
    assign P[73] = in1[31] ^ in2[31];
    assign G[74] = in1[30] & in2[30];
    assign P[74] = in1[30] ^ in2[30];
    assign G[75] = in1[29] & in2[29];
    assign P[75] = in1[29] ^ in2[29];
    assign G[76] = in1[28] & in2[28];
    assign P[76] = in1[28] ^ in2[28];
    assign G[77] = in1[27] & in2[27];
    assign P[77] = in1[27] ^ in2[27];
    assign G[78] = in1[26] & in2[26];
    assign P[78] = in1[26] ^ in2[26];
    assign G[79] = in1[25] & in2[25];
    assign P[79] = in1[25] ^ in2[25];
    assign G[80] = in1[24] & in2[24];
    assign P[80] = in1[24] ^ in2[24];
    assign G[81] = in1[23] & in2[23];
    assign P[81] = in1[23] ^ in2[23];
    assign G[82] = in1[22] & in2[22];
    assign P[82] = in1[22] ^ in2[22];
    assign G[83] = in1[21] & in2[21];
    assign P[83] = in1[21] ^ in2[21];
    assign G[84] = in1[20] & in2[20];
    assign P[84] = in1[20] ^ in2[20];
    assign G[85] = in1[19] & in2[19];
    assign P[85] = in1[19] ^ in2[19];
    assign G[86] = in1[18] & in2[18];
    assign P[86] = in1[18] ^ in2[18];
    assign G[87] = in1[17] & in2[17];
    assign P[87] = in1[17] ^ in2[17];
    assign G[88] = in1[16] & in2[16];
    assign P[88] = in1[16] ^ in2[16];
    assign G[89] = in1[15] & in2[15];
    assign P[89] = in1[15] ^ in2[15];
    assign G[90] = in1[14] & in2[14];
    assign P[90] = in1[14] ^ in2[14];
    assign G[91] = in1[13] & in2[13];
    assign P[91] = in1[13] ^ in2[13];
    assign G[92] = in1[12] & in2[12];
    assign P[92] = in1[12] ^ in2[12];
    assign G[93] = in1[11] & in2[11];
    assign P[93] = in1[11] ^ in2[11];
    assign G[94] = in1[10] & in2[10];
    assign P[94] = in1[10] ^ in2[10];
    assign G[95] = in1[9] & in2[9];
    assign P[95] = in1[9] ^ in2[9];
    assign G[96] = in1[8] & in2[8];
    assign P[96] = in1[8] ^ in2[8];
    assign G[97] = in1[7] & in2[7];
    assign P[97] = in1[7] ^ in2[7];
    assign G[98] = in1[6] & in2[6];
    assign P[98] = in1[6] ^ in2[6];
    assign G[99] = in1[5] & in2[5];
    assign P[99] = in1[5] ^ in2[5];
    assign G[100] = in1[4] & in2[4];
    assign P[100] = in1[4] ^ in2[4];
    assign G[101] = in1[3] & in2[3];
    assign P[101] = in1[3] ^ in2[3];
    assign G[102] = in1[2] & in2[2];
    assign P[102] = in1[2] ^ in2[2];
    assign G[103] = in1[1] & in2[1];
    assign P[103] = in1[1] ^ in2[1];
    assign G[104] = in1[0] & in2[0];
    assign P[104] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign cout = G[104] | (P[104] & C[104]);
    assign sum = P ^ C;
endmodule

module CLA_104(output [103:0] sum, output cout, input [103:0] in1, input [103:0] in2);

    wire[103:0] G;
    wire[103:0] C;
    wire[103:0] P;

    assign G[0] = in1[103] & in2[103];
    assign P[0] = in1[103] ^ in2[103];
    assign G[1] = in1[102] & in2[102];
    assign P[1] = in1[102] ^ in2[102];
    assign G[2] = in1[101] & in2[101];
    assign P[2] = in1[101] ^ in2[101];
    assign G[3] = in1[100] & in2[100];
    assign P[3] = in1[100] ^ in2[100];
    assign G[4] = in1[99] & in2[99];
    assign P[4] = in1[99] ^ in2[99];
    assign G[5] = in1[98] & in2[98];
    assign P[5] = in1[98] ^ in2[98];
    assign G[6] = in1[97] & in2[97];
    assign P[6] = in1[97] ^ in2[97];
    assign G[7] = in1[96] & in2[96];
    assign P[7] = in1[96] ^ in2[96];
    assign G[8] = in1[95] & in2[95];
    assign P[8] = in1[95] ^ in2[95];
    assign G[9] = in1[94] & in2[94];
    assign P[9] = in1[94] ^ in2[94];
    assign G[10] = in1[93] & in2[93];
    assign P[10] = in1[93] ^ in2[93];
    assign G[11] = in1[92] & in2[92];
    assign P[11] = in1[92] ^ in2[92];
    assign G[12] = in1[91] & in2[91];
    assign P[12] = in1[91] ^ in2[91];
    assign G[13] = in1[90] & in2[90];
    assign P[13] = in1[90] ^ in2[90];
    assign G[14] = in1[89] & in2[89];
    assign P[14] = in1[89] ^ in2[89];
    assign G[15] = in1[88] & in2[88];
    assign P[15] = in1[88] ^ in2[88];
    assign G[16] = in1[87] & in2[87];
    assign P[16] = in1[87] ^ in2[87];
    assign G[17] = in1[86] & in2[86];
    assign P[17] = in1[86] ^ in2[86];
    assign G[18] = in1[85] & in2[85];
    assign P[18] = in1[85] ^ in2[85];
    assign G[19] = in1[84] & in2[84];
    assign P[19] = in1[84] ^ in2[84];
    assign G[20] = in1[83] & in2[83];
    assign P[20] = in1[83] ^ in2[83];
    assign G[21] = in1[82] & in2[82];
    assign P[21] = in1[82] ^ in2[82];
    assign G[22] = in1[81] & in2[81];
    assign P[22] = in1[81] ^ in2[81];
    assign G[23] = in1[80] & in2[80];
    assign P[23] = in1[80] ^ in2[80];
    assign G[24] = in1[79] & in2[79];
    assign P[24] = in1[79] ^ in2[79];
    assign G[25] = in1[78] & in2[78];
    assign P[25] = in1[78] ^ in2[78];
    assign G[26] = in1[77] & in2[77];
    assign P[26] = in1[77] ^ in2[77];
    assign G[27] = in1[76] & in2[76];
    assign P[27] = in1[76] ^ in2[76];
    assign G[28] = in1[75] & in2[75];
    assign P[28] = in1[75] ^ in2[75];
    assign G[29] = in1[74] & in2[74];
    assign P[29] = in1[74] ^ in2[74];
    assign G[30] = in1[73] & in2[73];
    assign P[30] = in1[73] ^ in2[73];
    assign G[31] = in1[72] & in2[72];
    assign P[31] = in1[72] ^ in2[72];
    assign G[32] = in1[71] & in2[71];
    assign P[32] = in1[71] ^ in2[71];
    assign G[33] = in1[70] & in2[70];
    assign P[33] = in1[70] ^ in2[70];
    assign G[34] = in1[69] & in2[69];
    assign P[34] = in1[69] ^ in2[69];
    assign G[35] = in1[68] & in2[68];
    assign P[35] = in1[68] ^ in2[68];
    assign G[36] = in1[67] & in2[67];
    assign P[36] = in1[67] ^ in2[67];
    assign G[37] = in1[66] & in2[66];
    assign P[37] = in1[66] ^ in2[66];
    assign G[38] = in1[65] & in2[65];
    assign P[38] = in1[65] ^ in2[65];
    assign G[39] = in1[64] & in2[64];
    assign P[39] = in1[64] ^ in2[64];
    assign G[40] = in1[63] & in2[63];
    assign P[40] = in1[63] ^ in2[63];
    assign G[41] = in1[62] & in2[62];
    assign P[41] = in1[62] ^ in2[62];
    assign G[42] = in1[61] & in2[61];
    assign P[42] = in1[61] ^ in2[61];
    assign G[43] = in1[60] & in2[60];
    assign P[43] = in1[60] ^ in2[60];
    assign G[44] = in1[59] & in2[59];
    assign P[44] = in1[59] ^ in2[59];
    assign G[45] = in1[58] & in2[58];
    assign P[45] = in1[58] ^ in2[58];
    assign G[46] = in1[57] & in2[57];
    assign P[46] = in1[57] ^ in2[57];
    assign G[47] = in1[56] & in2[56];
    assign P[47] = in1[56] ^ in2[56];
    assign G[48] = in1[55] & in2[55];
    assign P[48] = in1[55] ^ in2[55];
    assign G[49] = in1[54] & in2[54];
    assign P[49] = in1[54] ^ in2[54];
    assign G[50] = in1[53] & in2[53];
    assign P[50] = in1[53] ^ in2[53];
    assign G[51] = in1[52] & in2[52];
    assign P[51] = in1[52] ^ in2[52];
    assign G[52] = in1[51] & in2[51];
    assign P[52] = in1[51] ^ in2[51];
    assign G[53] = in1[50] & in2[50];
    assign P[53] = in1[50] ^ in2[50];
    assign G[54] = in1[49] & in2[49];
    assign P[54] = in1[49] ^ in2[49];
    assign G[55] = in1[48] & in2[48];
    assign P[55] = in1[48] ^ in2[48];
    assign G[56] = in1[47] & in2[47];
    assign P[56] = in1[47] ^ in2[47];
    assign G[57] = in1[46] & in2[46];
    assign P[57] = in1[46] ^ in2[46];
    assign G[58] = in1[45] & in2[45];
    assign P[58] = in1[45] ^ in2[45];
    assign G[59] = in1[44] & in2[44];
    assign P[59] = in1[44] ^ in2[44];
    assign G[60] = in1[43] & in2[43];
    assign P[60] = in1[43] ^ in2[43];
    assign G[61] = in1[42] & in2[42];
    assign P[61] = in1[42] ^ in2[42];
    assign G[62] = in1[41] & in2[41];
    assign P[62] = in1[41] ^ in2[41];
    assign G[63] = in1[40] & in2[40];
    assign P[63] = in1[40] ^ in2[40];
    assign G[64] = in1[39] & in2[39];
    assign P[64] = in1[39] ^ in2[39];
    assign G[65] = in1[38] & in2[38];
    assign P[65] = in1[38] ^ in2[38];
    assign G[66] = in1[37] & in2[37];
    assign P[66] = in1[37] ^ in2[37];
    assign G[67] = in1[36] & in2[36];
    assign P[67] = in1[36] ^ in2[36];
    assign G[68] = in1[35] & in2[35];
    assign P[68] = in1[35] ^ in2[35];
    assign G[69] = in1[34] & in2[34];
    assign P[69] = in1[34] ^ in2[34];
    assign G[70] = in1[33] & in2[33];
    assign P[70] = in1[33] ^ in2[33];
    assign G[71] = in1[32] & in2[32];
    assign P[71] = in1[32] ^ in2[32];
    assign G[72] = in1[31] & in2[31];
    assign P[72] = in1[31] ^ in2[31];
    assign G[73] = in1[30] & in2[30];
    assign P[73] = in1[30] ^ in2[30];
    assign G[74] = in1[29] & in2[29];
    assign P[74] = in1[29] ^ in2[29];
    assign G[75] = in1[28] & in2[28];
    assign P[75] = in1[28] ^ in2[28];
    assign G[76] = in1[27] & in2[27];
    assign P[76] = in1[27] ^ in2[27];
    assign G[77] = in1[26] & in2[26];
    assign P[77] = in1[26] ^ in2[26];
    assign G[78] = in1[25] & in2[25];
    assign P[78] = in1[25] ^ in2[25];
    assign G[79] = in1[24] & in2[24];
    assign P[79] = in1[24] ^ in2[24];
    assign G[80] = in1[23] & in2[23];
    assign P[80] = in1[23] ^ in2[23];
    assign G[81] = in1[22] & in2[22];
    assign P[81] = in1[22] ^ in2[22];
    assign G[82] = in1[21] & in2[21];
    assign P[82] = in1[21] ^ in2[21];
    assign G[83] = in1[20] & in2[20];
    assign P[83] = in1[20] ^ in2[20];
    assign G[84] = in1[19] & in2[19];
    assign P[84] = in1[19] ^ in2[19];
    assign G[85] = in1[18] & in2[18];
    assign P[85] = in1[18] ^ in2[18];
    assign G[86] = in1[17] & in2[17];
    assign P[86] = in1[17] ^ in2[17];
    assign G[87] = in1[16] & in2[16];
    assign P[87] = in1[16] ^ in2[16];
    assign G[88] = in1[15] & in2[15];
    assign P[88] = in1[15] ^ in2[15];
    assign G[89] = in1[14] & in2[14];
    assign P[89] = in1[14] ^ in2[14];
    assign G[90] = in1[13] & in2[13];
    assign P[90] = in1[13] ^ in2[13];
    assign G[91] = in1[12] & in2[12];
    assign P[91] = in1[12] ^ in2[12];
    assign G[92] = in1[11] & in2[11];
    assign P[92] = in1[11] ^ in2[11];
    assign G[93] = in1[10] & in2[10];
    assign P[93] = in1[10] ^ in2[10];
    assign G[94] = in1[9] & in2[9];
    assign P[94] = in1[9] ^ in2[9];
    assign G[95] = in1[8] & in2[8];
    assign P[95] = in1[8] ^ in2[8];
    assign G[96] = in1[7] & in2[7];
    assign P[96] = in1[7] ^ in2[7];
    assign G[97] = in1[6] & in2[6];
    assign P[97] = in1[6] ^ in2[6];
    assign G[98] = in1[5] & in2[5];
    assign P[98] = in1[5] ^ in2[5];
    assign G[99] = in1[4] & in2[4];
    assign P[99] = in1[4] ^ in2[4];
    assign G[100] = in1[3] & in2[3];
    assign P[100] = in1[3] ^ in2[3];
    assign G[101] = in1[2] & in2[2];
    assign P[101] = in1[2] ^ in2[2];
    assign G[102] = in1[1] & in2[1];
    assign P[102] = in1[1] ^ in2[1];
    assign G[103] = in1[0] & in2[0];
    assign P[103] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign cout = G[103] | (P[103] & C[103]);
    assign sum = P ^ C;
endmodule

module CLA_103(output [102:0] sum, output cout, input [102:0] in1, input [102:0] in2);

    wire[102:0] G;
    wire[102:0] C;
    wire[102:0] P;

    assign G[0] = in1[102] & in2[102];
    assign P[0] = in1[102] ^ in2[102];
    assign G[1] = in1[101] & in2[101];
    assign P[1] = in1[101] ^ in2[101];
    assign G[2] = in1[100] & in2[100];
    assign P[2] = in1[100] ^ in2[100];
    assign G[3] = in1[99] & in2[99];
    assign P[3] = in1[99] ^ in2[99];
    assign G[4] = in1[98] & in2[98];
    assign P[4] = in1[98] ^ in2[98];
    assign G[5] = in1[97] & in2[97];
    assign P[5] = in1[97] ^ in2[97];
    assign G[6] = in1[96] & in2[96];
    assign P[6] = in1[96] ^ in2[96];
    assign G[7] = in1[95] & in2[95];
    assign P[7] = in1[95] ^ in2[95];
    assign G[8] = in1[94] & in2[94];
    assign P[8] = in1[94] ^ in2[94];
    assign G[9] = in1[93] & in2[93];
    assign P[9] = in1[93] ^ in2[93];
    assign G[10] = in1[92] & in2[92];
    assign P[10] = in1[92] ^ in2[92];
    assign G[11] = in1[91] & in2[91];
    assign P[11] = in1[91] ^ in2[91];
    assign G[12] = in1[90] & in2[90];
    assign P[12] = in1[90] ^ in2[90];
    assign G[13] = in1[89] & in2[89];
    assign P[13] = in1[89] ^ in2[89];
    assign G[14] = in1[88] & in2[88];
    assign P[14] = in1[88] ^ in2[88];
    assign G[15] = in1[87] & in2[87];
    assign P[15] = in1[87] ^ in2[87];
    assign G[16] = in1[86] & in2[86];
    assign P[16] = in1[86] ^ in2[86];
    assign G[17] = in1[85] & in2[85];
    assign P[17] = in1[85] ^ in2[85];
    assign G[18] = in1[84] & in2[84];
    assign P[18] = in1[84] ^ in2[84];
    assign G[19] = in1[83] & in2[83];
    assign P[19] = in1[83] ^ in2[83];
    assign G[20] = in1[82] & in2[82];
    assign P[20] = in1[82] ^ in2[82];
    assign G[21] = in1[81] & in2[81];
    assign P[21] = in1[81] ^ in2[81];
    assign G[22] = in1[80] & in2[80];
    assign P[22] = in1[80] ^ in2[80];
    assign G[23] = in1[79] & in2[79];
    assign P[23] = in1[79] ^ in2[79];
    assign G[24] = in1[78] & in2[78];
    assign P[24] = in1[78] ^ in2[78];
    assign G[25] = in1[77] & in2[77];
    assign P[25] = in1[77] ^ in2[77];
    assign G[26] = in1[76] & in2[76];
    assign P[26] = in1[76] ^ in2[76];
    assign G[27] = in1[75] & in2[75];
    assign P[27] = in1[75] ^ in2[75];
    assign G[28] = in1[74] & in2[74];
    assign P[28] = in1[74] ^ in2[74];
    assign G[29] = in1[73] & in2[73];
    assign P[29] = in1[73] ^ in2[73];
    assign G[30] = in1[72] & in2[72];
    assign P[30] = in1[72] ^ in2[72];
    assign G[31] = in1[71] & in2[71];
    assign P[31] = in1[71] ^ in2[71];
    assign G[32] = in1[70] & in2[70];
    assign P[32] = in1[70] ^ in2[70];
    assign G[33] = in1[69] & in2[69];
    assign P[33] = in1[69] ^ in2[69];
    assign G[34] = in1[68] & in2[68];
    assign P[34] = in1[68] ^ in2[68];
    assign G[35] = in1[67] & in2[67];
    assign P[35] = in1[67] ^ in2[67];
    assign G[36] = in1[66] & in2[66];
    assign P[36] = in1[66] ^ in2[66];
    assign G[37] = in1[65] & in2[65];
    assign P[37] = in1[65] ^ in2[65];
    assign G[38] = in1[64] & in2[64];
    assign P[38] = in1[64] ^ in2[64];
    assign G[39] = in1[63] & in2[63];
    assign P[39] = in1[63] ^ in2[63];
    assign G[40] = in1[62] & in2[62];
    assign P[40] = in1[62] ^ in2[62];
    assign G[41] = in1[61] & in2[61];
    assign P[41] = in1[61] ^ in2[61];
    assign G[42] = in1[60] & in2[60];
    assign P[42] = in1[60] ^ in2[60];
    assign G[43] = in1[59] & in2[59];
    assign P[43] = in1[59] ^ in2[59];
    assign G[44] = in1[58] & in2[58];
    assign P[44] = in1[58] ^ in2[58];
    assign G[45] = in1[57] & in2[57];
    assign P[45] = in1[57] ^ in2[57];
    assign G[46] = in1[56] & in2[56];
    assign P[46] = in1[56] ^ in2[56];
    assign G[47] = in1[55] & in2[55];
    assign P[47] = in1[55] ^ in2[55];
    assign G[48] = in1[54] & in2[54];
    assign P[48] = in1[54] ^ in2[54];
    assign G[49] = in1[53] & in2[53];
    assign P[49] = in1[53] ^ in2[53];
    assign G[50] = in1[52] & in2[52];
    assign P[50] = in1[52] ^ in2[52];
    assign G[51] = in1[51] & in2[51];
    assign P[51] = in1[51] ^ in2[51];
    assign G[52] = in1[50] & in2[50];
    assign P[52] = in1[50] ^ in2[50];
    assign G[53] = in1[49] & in2[49];
    assign P[53] = in1[49] ^ in2[49];
    assign G[54] = in1[48] & in2[48];
    assign P[54] = in1[48] ^ in2[48];
    assign G[55] = in1[47] & in2[47];
    assign P[55] = in1[47] ^ in2[47];
    assign G[56] = in1[46] & in2[46];
    assign P[56] = in1[46] ^ in2[46];
    assign G[57] = in1[45] & in2[45];
    assign P[57] = in1[45] ^ in2[45];
    assign G[58] = in1[44] & in2[44];
    assign P[58] = in1[44] ^ in2[44];
    assign G[59] = in1[43] & in2[43];
    assign P[59] = in1[43] ^ in2[43];
    assign G[60] = in1[42] & in2[42];
    assign P[60] = in1[42] ^ in2[42];
    assign G[61] = in1[41] & in2[41];
    assign P[61] = in1[41] ^ in2[41];
    assign G[62] = in1[40] & in2[40];
    assign P[62] = in1[40] ^ in2[40];
    assign G[63] = in1[39] & in2[39];
    assign P[63] = in1[39] ^ in2[39];
    assign G[64] = in1[38] & in2[38];
    assign P[64] = in1[38] ^ in2[38];
    assign G[65] = in1[37] & in2[37];
    assign P[65] = in1[37] ^ in2[37];
    assign G[66] = in1[36] & in2[36];
    assign P[66] = in1[36] ^ in2[36];
    assign G[67] = in1[35] & in2[35];
    assign P[67] = in1[35] ^ in2[35];
    assign G[68] = in1[34] & in2[34];
    assign P[68] = in1[34] ^ in2[34];
    assign G[69] = in1[33] & in2[33];
    assign P[69] = in1[33] ^ in2[33];
    assign G[70] = in1[32] & in2[32];
    assign P[70] = in1[32] ^ in2[32];
    assign G[71] = in1[31] & in2[31];
    assign P[71] = in1[31] ^ in2[31];
    assign G[72] = in1[30] & in2[30];
    assign P[72] = in1[30] ^ in2[30];
    assign G[73] = in1[29] & in2[29];
    assign P[73] = in1[29] ^ in2[29];
    assign G[74] = in1[28] & in2[28];
    assign P[74] = in1[28] ^ in2[28];
    assign G[75] = in1[27] & in2[27];
    assign P[75] = in1[27] ^ in2[27];
    assign G[76] = in1[26] & in2[26];
    assign P[76] = in1[26] ^ in2[26];
    assign G[77] = in1[25] & in2[25];
    assign P[77] = in1[25] ^ in2[25];
    assign G[78] = in1[24] & in2[24];
    assign P[78] = in1[24] ^ in2[24];
    assign G[79] = in1[23] & in2[23];
    assign P[79] = in1[23] ^ in2[23];
    assign G[80] = in1[22] & in2[22];
    assign P[80] = in1[22] ^ in2[22];
    assign G[81] = in1[21] & in2[21];
    assign P[81] = in1[21] ^ in2[21];
    assign G[82] = in1[20] & in2[20];
    assign P[82] = in1[20] ^ in2[20];
    assign G[83] = in1[19] & in2[19];
    assign P[83] = in1[19] ^ in2[19];
    assign G[84] = in1[18] & in2[18];
    assign P[84] = in1[18] ^ in2[18];
    assign G[85] = in1[17] & in2[17];
    assign P[85] = in1[17] ^ in2[17];
    assign G[86] = in1[16] & in2[16];
    assign P[86] = in1[16] ^ in2[16];
    assign G[87] = in1[15] & in2[15];
    assign P[87] = in1[15] ^ in2[15];
    assign G[88] = in1[14] & in2[14];
    assign P[88] = in1[14] ^ in2[14];
    assign G[89] = in1[13] & in2[13];
    assign P[89] = in1[13] ^ in2[13];
    assign G[90] = in1[12] & in2[12];
    assign P[90] = in1[12] ^ in2[12];
    assign G[91] = in1[11] & in2[11];
    assign P[91] = in1[11] ^ in2[11];
    assign G[92] = in1[10] & in2[10];
    assign P[92] = in1[10] ^ in2[10];
    assign G[93] = in1[9] & in2[9];
    assign P[93] = in1[9] ^ in2[9];
    assign G[94] = in1[8] & in2[8];
    assign P[94] = in1[8] ^ in2[8];
    assign G[95] = in1[7] & in2[7];
    assign P[95] = in1[7] ^ in2[7];
    assign G[96] = in1[6] & in2[6];
    assign P[96] = in1[6] ^ in2[6];
    assign G[97] = in1[5] & in2[5];
    assign P[97] = in1[5] ^ in2[5];
    assign G[98] = in1[4] & in2[4];
    assign P[98] = in1[4] ^ in2[4];
    assign G[99] = in1[3] & in2[3];
    assign P[99] = in1[3] ^ in2[3];
    assign G[100] = in1[2] & in2[2];
    assign P[100] = in1[2] ^ in2[2];
    assign G[101] = in1[1] & in2[1];
    assign P[101] = in1[1] ^ in2[1];
    assign G[102] = in1[0] & in2[0];
    assign P[102] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign cout = G[102] | (P[102] & C[102]);
    assign sum = P ^ C;
endmodule

module CLA_102(output [101:0] sum, output cout, input [101:0] in1, input [101:0] in2);

    wire[101:0] G;
    wire[101:0] C;
    wire[101:0] P;

    assign G[0] = in1[101] & in2[101];
    assign P[0] = in1[101] ^ in2[101];
    assign G[1] = in1[100] & in2[100];
    assign P[1] = in1[100] ^ in2[100];
    assign G[2] = in1[99] & in2[99];
    assign P[2] = in1[99] ^ in2[99];
    assign G[3] = in1[98] & in2[98];
    assign P[3] = in1[98] ^ in2[98];
    assign G[4] = in1[97] & in2[97];
    assign P[4] = in1[97] ^ in2[97];
    assign G[5] = in1[96] & in2[96];
    assign P[5] = in1[96] ^ in2[96];
    assign G[6] = in1[95] & in2[95];
    assign P[6] = in1[95] ^ in2[95];
    assign G[7] = in1[94] & in2[94];
    assign P[7] = in1[94] ^ in2[94];
    assign G[8] = in1[93] & in2[93];
    assign P[8] = in1[93] ^ in2[93];
    assign G[9] = in1[92] & in2[92];
    assign P[9] = in1[92] ^ in2[92];
    assign G[10] = in1[91] & in2[91];
    assign P[10] = in1[91] ^ in2[91];
    assign G[11] = in1[90] & in2[90];
    assign P[11] = in1[90] ^ in2[90];
    assign G[12] = in1[89] & in2[89];
    assign P[12] = in1[89] ^ in2[89];
    assign G[13] = in1[88] & in2[88];
    assign P[13] = in1[88] ^ in2[88];
    assign G[14] = in1[87] & in2[87];
    assign P[14] = in1[87] ^ in2[87];
    assign G[15] = in1[86] & in2[86];
    assign P[15] = in1[86] ^ in2[86];
    assign G[16] = in1[85] & in2[85];
    assign P[16] = in1[85] ^ in2[85];
    assign G[17] = in1[84] & in2[84];
    assign P[17] = in1[84] ^ in2[84];
    assign G[18] = in1[83] & in2[83];
    assign P[18] = in1[83] ^ in2[83];
    assign G[19] = in1[82] & in2[82];
    assign P[19] = in1[82] ^ in2[82];
    assign G[20] = in1[81] & in2[81];
    assign P[20] = in1[81] ^ in2[81];
    assign G[21] = in1[80] & in2[80];
    assign P[21] = in1[80] ^ in2[80];
    assign G[22] = in1[79] & in2[79];
    assign P[22] = in1[79] ^ in2[79];
    assign G[23] = in1[78] & in2[78];
    assign P[23] = in1[78] ^ in2[78];
    assign G[24] = in1[77] & in2[77];
    assign P[24] = in1[77] ^ in2[77];
    assign G[25] = in1[76] & in2[76];
    assign P[25] = in1[76] ^ in2[76];
    assign G[26] = in1[75] & in2[75];
    assign P[26] = in1[75] ^ in2[75];
    assign G[27] = in1[74] & in2[74];
    assign P[27] = in1[74] ^ in2[74];
    assign G[28] = in1[73] & in2[73];
    assign P[28] = in1[73] ^ in2[73];
    assign G[29] = in1[72] & in2[72];
    assign P[29] = in1[72] ^ in2[72];
    assign G[30] = in1[71] & in2[71];
    assign P[30] = in1[71] ^ in2[71];
    assign G[31] = in1[70] & in2[70];
    assign P[31] = in1[70] ^ in2[70];
    assign G[32] = in1[69] & in2[69];
    assign P[32] = in1[69] ^ in2[69];
    assign G[33] = in1[68] & in2[68];
    assign P[33] = in1[68] ^ in2[68];
    assign G[34] = in1[67] & in2[67];
    assign P[34] = in1[67] ^ in2[67];
    assign G[35] = in1[66] & in2[66];
    assign P[35] = in1[66] ^ in2[66];
    assign G[36] = in1[65] & in2[65];
    assign P[36] = in1[65] ^ in2[65];
    assign G[37] = in1[64] & in2[64];
    assign P[37] = in1[64] ^ in2[64];
    assign G[38] = in1[63] & in2[63];
    assign P[38] = in1[63] ^ in2[63];
    assign G[39] = in1[62] & in2[62];
    assign P[39] = in1[62] ^ in2[62];
    assign G[40] = in1[61] & in2[61];
    assign P[40] = in1[61] ^ in2[61];
    assign G[41] = in1[60] & in2[60];
    assign P[41] = in1[60] ^ in2[60];
    assign G[42] = in1[59] & in2[59];
    assign P[42] = in1[59] ^ in2[59];
    assign G[43] = in1[58] & in2[58];
    assign P[43] = in1[58] ^ in2[58];
    assign G[44] = in1[57] & in2[57];
    assign P[44] = in1[57] ^ in2[57];
    assign G[45] = in1[56] & in2[56];
    assign P[45] = in1[56] ^ in2[56];
    assign G[46] = in1[55] & in2[55];
    assign P[46] = in1[55] ^ in2[55];
    assign G[47] = in1[54] & in2[54];
    assign P[47] = in1[54] ^ in2[54];
    assign G[48] = in1[53] & in2[53];
    assign P[48] = in1[53] ^ in2[53];
    assign G[49] = in1[52] & in2[52];
    assign P[49] = in1[52] ^ in2[52];
    assign G[50] = in1[51] & in2[51];
    assign P[50] = in1[51] ^ in2[51];
    assign G[51] = in1[50] & in2[50];
    assign P[51] = in1[50] ^ in2[50];
    assign G[52] = in1[49] & in2[49];
    assign P[52] = in1[49] ^ in2[49];
    assign G[53] = in1[48] & in2[48];
    assign P[53] = in1[48] ^ in2[48];
    assign G[54] = in1[47] & in2[47];
    assign P[54] = in1[47] ^ in2[47];
    assign G[55] = in1[46] & in2[46];
    assign P[55] = in1[46] ^ in2[46];
    assign G[56] = in1[45] & in2[45];
    assign P[56] = in1[45] ^ in2[45];
    assign G[57] = in1[44] & in2[44];
    assign P[57] = in1[44] ^ in2[44];
    assign G[58] = in1[43] & in2[43];
    assign P[58] = in1[43] ^ in2[43];
    assign G[59] = in1[42] & in2[42];
    assign P[59] = in1[42] ^ in2[42];
    assign G[60] = in1[41] & in2[41];
    assign P[60] = in1[41] ^ in2[41];
    assign G[61] = in1[40] & in2[40];
    assign P[61] = in1[40] ^ in2[40];
    assign G[62] = in1[39] & in2[39];
    assign P[62] = in1[39] ^ in2[39];
    assign G[63] = in1[38] & in2[38];
    assign P[63] = in1[38] ^ in2[38];
    assign G[64] = in1[37] & in2[37];
    assign P[64] = in1[37] ^ in2[37];
    assign G[65] = in1[36] & in2[36];
    assign P[65] = in1[36] ^ in2[36];
    assign G[66] = in1[35] & in2[35];
    assign P[66] = in1[35] ^ in2[35];
    assign G[67] = in1[34] & in2[34];
    assign P[67] = in1[34] ^ in2[34];
    assign G[68] = in1[33] & in2[33];
    assign P[68] = in1[33] ^ in2[33];
    assign G[69] = in1[32] & in2[32];
    assign P[69] = in1[32] ^ in2[32];
    assign G[70] = in1[31] & in2[31];
    assign P[70] = in1[31] ^ in2[31];
    assign G[71] = in1[30] & in2[30];
    assign P[71] = in1[30] ^ in2[30];
    assign G[72] = in1[29] & in2[29];
    assign P[72] = in1[29] ^ in2[29];
    assign G[73] = in1[28] & in2[28];
    assign P[73] = in1[28] ^ in2[28];
    assign G[74] = in1[27] & in2[27];
    assign P[74] = in1[27] ^ in2[27];
    assign G[75] = in1[26] & in2[26];
    assign P[75] = in1[26] ^ in2[26];
    assign G[76] = in1[25] & in2[25];
    assign P[76] = in1[25] ^ in2[25];
    assign G[77] = in1[24] & in2[24];
    assign P[77] = in1[24] ^ in2[24];
    assign G[78] = in1[23] & in2[23];
    assign P[78] = in1[23] ^ in2[23];
    assign G[79] = in1[22] & in2[22];
    assign P[79] = in1[22] ^ in2[22];
    assign G[80] = in1[21] & in2[21];
    assign P[80] = in1[21] ^ in2[21];
    assign G[81] = in1[20] & in2[20];
    assign P[81] = in1[20] ^ in2[20];
    assign G[82] = in1[19] & in2[19];
    assign P[82] = in1[19] ^ in2[19];
    assign G[83] = in1[18] & in2[18];
    assign P[83] = in1[18] ^ in2[18];
    assign G[84] = in1[17] & in2[17];
    assign P[84] = in1[17] ^ in2[17];
    assign G[85] = in1[16] & in2[16];
    assign P[85] = in1[16] ^ in2[16];
    assign G[86] = in1[15] & in2[15];
    assign P[86] = in1[15] ^ in2[15];
    assign G[87] = in1[14] & in2[14];
    assign P[87] = in1[14] ^ in2[14];
    assign G[88] = in1[13] & in2[13];
    assign P[88] = in1[13] ^ in2[13];
    assign G[89] = in1[12] & in2[12];
    assign P[89] = in1[12] ^ in2[12];
    assign G[90] = in1[11] & in2[11];
    assign P[90] = in1[11] ^ in2[11];
    assign G[91] = in1[10] & in2[10];
    assign P[91] = in1[10] ^ in2[10];
    assign G[92] = in1[9] & in2[9];
    assign P[92] = in1[9] ^ in2[9];
    assign G[93] = in1[8] & in2[8];
    assign P[93] = in1[8] ^ in2[8];
    assign G[94] = in1[7] & in2[7];
    assign P[94] = in1[7] ^ in2[7];
    assign G[95] = in1[6] & in2[6];
    assign P[95] = in1[6] ^ in2[6];
    assign G[96] = in1[5] & in2[5];
    assign P[96] = in1[5] ^ in2[5];
    assign G[97] = in1[4] & in2[4];
    assign P[97] = in1[4] ^ in2[4];
    assign G[98] = in1[3] & in2[3];
    assign P[98] = in1[3] ^ in2[3];
    assign G[99] = in1[2] & in2[2];
    assign P[99] = in1[2] ^ in2[2];
    assign G[100] = in1[1] & in2[1];
    assign P[100] = in1[1] ^ in2[1];
    assign G[101] = in1[0] & in2[0];
    assign P[101] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign cout = G[101] | (P[101] & C[101]);
    assign sum = P ^ C;
endmodule

module CLA_101(output [100:0] sum, output cout, input [100:0] in1, input [100:0] in2);

    wire[100:0] G;
    wire[100:0] C;
    wire[100:0] P;

    assign G[0] = in1[100] & in2[100];
    assign P[0] = in1[100] ^ in2[100];
    assign G[1] = in1[99] & in2[99];
    assign P[1] = in1[99] ^ in2[99];
    assign G[2] = in1[98] & in2[98];
    assign P[2] = in1[98] ^ in2[98];
    assign G[3] = in1[97] & in2[97];
    assign P[3] = in1[97] ^ in2[97];
    assign G[4] = in1[96] & in2[96];
    assign P[4] = in1[96] ^ in2[96];
    assign G[5] = in1[95] & in2[95];
    assign P[5] = in1[95] ^ in2[95];
    assign G[6] = in1[94] & in2[94];
    assign P[6] = in1[94] ^ in2[94];
    assign G[7] = in1[93] & in2[93];
    assign P[7] = in1[93] ^ in2[93];
    assign G[8] = in1[92] & in2[92];
    assign P[8] = in1[92] ^ in2[92];
    assign G[9] = in1[91] & in2[91];
    assign P[9] = in1[91] ^ in2[91];
    assign G[10] = in1[90] & in2[90];
    assign P[10] = in1[90] ^ in2[90];
    assign G[11] = in1[89] & in2[89];
    assign P[11] = in1[89] ^ in2[89];
    assign G[12] = in1[88] & in2[88];
    assign P[12] = in1[88] ^ in2[88];
    assign G[13] = in1[87] & in2[87];
    assign P[13] = in1[87] ^ in2[87];
    assign G[14] = in1[86] & in2[86];
    assign P[14] = in1[86] ^ in2[86];
    assign G[15] = in1[85] & in2[85];
    assign P[15] = in1[85] ^ in2[85];
    assign G[16] = in1[84] & in2[84];
    assign P[16] = in1[84] ^ in2[84];
    assign G[17] = in1[83] & in2[83];
    assign P[17] = in1[83] ^ in2[83];
    assign G[18] = in1[82] & in2[82];
    assign P[18] = in1[82] ^ in2[82];
    assign G[19] = in1[81] & in2[81];
    assign P[19] = in1[81] ^ in2[81];
    assign G[20] = in1[80] & in2[80];
    assign P[20] = in1[80] ^ in2[80];
    assign G[21] = in1[79] & in2[79];
    assign P[21] = in1[79] ^ in2[79];
    assign G[22] = in1[78] & in2[78];
    assign P[22] = in1[78] ^ in2[78];
    assign G[23] = in1[77] & in2[77];
    assign P[23] = in1[77] ^ in2[77];
    assign G[24] = in1[76] & in2[76];
    assign P[24] = in1[76] ^ in2[76];
    assign G[25] = in1[75] & in2[75];
    assign P[25] = in1[75] ^ in2[75];
    assign G[26] = in1[74] & in2[74];
    assign P[26] = in1[74] ^ in2[74];
    assign G[27] = in1[73] & in2[73];
    assign P[27] = in1[73] ^ in2[73];
    assign G[28] = in1[72] & in2[72];
    assign P[28] = in1[72] ^ in2[72];
    assign G[29] = in1[71] & in2[71];
    assign P[29] = in1[71] ^ in2[71];
    assign G[30] = in1[70] & in2[70];
    assign P[30] = in1[70] ^ in2[70];
    assign G[31] = in1[69] & in2[69];
    assign P[31] = in1[69] ^ in2[69];
    assign G[32] = in1[68] & in2[68];
    assign P[32] = in1[68] ^ in2[68];
    assign G[33] = in1[67] & in2[67];
    assign P[33] = in1[67] ^ in2[67];
    assign G[34] = in1[66] & in2[66];
    assign P[34] = in1[66] ^ in2[66];
    assign G[35] = in1[65] & in2[65];
    assign P[35] = in1[65] ^ in2[65];
    assign G[36] = in1[64] & in2[64];
    assign P[36] = in1[64] ^ in2[64];
    assign G[37] = in1[63] & in2[63];
    assign P[37] = in1[63] ^ in2[63];
    assign G[38] = in1[62] & in2[62];
    assign P[38] = in1[62] ^ in2[62];
    assign G[39] = in1[61] & in2[61];
    assign P[39] = in1[61] ^ in2[61];
    assign G[40] = in1[60] & in2[60];
    assign P[40] = in1[60] ^ in2[60];
    assign G[41] = in1[59] & in2[59];
    assign P[41] = in1[59] ^ in2[59];
    assign G[42] = in1[58] & in2[58];
    assign P[42] = in1[58] ^ in2[58];
    assign G[43] = in1[57] & in2[57];
    assign P[43] = in1[57] ^ in2[57];
    assign G[44] = in1[56] & in2[56];
    assign P[44] = in1[56] ^ in2[56];
    assign G[45] = in1[55] & in2[55];
    assign P[45] = in1[55] ^ in2[55];
    assign G[46] = in1[54] & in2[54];
    assign P[46] = in1[54] ^ in2[54];
    assign G[47] = in1[53] & in2[53];
    assign P[47] = in1[53] ^ in2[53];
    assign G[48] = in1[52] & in2[52];
    assign P[48] = in1[52] ^ in2[52];
    assign G[49] = in1[51] & in2[51];
    assign P[49] = in1[51] ^ in2[51];
    assign G[50] = in1[50] & in2[50];
    assign P[50] = in1[50] ^ in2[50];
    assign G[51] = in1[49] & in2[49];
    assign P[51] = in1[49] ^ in2[49];
    assign G[52] = in1[48] & in2[48];
    assign P[52] = in1[48] ^ in2[48];
    assign G[53] = in1[47] & in2[47];
    assign P[53] = in1[47] ^ in2[47];
    assign G[54] = in1[46] & in2[46];
    assign P[54] = in1[46] ^ in2[46];
    assign G[55] = in1[45] & in2[45];
    assign P[55] = in1[45] ^ in2[45];
    assign G[56] = in1[44] & in2[44];
    assign P[56] = in1[44] ^ in2[44];
    assign G[57] = in1[43] & in2[43];
    assign P[57] = in1[43] ^ in2[43];
    assign G[58] = in1[42] & in2[42];
    assign P[58] = in1[42] ^ in2[42];
    assign G[59] = in1[41] & in2[41];
    assign P[59] = in1[41] ^ in2[41];
    assign G[60] = in1[40] & in2[40];
    assign P[60] = in1[40] ^ in2[40];
    assign G[61] = in1[39] & in2[39];
    assign P[61] = in1[39] ^ in2[39];
    assign G[62] = in1[38] & in2[38];
    assign P[62] = in1[38] ^ in2[38];
    assign G[63] = in1[37] & in2[37];
    assign P[63] = in1[37] ^ in2[37];
    assign G[64] = in1[36] & in2[36];
    assign P[64] = in1[36] ^ in2[36];
    assign G[65] = in1[35] & in2[35];
    assign P[65] = in1[35] ^ in2[35];
    assign G[66] = in1[34] & in2[34];
    assign P[66] = in1[34] ^ in2[34];
    assign G[67] = in1[33] & in2[33];
    assign P[67] = in1[33] ^ in2[33];
    assign G[68] = in1[32] & in2[32];
    assign P[68] = in1[32] ^ in2[32];
    assign G[69] = in1[31] & in2[31];
    assign P[69] = in1[31] ^ in2[31];
    assign G[70] = in1[30] & in2[30];
    assign P[70] = in1[30] ^ in2[30];
    assign G[71] = in1[29] & in2[29];
    assign P[71] = in1[29] ^ in2[29];
    assign G[72] = in1[28] & in2[28];
    assign P[72] = in1[28] ^ in2[28];
    assign G[73] = in1[27] & in2[27];
    assign P[73] = in1[27] ^ in2[27];
    assign G[74] = in1[26] & in2[26];
    assign P[74] = in1[26] ^ in2[26];
    assign G[75] = in1[25] & in2[25];
    assign P[75] = in1[25] ^ in2[25];
    assign G[76] = in1[24] & in2[24];
    assign P[76] = in1[24] ^ in2[24];
    assign G[77] = in1[23] & in2[23];
    assign P[77] = in1[23] ^ in2[23];
    assign G[78] = in1[22] & in2[22];
    assign P[78] = in1[22] ^ in2[22];
    assign G[79] = in1[21] & in2[21];
    assign P[79] = in1[21] ^ in2[21];
    assign G[80] = in1[20] & in2[20];
    assign P[80] = in1[20] ^ in2[20];
    assign G[81] = in1[19] & in2[19];
    assign P[81] = in1[19] ^ in2[19];
    assign G[82] = in1[18] & in2[18];
    assign P[82] = in1[18] ^ in2[18];
    assign G[83] = in1[17] & in2[17];
    assign P[83] = in1[17] ^ in2[17];
    assign G[84] = in1[16] & in2[16];
    assign P[84] = in1[16] ^ in2[16];
    assign G[85] = in1[15] & in2[15];
    assign P[85] = in1[15] ^ in2[15];
    assign G[86] = in1[14] & in2[14];
    assign P[86] = in1[14] ^ in2[14];
    assign G[87] = in1[13] & in2[13];
    assign P[87] = in1[13] ^ in2[13];
    assign G[88] = in1[12] & in2[12];
    assign P[88] = in1[12] ^ in2[12];
    assign G[89] = in1[11] & in2[11];
    assign P[89] = in1[11] ^ in2[11];
    assign G[90] = in1[10] & in2[10];
    assign P[90] = in1[10] ^ in2[10];
    assign G[91] = in1[9] & in2[9];
    assign P[91] = in1[9] ^ in2[9];
    assign G[92] = in1[8] & in2[8];
    assign P[92] = in1[8] ^ in2[8];
    assign G[93] = in1[7] & in2[7];
    assign P[93] = in1[7] ^ in2[7];
    assign G[94] = in1[6] & in2[6];
    assign P[94] = in1[6] ^ in2[6];
    assign G[95] = in1[5] & in2[5];
    assign P[95] = in1[5] ^ in2[5];
    assign G[96] = in1[4] & in2[4];
    assign P[96] = in1[4] ^ in2[4];
    assign G[97] = in1[3] & in2[3];
    assign P[97] = in1[3] ^ in2[3];
    assign G[98] = in1[2] & in2[2];
    assign P[98] = in1[2] ^ in2[2];
    assign G[99] = in1[1] & in2[1];
    assign P[99] = in1[1] ^ in2[1];
    assign G[100] = in1[0] & in2[0];
    assign P[100] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign cout = G[100] | (P[100] & C[100]);
    assign sum = P ^ C;
endmodule

module CLA_100(output [99:0] sum, output cout, input [99:0] in1, input [99:0] in2);

    wire[99:0] G;
    wire[99:0] C;
    wire[99:0] P;

    assign G[0] = in1[99] & in2[99];
    assign P[0] = in1[99] ^ in2[99];
    assign G[1] = in1[98] & in2[98];
    assign P[1] = in1[98] ^ in2[98];
    assign G[2] = in1[97] & in2[97];
    assign P[2] = in1[97] ^ in2[97];
    assign G[3] = in1[96] & in2[96];
    assign P[3] = in1[96] ^ in2[96];
    assign G[4] = in1[95] & in2[95];
    assign P[4] = in1[95] ^ in2[95];
    assign G[5] = in1[94] & in2[94];
    assign P[5] = in1[94] ^ in2[94];
    assign G[6] = in1[93] & in2[93];
    assign P[6] = in1[93] ^ in2[93];
    assign G[7] = in1[92] & in2[92];
    assign P[7] = in1[92] ^ in2[92];
    assign G[8] = in1[91] & in2[91];
    assign P[8] = in1[91] ^ in2[91];
    assign G[9] = in1[90] & in2[90];
    assign P[9] = in1[90] ^ in2[90];
    assign G[10] = in1[89] & in2[89];
    assign P[10] = in1[89] ^ in2[89];
    assign G[11] = in1[88] & in2[88];
    assign P[11] = in1[88] ^ in2[88];
    assign G[12] = in1[87] & in2[87];
    assign P[12] = in1[87] ^ in2[87];
    assign G[13] = in1[86] & in2[86];
    assign P[13] = in1[86] ^ in2[86];
    assign G[14] = in1[85] & in2[85];
    assign P[14] = in1[85] ^ in2[85];
    assign G[15] = in1[84] & in2[84];
    assign P[15] = in1[84] ^ in2[84];
    assign G[16] = in1[83] & in2[83];
    assign P[16] = in1[83] ^ in2[83];
    assign G[17] = in1[82] & in2[82];
    assign P[17] = in1[82] ^ in2[82];
    assign G[18] = in1[81] & in2[81];
    assign P[18] = in1[81] ^ in2[81];
    assign G[19] = in1[80] & in2[80];
    assign P[19] = in1[80] ^ in2[80];
    assign G[20] = in1[79] & in2[79];
    assign P[20] = in1[79] ^ in2[79];
    assign G[21] = in1[78] & in2[78];
    assign P[21] = in1[78] ^ in2[78];
    assign G[22] = in1[77] & in2[77];
    assign P[22] = in1[77] ^ in2[77];
    assign G[23] = in1[76] & in2[76];
    assign P[23] = in1[76] ^ in2[76];
    assign G[24] = in1[75] & in2[75];
    assign P[24] = in1[75] ^ in2[75];
    assign G[25] = in1[74] & in2[74];
    assign P[25] = in1[74] ^ in2[74];
    assign G[26] = in1[73] & in2[73];
    assign P[26] = in1[73] ^ in2[73];
    assign G[27] = in1[72] & in2[72];
    assign P[27] = in1[72] ^ in2[72];
    assign G[28] = in1[71] & in2[71];
    assign P[28] = in1[71] ^ in2[71];
    assign G[29] = in1[70] & in2[70];
    assign P[29] = in1[70] ^ in2[70];
    assign G[30] = in1[69] & in2[69];
    assign P[30] = in1[69] ^ in2[69];
    assign G[31] = in1[68] & in2[68];
    assign P[31] = in1[68] ^ in2[68];
    assign G[32] = in1[67] & in2[67];
    assign P[32] = in1[67] ^ in2[67];
    assign G[33] = in1[66] & in2[66];
    assign P[33] = in1[66] ^ in2[66];
    assign G[34] = in1[65] & in2[65];
    assign P[34] = in1[65] ^ in2[65];
    assign G[35] = in1[64] & in2[64];
    assign P[35] = in1[64] ^ in2[64];
    assign G[36] = in1[63] & in2[63];
    assign P[36] = in1[63] ^ in2[63];
    assign G[37] = in1[62] & in2[62];
    assign P[37] = in1[62] ^ in2[62];
    assign G[38] = in1[61] & in2[61];
    assign P[38] = in1[61] ^ in2[61];
    assign G[39] = in1[60] & in2[60];
    assign P[39] = in1[60] ^ in2[60];
    assign G[40] = in1[59] & in2[59];
    assign P[40] = in1[59] ^ in2[59];
    assign G[41] = in1[58] & in2[58];
    assign P[41] = in1[58] ^ in2[58];
    assign G[42] = in1[57] & in2[57];
    assign P[42] = in1[57] ^ in2[57];
    assign G[43] = in1[56] & in2[56];
    assign P[43] = in1[56] ^ in2[56];
    assign G[44] = in1[55] & in2[55];
    assign P[44] = in1[55] ^ in2[55];
    assign G[45] = in1[54] & in2[54];
    assign P[45] = in1[54] ^ in2[54];
    assign G[46] = in1[53] & in2[53];
    assign P[46] = in1[53] ^ in2[53];
    assign G[47] = in1[52] & in2[52];
    assign P[47] = in1[52] ^ in2[52];
    assign G[48] = in1[51] & in2[51];
    assign P[48] = in1[51] ^ in2[51];
    assign G[49] = in1[50] & in2[50];
    assign P[49] = in1[50] ^ in2[50];
    assign G[50] = in1[49] & in2[49];
    assign P[50] = in1[49] ^ in2[49];
    assign G[51] = in1[48] & in2[48];
    assign P[51] = in1[48] ^ in2[48];
    assign G[52] = in1[47] & in2[47];
    assign P[52] = in1[47] ^ in2[47];
    assign G[53] = in1[46] & in2[46];
    assign P[53] = in1[46] ^ in2[46];
    assign G[54] = in1[45] & in2[45];
    assign P[54] = in1[45] ^ in2[45];
    assign G[55] = in1[44] & in2[44];
    assign P[55] = in1[44] ^ in2[44];
    assign G[56] = in1[43] & in2[43];
    assign P[56] = in1[43] ^ in2[43];
    assign G[57] = in1[42] & in2[42];
    assign P[57] = in1[42] ^ in2[42];
    assign G[58] = in1[41] & in2[41];
    assign P[58] = in1[41] ^ in2[41];
    assign G[59] = in1[40] & in2[40];
    assign P[59] = in1[40] ^ in2[40];
    assign G[60] = in1[39] & in2[39];
    assign P[60] = in1[39] ^ in2[39];
    assign G[61] = in1[38] & in2[38];
    assign P[61] = in1[38] ^ in2[38];
    assign G[62] = in1[37] & in2[37];
    assign P[62] = in1[37] ^ in2[37];
    assign G[63] = in1[36] & in2[36];
    assign P[63] = in1[36] ^ in2[36];
    assign G[64] = in1[35] & in2[35];
    assign P[64] = in1[35] ^ in2[35];
    assign G[65] = in1[34] & in2[34];
    assign P[65] = in1[34] ^ in2[34];
    assign G[66] = in1[33] & in2[33];
    assign P[66] = in1[33] ^ in2[33];
    assign G[67] = in1[32] & in2[32];
    assign P[67] = in1[32] ^ in2[32];
    assign G[68] = in1[31] & in2[31];
    assign P[68] = in1[31] ^ in2[31];
    assign G[69] = in1[30] & in2[30];
    assign P[69] = in1[30] ^ in2[30];
    assign G[70] = in1[29] & in2[29];
    assign P[70] = in1[29] ^ in2[29];
    assign G[71] = in1[28] & in2[28];
    assign P[71] = in1[28] ^ in2[28];
    assign G[72] = in1[27] & in2[27];
    assign P[72] = in1[27] ^ in2[27];
    assign G[73] = in1[26] & in2[26];
    assign P[73] = in1[26] ^ in2[26];
    assign G[74] = in1[25] & in2[25];
    assign P[74] = in1[25] ^ in2[25];
    assign G[75] = in1[24] & in2[24];
    assign P[75] = in1[24] ^ in2[24];
    assign G[76] = in1[23] & in2[23];
    assign P[76] = in1[23] ^ in2[23];
    assign G[77] = in1[22] & in2[22];
    assign P[77] = in1[22] ^ in2[22];
    assign G[78] = in1[21] & in2[21];
    assign P[78] = in1[21] ^ in2[21];
    assign G[79] = in1[20] & in2[20];
    assign P[79] = in1[20] ^ in2[20];
    assign G[80] = in1[19] & in2[19];
    assign P[80] = in1[19] ^ in2[19];
    assign G[81] = in1[18] & in2[18];
    assign P[81] = in1[18] ^ in2[18];
    assign G[82] = in1[17] & in2[17];
    assign P[82] = in1[17] ^ in2[17];
    assign G[83] = in1[16] & in2[16];
    assign P[83] = in1[16] ^ in2[16];
    assign G[84] = in1[15] & in2[15];
    assign P[84] = in1[15] ^ in2[15];
    assign G[85] = in1[14] & in2[14];
    assign P[85] = in1[14] ^ in2[14];
    assign G[86] = in1[13] & in2[13];
    assign P[86] = in1[13] ^ in2[13];
    assign G[87] = in1[12] & in2[12];
    assign P[87] = in1[12] ^ in2[12];
    assign G[88] = in1[11] & in2[11];
    assign P[88] = in1[11] ^ in2[11];
    assign G[89] = in1[10] & in2[10];
    assign P[89] = in1[10] ^ in2[10];
    assign G[90] = in1[9] & in2[9];
    assign P[90] = in1[9] ^ in2[9];
    assign G[91] = in1[8] & in2[8];
    assign P[91] = in1[8] ^ in2[8];
    assign G[92] = in1[7] & in2[7];
    assign P[92] = in1[7] ^ in2[7];
    assign G[93] = in1[6] & in2[6];
    assign P[93] = in1[6] ^ in2[6];
    assign G[94] = in1[5] & in2[5];
    assign P[94] = in1[5] ^ in2[5];
    assign G[95] = in1[4] & in2[4];
    assign P[95] = in1[4] ^ in2[4];
    assign G[96] = in1[3] & in2[3];
    assign P[96] = in1[3] ^ in2[3];
    assign G[97] = in1[2] & in2[2];
    assign P[97] = in1[2] ^ in2[2];
    assign G[98] = in1[1] & in2[1];
    assign P[98] = in1[1] ^ in2[1];
    assign G[99] = in1[0] & in2[0];
    assign P[99] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign cout = G[99] | (P[99] & C[99]);
    assign sum = P ^ C;
endmodule

module CLA_99(output [98:0] sum, output cout, input [98:0] in1, input [98:0] in2);

    wire[98:0] G;
    wire[98:0] C;
    wire[98:0] P;

    assign G[0] = in1[98] & in2[98];
    assign P[0] = in1[98] ^ in2[98];
    assign G[1] = in1[97] & in2[97];
    assign P[1] = in1[97] ^ in2[97];
    assign G[2] = in1[96] & in2[96];
    assign P[2] = in1[96] ^ in2[96];
    assign G[3] = in1[95] & in2[95];
    assign P[3] = in1[95] ^ in2[95];
    assign G[4] = in1[94] & in2[94];
    assign P[4] = in1[94] ^ in2[94];
    assign G[5] = in1[93] & in2[93];
    assign P[5] = in1[93] ^ in2[93];
    assign G[6] = in1[92] & in2[92];
    assign P[6] = in1[92] ^ in2[92];
    assign G[7] = in1[91] & in2[91];
    assign P[7] = in1[91] ^ in2[91];
    assign G[8] = in1[90] & in2[90];
    assign P[8] = in1[90] ^ in2[90];
    assign G[9] = in1[89] & in2[89];
    assign P[9] = in1[89] ^ in2[89];
    assign G[10] = in1[88] & in2[88];
    assign P[10] = in1[88] ^ in2[88];
    assign G[11] = in1[87] & in2[87];
    assign P[11] = in1[87] ^ in2[87];
    assign G[12] = in1[86] & in2[86];
    assign P[12] = in1[86] ^ in2[86];
    assign G[13] = in1[85] & in2[85];
    assign P[13] = in1[85] ^ in2[85];
    assign G[14] = in1[84] & in2[84];
    assign P[14] = in1[84] ^ in2[84];
    assign G[15] = in1[83] & in2[83];
    assign P[15] = in1[83] ^ in2[83];
    assign G[16] = in1[82] & in2[82];
    assign P[16] = in1[82] ^ in2[82];
    assign G[17] = in1[81] & in2[81];
    assign P[17] = in1[81] ^ in2[81];
    assign G[18] = in1[80] & in2[80];
    assign P[18] = in1[80] ^ in2[80];
    assign G[19] = in1[79] & in2[79];
    assign P[19] = in1[79] ^ in2[79];
    assign G[20] = in1[78] & in2[78];
    assign P[20] = in1[78] ^ in2[78];
    assign G[21] = in1[77] & in2[77];
    assign P[21] = in1[77] ^ in2[77];
    assign G[22] = in1[76] & in2[76];
    assign P[22] = in1[76] ^ in2[76];
    assign G[23] = in1[75] & in2[75];
    assign P[23] = in1[75] ^ in2[75];
    assign G[24] = in1[74] & in2[74];
    assign P[24] = in1[74] ^ in2[74];
    assign G[25] = in1[73] & in2[73];
    assign P[25] = in1[73] ^ in2[73];
    assign G[26] = in1[72] & in2[72];
    assign P[26] = in1[72] ^ in2[72];
    assign G[27] = in1[71] & in2[71];
    assign P[27] = in1[71] ^ in2[71];
    assign G[28] = in1[70] & in2[70];
    assign P[28] = in1[70] ^ in2[70];
    assign G[29] = in1[69] & in2[69];
    assign P[29] = in1[69] ^ in2[69];
    assign G[30] = in1[68] & in2[68];
    assign P[30] = in1[68] ^ in2[68];
    assign G[31] = in1[67] & in2[67];
    assign P[31] = in1[67] ^ in2[67];
    assign G[32] = in1[66] & in2[66];
    assign P[32] = in1[66] ^ in2[66];
    assign G[33] = in1[65] & in2[65];
    assign P[33] = in1[65] ^ in2[65];
    assign G[34] = in1[64] & in2[64];
    assign P[34] = in1[64] ^ in2[64];
    assign G[35] = in1[63] & in2[63];
    assign P[35] = in1[63] ^ in2[63];
    assign G[36] = in1[62] & in2[62];
    assign P[36] = in1[62] ^ in2[62];
    assign G[37] = in1[61] & in2[61];
    assign P[37] = in1[61] ^ in2[61];
    assign G[38] = in1[60] & in2[60];
    assign P[38] = in1[60] ^ in2[60];
    assign G[39] = in1[59] & in2[59];
    assign P[39] = in1[59] ^ in2[59];
    assign G[40] = in1[58] & in2[58];
    assign P[40] = in1[58] ^ in2[58];
    assign G[41] = in1[57] & in2[57];
    assign P[41] = in1[57] ^ in2[57];
    assign G[42] = in1[56] & in2[56];
    assign P[42] = in1[56] ^ in2[56];
    assign G[43] = in1[55] & in2[55];
    assign P[43] = in1[55] ^ in2[55];
    assign G[44] = in1[54] & in2[54];
    assign P[44] = in1[54] ^ in2[54];
    assign G[45] = in1[53] & in2[53];
    assign P[45] = in1[53] ^ in2[53];
    assign G[46] = in1[52] & in2[52];
    assign P[46] = in1[52] ^ in2[52];
    assign G[47] = in1[51] & in2[51];
    assign P[47] = in1[51] ^ in2[51];
    assign G[48] = in1[50] & in2[50];
    assign P[48] = in1[50] ^ in2[50];
    assign G[49] = in1[49] & in2[49];
    assign P[49] = in1[49] ^ in2[49];
    assign G[50] = in1[48] & in2[48];
    assign P[50] = in1[48] ^ in2[48];
    assign G[51] = in1[47] & in2[47];
    assign P[51] = in1[47] ^ in2[47];
    assign G[52] = in1[46] & in2[46];
    assign P[52] = in1[46] ^ in2[46];
    assign G[53] = in1[45] & in2[45];
    assign P[53] = in1[45] ^ in2[45];
    assign G[54] = in1[44] & in2[44];
    assign P[54] = in1[44] ^ in2[44];
    assign G[55] = in1[43] & in2[43];
    assign P[55] = in1[43] ^ in2[43];
    assign G[56] = in1[42] & in2[42];
    assign P[56] = in1[42] ^ in2[42];
    assign G[57] = in1[41] & in2[41];
    assign P[57] = in1[41] ^ in2[41];
    assign G[58] = in1[40] & in2[40];
    assign P[58] = in1[40] ^ in2[40];
    assign G[59] = in1[39] & in2[39];
    assign P[59] = in1[39] ^ in2[39];
    assign G[60] = in1[38] & in2[38];
    assign P[60] = in1[38] ^ in2[38];
    assign G[61] = in1[37] & in2[37];
    assign P[61] = in1[37] ^ in2[37];
    assign G[62] = in1[36] & in2[36];
    assign P[62] = in1[36] ^ in2[36];
    assign G[63] = in1[35] & in2[35];
    assign P[63] = in1[35] ^ in2[35];
    assign G[64] = in1[34] & in2[34];
    assign P[64] = in1[34] ^ in2[34];
    assign G[65] = in1[33] & in2[33];
    assign P[65] = in1[33] ^ in2[33];
    assign G[66] = in1[32] & in2[32];
    assign P[66] = in1[32] ^ in2[32];
    assign G[67] = in1[31] & in2[31];
    assign P[67] = in1[31] ^ in2[31];
    assign G[68] = in1[30] & in2[30];
    assign P[68] = in1[30] ^ in2[30];
    assign G[69] = in1[29] & in2[29];
    assign P[69] = in1[29] ^ in2[29];
    assign G[70] = in1[28] & in2[28];
    assign P[70] = in1[28] ^ in2[28];
    assign G[71] = in1[27] & in2[27];
    assign P[71] = in1[27] ^ in2[27];
    assign G[72] = in1[26] & in2[26];
    assign P[72] = in1[26] ^ in2[26];
    assign G[73] = in1[25] & in2[25];
    assign P[73] = in1[25] ^ in2[25];
    assign G[74] = in1[24] & in2[24];
    assign P[74] = in1[24] ^ in2[24];
    assign G[75] = in1[23] & in2[23];
    assign P[75] = in1[23] ^ in2[23];
    assign G[76] = in1[22] & in2[22];
    assign P[76] = in1[22] ^ in2[22];
    assign G[77] = in1[21] & in2[21];
    assign P[77] = in1[21] ^ in2[21];
    assign G[78] = in1[20] & in2[20];
    assign P[78] = in1[20] ^ in2[20];
    assign G[79] = in1[19] & in2[19];
    assign P[79] = in1[19] ^ in2[19];
    assign G[80] = in1[18] & in2[18];
    assign P[80] = in1[18] ^ in2[18];
    assign G[81] = in1[17] & in2[17];
    assign P[81] = in1[17] ^ in2[17];
    assign G[82] = in1[16] & in2[16];
    assign P[82] = in1[16] ^ in2[16];
    assign G[83] = in1[15] & in2[15];
    assign P[83] = in1[15] ^ in2[15];
    assign G[84] = in1[14] & in2[14];
    assign P[84] = in1[14] ^ in2[14];
    assign G[85] = in1[13] & in2[13];
    assign P[85] = in1[13] ^ in2[13];
    assign G[86] = in1[12] & in2[12];
    assign P[86] = in1[12] ^ in2[12];
    assign G[87] = in1[11] & in2[11];
    assign P[87] = in1[11] ^ in2[11];
    assign G[88] = in1[10] & in2[10];
    assign P[88] = in1[10] ^ in2[10];
    assign G[89] = in1[9] & in2[9];
    assign P[89] = in1[9] ^ in2[9];
    assign G[90] = in1[8] & in2[8];
    assign P[90] = in1[8] ^ in2[8];
    assign G[91] = in1[7] & in2[7];
    assign P[91] = in1[7] ^ in2[7];
    assign G[92] = in1[6] & in2[6];
    assign P[92] = in1[6] ^ in2[6];
    assign G[93] = in1[5] & in2[5];
    assign P[93] = in1[5] ^ in2[5];
    assign G[94] = in1[4] & in2[4];
    assign P[94] = in1[4] ^ in2[4];
    assign G[95] = in1[3] & in2[3];
    assign P[95] = in1[3] ^ in2[3];
    assign G[96] = in1[2] & in2[2];
    assign P[96] = in1[2] ^ in2[2];
    assign G[97] = in1[1] & in2[1];
    assign P[97] = in1[1] ^ in2[1];
    assign G[98] = in1[0] & in2[0];
    assign P[98] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign cout = G[98] | (P[98] & C[98]);
    assign sum = P ^ C;
endmodule

module CLA_98(output [97:0] sum, output cout, input [97:0] in1, input [97:0] in2);

    wire[97:0] G;
    wire[97:0] C;
    wire[97:0] P;

    assign G[0] = in1[97] & in2[97];
    assign P[0] = in1[97] ^ in2[97];
    assign G[1] = in1[96] & in2[96];
    assign P[1] = in1[96] ^ in2[96];
    assign G[2] = in1[95] & in2[95];
    assign P[2] = in1[95] ^ in2[95];
    assign G[3] = in1[94] & in2[94];
    assign P[3] = in1[94] ^ in2[94];
    assign G[4] = in1[93] & in2[93];
    assign P[4] = in1[93] ^ in2[93];
    assign G[5] = in1[92] & in2[92];
    assign P[5] = in1[92] ^ in2[92];
    assign G[6] = in1[91] & in2[91];
    assign P[6] = in1[91] ^ in2[91];
    assign G[7] = in1[90] & in2[90];
    assign P[7] = in1[90] ^ in2[90];
    assign G[8] = in1[89] & in2[89];
    assign P[8] = in1[89] ^ in2[89];
    assign G[9] = in1[88] & in2[88];
    assign P[9] = in1[88] ^ in2[88];
    assign G[10] = in1[87] & in2[87];
    assign P[10] = in1[87] ^ in2[87];
    assign G[11] = in1[86] & in2[86];
    assign P[11] = in1[86] ^ in2[86];
    assign G[12] = in1[85] & in2[85];
    assign P[12] = in1[85] ^ in2[85];
    assign G[13] = in1[84] & in2[84];
    assign P[13] = in1[84] ^ in2[84];
    assign G[14] = in1[83] & in2[83];
    assign P[14] = in1[83] ^ in2[83];
    assign G[15] = in1[82] & in2[82];
    assign P[15] = in1[82] ^ in2[82];
    assign G[16] = in1[81] & in2[81];
    assign P[16] = in1[81] ^ in2[81];
    assign G[17] = in1[80] & in2[80];
    assign P[17] = in1[80] ^ in2[80];
    assign G[18] = in1[79] & in2[79];
    assign P[18] = in1[79] ^ in2[79];
    assign G[19] = in1[78] & in2[78];
    assign P[19] = in1[78] ^ in2[78];
    assign G[20] = in1[77] & in2[77];
    assign P[20] = in1[77] ^ in2[77];
    assign G[21] = in1[76] & in2[76];
    assign P[21] = in1[76] ^ in2[76];
    assign G[22] = in1[75] & in2[75];
    assign P[22] = in1[75] ^ in2[75];
    assign G[23] = in1[74] & in2[74];
    assign P[23] = in1[74] ^ in2[74];
    assign G[24] = in1[73] & in2[73];
    assign P[24] = in1[73] ^ in2[73];
    assign G[25] = in1[72] & in2[72];
    assign P[25] = in1[72] ^ in2[72];
    assign G[26] = in1[71] & in2[71];
    assign P[26] = in1[71] ^ in2[71];
    assign G[27] = in1[70] & in2[70];
    assign P[27] = in1[70] ^ in2[70];
    assign G[28] = in1[69] & in2[69];
    assign P[28] = in1[69] ^ in2[69];
    assign G[29] = in1[68] & in2[68];
    assign P[29] = in1[68] ^ in2[68];
    assign G[30] = in1[67] & in2[67];
    assign P[30] = in1[67] ^ in2[67];
    assign G[31] = in1[66] & in2[66];
    assign P[31] = in1[66] ^ in2[66];
    assign G[32] = in1[65] & in2[65];
    assign P[32] = in1[65] ^ in2[65];
    assign G[33] = in1[64] & in2[64];
    assign P[33] = in1[64] ^ in2[64];
    assign G[34] = in1[63] & in2[63];
    assign P[34] = in1[63] ^ in2[63];
    assign G[35] = in1[62] & in2[62];
    assign P[35] = in1[62] ^ in2[62];
    assign G[36] = in1[61] & in2[61];
    assign P[36] = in1[61] ^ in2[61];
    assign G[37] = in1[60] & in2[60];
    assign P[37] = in1[60] ^ in2[60];
    assign G[38] = in1[59] & in2[59];
    assign P[38] = in1[59] ^ in2[59];
    assign G[39] = in1[58] & in2[58];
    assign P[39] = in1[58] ^ in2[58];
    assign G[40] = in1[57] & in2[57];
    assign P[40] = in1[57] ^ in2[57];
    assign G[41] = in1[56] & in2[56];
    assign P[41] = in1[56] ^ in2[56];
    assign G[42] = in1[55] & in2[55];
    assign P[42] = in1[55] ^ in2[55];
    assign G[43] = in1[54] & in2[54];
    assign P[43] = in1[54] ^ in2[54];
    assign G[44] = in1[53] & in2[53];
    assign P[44] = in1[53] ^ in2[53];
    assign G[45] = in1[52] & in2[52];
    assign P[45] = in1[52] ^ in2[52];
    assign G[46] = in1[51] & in2[51];
    assign P[46] = in1[51] ^ in2[51];
    assign G[47] = in1[50] & in2[50];
    assign P[47] = in1[50] ^ in2[50];
    assign G[48] = in1[49] & in2[49];
    assign P[48] = in1[49] ^ in2[49];
    assign G[49] = in1[48] & in2[48];
    assign P[49] = in1[48] ^ in2[48];
    assign G[50] = in1[47] & in2[47];
    assign P[50] = in1[47] ^ in2[47];
    assign G[51] = in1[46] & in2[46];
    assign P[51] = in1[46] ^ in2[46];
    assign G[52] = in1[45] & in2[45];
    assign P[52] = in1[45] ^ in2[45];
    assign G[53] = in1[44] & in2[44];
    assign P[53] = in1[44] ^ in2[44];
    assign G[54] = in1[43] & in2[43];
    assign P[54] = in1[43] ^ in2[43];
    assign G[55] = in1[42] & in2[42];
    assign P[55] = in1[42] ^ in2[42];
    assign G[56] = in1[41] & in2[41];
    assign P[56] = in1[41] ^ in2[41];
    assign G[57] = in1[40] & in2[40];
    assign P[57] = in1[40] ^ in2[40];
    assign G[58] = in1[39] & in2[39];
    assign P[58] = in1[39] ^ in2[39];
    assign G[59] = in1[38] & in2[38];
    assign P[59] = in1[38] ^ in2[38];
    assign G[60] = in1[37] & in2[37];
    assign P[60] = in1[37] ^ in2[37];
    assign G[61] = in1[36] & in2[36];
    assign P[61] = in1[36] ^ in2[36];
    assign G[62] = in1[35] & in2[35];
    assign P[62] = in1[35] ^ in2[35];
    assign G[63] = in1[34] & in2[34];
    assign P[63] = in1[34] ^ in2[34];
    assign G[64] = in1[33] & in2[33];
    assign P[64] = in1[33] ^ in2[33];
    assign G[65] = in1[32] & in2[32];
    assign P[65] = in1[32] ^ in2[32];
    assign G[66] = in1[31] & in2[31];
    assign P[66] = in1[31] ^ in2[31];
    assign G[67] = in1[30] & in2[30];
    assign P[67] = in1[30] ^ in2[30];
    assign G[68] = in1[29] & in2[29];
    assign P[68] = in1[29] ^ in2[29];
    assign G[69] = in1[28] & in2[28];
    assign P[69] = in1[28] ^ in2[28];
    assign G[70] = in1[27] & in2[27];
    assign P[70] = in1[27] ^ in2[27];
    assign G[71] = in1[26] & in2[26];
    assign P[71] = in1[26] ^ in2[26];
    assign G[72] = in1[25] & in2[25];
    assign P[72] = in1[25] ^ in2[25];
    assign G[73] = in1[24] & in2[24];
    assign P[73] = in1[24] ^ in2[24];
    assign G[74] = in1[23] & in2[23];
    assign P[74] = in1[23] ^ in2[23];
    assign G[75] = in1[22] & in2[22];
    assign P[75] = in1[22] ^ in2[22];
    assign G[76] = in1[21] & in2[21];
    assign P[76] = in1[21] ^ in2[21];
    assign G[77] = in1[20] & in2[20];
    assign P[77] = in1[20] ^ in2[20];
    assign G[78] = in1[19] & in2[19];
    assign P[78] = in1[19] ^ in2[19];
    assign G[79] = in1[18] & in2[18];
    assign P[79] = in1[18] ^ in2[18];
    assign G[80] = in1[17] & in2[17];
    assign P[80] = in1[17] ^ in2[17];
    assign G[81] = in1[16] & in2[16];
    assign P[81] = in1[16] ^ in2[16];
    assign G[82] = in1[15] & in2[15];
    assign P[82] = in1[15] ^ in2[15];
    assign G[83] = in1[14] & in2[14];
    assign P[83] = in1[14] ^ in2[14];
    assign G[84] = in1[13] & in2[13];
    assign P[84] = in1[13] ^ in2[13];
    assign G[85] = in1[12] & in2[12];
    assign P[85] = in1[12] ^ in2[12];
    assign G[86] = in1[11] & in2[11];
    assign P[86] = in1[11] ^ in2[11];
    assign G[87] = in1[10] & in2[10];
    assign P[87] = in1[10] ^ in2[10];
    assign G[88] = in1[9] & in2[9];
    assign P[88] = in1[9] ^ in2[9];
    assign G[89] = in1[8] & in2[8];
    assign P[89] = in1[8] ^ in2[8];
    assign G[90] = in1[7] & in2[7];
    assign P[90] = in1[7] ^ in2[7];
    assign G[91] = in1[6] & in2[6];
    assign P[91] = in1[6] ^ in2[6];
    assign G[92] = in1[5] & in2[5];
    assign P[92] = in1[5] ^ in2[5];
    assign G[93] = in1[4] & in2[4];
    assign P[93] = in1[4] ^ in2[4];
    assign G[94] = in1[3] & in2[3];
    assign P[94] = in1[3] ^ in2[3];
    assign G[95] = in1[2] & in2[2];
    assign P[95] = in1[2] ^ in2[2];
    assign G[96] = in1[1] & in2[1];
    assign P[96] = in1[1] ^ in2[1];
    assign G[97] = in1[0] & in2[0];
    assign P[97] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign cout = G[97] | (P[97] & C[97]);
    assign sum = P ^ C;
endmodule

module CLA_97(output [96:0] sum, output cout, input [96:0] in1, input [96:0] in2);

    wire[96:0] G;
    wire[96:0] C;
    wire[96:0] P;

    assign G[0] = in1[96] & in2[96];
    assign P[0] = in1[96] ^ in2[96];
    assign G[1] = in1[95] & in2[95];
    assign P[1] = in1[95] ^ in2[95];
    assign G[2] = in1[94] & in2[94];
    assign P[2] = in1[94] ^ in2[94];
    assign G[3] = in1[93] & in2[93];
    assign P[3] = in1[93] ^ in2[93];
    assign G[4] = in1[92] & in2[92];
    assign P[4] = in1[92] ^ in2[92];
    assign G[5] = in1[91] & in2[91];
    assign P[5] = in1[91] ^ in2[91];
    assign G[6] = in1[90] & in2[90];
    assign P[6] = in1[90] ^ in2[90];
    assign G[7] = in1[89] & in2[89];
    assign P[7] = in1[89] ^ in2[89];
    assign G[8] = in1[88] & in2[88];
    assign P[8] = in1[88] ^ in2[88];
    assign G[9] = in1[87] & in2[87];
    assign P[9] = in1[87] ^ in2[87];
    assign G[10] = in1[86] & in2[86];
    assign P[10] = in1[86] ^ in2[86];
    assign G[11] = in1[85] & in2[85];
    assign P[11] = in1[85] ^ in2[85];
    assign G[12] = in1[84] & in2[84];
    assign P[12] = in1[84] ^ in2[84];
    assign G[13] = in1[83] & in2[83];
    assign P[13] = in1[83] ^ in2[83];
    assign G[14] = in1[82] & in2[82];
    assign P[14] = in1[82] ^ in2[82];
    assign G[15] = in1[81] & in2[81];
    assign P[15] = in1[81] ^ in2[81];
    assign G[16] = in1[80] & in2[80];
    assign P[16] = in1[80] ^ in2[80];
    assign G[17] = in1[79] & in2[79];
    assign P[17] = in1[79] ^ in2[79];
    assign G[18] = in1[78] & in2[78];
    assign P[18] = in1[78] ^ in2[78];
    assign G[19] = in1[77] & in2[77];
    assign P[19] = in1[77] ^ in2[77];
    assign G[20] = in1[76] & in2[76];
    assign P[20] = in1[76] ^ in2[76];
    assign G[21] = in1[75] & in2[75];
    assign P[21] = in1[75] ^ in2[75];
    assign G[22] = in1[74] & in2[74];
    assign P[22] = in1[74] ^ in2[74];
    assign G[23] = in1[73] & in2[73];
    assign P[23] = in1[73] ^ in2[73];
    assign G[24] = in1[72] & in2[72];
    assign P[24] = in1[72] ^ in2[72];
    assign G[25] = in1[71] & in2[71];
    assign P[25] = in1[71] ^ in2[71];
    assign G[26] = in1[70] & in2[70];
    assign P[26] = in1[70] ^ in2[70];
    assign G[27] = in1[69] & in2[69];
    assign P[27] = in1[69] ^ in2[69];
    assign G[28] = in1[68] & in2[68];
    assign P[28] = in1[68] ^ in2[68];
    assign G[29] = in1[67] & in2[67];
    assign P[29] = in1[67] ^ in2[67];
    assign G[30] = in1[66] & in2[66];
    assign P[30] = in1[66] ^ in2[66];
    assign G[31] = in1[65] & in2[65];
    assign P[31] = in1[65] ^ in2[65];
    assign G[32] = in1[64] & in2[64];
    assign P[32] = in1[64] ^ in2[64];
    assign G[33] = in1[63] & in2[63];
    assign P[33] = in1[63] ^ in2[63];
    assign G[34] = in1[62] & in2[62];
    assign P[34] = in1[62] ^ in2[62];
    assign G[35] = in1[61] & in2[61];
    assign P[35] = in1[61] ^ in2[61];
    assign G[36] = in1[60] & in2[60];
    assign P[36] = in1[60] ^ in2[60];
    assign G[37] = in1[59] & in2[59];
    assign P[37] = in1[59] ^ in2[59];
    assign G[38] = in1[58] & in2[58];
    assign P[38] = in1[58] ^ in2[58];
    assign G[39] = in1[57] & in2[57];
    assign P[39] = in1[57] ^ in2[57];
    assign G[40] = in1[56] & in2[56];
    assign P[40] = in1[56] ^ in2[56];
    assign G[41] = in1[55] & in2[55];
    assign P[41] = in1[55] ^ in2[55];
    assign G[42] = in1[54] & in2[54];
    assign P[42] = in1[54] ^ in2[54];
    assign G[43] = in1[53] & in2[53];
    assign P[43] = in1[53] ^ in2[53];
    assign G[44] = in1[52] & in2[52];
    assign P[44] = in1[52] ^ in2[52];
    assign G[45] = in1[51] & in2[51];
    assign P[45] = in1[51] ^ in2[51];
    assign G[46] = in1[50] & in2[50];
    assign P[46] = in1[50] ^ in2[50];
    assign G[47] = in1[49] & in2[49];
    assign P[47] = in1[49] ^ in2[49];
    assign G[48] = in1[48] & in2[48];
    assign P[48] = in1[48] ^ in2[48];
    assign G[49] = in1[47] & in2[47];
    assign P[49] = in1[47] ^ in2[47];
    assign G[50] = in1[46] & in2[46];
    assign P[50] = in1[46] ^ in2[46];
    assign G[51] = in1[45] & in2[45];
    assign P[51] = in1[45] ^ in2[45];
    assign G[52] = in1[44] & in2[44];
    assign P[52] = in1[44] ^ in2[44];
    assign G[53] = in1[43] & in2[43];
    assign P[53] = in1[43] ^ in2[43];
    assign G[54] = in1[42] & in2[42];
    assign P[54] = in1[42] ^ in2[42];
    assign G[55] = in1[41] & in2[41];
    assign P[55] = in1[41] ^ in2[41];
    assign G[56] = in1[40] & in2[40];
    assign P[56] = in1[40] ^ in2[40];
    assign G[57] = in1[39] & in2[39];
    assign P[57] = in1[39] ^ in2[39];
    assign G[58] = in1[38] & in2[38];
    assign P[58] = in1[38] ^ in2[38];
    assign G[59] = in1[37] & in2[37];
    assign P[59] = in1[37] ^ in2[37];
    assign G[60] = in1[36] & in2[36];
    assign P[60] = in1[36] ^ in2[36];
    assign G[61] = in1[35] & in2[35];
    assign P[61] = in1[35] ^ in2[35];
    assign G[62] = in1[34] & in2[34];
    assign P[62] = in1[34] ^ in2[34];
    assign G[63] = in1[33] & in2[33];
    assign P[63] = in1[33] ^ in2[33];
    assign G[64] = in1[32] & in2[32];
    assign P[64] = in1[32] ^ in2[32];
    assign G[65] = in1[31] & in2[31];
    assign P[65] = in1[31] ^ in2[31];
    assign G[66] = in1[30] & in2[30];
    assign P[66] = in1[30] ^ in2[30];
    assign G[67] = in1[29] & in2[29];
    assign P[67] = in1[29] ^ in2[29];
    assign G[68] = in1[28] & in2[28];
    assign P[68] = in1[28] ^ in2[28];
    assign G[69] = in1[27] & in2[27];
    assign P[69] = in1[27] ^ in2[27];
    assign G[70] = in1[26] & in2[26];
    assign P[70] = in1[26] ^ in2[26];
    assign G[71] = in1[25] & in2[25];
    assign P[71] = in1[25] ^ in2[25];
    assign G[72] = in1[24] & in2[24];
    assign P[72] = in1[24] ^ in2[24];
    assign G[73] = in1[23] & in2[23];
    assign P[73] = in1[23] ^ in2[23];
    assign G[74] = in1[22] & in2[22];
    assign P[74] = in1[22] ^ in2[22];
    assign G[75] = in1[21] & in2[21];
    assign P[75] = in1[21] ^ in2[21];
    assign G[76] = in1[20] & in2[20];
    assign P[76] = in1[20] ^ in2[20];
    assign G[77] = in1[19] & in2[19];
    assign P[77] = in1[19] ^ in2[19];
    assign G[78] = in1[18] & in2[18];
    assign P[78] = in1[18] ^ in2[18];
    assign G[79] = in1[17] & in2[17];
    assign P[79] = in1[17] ^ in2[17];
    assign G[80] = in1[16] & in2[16];
    assign P[80] = in1[16] ^ in2[16];
    assign G[81] = in1[15] & in2[15];
    assign P[81] = in1[15] ^ in2[15];
    assign G[82] = in1[14] & in2[14];
    assign P[82] = in1[14] ^ in2[14];
    assign G[83] = in1[13] & in2[13];
    assign P[83] = in1[13] ^ in2[13];
    assign G[84] = in1[12] & in2[12];
    assign P[84] = in1[12] ^ in2[12];
    assign G[85] = in1[11] & in2[11];
    assign P[85] = in1[11] ^ in2[11];
    assign G[86] = in1[10] & in2[10];
    assign P[86] = in1[10] ^ in2[10];
    assign G[87] = in1[9] & in2[9];
    assign P[87] = in1[9] ^ in2[9];
    assign G[88] = in1[8] & in2[8];
    assign P[88] = in1[8] ^ in2[8];
    assign G[89] = in1[7] & in2[7];
    assign P[89] = in1[7] ^ in2[7];
    assign G[90] = in1[6] & in2[6];
    assign P[90] = in1[6] ^ in2[6];
    assign G[91] = in1[5] & in2[5];
    assign P[91] = in1[5] ^ in2[5];
    assign G[92] = in1[4] & in2[4];
    assign P[92] = in1[4] ^ in2[4];
    assign G[93] = in1[3] & in2[3];
    assign P[93] = in1[3] ^ in2[3];
    assign G[94] = in1[2] & in2[2];
    assign P[94] = in1[2] ^ in2[2];
    assign G[95] = in1[1] & in2[1];
    assign P[95] = in1[1] ^ in2[1];
    assign G[96] = in1[0] & in2[0];
    assign P[96] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign cout = G[96] | (P[96] & C[96]);
    assign sum = P ^ C;
endmodule

module CLA_96(output [95:0] sum, output cout, input [95:0] in1, input [95:0] in2);

    wire[95:0] G;
    wire[95:0] C;
    wire[95:0] P;

    assign G[0] = in1[95] & in2[95];
    assign P[0] = in1[95] ^ in2[95];
    assign G[1] = in1[94] & in2[94];
    assign P[1] = in1[94] ^ in2[94];
    assign G[2] = in1[93] & in2[93];
    assign P[2] = in1[93] ^ in2[93];
    assign G[3] = in1[92] & in2[92];
    assign P[3] = in1[92] ^ in2[92];
    assign G[4] = in1[91] & in2[91];
    assign P[4] = in1[91] ^ in2[91];
    assign G[5] = in1[90] & in2[90];
    assign P[5] = in1[90] ^ in2[90];
    assign G[6] = in1[89] & in2[89];
    assign P[6] = in1[89] ^ in2[89];
    assign G[7] = in1[88] & in2[88];
    assign P[7] = in1[88] ^ in2[88];
    assign G[8] = in1[87] & in2[87];
    assign P[8] = in1[87] ^ in2[87];
    assign G[9] = in1[86] & in2[86];
    assign P[9] = in1[86] ^ in2[86];
    assign G[10] = in1[85] & in2[85];
    assign P[10] = in1[85] ^ in2[85];
    assign G[11] = in1[84] & in2[84];
    assign P[11] = in1[84] ^ in2[84];
    assign G[12] = in1[83] & in2[83];
    assign P[12] = in1[83] ^ in2[83];
    assign G[13] = in1[82] & in2[82];
    assign P[13] = in1[82] ^ in2[82];
    assign G[14] = in1[81] & in2[81];
    assign P[14] = in1[81] ^ in2[81];
    assign G[15] = in1[80] & in2[80];
    assign P[15] = in1[80] ^ in2[80];
    assign G[16] = in1[79] & in2[79];
    assign P[16] = in1[79] ^ in2[79];
    assign G[17] = in1[78] & in2[78];
    assign P[17] = in1[78] ^ in2[78];
    assign G[18] = in1[77] & in2[77];
    assign P[18] = in1[77] ^ in2[77];
    assign G[19] = in1[76] & in2[76];
    assign P[19] = in1[76] ^ in2[76];
    assign G[20] = in1[75] & in2[75];
    assign P[20] = in1[75] ^ in2[75];
    assign G[21] = in1[74] & in2[74];
    assign P[21] = in1[74] ^ in2[74];
    assign G[22] = in1[73] & in2[73];
    assign P[22] = in1[73] ^ in2[73];
    assign G[23] = in1[72] & in2[72];
    assign P[23] = in1[72] ^ in2[72];
    assign G[24] = in1[71] & in2[71];
    assign P[24] = in1[71] ^ in2[71];
    assign G[25] = in1[70] & in2[70];
    assign P[25] = in1[70] ^ in2[70];
    assign G[26] = in1[69] & in2[69];
    assign P[26] = in1[69] ^ in2[69];
    assign G[27] = in1[68] & in2[68];
    assign P[27] = in1[68] ^ in2[68];
    assign G[28] = in1[67] & in2[67];
    assign P[28] = in1[67] ^ in2[67];
    assign G[29] = in1[66] & in2[66];
    assign P[29] = in1[66] ^ in2[66];
    assign G[30] = in1[65] & in2[65];
    assign P[30] = in1[65] ^ in2[65];
    assign G[31] = in1[64] & in2[64];
    assign P[31] = in1[64] ^ in2[64];
    assign G[32] = in1[63] & in2[63];
    assign P[32] = in1[63] ^ in2[63];
    assign G[33] = in1[62] & in2[62];
    assign P[33] = in1[62] ^ in2[62];
    assign G[34] = in1[61] & in2[61];
    assign P[34] = in1[61] ^ in2[61];
    assign G[35] = in1[60] & in2[60];
    assign P[35] = in1[60] ^ in2[60];
    assign G[36] = in1[59] & in2[59];
    assign P[36] = in1[59] ^ in2[59];
    assign G[37] = in1[58] & in2[58];
    assign P[37] = in1[58] ^ in2[58];
    assign G[38] = in1[57] & in2[57];
    assign P[38] = in1[57] ^ in2[57];
    assign G[39] = in1[56] & in2[56];
    assign P[39] = in1[56] ^ in2[56];
    assign G[40] = in1[55] & in2[55];
    assign P[40] = in1[55] ^ in2[55];
    assign G[41] = in1[54] & in2[54];
    assign P[41] = in1[54] ^ in2[54];
    assign G[42] = in1[53] & in2[53];
    assign P[42] = in1[53] ^ in2[53];
    assign G[43] = in1[52] & in2[52];
    assign P[43] = in1[52] ^ in2[52];
    assign G[44] = in1[51] & in2[51];
    assign P[44] = in1[51] ^ in2[51];
    assign G[45] = in1[50] & in2[50];
    assign P[45] = in1[50] ^ in2[50];
    assign G[46] = in1[49] & in2[49];
    assign P[46] = in1[49] ^ in2[49];
    assign G[47] = in1[48] & in2[48];
    assign P[47] = in1[48] ^ in2[48];
    assign G[48] = in1[47] & in2[47];
    assign P[48] = in1[47] ^ in2[47];
    assign G[49] = in1[46] & in2[46];
    assign P[49] = in1[46] ^ in2[46];
    assign G[50] = in1[45] & in2[45];
    assign P[50] = in1[45] ^ in2[45];
    assign G[51] = in1[44] & in2[44];
    assign P[51] = in1[44] ^ in2[44];
    assign G[52] = in1[43] & in2[43];
    assign P[52] = in1[43] ^ in2[43];
    assign G[53] = in1[42] & in2[42];
    assign P[53] = in1[42] ^ in2[42];
    assign G[54] = in1[41] & in2[41];
    assign P[54] = in1[41] ^ in2[41];
    assign G[55] = in1[40] & in2[40];
    assign P[55] = in1[40] ^ in2[40];
    assign G[56] = in1[39] & in2[39];
    assign P[56] = in1[39] ^ in2[39];
    assign G[57] = in1[38] & in2[38];
    assign P[57] = in1[38] ^ in2[38];
    assign G[58] = in1[37] & in2[37];
    assign P[58] = in1[37] ^ in2[37];
    assign G[59] = in1[36] & in2[36];
    assign P[59] = in1[36] ^ in2[36];
    assign G[60] = in1[35] & in2[35];
    assign P[60] = in1[35] ^ in2[35];
    assign G[61] = in1[34] & in2[34];
    assign P[61] = in1[34] ^ in2[34];
    assign G[62] = in1[33] & in2[33];
    assign P[62] = in1[33] ^ in2[33];
    assign G[63] = in1[32] & in2[32];
    assign P[63] = in1[32] ^ in2[32];
    assign G[64] = in1[31] & in2[31];
    assign P[64] = in1[31] ^ in2[31];
    assign G[65] = in1[30] & in2[30];
    assign P[65] = in1[30] ^ in2[30];
    assign G[66] = in1[29] & in2[29];
    assign P[66] = in1[29] ^ in2[29];
    assign G[67] = in1[28] & in2[28];
    assign P[67] = in1[28] ^ in2[28];
    assign G[68] = in1[27] & in2[27];
    assign P[68] = in1[27] ^ in2[27];
    assign G[69] = in1[26] & in2[26];
    assign P[69] = in1[26] ^ in2[26];
    assign G[70] = in1[25] & in2[25];
    assign P[70] = in1[25] ^ in2[25];
    assign G[71] = in1[24] & in2[24];
    assign P[71] = in1[24] ^ in2[24];
    assign G[72] = in1[23] & in2[23];
    assign P[72] = in1[23] ^ in2[23];
    assign G[73] = in1[22] & in2[22];
    assign P[73] = in1[22] ^ in2[22];
    assign G[74] = in1[21] & in2[21];
    assign P[74] = in1[21] ^ in2[21];
    assign G[75] = in1[20] & in2[20];
    assign P[75] = in1[20] ^ in2[20];
    assign G[76] = in1[19] & in2[19];
    assign P[76] = in1[19] ^ in2[19];
    assign G[77] = in1[18] & in2[18];
    assign P[77] = in1[18] ^ in2[18];
    assign G[78] = in1[17] & in2[17];
    assign P[78] = in1[17] ^ in2[17];
    assign G[79] = in1[16] & in2[16];
    assign P[79] = in1[16] ^ in2[16];
    assign G[80] = in1[15] & in2[15];
    assign P[80] = in1[15] ^ in2[15];
    assign G[81] = in1[14] & in2[14];
    assign P[81] = in1[14] ^ in2[14];
    assign G[82] = in1[13] & in2[13];
    assign P[82] = in1[13] ^ in2[13];
    assign G[83] = in1[12] & in2[12];
    assign P[83] = in1[12] ^ in2[12];
    assign G[84] = in1[11] & in2[11];
    assign P[84] = in1[11] ^ in2[11];
    assign G[85] = in1[10] & in2[10];
    assign P[85] = in1[10] ^ in2[10];
    assign G[86] = in1[9] & in2[9];
    assign P[86] = in1[9] ^ in2[9];
    assign G[87] = in1[8] & in2[8];
    assign P[87] = in1[8] ^ in2[8];
    assign G[88] = in1[7] & in2[7];
    assign P[88] = in1[7] ^ in2[7];
    assign G[89] = in1[6] & in2[6];
    assign P[89] = in1[6] ^ in2[6];
    assign G[90] = in1[5] & in2[5];
    assign P[90] = in1[5] ^ in2[5];
    assign G[91] = in1[4] & in2[4];
    assign P[91] = in1[4] ^ in2[4];
    assign G[92] = in1[3] & in2[3];
    assign P[92] = in1[3] ^ in2[3];
    assign G[93] = in1[2] & in2[2];
    assign P[93] = in1[2] ^ in2[2];
    assign G[94] = in1[1] & in2[1];
    assign P[94] = in1[1] ^ in2[1];
    assign G[95] = in1[0] & in2[0];
    assign P[95] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign cout = G[95] | (P[95] & C[95]);
    assign sum = P ^ C;
endmodule

module CLA_95(output [94:0] sum, output cout, input [94:0] in1, input [94:0] in2);

    wire[94:0] G;
    wire[94:0] C;
    wire[94:0] P;

    assign G[0] = in1[94] & in2[94];
    assign P[0] = in1[94] ^ in2[94];
    assign G[1] = in1[93] & in2[93];
    assign P[1] = in1[93] ^ in2[93];
    assign G[2] = in1[92] & in2[92];
    assign P[2] = in1[92] ^ in2[92];
    assign G[3] = in1[91] & in2[91];
    assign P[3] = in1[91] ^ in2[91];
    assign G[4] = in1[90] & in2[90];
    assign P[4] = in1[90] ^ in2[90];
    assign G[5] = in1[89] & in2[89];
    assign P[5] = in1[89] ^ in2[89];
    assign G[6] = in1[88] & in2[88];
    assign P[6] = in1[88] ^ in2[88];
    assign G[7] = in1[87] & in2[87];
    assign P[7] = in1[87] ^ in2[87];
    assign G[8] = in1[86] & in2[86];
    assign P[8] = in1[86] ^ in2[86];
    assign G[9] = in1[85] & in2[85];
    assign P[9] = in1[85] ^ in2[85];
    assign G[10] = in1[84] & in2[84];
    assign P[10] = in1[84] ^ in2[84];
    assign G[11] = in1[83] & in2[83];
    assign P[11] = in1[83] ^ in2[83];
    assign G[12] = in1[82] & in2[82];
    assign P[12] = in1[82] ^ in2[82];
    assign G[13] = in1[81] & in2[81];
    assign P[13] = in1[81] ^ in2[81];
    assign G[14] = in1[80] & in2[80];
    assign P[14] = in1[80] ^ in2[80];
    assign G[15] = in1[79] & in2[79];
    assign P[15] = in1[79] ^ in2[79];
    assign G[16] = in1[78] & in2[78];
    assign P[16] = in1[78] ^ in2[78];
    assign G[17] = in1[77] & in2[77];
    assign P[17] = in1[77] ^ in2[77];
    assign G[18] = in1[76] & in2[76];
    assign P[18] = in1[76] ^ in2[76];
    assign G[19] = in1[75] & in2[75];
    assign P[19] = in1[75] ^ in2[75];
    assign G[20] = in1[74] & in2[74];
    assign P[20] = in1[74] ^ in2[74];
    assign G[21] = in1[73] & in2[73];
    assign P[21] = in1[73] ^ in2[73];
    assign G[22] = in1[72] & in2[72];
    assign P[22] = in1[72] ^ in2[72];
    assign G[23] = in1[71] & in2[71];
    assign P[23] = in1[71] ^ in2[71];
    assign G[24] = in1[70] & in2[70];
    assign P[24] = in1[70] ^ in2[70];
    assign G[25] = in1[69] & in2[69];
    assign P[25] = in1[69] ^ in2[69];
    assign G[26] = in1[68] & in2[68];
    assign P[26] = in1[68] ^ in2[68];
    assign G[27] = in1[67] & in2[67];
    assign P[27] = in1[67] ^ in2[67];
    assign G[28] = in1[66] & in2[66];
    assign P[28] = in1[66] ^ in2[66];
    assign G[29] = in1[65] & in2[65];
    assign P[29] = in1[65] ^ in2[65];
    assign G[30] = in1[64] & in2[64];
    assign P[30] = in1[64] ^ in2[64];
    assign G[31] = in1[63] & in2[63];
    assign P[31] = in1[63] ^ in2[63];
    assign G[32] = in1[62] & in2[62];
    assign P[32] = in1[62] ^ in2[62];
    assign G[33] = in1[61] & in2[61];
    assign P[33] = in1[61] ^ in2[61];
    assign G[34] = in1[60] & in2[60];
    assign P[34] = in1[60] ^ in2[60];
    assign G[35] = in1[59] & in2[59];
    assign P[35] = in1[59] ^ in2[59];
    assign G[36] = in1[58] & in2[58];
    assign P[36] = in1[58] ^ in2[58];
    assign G[37] = in1[57] & in2[57];
    assign P[37] = in1[57] ^ in2[57];
    assign G[38] = in1[56] & in2[56];
    assign P[38] = in1[56] ^ in2[56];
    assign G[39] = in1[55] & in2[55];
    assign P[39] = in1[55] ^ in2[55];
    assign G[40] = in1[54] & in2[54];
    assign P[40] = in1[54] ^ in2[54];
    assign G[41] = in1[53] & in2[53];
    assign P[41] = in1[53] ^ in2[53];
    assign G[42] = in1[52] & in2[52];
    assign P[42] = in1[52] ^ in2[52];
    assign G[43] = in1[51] & in2[51];
    assign P[43] = in1[51] ^ in2[51];
    assign G[44] = in1[50] & in2[50];
    assign P[44] = in1[50] ^ in2[50];
    assign G[45] = in1[49] & in2[49];
    assign P[45] = in1[49] ^ in2[49];
    assign G[46] = in1[48] & in2[48];
    assign P[46] = in1[48] ^ in2[48];
    assign G[47] = in1[47] & in2[47];
    assign P[47] = in1[47] ^ in2[47];
    assign G[48] = in1[46] & in2[46];
    assign P[48] = in1[46] ^ in2[46];
    assign G[49] = in1[45] & in2[45];
    assign P[49] = in1[45] ^ in2[45];
    assign G[50] = in1[44] & in2[44];
    assign P[50] = in1[44] ^ in2[44];
    assign G[51] = in1[43] & in2[43];
    assign P[51] = in1[43] ^ in2[43];
    assign G[52] = in1[42] & in2[42];
    assign P[52] = in1[42] ^ in2[42];
    assign G[53] = in1[41] & in2[41];
    assign P[53] = in1[41] ^ in2[41];
    assign G[54] = in1[40] & in2[40];
    assign P[54] = in1[40] ^ in2[40];
    assign G[55] = in1[39] & in2[39];
    assign P[55] = in1[39] ^ in2[39];
    assign G[56] = in1[38] & in2[38];
    assign P[56] = in1[38] ^ in2[38];
    assign G[57] = in1[37] & in2[37];
    assign P[57] = in1[37] ^ in2[37];
    assign G[58] = in1[36] & in2[36];
    assign P[58] = in1[36] ^ in2[36];
    assign G[59] = in1[35] & in2[35];
    assign P[59] = in1[35] ^ in2[35];
    assign G[60] = in1[34] & in2[34];
    assign P[60] = in1[34] ^ in2[34];
    assign G[61] = in1[33] & in2[33];
    assign P[61] = in1[33] ^ in2[33];
    assign G[62] = in1[32] & in2[32];
    assign P[62] = in1[32] ^ in2[32];
    assign G[63] = in1[31] & in2[31];
    assign P[63] = in1[31] ^ in2[31];
    assign G[64] = in1[30] & in2[30];
    assign P[64] = in1[30] ^ in2[30];
    assign G[65] = in1[29] & in2[29];
    assign P[65] = in1[29] ^ in2[29];
    assign G[66] = in1[28] & in2[28];
    assign P[66] = in1[28] ^ in2[28];
    assign G[67] = in1[27] & in2[27];
    assign P[67] = in1[27] ^ in2[27];
    assign G[68] = in1[26] & in2[26];
    assign P[68] = in1[26] ^ in2[26];
    assign G[69] = in1[25] & in2[25];
    assign P[69] = in1[25] ^ in2[25];
    assign G[70] = in1[24] & in2[24];
    assign P[70] = in1[24] ^ in2[24];
    assign G[71] = in1[23] & in2[23];
    assign P[71] = in1[23] ^ in2[23];
    assign G[72] = in1[22] & in2[22];
    assign P[72] = in1[22] ^ in2[22];
    assign G[73] = in1[21] & in2[21];
    assign P[73] = in1[21] ^ in2[21];
    assign G[74] = in1[20] & in2[20];
    assign P[74] = in1[20] ^ in2[20];
    assign G[75] = in1[19] & in2[19];
    assign P[75] = in1[19] ^ in2[19];
    assign G[76] = in1[18] & in2[18];
    assign P[76] = in1[18] ^ in2[18];
    assign G[77] = in1[17] & in2[17];
    assign P[77] = in1[17] ^ in2[17];
    assign G[78] = in1[16] & in2[16];
    assign P[78] = in1[16] ^ in2[16];
    assign G[79] = in1[15] & in2[15];
    assign P[79] = in1[15] ^ in2[15];
    assign G[80] = in1[14] & in2[14];
    assign P[80] = in1[14] ^ in2[14];
    assign G[81] = in1[13] & in2[13];
    assign P[81] = in1[13] ^ in2[13];
    assign G[82] = in1[12] & in2[12];
    assign P[82] = in1[12] ^ in2[12];
    assign G[83] = in1[11] & in2[11];
    assign P[83] = in1[11] ^ in2[11];
    assign G[84] = in1[10] & in2[10];
    assign P[84] = in1[10] ^ in2[10];
    assign G[85] = in1[9] & in2[9];
    assign P[85] = in1[9] ^ in2[9];
    assign G[86] = in1[8] & in2[8];
    assign P[86] = in1[8] ^ in2[8];
    assign G[87] = in1[7] & in2[7];
    assign P[87] = in1[7] ^ in2[7];
    assign G[88] = in1[6] & in2[6];
    assign P[88] = in1[6] ^ in2[6];
    assign G[89] = in1[5] & in2[5];
    assign P[89] = in1[5] ^ in2[5];
    assign G[90] = in1[4] & in2[4];
    assign P[90] = in1[4] ^ in2[4];
    assign G[91] = in1[3] & in2[3];
    assign P[91] = in1[3] ^ in2[3];
    assign G[92] = in1[2] & in2[2];
    assign P[92] = in1[2] ^ in2[2];
    assign G[93] = in1[1] & in2[1];
    assign P[93] = in1[1] ^ in2[1];
    assign G[94] = in1[0] & in2[0];
    assign P[94] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign cout = G[94] | (P[94] & C[94]);
    assign sum = P ^ C;
endmodule

module CLA_94(output [93:0] sum, output cout, input [93:0] in1, input [93:0] in2);

    wire[93:0] G;
    wire[93:0] C;
    wire[93:0] P;

    assign G[0] = in1[93] & in2[93];
    assign P[0] = in1[93] ^ in2[93];
    assign G[1] = in1[92] & in2[92];
    assign P[1] = in1[92] ^ in2[92];
    assign G[2] = in1[91] & in2[91];
    assign P[2] = in1[91] ^ in2[91];
    assign G[3] = in1[90] & in2[90];
    assign P[3] = in1[90] ^ in2[90];
    assign G[4] = in1[89] & in2[89];
    assign P[4] = in1[89] ^ in2[89];
    assign G[5] = in1[88] & in2[88];
    assign P[5] = in1[88] ^ in2[88];
    assign G[6] = in1[87] & in2[87];
    assign P[6] = in1[87] ^ in2[87];
    assign G[7] = in1[86] & in2[86];
    assign P[7] = in1[86] ^ in2[86];
    assign G[8] = in1[85] & in2[85];
    assign P[8] = in1[85] ^ in2[85];
    assign G[9] = in1[84] & in2[84];
    assign P[9] = in1[84] ^ in2[84];
    assign G[10] = in1[83] & in2[83];
    assign P[10] = in1[83] ^ in2[83];
    assign G[11] = in1[82] & in2[82];
    assign P[11] = in1[82] ^ in2[82];
    assign G[12] = in1[81] & in2[81];
    assign P[12] = in1[81] ^ in2[81];
    assign G[13] = in1[80] & in2[80];
    assign P[13] = in1[80] ^ in2[80];
    assign G[14] = in1[79] & in2[79];
    assign P[14] = in1[79] ^ in2[79];
    assign G[15] = in1[78] & in2[78];
    assign P[15] = in1[78] ^ in2[78];
    assign G[16] = in1[77] & in2[77];
    assign P[16] = in1[77] ^ in2[77];
    assign G[17] = in1[76] & in2[76];
    assign P[17] = in1[76] ^ in2[76];
    assign G[18] = in1[75] & in2[75];
    assign P[18] = in1[75] ^ in2[75];
    assign G[19] = in1[74] & in2[74];
    assign P[19] = in1[74] ^ in2[74];
    assign G[20] = in1[73] & in2[73];
    assign P[20] = in1[73] ^ in2[73];
    assign G[21] = in1[72] & in2[72];
    assign P[21] = in1[72] ^ in2[72];
    assign G[22] = in1[71] & in2[71];
    assign P[22] = in1[71] ^ in2[71];
    assign G[23] = in1[70] & in2[70];
    assign P[23] = in1[70] ^ in2[70];
    assign G[24] = in1[69] & in2[69];
    assign P[24] = in1[69] ^ in2[69];
    assign G[25] = in1[68] & in2[68];
    assign P[25] = in1[68] ^ in2[68];
    assign G[26] = in1[67] & in2[67];
    assign P[26] = in1[67] ^ in2[67];
    assign G[27] = in1[66] & in2[66];
    assign P[27] = in1[66] ^ in2[66];
    assign G[28] = in1[65] & in2[65];
    assign P[28] = in1[65] ^ in2[65];
    assign G[29] = in1[64] & in2[64];
    assign P[29] = in1[64] ^ in2[64];
    assign G[30] = in1[63] & in2[63];
    assign P[30] = in1[63] ^ in2[63];
    assign G[31] = in1[62] & in2[62];
    assign P[31] = in1[62] ^ in2[62];
    assign G[32] = in1[61] & in2[61];
    assign P[32] = in1[61] ^ in2[61];
    assign G[33] = in1[60] & in2[60];
    assign P[33] = in1[60] ^ in2[60];
    assign G[34] = in1[59] & in2[59];
    assign P[34] = in1[59] ^ in2[59];
    assign G[35] = in1[58] & in2[58];
    assign P[35] = in1[58] ^ in2[58];
    assign G[36] = in1[57] & in2[57];
    assign P[36] = in1[57] ^ in2[57];
    assign G[37] = in1[56] & in2[56];
    assign P[37] = in1[56] ^ in2[56];
    assign G[38] = in1[55] & in2[55];
    assign P[38] = in1[55] ^ in2[55];
    assign G[39] = in1[54] & in2[54];
    assign P[39] = in1[54] ^ in2[54];
    assign G[40] = in1[53] & in2[53];
    assign P[40] = in1[53] ^ in2[53];
    assign G[41] = in1[52] & in2[52];
    assign P[41] = in1[52] ^ in2[52];
    assign G[42] = in1[51] & in2[51];
    assign P[42] = in1[51] ^ in2[51];
    assign G[43] = in1[50] & in2[50];
    assign P[43] = in1[50] ^ in2[50];
    assign G[44] = in1[49] & in2[49];
    assign P[44] = in1[49] ^ in2[49];
    assign G[45] = in1[48] & in2[48];
    assign P[45] = in1[48] ^ in2[48];
    assign G[46] = in1[47] & in2[47];
    assign P[46] = in1[47] ^ in2[47];
    assign G[47] = in1[46] & in2[46];
    assign P[47] = in1[46] ^ in2[46];
    assign G[48] = in1[45] & in2[45];
    assign P[48] = in1[45] ^ in2[45];
    assign G[49] = in1[44] & in2[44];
    assign P[49] = in1[44] ^ in2[44];
    assign G[50] = in1[43] & in2[43];
    assign P[50] = in1[43] ^ in2[43];
    assign G[51] = in1[42] & in2[42];
    assign P[51] = in1[42] ^ in2[42];
    assign G[52] = in1[41] & in2[41];
    assign P[52] = in1[41] ^ in2[41];
    assign G[53] = in1[40] & in2[40];
    assign P[53] = in1[40] ^ in2[40];
    assign G[54] = in1[39] & in2[39];
    assign P[54] = in1[39] ^ in2[39];
    assign G[55] = in1[38] & in2[38];
    assign P[55] = in1[38] ^ in2[38];
    assign G[56] = in1[37] & in2[37];
    assign P[56] = in1[37] ^ in2[37];
    assign G[57] = in1[36] & in2[36];
    assign P[57] = in1[36] ^ in2[36];
    assign G[58] = in1[35] & in2[35];
    assign P[58] = in1[35] ^ in2[35];
    assign G[59] = in1[34] & in2[34];
    assign P[59] = in1[34] ^ in2[34];
    assign G[60] = in1[33] & in2[33];
    assign P[60] = in1[33] ^ in2[33];
    assign G[61] = in1[32] & in2[32];
    assign P[61] = in1[32] ^ in2[32];
    assign G[62] = in1[31] & in2[31];
    assign P[62] = in1[31] ^ in2[31];
    assign G[63] = in1[30] & in2[30];
    assign P[63] = in1[30] ^ in2[30];
    assign G[64] = in1[29] & in2[29];
    assign P[64] = in1[29] ^ in2[29];
    assign G[65] = in1[28] & in2[28];
    assign P[65] = in1[28] ^ in2[28];
    assign G[66] = in1[27] & in2[27];
    assign P[66] = in1[27] ^ in2[27];
    assign G[67] = in1[26] & in2[26];
    assign P[67] = in1[26] ^ in2[26];
    assign G[68] = in1[25] & in2[25];
    assign P[68] = in1[25] ^ in2[25];
    assign G[69] = in1[24] & in2[24];
    assign P[69] = in1[24] ^ in2[24];
    assign G[70] = in1[23] & in2[23];
    assign P[70] = in1[23] ^ in2[23];
    assign G[71] = in1[22] & in2[22];
    assign P[71] = in1[22] ^ in2[22];
    assign G[72] = in1[21] & in2[21];
    assign P[72] = in1[21] ^ in2[21];
    assign G[73] = in1[20] & in2[20];
    assign P[73] = in1[20] ^ in2[20];
    assign G[74] = in1[19] & in2[19];
    assign P[74] = in1[19] ^ in2[19];
    assign G[75] = in1[18] & in2[18];
    assign P[75] = in1[18] ^ in2[18];
    assign G[76] = in1[17] & in2[17];
    assign P[76] = in1[17] ^ in2[17];
    assign G[77] = in1[16] & in2[16];
    assign P[77] = in1[16] ^ in2[16];
    assign G[78] = in1[15] & in2[15];
    assign P[78] = in1[15] ^ in2[15];
    assign G[79] = in1[14] & in2[14];
    assign P[79] = in1[14] ^ in2[14];
    assign G[80] = in1[13] & in2[13];
    assign P[80] = in1[13] ^ in2[13];
    assign G[81] = in1[12] & in2[12];
    assign P[81] = in1[12] ^ in2[12];
    assign G[82] = in1[11] & in2[11];
    assign P[82] = in1[11] ^ in2[11];
    assign G[83] = in1[10] & in2[10];
    assign P[83] = in1[10] ^ in2[10];
    assign G[84] = in1[9] & in2[9];
    assign P[84] = in1[9] ^ in2[9];
    assign G[85] = in1[8] & in2[8];
    assign P[85] = in1[8] ^ in2[8];
    assign G[86] = in1[7] & in2[7];
    assign P[86] = in1[7] ^ in2[7];
    assign G[87] = in1[6] & in2[6];
    assign P[87] = in1[6] ^ in2[6];
    assign G[88] = in1[5] & in2[5];
    assign P[88] = in1[5] ^ in2[5];
    assign G[89] = in1[4] & in2[4];
    assign P[89] = in1[4] ^ in2[4];
    assign G[90] = in1[3] & in2[3];
    assign P[90] = in1[3] ^ in2[3];
    assign G[91] = in1[2] & in2[2];
    assign P[91] = in1[2] ^ in2[2];
    assign G[92] = in1[1] & in2[1];
    assign P[92] = in1[1] ^ in2[1];
    assign G[93] = in1[0] & in2[0];
    assign P[93] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign cout = G[93] | (P[93] & C[93]);
    assign sum = P ^ C;
endmodule

module CLA_93(output [92:0] sum, output cout, input [92:0] in1, input [92:0] in2);

    wire[92:0] G;
    wire[92:0] C;
    wire[92:0] P;

    assign G[0] = in1[92] & in2[92];
    assign P[0] = in1[92] ^ in2[92];
    assign G[1] = in1[91] & in2[91];
    assign P[1] = in1[91] ^ in2[91];
    assign G[2] = in1[90] & in2[90];
    assign P[2] = in1[90] ^ in2[90];
    assign G[3] = in1[89] & in2[89];
    assign P[3] = in1[89] ^ in2[89];
    assign G[4] = in1[88] & in2[88];
    assign P[4] = in1[88] ^ in2[88];
    assign G[5] = in1[87] & in2[87];
    assign P[5] = in1[87] ^ in2[87];
    assign G[6] = in1[86] & in2[86];
    assign P[6] = in1[86] ^ in2[86];
    assign G[7] = in1[85] & in2[85];
    assign P[7] = in1[85] ^ in2[85];
    assign G[8] = in1[84] & in2[84];
    assign P[8] = in1[84] ^ in2[84];
    assign G[9] = in1[83] & in2[83];
    assign P[9] = in1[83] ^ in2[83];
    assign G[10] = in1[82] & in2[82];
    assign P[10] = in1[82] ^ in2[82];
    assign G[11] = in1[81] & in2[81];
    assign P[11] = in1[81] ^ in2[81];
    assign G[12] = in1[80] & in2[80];
    assign P[12] = in1[80] ^ in2[80];
    assign G[13] = in1[79] & in2[79];
    assign P[13] = in1[79] ^ in2[79];
    assign G[14] = in1[78] & in2[78];
    assign P[14] = in1[78] ^ in2[78];
    assign G[15] = in1[77] & in2[77];
    assign P[15] = in1[77] ^ in2[77];
    assign G[16] = in1[76] & in2[76];
    assign P[16] = in1[76] ^ in2[76];
    assign G[17] = in1[75] & in2[75];
    assign P[17] = in1[75] ^ in2[75];
    assign G[18] = in1[74] & in2[74];
    assign P[18] = in1[74] ^ in2[74];
    assign G[19] = in1[73] & in2[73];
    assign P[19] = in1[73] ^ in2[73];
    assign G[20] = in1[72] & in2[72];
    assign P[20] = in1[72] ^ in2[72];
    assign G[21] = in1[71] & in2[71];
    assign P[21] = in1[71] ^ in2[71];
    assign G[22] = in1[70] & in2[70];
    assign P[22] = in1[70] ^ in2[70];
    assign G[23] = in1[69] & in2[69];
    assign P[23] = in1[69] ^ in2[69];
    assign G[24] = in1[68] & in2[68];
    assign P[24] = in1[68] ^ in2[68];
    assign G[25] = in1[67] & in2[67];
    assign P[25] = in1[67] ^ in2[67];
    assign G[26] = in1[66] & in2[66];
    assign P[26] = in1[66] ^ in2[66];
    assign G[27] = in1[65] & in2[65];
    assign P[27] = in1[65] ^ in2[65];
    assign G[28] = in1[64] & in2[64];
    assign P[28] = in1[64] ^ in2[64];
    assign G[29] = in1[63] & in2[63];
    assign P[29] = in1[63] ^ in2[63];
    assign G[30] = in1[62] & in2[62];
    assign P[30] = in1[62] ^ in2[62];
    assign G[31] = in1[61] & in2[61];
    assign P[31] = in1[61] ^ in2[61];
    assign G[32] = in1[60] & in2[60];
    assign P[32] = in1[60] ^ in2[60];
    assign G[33] = in1[59] & in2[59];
    assign P[33] = in1[59] ^ in2[59];
    assign G[34] = in1[58] & in2[58];
    assign P[34] = in1[58] ^ in2[58];
    assign G[35] = in1[57] & in2[57];
    assign P[35] = in1[57] ^ in2[57];
    assign G[36] = in1[56] & in2[56];
    assign P[36] = in1[56] ^ in2[56];
    assign G[37] = in1[55] & in2[55];
    assign P[37] = in1[55] ^ in2[55];
    assign G[38] = in1[54] & in2[54];
    assign P[38] = in1[54] ^ in2[54];
    assign G[39] = in1[53] & in2[53];
    assign P[39] = in1[53] ^ in2[53];
    assign G[40] = in1[52] & in2[52];
    assign P[40] = in1[52] ^ in2[52];
    assign G[41] = in1[51] & in2[51];
    assign P[41] = in1[51] ^ in2[51];
    assign G[42] = in1[50] & in2[50];
    assign P[42] = in1[50] ^ in2[50];
    assign G[43] = in1[49] & in2[49];
    assign P[43] = in1[49] ^ in2[49];
    assign G[44] = in1[48] & in2[48];
    assign P[44] = in1[48] ^ in2[48];
    assign G[45] = in1[47] & in2[47];
    assign P[45] = in1[47] ^ in2[47];
    assign G[46] = in1[46] & in2[46];
    assign P[46] = in1[46] ^ in2[46];
    assign G[47] = in1[45] & in2[45];
    assign P[47] = in1[45] ^ in2[45];
    assign G[48] = in1[44] & in2[44];
    assign P[48] = in1[44] ^ in2[44];
    assign G[49] = in1[43] & in2[43];
    assign P[49] = in1[43] ^ in2[43];
    assign G[50] = in1[42] & in2[42];
    assign P[50] = in1[42] ^ in2[42];
    assign G[51] = in1[41] & in2[41];
    assign P[51] = in1[41] ^ in2[41];
    assign G[52] = in1[40] & in2[40];
    assign P[52] = in1[40] ^ in2[40];
    assign G[53] = in1[39] & in2[39];
    assign P[53] = in1[39] ^ in2[39];
    assign G[54] = in1[38] & in2[38];
    assign P[54] = in1[38] ^ in2[38];
    assign G[55] = in1[37] & in2[37];
    assign P[55] = in1[37] ^ in2[37];
    assign G[56] = in1[36] & in2[36];
    assign P[56] = in1[36] ^ in2[36];
    assign G[57] = in1[35] & in2[35];
    assign P[57] = in1[35] ^ in2[35];
    assign G[58] = in1[34] & in2[34];
    assign P[58] = in1[34] ^ in2[34];
    assign G[59] = in1[33] & in2[33];
    assign P[59] = in1[33] ^ in2[33];
    assign G[60] = in1[32] & in2[32];
    assign P[60] = in1[32] ^ in2[32];
    assign G[61] = in1[31] & in2[31];
    assign P[61] = in1[31] ^ in2[31];
    assign G[62] = in1[30] & in2[30];
    assign P[62] = in1[30] ^ in2[30];
    assign G[63] = in1[29] & in2[29];
    assign P[63] = in1[29] ^ in2[29];
    assign G[64] = in1[28] & in2[28];
    assign P[64] = in1[28] ^ in2[28];
    assign G[65] = in1[27] & in2[27];
    assign P[65] = in1[27] ^ in2[27];
    assign G[66] = in1[26] & in2[26];
    assign P[66] = in1[26] ^ in2[26];
    assign G[67] = in1[25] & in2[25];
    assign P[67] = in1[25] ^ in2[25];
    assign G[68] = in1[24] & in2[24];
    assign P[68] = in1[24] ^ in2[24];
    assign G[69] = in1[23] & in2[23];
    assign P[69] = in1[23] ^ in2[23];
    assign G[70] = in1[22] & in2[22];
    assign P[70] = in1[22] ^ in2[22];
    assign G[71] = in1[21] & in2[21];
    assign P[71] = in1[21] ^ in2[21];
    assign G[72] = in1[20] & in2[20];
    assign P[72] = in1[20] ^ in2[20];
    assign G[73] = in1[19] & in2[19];
    assign P[73] = in1[19] ^ in2[19];
    assign G[74] = in1[18] & in2[18];
    assign P[74] = in1[18] ^ in2[18];
    assign G[75] = in1[17] & in2[17];
    assign P[75] = in1[17] ^ in2[17];
    assign G[76] = in1[16] & in2[16];
    assign P[76] = in1[16] ^ in2[16];
    assign G[77] = in1[15] & in2[15];
    assign P[77] = in1[15] ^ in2[15];
    assign G[78] = in1[14] & in2[14];
    assign P[78] = in1[14] ^ in2[14];
    assign G[79] = in1[13] & in2[13];
    assign P[79] = in1[13] ^ in2[13];
    assign G[80] = in1[12] & in2[12];
    assign P[80] = in1[12] ^ in2[12];
    assign G[81] = in1[11] & in2[11];
    assign P[81] = in1[11] ^ in2[11];
    assign G[82] = in1[10] & in2[10];
    assign P[82] = in1[10] ^ in2[10];
    assign G[83] = in1[9] & in2[9];
    assign P[83] = in1[9] ^ in2[9];
    assign G[84] = in1[8] & in2[8];
    assign P[84] = in1[8] ^ in2[8];
    assign G[85] = in1[7] & in2[7];
    assign P[85] = in1[7] ^ in2[7];
    assign G[86] = in1[6] & in2[6];
    assign P[86] = in1[6] ^ in2[6];
    assign G[87] = in1[5] & in2[5];
    assign P[87] = in1[5] ^ in2[5];
    assign G[88] = in1[4] & in2[4];
    assign P[88] = in1[4] ^ in2[4];
    assign G[89] = in1[3] & in2[3];
    assign P[89] = in1[3] ^ in2[3];
    assign G[90] = in1[2] & in2[2];
    assign P[90] = in1[2] ^ in2[2];
    assign G[91] = in1[1] & in2[1];
    assign P[91] = in1[1] ^ in2[1];
    assign G[92] = in1[0] & in2[0];
    assign P[92] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign cout = G[92] | (P[92] & C[92]);
    assign sum = P ^ C;
endmodule

module CLA_92(output [91:0] sum, output cout, input [91:0] in1, input [91:0] in2);

    wire[91:0] G;
    wire[91:0] C;
    wire[91:0] P;

    assign G[0] = in1[91] & in2[91];
    assign P[0] = in1[91] ^ in2[91];
    assign G[1] = in1[90] & in2[90];
    assign P[1] = in1[90] ^ in2[90];
    assign G[2] = in1[89] & in2[89];
    assign P[2] = in1[89] ^ in2[89];
    assign G[3] = in1[88] & in2[88];
    assign P[3] = in1[88] ^ in2[88];
    assign G[4] = in1[87] & in2[87];
    assign P[4] = in1[87] ^ in2[87];
    assign G[5] = in1[86] & in2[86];
    assign P[5] = in1[86] ^ in2[86];
    assign G[6] = in1[85] & in2[85];
    assign P[6] = in1[85] ^ in2[85];
    assign G[7] = in1[84] & in2[84];
    assign P[7] = in1[84] ^ in2[84];
    assign G[8] = in1[83] & in2[83];
    assign P[8] = in1[83] ^ in2[83];
    assign G[9] = in1[82] & in2[82];
    assign P[9] = in1[82] ^ in2[82];
    assign G[10] = in1[81] & in2[81];
    assign P[10] = in1[81] ^ in2[81];
    assign G[11] = in1[80] & in2[80];
    assign P[11] = in1[80] ^ in2[80];
    assign G[12] = in1[79] & in2[79];
    assign P[12] = in1[79] ^ in2[79];
    assign G[13] = in1[78] & in2[78];
    assign P[13] = in1[78] ^ in2[78];
    assign G[14] = in1[77] & in2[77];
    assign P[14] = in1[77] ^ in2[77];
    assign G[15] = in1[76] & in2[76];
    assign P[15] = in1[76] ^ in2[76];
    assign G[16] = in1[75] & in2[75];
    assign P[16] = in1[75] ^ in2[75];
    assign G[17] = in1[74] & in2[74];
    assign P[17] = in1[74] ^ in2[74];
    assign G[18] = in1[73] & in2[73];
    assign P[18] = in1[73] ^ in2[73];
    assign G[19] = in1[72] & in2[72];
    assign P[19] = in1[72] ^ in2[72];
    assign G[20] = in1[71] & in2[71];
    assign P[20] = in1[71] ^ in2[71];
    assign G[21] = in1[70] & in2[70];
    assign P[21] = in1[70] ^ in2[70];
    assign G[22] = in1[69] & in2[69];
    assign P[22] = in1[69] ^ in2[69];
    assign G[23] = in1[68] & in2[68];
    assign P[23] = in1[68] ^ in2[68];
    assign G[24] = in1[67] & in2[67];
    assign P[24] = in1[67] ^ in2[67];
    assign G[25] = in1[66] & in2[66];
    assign P[25] = in1[66] ^ in2[66];
    assign G[26] = in1[65] & in2[65];
    assign P[26] = in1[65] ^ in2[65];
    assign G[27] = in1[64] & in2[64];
    assign P[27] = in1[64] ^ in2[64];
    assign G[28] = in1[63] & in2[63];
    assign P[28] = in1[63] ^ in2[63];
    assign G[29] = in1[62] & in2[62];
    assign P[29] = in1[62] ^ in2[62];
    assign G[30] = in1[61] & in2[61];
    assign P[30] = in1[61] ^ in2[61];
    assign G[31] = in1[60] & in2[60];
    assign P[31] = in1[60] ^ in2[60];
    assign G[32] = in1[59] & in2[59];
    assign P[32] = in1[59] ^ in2[59];
    assign G[33] = in1[58] & in2[58];
    assign P[33] = in1[58] ^ in2[58];
    assign G[34] = in1[57] & in2[57];
    assign P[34] = in1[57] ^ in2[57];
    assign G[35] = in1[56] & in2[56];
    assign P[35] = in1[56] ^ in2[56];
    assign G[36] = in1[55] & in2[55];
    assign P[36] = in1[55] ^ in2[55];
    assign G[37] = in1[54] & in2[54];
    assign P[37] = in1[54] ^ in2[54];
    assign G[38] = in1[53] & in2[53];
    assign P[38] = in1[53] ^ in2[53];
    assign G[39] = in1[52] & in2[52];
    assign P[39] = in1[52] ^ in2[52];
    assign G[40] = in1[51] & in2[51];
    assign P[40] = in1[51] ^ in2[51];
    assign G[41] = in1[50] & in2[50];
    assign P[41] = in1[50] ^ in2[50];
    assign G[42] = in1[49] & in2[49];
    assign P[42] = in1[49] ^ in2[49];
    assign G[43] = in1[48] & in2[48];
    assign P[43] = in1[48] ^ in2[48];
    assign G[44] = in1[47] & in2[47];
    assign P[44] = in1[47] ^ in2[47];
    assign G[45] = in1[46] & in2[46];
    assign P[45] = in1[46] ^ in2[46];
    assign G[46] = in1[45] & in2[45];
    assign P[46] = in1[45] ^ in2[45];
    assign G[47] = in1[44] & in2[44];
    assign P[47] = in1[44] ^ in2[44];
    assign G[48] = in1[43] & in2[43];
    assign P[48] = in1[43] ^ in2[43];
    assign G[49] = in1[42] & in2[42];
    assign P[49] = in1[42] ^ in2[42];
    assign G[50] = in1[41] & in2[41];
    assign P[50] = in1[41] ^ in2[41];
    assign G[51] = in1[40] & in2[40];
    assign P[51] = in1[40] ^ in2[40];
    assign G[52] = in1[39] & in2[39];
    assign P[52] = in1[39] ^ in2[39];
    assign G[53] = in1[38] & in2[38];
    assign P[53] = in1[38] ^ in2[38];
    assign G[54] = in1[37] & in2[37];
    assign P[54] = in1[37] ^ in2[37];
    assign G[55] = in1[36] & in2[36];
    assign P[55] = in1[36] ^ in2[36];
    assign G[56] = in1[35] & in2[35];
    assign P[56] = in1[35] ^ in2[35];
    assign G[57] = in1[34] & in2[34];
    assign P[57] = in1[34] ^ in2[34];
    assign G[58] = in1[33] & in2[33];
    assign P[58] = in1[33] ^ in2[33];
    assign G[59] = in1[32] & in2[32];
    assign P[59] = in1[32] ^ in2[32];
    assign G[60] = in1[31] & in2[31];
    assign P[60] = in1[31] ^ in2[31];
    assign G[61] = in1[30] & in2[30];
    assign P[61] = in1[30] ^ in2[30];
    assign G[62] = in1[29] & in2[29];
    assign P[62] = in1[29] ^ in2[29];
    assign G[63] = in1[28] & in2[28];
    assign P[63] = in1[28] ^ in2[28];
    assign G[64] = in1[27] & in2[27];
    assign P[64] = in1[27] ^ in2[27];
    assign G[65] = in1[26] & in2[26];
    assign P[65] = in1[26] ^ in2[26];
    assign G[66] = in1[25] & in2[25];
    assign P[66] = in1[25] ^ in2[25];
    assign G[67] = in1[24] & in2[24];
    assign P[67] = in1[24] ^ in2[24];
    assign G[68] = in1[23] & in2[23];
    assign P[68] = in1[23] ^ in2[23];
    assign G[69] = in1[22] & in2[22];
    assign P[69] = in1[22] ^ in2[22];
    assign G[70] = in1[21] & in2[21];
    assign P[70] = in1[21] ^ in2[21];
    assign G[71] = in1[20] & in2[20];
    assign P[71] = in1[20] ^ in2[20];
    assign G[72] = in1[19] & in2[19];
    assign P[72] = in1[19] ^ in2[19];
    assign G[73] = in1[18] & in2[18];
    assign P[73] = in1[18] ^ in2[18];
    assign G[74] = in1[17] & in2[17];
    assign P[74] = in1[17] ^ in2[17];
    assign G[75] = in1[16] & in2[16];
    assign P[75] = in1[16] ^ in2[16];
    assign G[76] = in1[15] & in2[15];
    assign P[76] = in1[15] ^ in2[15];
    assign G[77] = in1[14] & in2[14];
    assign P[77] = in1[14] ^ in2[14];
    assign G[78] = in1[13] & in2[13];
    assign P[78] = in1[13] ^ in2[13];
    assign G[79] = in1[12] & in2[12];
    assign P[79] = in1[12] ^ in2[12];
    assign G[80] = in1[11] & in2[11];
    assign P[80] = in1[11] ^ in2[11];
    assign G[81] = in1[10] & in2[10];
    assign P[81] = in1[10] ^ in2[10];
    assign G[82] = in1[9] & in2[9];
    assign P[82] = in1[9] ^ in2[9];
    assign G[83] = in1[8] & in2[8];
    assign P[83] = in1[8] ^ in2[8];
    assign G[84] = in1[7] & in2[7];
    assign P[84] = in1[7] ^ in2[7];
    assign G[85] = in1[6] & in2[6];
    assign P[85] = in1[6] ^ in2[6];
    assign G[86] = in1[5] & in2[5];
    assign P[86] = in1[5] ^ in2[5];
    assign G[87] = in1[4] & in2[4];
    assign P[87] = in1[4] ^ in2[4];
    assign G[88] = in1[3] & in2[3];
    assign P[88] = in1[3] ^ in2[3];
    assign G[89] = in1[2] & in2[2];
    assign P[89] = in1[2] ^ in2[2];
    assign G[90] = in1[1] & in2[1];
    assign P[90] = in1[1] ^ in2[1];
    assign G[91] = in1[0] & in2[0];
    assign P[91] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign cout = G[91] | (P[91] & C[91]);
    assign sum = P ^ C;
endmodule

module CLA_91(output [90:0] sum, output cout, input [90:0] in1, input [90:0] in2);

    wire[90:0] G;
    wire[90:0] C;
    wire[90:0] P;

    assign G[0] = in1[90] & in2[90];
    assign P[0] = in1[90] ^ in2[90];
    assign G[1] = in1[89] & in2[89];
    assign P[1] = in1[89] ^ in2[89];
    assign G[2] = in1[88] & in2[88];
    assign P[2] = in1[88] ^ in2[88];
    assign G[3] = in1[87] & in2[87];
    assign P[3] = in1[87] ^ in2[87];
    assign G[4] = in1[86] & in2[86];
    assign P[4] = in1[86] ^ in2[86];
    assign G[5] = in1[85] & in2[85];
    assign P[5] = in1[85] ^ in2[85];
    assign G[6] = in1[84] & in2[84];
    assign P[6] = in1[84] ^ in2[84];
    assign G[7] = in1[83] & in2[83];
    assign P[7] = in1[83] ^ in2[83];
    assign G[8] = in1[82] & in2[82];
    assign P[8] = in1[82] ^ in2[82];
    assign G[9] = in1[81] & in2[81];
    assign P[9] = in1[81] ^ in2[81];
    assign G[10] = in1[80] & in2[80];
    assign P[10] = in1[80] ^ in2[80];
    assign G[11] = in1[79] & in2[79];
    assign P[11] = in1[79] ^ in2[79];
    assign G[12] = in1[78] & in2[78];
    assign P[12] = in1[78] ^ in2[78];
    assign G[13] = in1[77] & in2[77];
    assign P[13] = in1[77] ^ in2[77];
    assign G[14] = in1[76] & in2[76];
    assign P[14] = in1[76] ^ in2[76];
    assign G[15] = in1[75] & in2[75];
    assign P[15] = in1[75] ^ in2[75];
    assign G[16] = in1[74] & in2[74];
    assign P[16] = in1[74] ^ in2[74];
    assign G[17] = in1[73] & in2[73];
    assign P[17] = in1[73] ^ in2[73];
    assign G[18] = in1[72] & in2[72];
    assign P[18] = in1[72] ^ in2[72];
    assign G[19] = in1[71] & in2[71];
    assign P[19] = in1[71] ^ in2[71];
    assign G[20] = in1[70] & in2[70];
    assign P[20] = in1[70] ^ in2[70];
    assign G[21] = in1[69] & in2[69];
    assign P[21] = in1[69] ^ in2[69];
    assign G[22] = in1[68] & in2[68];
    assign P[22] = in1[68] ^ in2[68];
    assign G[23] = in1[67] & in2[67];
    assign P[23] = in1[67] ^ in2[67];
    assign G[24] = in1[66] & in2[66];
    assign P[24] = in1[66] ^ in2[66];
    assign G[25] = in1[65] & in2[65];
    assign P[25] = in1[65] ^ in2[65];
    assign G[26] = in1[64] & in2[64];
    assign P[26] = in1[64] ^ in2[64];
    assign G[27] = in1[63] & in2[63];
    assign P[27] = in1[63] ^ in2[63];
    assign G[28] = in1[62] & in2[62];
    assign P[28] = in1[62] ^ in2[62];
    assign G[29] = in1[61] & in2[61];
    assign P[29] = in1[61] ^ in2[61];
    assign G[30] = in1[60] & in2[60];
    assign P[30] = in1[60] ^ in2[60];
    assign G[31] = in1[59] & in2[59];
    assign P[31] = in1[59] ^ in2[59];
    assign G[32] = in1[58] & in2[58];
    assign P[32] = in1[58] ^ in2[58];
    assign G[33] = in1[57] & in2[57];
    assign P[33] = in1[57] ^ in2[57];
    assign G[34] = in1[56] & in2[56];
    assign P[34] = in1[56] ^ in2[56];
    assign G[35] = in1[55] & in2[55];
    assign P[35] = in1[55] ^ in2[55];
    assign G[36] = in1[54] & in2[54];
    assign P[36] = in1[54] ^ in2[54];
    assign G[37] = in1[53] & in2[53];
    assign P[37] = in1[53] ^ in2[53];
    assign G[38] = in1[52] & in2[52];
    assign P[38] = in1[52] ^ in2[52];
    assign G[39] = in1[51] & in2[51];
    assign P[39] = in1[51] ^ in2[51];
    assign G[40] = in1[50] & in2[50];
    assign P[40] = in1[50] ^ in2[50];
    assign G[41] = in1[49] & in2[49];
    assign P[41] = in1[49] ^ in2[49];
    assign G[42] = in1[48] & in2[48];
    assign P[42] = in1[48] ^ in2[48];
    assign G[43] = in1[47] & in2[47];
    assign P[43] = in1[47] ^ in2[47];
    assign G[44] = in1[46] & in2[46];
    assign P[44] = in1[46] ^ in2[46];
    assign G[45] = in1[45] & in2[45];
    assign P[45] = in1[45] ^ in2[45];
    assign G[46] = in1[44] & in2[44];
    assign P[46] = in1[44] ^ in2[44];
    assign G[47] = in1[43] & in2[43];
    assign P[47] = in1[43] ^ in2[43];
    assign G[48] = in1[42] & in2[42];
    assign P[48] = in1[42] ^ in2[42];
    assign G[49] = in1[41] & in2[41];
    assign P[49] = in1[41] ^ in2[41];
    assign G[50] = in1[40] & in2[40];
    assign P[50] = in1[40] ^ in2[40];
    assign G[51] = in1[39] & in2[39];
    assign P[51] = in1[39] ^ in2[39];
    assign G[52] = in1[38] & in2[38];
    assign P[52] = in1[38] ^ in2[38];
    assign G[53] = in1[37] & in2[37];
    assign P[53] = in1[37] ^ in2[37];
    assign G[54] = in1[36] & in2[36];
    assign P[54] = in1[36] ^ in2[36];
    assign G[55] = in1[35] & in2[35];
    assign P[55] = in1[35] ^ in2[35];
    assign G[56] = in1[34] & in2[34];
    assign P[56] = in1[34] ^ in2[34];
    assign G[57] = in1[33] & in2[33];
    assign P[57] = in1[33] ^ in2[33];
    assign G[58] = in1[32] & in2[32];
    assign P[58] = in1[32] ^ in2[32];
    assign G[59] = in1[31] & in2[31];
    assign P[59] = in1[31] ^ in2[31];
    assign G[60] = in1[30] & in2[30];
    assign P[60] = in1[30] ^ in2[30];
    assign G[61] = in1[29] & in2[29];
    assign P[61] = in1[29] ^ in2[29];
    assign G[62] = in1[28] & in2[28];
    assign P[62] = in1[28] ^ in2[28];
    assign G[63] = in1[27] & in2[27];
    assign P[63] = in1[27] ^ in2[27];
    assign G[64] = in1[26] & in2[26];
    assign P[64] = in1[26] ^ in2[26];
    assign G[65] = in1[25] & in2[25];
    assign P[65] = in1[25] ^ in2[25];
    assign G[66] = in1[24] & in2[24];
    assign P[66] = in1[24] ^ in2[24];
    assign G[67] = in1[23] & in2[23];
    assign P[67] = in1[23] ^ in2[23];
    assign G[68] = in1[22] & in2[22];
    assign P[68] = in1[22] ^ in2[22];
    assign G[69] = in1[21] & in2[21];
    assign P[69] = in1[21] ^ in2[21];
    assign G[70] = in1[20] & in2[20];
    assign P[70] = in1[20] ^ in2[20];
    assign G[71] = in1[19] & in2[19];
    assign P[71] = in1[19] ^ in2[19];
    assign G[72] = in1[18] & in2[18];
    assign P[72] = in1[18] ^ in2[18];
    assign G[73] = in1[17] & in2[17];
    assign P[73] = in1[17] ^ in2[17];
    assign G[74] = in1[16] & in2[16];
    assign P[74] = in1[16] ^ in2[16];
    assign G[75] = in1[15] & in2[15];
    assign P[75] = in1[15] ^ in2[15];
    assign G[76] = in1[14] & in2[14];
    assign P[76] = in1[14] ^ in2[14];
    assign G[77] = in1[13] & in2[13];
    assign P[77] = in1[13] ^ in2[13];
    assign G[78] = in1[12] & in2[12];
    assign P[78] = in1[12] ^ in2[12];
    assign G[79] = in1[11] & in2[11];
    assign P[79] = in1[11] ^ in2[11];
    assign G[80] = in1[10] & in2[10];
    assign P[80] = in1[10] ^ in2[10];
    assign G[81] = in1[9] & in2[9];
    assign P[81] = in1[9] ^ in2[9];
    assign G[82] = in1[8] & in2[8];
    assign P[82] = in1[8] ^ in2[8];
    assign G[83] = in1[7] & in2[7];
    assign P[83] = in1[7] ^ in2[7];
    assign G[84] = in1[6] & in2[6];
    assign P[84] = in1[6] ^ in2[6];
    assign G[85] = in1[5] & in2[5];
    assign P[85] = in1[5] ^ in2[5];
    assign G[86] = in1[4] & in2[4];
    assign P[86] = in1[4] ^ in2[4];
    assign G[87] = in1[3] & in2[3];
    assign P[87] = in1[3] ^ in2[3];
    assign G[88] = in1[2] & in2[2];
    assign P[88] = in1[2] ^ in2[2];
    assign G[89] = in1[1] & in2[1];
    assign P[89] = in1[1] ^ in2[1];
    assign G[90] = in1[0] & in2[0];
    assign P[90] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign cout = G[90] | (P[90] & C[90]);
    assign sum = P ^ C;
endmodule

module CLA_90(output [89:0] sum, output cout, input [89:0] in1, input [89:0] in2);

    wire[89:0] G;
    wire[89:0] C;
    wire[89:0] P;

    assign G[0] = in1[89] & in2[89];
    assign P[0] = in1[89] ^ in2[89];
    assign G[1] = in1[88] & in2[88];
    assign P[1] = in1[88] ^ in2[88];
    assign G[2] = in1[87] & in2[87];
    assign P[2] = in1[87] ^ in2[87];
    assign G[3] = in1[86] & in2[86];
    assign P[3] = in1[86] ^ in2[86];
    assign G[4] = in1[85] & in2[85];
    assign P[4] = in1[85] ^ in2[85];
    assign G[5] = in1[84] & in2[84];
    assign P[5] = in1[84] ^ in2[84];
    assign G[6] = in1[83] & in2[83];
    assign P[6] = in1[83] ^ in2[83];
    assign G[7] = in1[82] & in2[82];
    assign P[7] = in1[82] ^ in2[82];
    assign G[8] = in1[81] & in2[81];
    assign P[8] = in1[81] ^ in2[81];
    assign G[9] = in1[80] & in2[80];
    assign P[9] = in1[80] ^ in2[80];
    assign G[10] = in1[79] & in2[79];
    assign P[10] = in1[79] ^ in2[79];
    assign G[11] = in1[78] & in2[78];
    assign P[11] = in1[78] ^ in2[78];
    assign G[12] = in1[77] & in2[77];
    assign P[12] = in1[77] ^ in2[77];
    assign G[13] = in1[76] & in2[76];
    assign P[13] = in1[76] ^ in2[76];
    assign G[14] = in1[75] & in2[75];
    assign P[14] = in1[75] ^ in2[75];
    assign G[15] = in1[74] & in2[74];
    assign P[15] = in1[74] ^ in2[74];
    assign G[16] = in1[73] & in2[73];
    assign P[16] = in1[73] ^ in2[73];
    assign G[17] = in1[72] & in2[72];
    assign P[17] = in1[72] ^ in2[72];
    assign G[18] = in1[71] & in2[71];
    assign P[18] = in1[71] ^ in2[71];
    assign G[19] = in1[70] & in2[70];
    assign P[19] = in1[70] ^ in2[70];
    assign G[20] = in1[69] & in2[69];
    assign P[20] = in1[69] ^ in2[69];
    assign G[21] = in1[68] & in2[68];
    assign P[21] = in1[68] ^ in2[68];
    assign G[22] = in1[67] & in2[67];
    assign P[22] = in1[67] ^ in2[67];
    assign G[23] = in1[66] & in2[66];
    assign P[23] = in1[66] ^ in2[66];
    assign G[24] = in1[65] & in2[65];
    assign P[24] = in1[65] ^ in2[65];
    assign G[25] = in1[64] & in2[64];
    assign P[25] = in1[64] ^ in2[64];
    assign G[26] = in1[63] & in2[63];
    assign P[26] = in1[63] ^ in2[63];
    assign G[27] = in1[62] & in2[62];
    assign P[27] = in1[62] ^ in2[62];
    assign G[28] = in1[61] & in2[61];
    assign P[28] = in1[61] ^ in2[61];
    assign G[29] = in1[60] & in2[60];
    assign P[29] = in1[60] ^ in2[60];
    assign G[30] = in1[59] & in2[59];
    assign P[30] = in1[59] ^ in2[59];
    assign G[31] = in1[58] & in2[58];
    assign P[31] = in1[58] ^ in2[58];
    assign G[32] = in1[57] & in2[57];
    assign P[32] = in1[57] ^ in2[57];
    assign G[33] = in1[56] & in2[56];
    assign P[33] = in1[56] ^ in2[56];
    assign G[34] = in1[55] & in2[55];
    assign P[34] = in1[55] ^ in2[55];
    assign G[35] = in1[54] & in2[54];
    assign P[35] = in1[54] ^ in2[54];
    assign G[36] = in1[53] & in2[53];
    assign P[36] = in1[53] ^ in2[53];
    assign G[37] = in1[52] & in2[52];
    assign P[37] = in1[52] ^ in2[52];
    assign G[38] = in1[51] & in2[51];
    assign P[38] = in1[51] ^ in2[51];
    assign G[39] = in1[50] & in2[50];
    assign P[39] = in1[50] ^ in2[50];
    assign G[40] = in1[49] & in2[49];
    assign P[40] = in1[49] ^ in2[49];
    assign G[41] = in1[48] & in2[48];
    assign P[41] = in1[48] ^ in2[48];
    assign G[42] = in1[47] & in2[47];
    assign P[42] = in1[47] ^ in2[47];
    assign G[43] = in1[46] & in2[46];
    assign P[43] = in1[46] ^ in2[46];
    assign G[44] = in1[45] & in2[45];
    assign P[44] = in1[45] ^ in2[45];
    assign G[45] = in1[44] & in2[44];
    assign P[45] = in1[44] ^ in2[44];
    assign G[46] = in1[43] & in2[43];
    assign P[46] = in1[43] ^ in2[43];
    assign G[47] = in1[42] & in2[42];
    assign P[47] = in1[42] ^ in2[42];
    assign G[48] = in1[41] & in2[41];
    assign P[48] = in1[41] ^ in2[41];
    assign G[49] = in1[40] & in2[40];
    assign P[49] = in1[40] ^ in2[40];
    assign G[50] = in1[39] & in2[39];
    assign P[50] = in1[39] ^ in2[39];
    assign G[51] = in1[38] & in2[38];
    assign P[51] = in1[38] ^ in2[38];
    assign G[52] = in1[37] & in2[37];
    assign P[52] = in1[37] ^ in2[37];
    assign G[53] = in1[36] & in2[36];
    assign P[53] = in1[36] ^ in2[36];
    assign G[54] = in1[35] & in2[35];
    assign P[54] = in1[35] ^ in2[35];
    assign G[55] = in1[34] & in2[34];
    assign P[55] = in1[34] ^ in2[34];
    assign G[56] = in1[33] & in2[33];
    assign P[56] = in1[33] ^ in2[33];
    assign G[57] = in1[32] & in2[32];
    assign P[57] = in1[32] ^ in2[32];
    assign G[58] = in1[31] & in2[31];
    assign P[58] = in1[31] ^ in2[31];
    assign G[59] = in1[30] & in2[30];
    assign P[59] = in1[30] ^ in2[30];
    assign G[60] = in1[29] & in2[29];
    assign P[60] = in1[29] ^ in2[29];
    assign G[61] = in1[28] & in2[28];
    assign P[61] = in1[28] ^ in2[28];
    assign G[62] = in1[27] & in2[27];
    assign P[62] = in1[27] ^ in2[27];
    assign G[63] = in1[26] & in2[26];
    assign P[63] = in1[26] ^ in2[26];
    assign G[64] = in1[25] & in2[25];
    assign P[64] = in1[25] ^ in2[25];
    assign G[65] = in1[24] & in2[24];
    assign P[65] = in1[24] ^ in2[24];
    assign G[66] = in1[23] & in2[23];
    assign P[66] = in1[23] ^ in2[23];
    assign G[67] = in1[22] & in2[22];
    assign P[67] = in1[22] ^ in2[22];
    assign G[68] = in1[21] & in2[21];
    assign P[68] = in1[21] ^ in2[21];
    assign G[69] = in1[20] & in2[20];
    assign P[69] = in1[20] ^ in2[20];
    assign G[70] = in1[19] & in2[19];
    assign P[70] = in1[19] ^ in2[19];
    assign G[71] = in1[18] & in2[18];
    assign P[71] = in1[18] ^ in2[18];
    assign G[72] = in1[17] & in2[17];
    assign P[72] = in1[17] ^ in2[17];
    assign G[73] = in1[16] & in2[16];
    assign P[73] = in1[16] ^ in2[16];
    assign G[74] = in1[15] & in2[15];
    assign P[74] = in1[15] ^ in2[15];
    assign G[75] = in1[14] & in2[14];
    assign P[75] = in1[14] ^ in2[14];
    assign G[76] = in1[13] & in2[13];
    assign P[76] = in1[13] ^ in2[13];
    assign G[77] = in1[12] & in2[12];
    assign P[77] = in1[12] ^ in2[12];
    assign G[78] = in1[11] & in2[11];
    assign P[78] = in1[11] ^ in2[11];
    assign G[79] = in1[10] & in2[10];
    assign P[79] = in1[10] ^ in2[10];
    assign G[80] = in1[9] & in2[9];
    assign P[80] = in1[9] ^ in2[9];
    assign G[81] = in1[8] & in2[8];
    assign P[81] = in1[8] ^ in2[8];
    assign G[82] = in1[7] & in2[7];
    assign P[82] = in1[7] ^ in2[7];
    assign G[83] = in1[6] & in2[6];
    assign P[83] = in1[6] ^ in2[6];
    assign G[84] = in1[5] & in2[5];
    assign P[84] = in1[5] ^ in2[5];
    assign G[85] = in1[4] & in2[4];
    assign P[85] = in1[4] ^ in2[4];
    assign G[86] = in1[3] & in2[3];
    assign P[86] = in1[3] ^ in2[3];
    assign G[87] = in1[2] & in2[2];
    assign P[87] = in1[2] ^ in2[2];
    assign G[88] = in1[1] & in2[1];
    assign P[88] = in1[1] ^ in2[1];
    assign G[89] = in1[0] & in2[0];
    assign P[89] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign cout = G[89] | (P[89] & C[89]);
    assign sum = P ^ C;
endmodule

module CLA_89(output [88:0] sum, output cout, input [88:0] in1, input [88:0] in2);

    wire[88:0] G;
    wire[88:0] C;
    wire[88:0] P;

    assign G[0] = in1[88] & in2[88];
    assign P[0] = in1[88] ^ in2[88];
    assign G[1] = in1[87] & in2[87];
    assign P[1] = in1[87] ^ in2[87];
    assign G[2] = in1[86] & in2[86];
    assign P[2] = in1[86] ^ in2[86];
    assign G[3] = in1[85] & in2[85];
    assign P[3] = in1[85] ^ in2[85];
    assign G[4] = in1[84] & in2[84];
    assign P[4] = in1[84] ^ in2[84];
    assign G[5] = in1[83] & in2[83];
    assign P[5] = in1[83] ^ in2[83];
    assign G[6] = in1[82] & in2[82];
    assign P[6] = in1[82] ^ in2[82];
    assign G[7] = in1[81] & in2[81];
    assign P[7] = in1[81] ^ in2[81];
    assign G[8] = in1[80] & in2[80];
    assign P[8] = in1[80] ^ in2[80];
    assign G[9] = in1[79] & in2[79];
    assign P[9] = in1[79] ^ in2[79];
    assign G[10] = in1[78] & in2[78];
    assign P[10] = in1[78] ^ in2[78];
    assign G[11] = in1[77] & in2[77];
    assign P[11] = in1[77] ^ in2[77];
    assign G[12] = in1[76] & in2[76];
    assign P[12] = in1[76] ^ in2[76];
    assign G[13] = in1[75] & in2[75];
    assign P[13] = in1[75] ^ in2[75];
    assign G[14] = in1[74] & in2[74];
    assign P[14] = in1[74] ^ in2[74];
    assign G[15] = in1[73] & in2[73];
    assign P[15] = in1[73] ^ in2[73];
    assign G[16] = in1[72] & in2[72];
    assign P[16] = in1[72] ^ in2[72];
    assign G[17] = in1[71] & in2[71];
    assign P[17] = in1[71] ^ in2[71];
    assign G[18] = in1[70] & in2[70];
    assign P[18] = in1[70] ^ in2[70];
    assign G[19] = in1[69] & in2[69];
    assign P[19] = in1[69] ^ in2[69];
    assign G[20] = in1[68] & in2[68];
    assign P[20] = in1[68] ^ in2[68];
    assign G[21] = in1[67] & in2[67];
    assign P[21] = in1[67] ^ in2[67];
    assign G[22] = in1[66] & in2[66];
    assign P[22] = in1[66] ^ in2[66];
    assign G[23] = in1[65] & in2[65];
    assign P[23] = in1[65] ^ in2[65];
    assign G[24] = in1[64] & in2[64];
    assign P[24] = in1[64] ^ in2[64];
    assign G[25] = in1[63] & in2[63];
    assign P[25] = in1[63] ^ in2[63];
    assign G[26] = in1[62] & in2[62];
    assign P[26] = in1[62] ^ in2[62];
    assign G[27] = in1[61] & in2[61];
    assign P[27] = in1[61] ^ in2[61];
    assign G[28] = in1[60] & in2[60];
    assign P[28] = in1[60] ^ in2[60];
    assign G[29] = in1[59] & in2[59];
    assign P[29] = in1[59] ^ in2[59];
    assign G[30] = in1[58] & in2[58];
    assign P[30] = in1[58] ^ in2[58];
    assign G[31] = in1[57] & in2[57];
    assign P[31] = in1[57] ^ in2[57];
    assign G[32] = in1[56] & in2[56];
    assign P[32] = in1[56] ^ in2[56];
    assign G[33] = in1[55] & in2[55];
    assign P[33] = in1[55] ^ in2[55];
    assign G[34] = in1[54] & in2[54];
    assign P[34] = in1[54] ^ in2[54];
    assign G[35] = in1[53] & in2[53];
    assign P[35] = in1[53] ^ in2[53];
    assign G[36] = in1[52] & in2[52];
    assign P[36] = in1[52] ^ in2[52];
    assign G[37] = in1[51] & in2[51];
    assign P[37] = in1[51] ^ in2[51];
    assign G[38] = in1[50] & in2[50];
    assign P[38] = in1[50] ^ in2[50];
    assign G[39] = in1[49] & in2[49];
    assign P[39] = in1[49] ^ in2[49];
    assign G[40] = in1[48] & in2[48];
    assign P[40] = in1[48] ^ in2[48];
    assign G[41] = in1[47] & in2[47];
    assign P[41] = in1[47] ^ in2[47];
    assign G[42] = in1[46] & in2[46];
    assign P[42] = in1[46] ^ in2[46];
    assign G[43] = in1[45] & in2[45];
    assign P[43] = in1[45] ^ in2[45];
    assign G[44] = in1[44] & in2[44];
    assign P[44] = in1[44] ^ in2[44];
    assign G[45] = in1[43] & in2[43];
    assign P[45] = in1[43] ^ in2[43];
    assign G[46] = in1[42] & in2[42];
    assign P[46] = in1[42] ^ in2[42];
    assign G[47] = in1[41] & in2[41];
    assign P[47] = in1[41] ^ in2[41];
    assign G[48] = in1[40] & in2[40];
    assign P[48] = in1[40] ^ in2[40];
    assign G[49] = in1[39] & in2[39];
    assign P[49] = in1[39] ^ in2[39];
    assign G[50] = in1[38] & in2[38];
    assign P[50] = in1[38] ^ in2[38];
    assign G[51] = in1[37] & in2[37];
    assign P[51] = in1[37] ^ in2[37];
    assign G[52] = in1[36] & in2[36];
    assign P[52] = in1[36] ^ in2[36];
    assign G[53] = in1[35] & in2[35];
    assign P[53] = in1[35] ^ in2[35];
    assign G[54] = in1[34] & in2[34];
    assign P[54] = in1[34] ^ in2[34];
    assign G[55] = in1[33] & in2[33];
    assign P[55] = in1[33] ^ in2[33];
    assign G[56] = in1[32] & in2[32];
    assign P[56] = in1[32] ^ in2[32];
    assign G[57] = in1[31] & in2[31];
    assign P[57] = in1[31] ^ in2[31];
    assign G[58] = in1[30] & in2[30];
    assign P[58] = in1[30] ^ in2[30];
    assign G[59] = in1[29] & in2[29];
    assign P[59] = in1[29] ^ in2[29];
    assign G[60] = in1[28] & in2[28];
    assign P[60] = in1[28] ^ in2[28];
    assign G[61] = in1[27] & in2[27];
    assign P[61] = in1[27] ^ in2[27];
    assign G[62] = in1[26] & in2[26];
    assign P[62] = in1[26] ^ in2[26];
    assign G[63] = in1[25] & in2[25];
    assign P[63] = in1[25] ^ in2[25];
    assign G[64] = in1[24] & in2[24];
    assign P[64] = in1[24] ^ in2[24];
    assign G[65] = in1[23] & in2[23];
    assign P[65] = in1[23] ^ in2[23];
    assign G[66] = in1[22] & in2[22];
    assign P[66] = in1[22] ^ in2[22];
    assign G[67] = in1[21] & in2[21];
    assign P[67] = in1[21] ^ in2[21];
    assign G[68] = in1[20] & in2[20];
    assign P[68] = in1[20] ^ in2[20];
    assign G[69] = in1[19] & in2[19];
    assign P[69] = in1[19] ^ in2[19];
    assign G[70] = in1[18] & in2[18];
    assign P[70] = in1[18] ^ in2[18];
    assign G[71] = in1[17] & in2[17];
    assign P[71] = in1[17] ^ in2[17];
    assign G[72] = in1[16] & in2[16];
    assign P[72] = in1[16] ^ in2[16];
    assign G[73] = in1[15] & in2[15];
    assign P[73] = in1[15] ^ in2[15];
    assign G[74] = in1[14] & in2[14];
    assign P[74] = in1[14] ^ in2[14];
    assign G[75] = in1[13] & in2[13];
    assign P[75] = in1[13] ^ in2[13];
    assign G[76] = in1[12] & in2[12];
    assign P[76] = in1[12] ^ in2[12];
    assign G[77] = in1[11] & in2[11];
    assign P[77] = in1[11] ^ in2[11];
    assign G[78] = in1[10] & in2[10];
    assign P[78] = in1[10] ^ in2[10];
    assign G[79] = in1[9] & in2[9];
    assign P[79] = in1[9] ^ in2[9];
    assign G[80] = in1[8] & in2[8];
    assign P[80] = in1[8] ^ in2[8];
    assign G[81] = in1[7] & in2[7];
    assign P[81] = in1[7] ^ in2[7];
    assign G[82] = in1[6] & in2[6];
    assign P[82] = in1[6] ^ in2[6];
    assign G[83] = in1[5] & in2[5];
    assign P[83] = in1[5] ^ in2[5];
    assign G[84] = in1[4] & in2[4];
    assign P[84] = in1[4] ^ in2[4];
    assign G[85] = in1[3] & in2[3];
    assign P[85] = in1[3] ^ in2[3];
    assign G[86] = in1[2] & in2[2];
    assign P[86] = in1[2] ^ in2[2];
    assign G[87] = in1[1] & in2[1];
    assign P[87] = in1[1] ^ in2[1];
    assign G[88] = in1[0] & in2[0];
    assign P[88] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign cout = G[88] | (P[88] & C[88]);
    assign sum = P ^ C;
endmodule

module CLA_88(output [87:0] sum, output cout, input [87:0] in1, input [87:0] in2);

    wire[87:0] G;
    wire[87:0] C;
    wire[87:0] P;

    assign G[0] = in1[87] & in2[87];
    assign P[0] = in1[87] ^ in2[87];
    assign G[1] = in1[86] & in2[86];
    assign P[1] = in1[86] ^ in2[86];
    assign G[2] = in1[85] & in2[85];
    assign P[2] = in1[85] ^ in2[85];
    assign G[3] = in1[84] & in2[84];
    assign P[3] = in1[84] ^ in2[84];
    assign G[4] = in1[83] & in2[83];
    assign P[4] = in1[83] ^ in2[83];
    assign G[5] = in1[82] & in2[82];
    assign P[5] = in1[82] ^ in2[82];
    assign G[6] = in1[81] & in2[81];
    assign P[6] = in1[81] ^ in2[81];
    assign G[7] = in1[80] & in2[80];
    assign P[7] = in1[80] ^ in2[80];
    assign G[8] = in1[79] & in2[79];
    assign P[8] = in1[79] ^ in2[79];
    assign G[9] = in1[78] & in2[78];
    assign P[9] = in1[78] ^ in2[78];
    assign G[10] = in1[77] & in2[77];
    assign P[10] = in1[77] ^ in2[77];
    assign G[11] = in1[76] & in2[76];
    assign P[11] = in1[76] ^ in2[76];
    assign G[12] = in1[75] & in2[75];
    assign P[12] = in1[75] ^ in2[75];
    assign G[13] = in1[74] & in2[74];
    assign P[13] = in1[74] ^ in2[74];
    assign G[14] = in1[73] & in2[73];
    assign P[14] = in1[73] ^ in2[73];
    assign G[15] = in1[72] & in2[72];
    assign P[15] = in1[72] ^ in2[72];
    assign G[16] = in1[71] & in2[71];
    assign P[16] = in1[71] ^ in2[71];
    assign G[17] = in1[70] & in2[70];
    assign P[17] = in1[70] ^ in2[70];
    assign G[18] = in1[69] & in2[69];
    assign P[18] = in1[69] ^ in2[69];
    assign G[19] = in1[68] & in2[68];
    assign P[19] = in1[68] ^ in2[68];
    assign G[20] = in1[67] & in2[67];
    assign P[20] = in1[67] ^ in2[67];
    assign G[21] = in1[66] & in2[66];
    assign P[21] = in1[66] ^ in2[66];
    assign G[22] = in1[65] & in2[65];
    assign P[22] = in1[65] ^ in2[65];
    assign G[23] = in1[64] & in2[64];
    assign P[23] = in1[64] ^ in2[64];
    assign G[24] = in1[63] & in2[63];
    assign P[24] = in1[63] ^ in2[63];
    assign G[25] = in1[62] & in2[62];
    assign P[25] = in1[62] ^ in2[62];
    assign G[26] = in1[61] & in2[61];
    assign P[26] = in1[61] ^ in2[61];
    assign G[27] = in1[60] & in2[60];
    assign P[27] = in1[60] ^ in2[60];
    assign G[28] = in1[59] & in2[59];
    assign P[28] = in1[59] ^ in2[59];
    assign G[29] = in1[58] & in2[58];
    assign P[29] = in1[58] ^ in2[58];
    assign G[30] = in1[57] & in2[57];
    assign P[30] = in1[57] ^ in2[57];
    assign G[31] = in1[56] & in2[56];
    assign P[31] = in1[56] ^ in2[56];
    assign G[32] = in1[55] & in2[55];
    assign P[32] = in1[55] ^ in2[55];
    assign G[33] = in1[54] & in2[54];
    assign P[33] = in1[54] ^ in2[54];
    assign G[34] = in1[53] & in2[53];
    assign P[34] = in1[53] ^ in2[53];
    assign G[35] = in1[52] & in2[52];
    assign P[35] = in1[52] ^ in2[52];
    assign G[36] = in1[51] & in2[51];
    assign P[36] = in1[51] ^ in2[51];
    assign G[37] = in1[50] & in2[50];
    assign P[37] = in1[50] ^ in2[50];
    assign G[38] = in1[49] & in2[49];
    assign P[38] = in1[49] ^ in2[49];
    assign G[39] = in1[48] & in2[48];
    assign P[39] = in1[48] ^ in2[48];
    assign G[40] = in1[47] & in2[47];
    assign P[40] = in1[47] ^ in2[47];
    assign G[41] = in1[46] & in2[46];
    assign P[41] = in1[46] ^ in2[46];
    assign G[42] = in1[45] & in2[45];
    assign P[42] = in1[45] ^ in2[45];
    assign G[43] = in1[44] & in2[44];
    assign P[43] = in1[44] ^ in2[44];
    assign G[44] = in1[43] & in2[43];
    assign P[44] = in1[43] ^ in2[43];
    assign G[45] = in1[42] & in2[42];
    assign P[45] = in1[42] ^ in2[42];
    assign G[46] = in1[41] & in2[41];
    assign P[46] = in1[41] ^ in2[41];
    assign G[47] = in1[40] & in2[40];
    assign P[47] = in1[40] ^ in2[40];
    assign G[48] = in1[39] & in2[39];
    assign P[48] = in1[39] ^ in2[39];
    assign G[49] = in1[38] & in2[38];
    assign P[49] = in1[38] ^ in2[38];
    assign G[50] = in1[37] & in2[37];
    assign P[50] = in1[37] ^ in2[37];
    assign G[51] = in1[36] & in2[36];
    assign P[51] = in1[36] ^ in2[36];
    assign G[52] = in1[35] & in2[35];
    assign P[52] = in1[35] ^ in2[35];
    assign G[53] = in1[34] & in2[34];
    assign P[53] = in1[34] ^ in2[34];
    assign G[54] = in1[33] & in2[33];
    assign P[54] = in1[33] ^ in2[33];
    assign G[55] = in1[32] & in2[32];
    assign P[55] = in1[32] ^ in2[32];
    assign G[56] = in1[31] & in2[31];
    assign P[56] = in1[31] ^ in2[31];
    assign G[57] = in1[30] & in2[30];
    assign P[57] = in1[30] ^ in2[30];
    assign G[58] = in1[29] & in2[29];
    assign P[58] = in1[29] ^ in2[29];
    assign G[59] = in1[28] & in2[28];
    assign P[59] = in1[28] ^ in2[28];
    assign G[60] = in1[27] & in2[27];
    assign P[60] = in1[27] ^ in2[27];
    assign G[61] = in1[26] & in2[26];
    assign P[61] = in1[26] ^ in2[26];
    assign G[62] = in1[25] & in2[25];
    assign P[62] = in1[25] ^ in2[25];
    assign G[63] = in1[24] & in2[24];
    assign P[63] = in1[24] ^ in2[24];
    assign G[64] = in1[23] & in2[23];
    assign P[64] = in1[23] ^ in2[23];
    assign G[65] = in1[22] & in2[22];
    assign P[65] = in1[22] ^ in2[22];
    assign G[66] = in1[21] & in2[21];
    assign P[66] = in1[21] ^ in2[21];
    assign G[67] = in1[20] & in2[20];
    assign P[67] = in1[20] ^ in2[20];
    assign G[68] = in1[19] & in2[19];
    assign P[68] = in1[19] ^ in2[19];
    assign G[69] = in1[18] & in2[18];
    assign P[69] = in1[18] ^ in2[18];
    assign G[70] = in1[17] & in2[17];
    assign P[70] = in1[17] ^ in2[17];
    assign G[71] = in1[16] & in2[16];
    assign P[71] = in1[16] ^ in2[16];
    assign G[72] = in1[15] & in2[15];
    assign P[72] = in1[15] ^ in2[15];
    assign G[73] = in1[14] & in2[14];
    assign P[73] = in1[14] ^ in2[14];
    assign G[74] = in1[13] & in2[13];
    assign P[74] = in1[13] ^ in2[13];
    assign G[75] = in1[12] & in2[12];
    assign P[75] = in1[12] ^ in2[12];
    assign G[76] = in1[11] & in2[11];
    assign P[76] = in1[11] ^ in2[11];
    assign G[77] = in1[10] & in2[10];
    assign P[77] = in1[10] ^ in2[10];
    assign G[78] = in1[9] & in2[9];
    assign P[78] = in1[9] ^ in2[9];
    assign G[79] = in1[8] & in2[8];
    assign P[79] = in1[8] ^ in2[8];
    assign G[80] = in1[7] & in2[7];
    assign P[80] = in1[7] ^ in2[7];
    assign G[81] = in1[6] & in2[6];
    assign P[81] = in1[6] ^ in2[6];
    assign G[82] = in1[5] & in2[5];
    assign P[82] = in1[5] ^ in2[5];
    assign G[83] = in1[4] & in2[4];
    assign P[83] = in1[4] ^ in2[4];
    assign G[84] = in1[3] & in2[3];
    assign P[84] = in1[3] ^ in2[3];
    assign G[85] = in1[2] & in2[2];
    assign P[85] = in1[2] ^ in2[2];
    assign G[86] = in1[1] & in2[1];
    assign P[86] = in1[1] ^ in2[1];
    assign G[87] = in1[0] & in2[0];
    assign P[87] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign cout = G[87] | (P[87] & C[87]);
    assign sum = P ^ C;
endmodule

module CLA_87(output [86:0] sum, output cout, input [86:0] in1, input [86:0] in2);

    wire[86:0] G;
    wire[86:0] C;
    wire[86:0] P;

    assign G[0] = in1[86] & in2[86];
    assign P[0] = in1[86] ^ in2[86];
    assign G[1] = in1[85] & in2[85];
    assign P[1] = in1[85] ^ in2[85];
    assign G[2] = in1[84] & in2[84];
    assign P[2] = in1[84] ^ in2[84];
    assign G[3] = in1[83] & in2[83];
    assign P[3] = in1[83] ^ in2[83];
    assign G[4] = in1[82] & in2[82];
    assign P[4] = in1[82] ^ in2[82];
    assign G[5] = in1[81] & in2[81];
    assign P[5] = in1[81] ^ in2[81];
    assign G[6] = in1[80] & in2[80];
    assign P[6] = in1[80] ^ in2[80];
    assign G[7] = in1[79] & in2[79];
    assign P[7] = in1[79] ^ in2[79];
    assign G[8] = in1[78] & in2[78];
    assign P[8] = in1[78] ^ in2[78];
    assign G[9] = in1[77] & in2[77];
    assign P[9] = in1[77] ^ in2[77];
    assign G[10] = in1[76] & in2[76];
    assign P[10] = in1[76] ^ in2[76];
    assign G[11] = in1[75] & in2[75];
    assign P[11] = in1[75] ^ in2[75];
    assign G[12] = in1[74] & in2[74];
    assign P[12] = in1[74] ^ in2[74];
    assign G[13] = in1[73] & in2[73];
    assign P[13] = in1[73] ^ in2[73];
    assign G[14] = in1[72] & in2[72];
    assign P[14] = in1[72] ^ in2[72];
    assign G[15] = in1[71] & in2[71];
    assign P[15] = in1[71] ^ in2[71];
    assign G[16] = in1[70] & in2[70];
    assign P[16] = in1[70] ^ in2[70];
    assign G[17] = in1[69] & in2[69];
    assign P[17] = in1[69] ^ in2[69];
    assign G[18] = in1[68] & in2[68];
    assign P[18] = in1[68] ^ in2[68];
    assign G[19] = in1[67] & in2[67];
    assign P[19] = in1[67] ^ in2[67];
    assign G[20] = in1[66] & in2[66];
    assign P[20] = in1[66] ^ in2[66];
    assign G[21] = in1[65] & in2[65];
    assign P[21] = in1[65] ^ in2[65];
    assign G[22] = in1[64] & in2[64];
    assign P[22] = in1[64] ^ in2[64];
    assign G[23] = in1[63] & in2[63];
    assign P[23] = in1[63] ^ in2[63];
    assign G[24] = in1[62] & in2[62];
    assign P[24] = in1[62] ^ in2[62];
    assign G[25] = in1[61] & in2[61];
    assign P[25] = in1[61] ^ in2[61];
    assign G[26] = in1[60] & in2[60];
    assign P[26] = in1[60] ^ in2[60];
    assign G[27] = in1[59] & in2[59];
    assign P[27] = in1[59] ^ in2[59];
    assign G[28] = in1[58] & in2[58];
    assign P[28] = in1[58] ^ in2[58];
    assign G[29] = in1[57] & in2[57];
    assign P[29] = in1[57] ^ in2[57];
    assign G[30] = in1[56] & in2[56];
    assign P[30] = in1[56] ^ in2[56];
    assign G[31] = in1[55] & in2[55];
    assign P[31] = in1[55] ^ in2[55];
    assign G[32] = in1[54] & in2[54];
    assign P[32] = in1[54] ^ in2[54];
    assign G[33] = in1[53] & in2[53];
    assign P[33] = in1[53] ^ in2[53];
    assign G[34] = in1[52] & in2[52];
    assign P[34] = in1[52] ^ in2[52];
    assign G[35] = in1[51] & in2[51];
    assign P[35] = in1[51] ^ in2[51];
    assign G[36] = in1[50] & in2[50];
    assign P[36] = in1[50] ^ in2[50];
    assign G[37] = in1[49] & in2[49];
    assign P[37] = in1[49] ^ in2[49];
    assign G[38] = in1[48] & in2[48];
    assign P[38] = in1[48] ^ in2[48];
    assign G[39] = in1[47] & in2[47];
    assign P[39] = in1[47] ^ in2[47];
    assign G[40] = in1[46] & in2[46];
    assign P[40] = in1[46] ^ in2[46];
    assign G[41] = in1[45] & in2[45];
    assign P[41] = in1[45] ^ in2[45];
    assign G[42] = in1[44] & in2[44];
    assign P[42] = in1[44] ^ in2[44];
    assign G[43] = in1[43] & in2[43];
    assign P[43] = in1[43] ^ in2[43];
    assign G[44] = in1[42] & in2[42];
    assign P[44] = in1[42] ^ in2[42];
    assign G[45] = in1[41] & in2[41];
    assign P[45] = in1[41] ^ in2[41];
    assign G[46] = in1[40] & in2[40];
    assign P[46] = in1[40] ^ in2[40];
    assign G[47] = in1[39] & in2[39];
    assign P[47] = in1[39] ^ in2[39];
    assign G[48] = in1[38] & in2[38];
    assign P[48] = in1[38] ^ in2[38];
    assign G[49] = in1[37] & in2[37];
    assign P[49] = in1[37] ^ in2[37];
    assign G[50] = in1[36] & in2[36];
    assign P[50] = in1[36] ^ in2[36];
    assign G[51] = in1[35] & in2[35];
    assign P[51] = in1[35] ^ in2[35];
    assign G[52] = in1[34] & in2[34];
    assign P[52] = in1[34] ^ in2[34];
    assign G[53] = in1[33] & in2[33];
    assign P[53] = in1[33] ^ in2[33];
    assign G[54] = in1[32] & in2[32];
    assign P[54] = in1[32] ^ in2[32];
    assign G[55] = in1[31] & in2[31];
    assign P[55] = in1[31] ^ in2[31];
    assign G[56] = in1[30] & in2[30];
    assign P[56] = in1[30] ^ in2[30];
    assign G[57] = in1[29] & in2[29];
    assign P[57] = in1[29] ^ in2[29];
    assign G[58] = in1[28] & in2[28];
    assign P[58] = in1[28] ^ in2[28];
    assign G[59] = in1[27] & in2[27];
    assign P[59] = in1[27] ^ in2[27];
    assign G[60] = in1[26] & in2[26];
    assign P[60] = in1[26] ^ in2[26];
    assign G[61] = in1[25] & in2[25];
    assign P[61] = in1[25] ^ in2[25];
    assign G[62] = in1[24] & in2[24];
    assign P[62] = in1[24] ^ in2[24];
    assign G[63] = in1[23] & in2[23];
    assign P[63] = in1[23] ^ in2[23];
    assign G[64] = in1[22] & in2[22];
    assign P[64] = in1[22] ^ in2[22];
    assign G[65] = in1[21] & in2[21];
    assign P[65] = in1[21] ^ in2[21];
    assign G[66] = in1[20] & in2[20];
    assign P[66] = in1[20] ^ in2[20];
    assign G[67] = in1[19] & in2[19];
    assign P[67] = in1[19] ^ in2[19];
    assign G[68] = in1[18] & in2[18];
    assign P[68] = in1[18] ^ in2[18];
    assign G[69] = in1[17] & in2[17];
    assign P[69] = in1[17] ^ in2[17];
    assign G[70] = in1[16] & in2[16];
    assign P[70] = in1[16] ^ in2[16];
    assign G[71] = in1[15] & in2[15];
    assign P[71] = in1[15] ^ in2[15];
    assign G[72] = in1[14] & in2[14];
    assign P[72] = in1[14] ^ in2[14];
    assign G[73] = in1[13] & in2[13];
    assign P[73] = in1[13] ^ in2[13];
    assign G[74] = in1[12] & in2[12];
    assign P[74] = in1[12] ^ in2[12];
    assign G[75] = in1[11] & in2[11];
    assign P[75] = in1[11] ^ in2[11];
    assign G[76] = in1[10] & in2[10];
    assign P[76] = in1[10] ^ in2[10];
    assign G[77] = in1[9] & in2[9];
    assign P[77] = in1[9] ^ in2[9];
    assign G[78] = in1[8] & in2[8];
    assign P[78] = in1[8] ^ in2[8];
    assign G[79] = in1[7] & in2[7];
    assign P[79] = in1[7] ^ in2[7];
    assign G[80] = in1[6] & in2[6];
    assign P[80] = in1[6] ^ in2[6];
    assign G[81] = in1[5] & in2[5];
    assign P[81] = in1[5] ^ in2[5];
    assign G[82] = in1[4] & in2[4];
    assign P[82] = in1[4] ^ in2[4];
    assign G[83] = in1[3] & in2[3];
    assign P[83] = in1[3] ^ in2[3];
    assign G[84] = in1[2] & in2[2];
    assign P[84] = in1[2] ^ in2[2];
    assign G[85] = in1[1] & in2[1];
    assign P[85] = in1[1] ^ in2[1];
    assign G[86] = in1[0] & in2[0];
    assign P[86] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign cout = G[86] | (P[86] & C[86]);
    assign sum = P ^ C;
endmodule

module CLA_86(output [85:0] sum, output cout, input [85:0] in1, input [85:0] in2);

    wire[85:0] G;
    wire[85:0] C;
    wire[85:0] P;

    assign G[0] = in1[85] & in2[85];
    assign P[0] = in1[85] ^ in2[85];
    assign G[1] = in1[84] & in2[84];
    assign P[1] = in1[84] ^ in2[84];
    assign G[2] = in1[83] & in2[83];
    assign P[2] = in1[83] ^ in2[83];
    assign G[3] = in1[82] & in2[82];
    assign P[3] = in1[82] ^ in2[82];
    assign G[4] = in1[81] & in2[81];
    assign P[4] = in1[81] ^ in2[81];
    assign G[5] = in1[80] & in2[80];
    assign P[5] = in1[80] ^ in2[80];
    assign G[6] = in1[79] & in2[79];
    assign P[6] = in1[79] ^ in2[79];
    assign G[7] = in1[78] & in2[78];
    assign P[7] = in1[78] ^ in2[78];
    assign G[8] = in1[77] & in2[77];
    assign P[8] = in1[77] ^ in2[77];
    assign G[9] = in1[76] & in2[76];
    assign P[9] = in1[76] ^ in2[76];
    assign G[10] = in1[75] & in2[75];
    assign P[10] = in1[75] ^ in2[75];
    assign G[11] = in1[74] & in2[74];
    assign P[11] = in1[74] ^ in2[74];
    assign G[12] = in1[73] & in2[73];
    assign P[12] = in1[73] ^ in2[73];
    assign G[13] = in1[72] & in2[72];
    assign P[13] = in1[72] ^ in2[72];
    assign G[14] = in1[71] & in2[71];
    assign P[14] = in1[71] ^ in2[71];
    assign G[15] = in1[70] & in2[70];
    assign P[15] = in1[70] ^ in2[70];
    assign G[16] = in1[69] & in2[69];
    assign P[16] = in1[69] ^ in2[69];
    assign G[17] = in1[68] & in2[68];
    assign P[17] = in1[68] ^ in2[68];
    assign G[18] = in1[67] & in2[67];
    assign P[18] = in1[67] ^ in2[67];
    assign G[19] = in1[66] & in2[66];
    assign P[19] = in1[66] ^ in2[66];
    assign G[20] = in1[65] & in2[65];
    assign P[20] = in1[65] ^ in2[65];
    assign G[21] = in1[64] & in2[64];
    assign P[21] = in1[64] ^ in2[64];
    assign G[22] = in1[63] & in2[63];
    assign P[22] = in1[63] ^ in2[63];
    assign G[23] = in1[62] & in2[62];
    assign P[23] = in1[62] ^ in2[62];
    assign G[24] = in1[61] & in2[61];
    assign P[24] = in1[61] ^ in2[61];
    assign G[25] = in1[60] & in2[60];
    assign P[25] = in1[60] ^ in2[60];
    assign G[26] = in1[59] & in2[59];
    assign P[26] = in1[59] ^ in2[59];
    assign G[27] = in1[58] & in2[58];
    assign P[27] = in1[58] ^ in2[58];
    assign G[28] = in1[57] & in2[57];
    assign P[28] = in1[57] ^ in2[57];
    assign G[29] = in1[56] & in2[56];
    assign P[29] = in1[56] ^ in2[56];
    assign G[30] = in1[55] & in2[55];
    assign P[30] = in1[55] ^ in2[55];
    assign G[31] = in1[54] & in2[54];
    assign P[31] = in1[54] ^ in2[54];
    assign G[32] = in1[53] & in2[53];
    assign P[32] = in1[53] ^ in2[53];
    assign G[33] = in1[52] & in2[52];
    assign P[33] = in1[52] ^ in2[52];
    assign G[34] = in1[51] & in2[51];
    assign P[34] = in1[51] ^ in2[51];
    assign G[35] = in1[50] & in2[50];
    assign P[35] = in1[50] ^ in2[50];
    assign G[36] = in1[49] & in2[49];
    assign P[36] = in1[49] ^ in2[49];
    assign G[37] = in1[48] & in2[48];
    assign P[37] = in1[48] ^ in2[48];
    assign G[38] = in1[47] & in2[47];
    assign P[38] = in1[47] ^ in2[47];
    assign G[39] = in1[46] & in2[46];
    assign P[39] = in1[46] ^ in2[46];
    assign G[40] = in1[45] & in2[45];
    assign P[40] = in1[45] ^ in2[45];
    assign G[41] = in1[44] & in2[44];
    assign P[41] = in1[44] ^ in2[44];
    assign G[42] = in1[43] & in2[43];
    assign P[42] = in1[43] ^ in2[43];
    assign G[43] = in1[42] & in2[42];
    assign P[43] = in1[42] ^ in2[42];
    assign G[44] = in1[41] & in2[41];
    assign P[44] = in1[41] ^ in2[41];
    assign G[45] = in1[40] & in2[40];
    assign P[45] = in1[40] ^ in2[40];
    assign G[46] = in1[39] & in2[39];
    assign P[46] = in1[39] ^ in2[39];
    assign G[47] = in1[38] & in2[38];
    assign P[47] = in1[38] ^ in2[38];
    assign G[48] = in1[37] & in2[37];
    assign P[48] = in1[37] ^ in2[37];
    assign G[49] = in1[36] & in2[36];
    assign P[49] = in1[36] ^ in2[36];
    assign G[50] = in1[35] & in2[35];
    assign P[50] = in1[35] ^ in2[35];
    assign G[51] = in1[34] & in2[34];
    assign P[51] = in1[34] ^ in2[34];
    assign G[52] = in1[33] & in2[33];
    assign P[52] = in1[33] ^ in2[33];
    assign G[53] = in1[32] & in2[32];
    assign P[53] = in1[32] ^ in2[32];
    assign G[54] = in1[31] & in2[31];
    assign P[54] = in1[31] ^ in2[31];
    assign G[55] = in1[30] & in2[30];
    assign P[55] = in1[30] ^ in2[30];
    assign G[56] = in1[29] & in2[29];
    assign P[56] = in1[29] ^ in2[29];
    assign G[57] = in1[28] & in2[28];
    assign P[57] = in1[28] ^ in2[28];
    assign G[58] = in1[27] & in2[27];
    assign P[58] = in1[27] ^ in2[27];
    assign G[59] = in1[26] & in2[26];
    assign P[59] = in1[26] ^ in2[26];
    assign G[60] = in1[25] & in2[25];
    assign P[60] = in1[25] ^ in2[25];
    assign G[61] = in1[24] & in2[24];
    assign P[61] = in1[24] ^ in2[24];
    assign G[62] = in1[23] & in2[23];
    assign P[62] = in1[23] ^ in2[23];
    assign G[63] = in1[22] & in2[22];
    assign P[63] = in1[22] ^ in2[22];
    assign G[64] = in1[21] & in2[21];
    assign P[64] = in1[21] ^ in2[21];
    assign G[65] = in1[20] & in2[20];
    assign P[65] = in1[20] ^ in2[20];
    assign G[66] = in1[19] & in2[19];
    assign P[66] = in1[19] ^ in2[19];
    assign G[67] = in1[18] & in2[18];
    assign P[67] = in1[18] ^ in2[18];
    assign G[68] = in1[17] & in2[17];
    assign P[68] = in1[17] ^ in2[17];
    assign G[69] = in1[16] & in2[16];
    assign P[69] = in1[16] ^ in2[16];
    assign G[70] = in1[15] & in2[15];
    assign P[70] = in1[15] ^ in2[15];
    assign G[71] = in1[14] & in2[14];
    assign P[71] = in1[14] ^ in2[14];
    assign G[72] = in1[13] & in2[13];
    assign P[72] = in1[13] ^ in2[13];
    assign G[73] = in1[12] & in2[12];
    assign P[73] = in1[12] ^ in2[12];
    assign G[74] = in1[11] & in2[11];
    assign P[74] = in1[11] ^ in2[11];
    assign G[75] = in1[10] & in2[10];
    assign P[75] = in1[10] ^ in2[10];
    assign G[76] = in1[9] & in2[9];
    assign P[76] = in1[9] ^ in2[9];
    assign G[77] = in1[8] & in2[8];
    assign P[77] = in1[8] ^ in2[8];
    assign G[78] = in1[7] & in2[7];
    assign P[78] = in1[7] ^ in2[7];
    assign G[79] = in1[6] & in2[6];
    assign P[79] = in1[6] ^ in2[6];
    assign G[80] = in1[5] & in2[5];
    assign P[80] = in1[5] ^ in2[5];
    assign G[81] = in1[4] & in2[4];
    assign P[81] = in1[4] ^ in2[4];
    assign G[82] = in1[3] & in2[3];
    assign P[82] = in1[3] ^ in2[3];
    assign G[83] = in1[2] & in2[2];
    assign P[83] = in1[2] ^ in2[2];
    assign G[84] = in1[1] & in2[1];
    assign P[84] = in1[1] ^ in2[1];
    assign G[85] = in1[0] & in2[0];
    assign P[85] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign cout = G[85] | (P[85] & C[85]);
    assign sum = P ^ C;
endmodule

module CLA_85(output [84:0] sum, output cout, input [84:0] in1, input [84:0] in2);

    wire[84:0] G;
    wire[84:0] C;
    wire[84:0] P;

    assign G[0] = in1[84] & in2[84];
    assign P[0] = in1[84] ^ in2[84];
    assign G[1] = in1[83] & in2[83];
    assign P[1] = in1[83] ^ in2[83];
    assign G[2] = in1[82] & in2[82];
    assign P[2] = in1[82] ^ in2[82];
    assign G[3] = in1[81] & in2[81];
    assign P[3] = in1[81] ^ in2[81];
    assign G[4] = in1[80] & in2[80];
    assign P[4] = in1[80] ^ in2[80];
    assign G[5] = in1[79] & in2[79];
    assign P[5] = in1[79] ^ in2[79];
    assign G[6] = in1[78] & in2[78];
    assign P[6] = in1[78] ^ in2[78];
    assign G[7] = in1[77] & in2[77];
    assign P[7] = in1[77] ^ in2[77];
    assign G[8] = in1[76] & in2[76];
    assign P[8] = in1[76] ^ in2[76];
    assign G[9] = in1[75] & in2[75];
    assign P[9] = in1[75] ^ in2[75];
    assign G[10] = in1[74] & in2[74];
    assign P[10] = in1[74] ^ in2[74];
    assign G[11] = in1[73] & in2[73];
    assign P[11] = in1[73] ^ in2[73];
    assign G[12] = in1[72] & in2[72];
    assign P[12] = in1[72] ^ in2[72];
    assign G[13] = in1[71] & in2[71];
    assign P[13] = in1[71] ^ in2[71];
    assign G[14] = in1[70] & in2[70];
    assign P[14] = in1[70] ^ in2[70];
    assign G[15] = in1[69] & in2[69];
    assign P[15] = in1[69] ^ in2[69];
    assign G[16] = in1[68] & in2[68];
    assign P[16] = in1[68] ^ in2[68];
    assign G[17] = in1[67] & in2[67];
    assign P[17] = in1[67] ^ in2[67];
    assign G[18] = in1[66] & in2[66];
    assign P[18] = in1[66] ^ in2[66];
    assign G[19] = in1[65] & in2[65];
    assign P[19] = in1[65] ^ in2[65];
    assign G[20] = in1[64] & in2[64];
    assign P[20] = in1[64] ^ in2[64];
    assign G[21] = in1[63] & in2[63];
    assign P[21] = in1[63] ^ in2[63];
    assign G[22] = in1[62] & in2[62];
    assign P[22] = in1[62] ^ in2[62];
    assign G[23] = in1[61] & in2[61];
    assign P[23] = in1[61] ^ in2[61];
    assign G[24] = in1[60] & in2[60];
    assign P[24] = in1[60] ^ in2[60];
    assign G[25] = in1[59] & in2[59];
    assign P[25] = in1[59] ^ in2[59];
    assign G[26] = in1[58] & in2[58];
    assign P[26] = in1[58] ^ in2[58];
    assign G[27] = in1[57] & in2[57];
    assign P[27] = in1[57] ^ in2[57];
    assign G[28] = in1[56] & in2[56];
    assign P[28] = in1[56] ^ in2[56];
    assign G[29] = in1[55] & in2[55];
    assign P[29] = in1[55] ^ in2[55];
    assign G[30] = in1[54] & in2[54];
    assign P[30] = in1[54] ^ in2[54];
    assign G[31] = in1[53] & in2[53];
    assign P[31] = in1[53] ^ in2[53];
    assign G[32] = in1[52] & in2[52];
    assign P[32] = in1[52] ^ in2[52];
    assign G[33] = in1[51] & in2[51];
    assign P[33] = in1[51] ^ in2[51];
    assign G[34] = in1[50] & in2[50];
    assign P[34] = in1[50] ^ in2[50];
    assign G[35] = in1[49] & in2[49];
    assign P[35] = in1[49] ^ in2[49];
    assign G[36] = in1[48] & in2[48];
    assign P[36] = in1[48] ^ in2[48];
    assign G[37] = in1[47] & in2[47];
    assign P[37] = in1[47] ^ in2[47];
    assign G[38] = in1[46] & in2[46];
    assign P[38] = in1[46] ^ in2[46];
    assign G[39] = in1[45] & in2[45];
    assign P[39] = in1[45] ^ in2[45];
    assign G[40] = in1[44] & in2[44];
    assign P[40] = in1[44] ^ in2[44];
    assign G[41] = in1[43] & in2[43];
    assign P[41] = in1[43] ^ in2[43];
    assign G[42] = in1[42] & in2[42];
    assign P[42] = in1[42] ^ in2[42];
    assign G[43] = in1[41] & in2[41];
    assign P[43] = in1[41] ^ in2[41];
    assign G[44] = in1[40] & in2[40];
    assign P[44] = in1[40] ^ in2[40];
    assign G[45] = in1[39] & in2[39];
    assign P[45] = in1[39] ^ in2[39];
    assign G[46] = in1[38] & in2[38];
    assign P[46] = in1[38] ^ in2[38];
    assign G[47] = in1[37] & in2[37];
    assign P[47] = in1[37] ^ in2[37];
    assign G[48] = in1[36] & in2[36];
    assign P[48] = in1[36] ^ in2[36];
    assign G[49] = in1[35] & in2[35];
    assign P[49] = in1[35] ^ in2[35];
    assign G[50] = in1[34] & in2[34];
    assign P[50] = in1[34] ^ in2[34];
    assign G[51] = in1[33] & in2[33];
    assign P[51] = in1[33] ^ in2[33];
    assign G[52] = in1[32] & in2[32];
    assign P[52] = in1[32] ^ in2[32];
    assign G[53] = in1[31] & in2[31];
    assign P[53] = in1[31] ^ in2[31];
    assign G[54] = in1[30] & in2[30];
    assign P[54] = in1[30] ^ in2[30];
    assign G[55] = in1[29] & in2[29];
    assign P[55] = in1[29] ^ in2[29];
    assign G[56] = in1[28] & in2[28];
    assign P[56] = in1[28] ^ in2[28];
    assign G[57] = in1[27] & in2[27];
    assign P[57] = in1[27] ^ in2[27];
    assign G[58] = in1[26] & in2[26];
    assign P[58] = in1[26] ^ in2[26];
    assign G[59] = in1[25] & in2[25];
    assign P[59] = in1[25] ^ in2[25];
    assign G[60] = in1[24] & in2[24];
    assign P[60] = in1[24] ^ in2[24];
    assign G[61] = in1[23] & in2[23];
    assign P[61] = in1[23] ^ in2[23];
    assign G[62] = in1[22] & in2[22];
    assign P[62] = in1[22] ^ in2[22];
    assign G[63] = in1[21] & in2[21];
    assign P[63] = in1[21] ^ in2[21];
    assign G[64] = in1[20] & in2[20];
    assign P[64] = in1[20] ^ in2[20];
    assign G[65] = in1[19] & in2[19];
    assign P[65] = in1[19] ^ in2[19];
    assign G[66] = in1[18] & in2[18];
    assign P[66] = in1[18] ^ in2[18];
    assign G[67] = in1[17] & in2[17];
    assign P[67] = in1[17] ^ in2[17];
    assign G[68] = in1[16] & in2[16];
    assign P[68] = in1[16] ^ in2[16];
    assign G[69] = in1[15] & in2[15];
    assign P[69] = in1[15] ^ in2[15];
    assign G[70] = in1[14] & in2[14];
    assign P[70] = in1[14] ^ in2[14];
    assign G[71] = in1[13] & in2[13];
    assign P[71] = in1[13] ^ in2[13];
    assign G[72] = in1[12] & in2[12];
    assign P[72] = in1[12] ^ in2[12];
    assign G[73] = in1[11] & in2[11];
    assign P[73] = in1[11] ^ in2[11];
    assign G[74] = in1[10] & in2[10];
    assign P[74] = in1[10] ^ in2[10];
    assign G[75] = in1[9] & in2[9];
    assign P[75] = in1[9] ^ in2[9];
    assign G[76] = in1[8] & in2[8];
    assign P[76] = in1[8] ^ in2[8];
    assign G[77] = in1[7] & in2[7];
    assign P[77] = in1[7] ^ in2[7];
    assign G[78] = in1[6] & in2[6];
    assign P[78] = in1[6] ^ in2[6];
    assign G[79] = in1[5] & in2[5];
    assign P[79] = in1[5] ^ in2[5];
    assign G[80] = in1[4] & in2[4];
    assign P[80] = in1[4] ^ in2[4];
    assign G[81] = in1[3] & in2[3];
    assign P[81] = in1[3] ^ in2[3];
    assign G[82] = in1[2] & in2[2];
    assign P[82] = in1[2] ^ in2[2];
    assign G[83] = in1[1] & in2[1];
    assign P[83] = in1[1] ^ in2[1];
    assign G[84] = in1[0] & in2[0];
    assign P[84] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign cout = G[84] | (P[84] & C[84]);
    assign sum = P ^ C;
endmodule

module CLA_84(output [83:0] sum, output cout, input [83:0] in1, input [83:0] in2);

    wire[83:0] G;
    wire[83:0] C;
    wire[83:0] P;

    assign G[0] = in1[83] & in2[83];
    assign P[0] = in1[83] ^ in2[83];
    assign G[1] = in1[82] & in2[82];
    assign P[1] = in1[82] ^ in2[82];
    assign G[2] = in1[81] & in2[81];
    assign P[2] = in1[81] ^ in2[81];
    assign G[3] = in1[80] & in2[80];
    assign P[3] = in1[80] ^ in2[80];
    assign G[4] = in1[79] & in2[79];
    assign P[4] = in1[79] ^ in2[79];
    assign G[5] = in1[78] & in2[78];
    assign P[5] = in1[78] ^ in2[78];
    assign G[6] = in1[77] & in2[77];
    assign P[6] = in1[77] ^ in2[77];
    assign G[7] = in1[76] & in2[76];
    assign P[7] = in1[76] ^ in2[76];
    assign G[8] = in1[75] & in2[75];
    assign P[8] = in1[75] ^ in2[75];
    assign G[9] = in1[74] & in2[74];
    assign P[9] = in1[74] ^ in2[74];
    assign G[10] = in1[73] & in2[73];
    assign P[10] = in1[73] ^ in2[73];
    assign G[11] = in1[72] & in2[72];
    assign P[11] = in1[72] ^ in2[72];
    assign G[12] = in1[71] & in2[71];
    assign P[12] = in1[71] ^ in2[71];
    assign G[13] = in1[70] & in2[70];
    assign P[13] = in1[70] ^ in2[70];
    assign G[14] = in1[69] & in2[69];
    assign P[14] = in1[69] ^ in2[69];
    assign G[15] = in1[68] & in2[68];
    assign P[15] = in1[68] ^ in2[68];
    assign G[16] = in1[67] & in2[67];
    assign P[16] = in1[67] ^ in2[67];
    assign G[17] = in1[66] & in2[66];
    assign P[17] = in1[66] ^ in2[66];
    assign G[18] = in1[65] & in2[65];
    assign P[18] = in1[65] ^ in2[65];
    assign G[19] = in1[64] & in2[64];
    assign P[19] = in1[64] ^ in2[64];
    assign G[20] = in1[63] & in2[63];
    assign P[20] = in1[63] ^ in2[63];
    assign G[21] = in1[62] & in2[62];
    assign P[21] = in1[62] ^ in2[62];
    assign G[22] = in1[61] & in2[61];
    assign P[22] = in1[61] ^ in2[61];
    assign G[23] = in1[60] & in2[60];
    assign P[23] = in1[60] ^ in2[60];
    assign G[24] = in1[59] & in2[59];
    assign P[24] = in1[59] ^ in2[59];
    assign G[25] = in1[58] & in2[58];
    assign P[25] = in1[58] ^ in2[58];
    assign G[26] = in1[57] & in2[57];
    assign P[26] = in1[57] ^ in2[57];
    assign G[27] = in1[56] & in2[56];
    assign P[27] = in1[56] ^ in2[56];
    assign G[28] = in1[55] & in2[55];
    assign P[28] = in1[55] ^ in2[55];
    assign G[29] = in1[54] & in2[54];
    assign P[29] = in1[54] ^ in2[54];
    assign G[30] = in1[53] & in2[53];
    assign P[30] = in1[53] ^ in2[53];
    assign G[31] = in1[52] & in2[52];
    assign P[31] = in1[52] ^ in2[52];
    assign G[32] = in1[51] & in2[51];
    assign P[32] = in1[51] ^ in2[51];
    assign G[33] = in1[50] & in2[50];
    assign P[33] = in1[50] ^ in2[50];
    assign G[34] = in1[49] & in2[49];
    assign P[34] = in1[49] ^ in2[49];
    assign G[35] = in1[48] & in2[48];
    assign P[35] = in1[48] ^ in2[48];
    assign G[36] = in1[47] & in2[47];
    assign P[36] = in1[47] ^ in2[47];
    assign G[37] = in1[46] & in2[46];
    assign P[37] = in1[46] ^ in2[46];
    assign G[38] = in1[45] & in2[45];
    assign P[38] = in1[45] ^ in2[45];
    assign G[39] = in1[44] & in2[44];
    assign P[39] = in1[44] ^ in2[44];
    assign G[40] = in1[43] & in2[43];
    assign P[40] = in1[43] ^ in2[43];
    assign G[41] = in1[42] & in2[42];
    assign P[41] = in1[42] ^ in2[42];
    assign G[42] = in1[41] & in2[41];
    assign P[42] = in1[41] ^ in2[41];
    assign G[43] = in1[40] & in2[40];
    assign P[43] = in1[40] ^ in2[40];
    assign G[44] = in1[39] & in2[39];
    assign P[44] = in1[39] ^ in2[39];
    assign G[45] = in1[38] & in2[38];
    assign P[45] = in1[38] ^ in2[38];
    assign G[46] = in1[37] & in2[37];
    assign P[46] = in1[37] ^ in2[37];
    assign G[47] = in1[36] & in2[36];
    assign P[47] = in1[36] ^ in2[36];
    assign G[48] = in1[35] & in2[35];
    assign P[48] = in1[35] ^ in2[35];
    assign G[49] = in1[34] & in2[34];
    assign P[49] = in1[34] ^ in2[34];
    assign G[50] = in1[33] & in2[33];
    assign P[50] = in1[33] ^ in2[33];
    assign G[51] = in1[32] & in2[32];
    assign P[51] = in1[32] ^ in2[32];
    assign G[52] = in1[31] & in2[31];
    assign P[52] = in1[31] ^ in2[31];
    assign G[53] = in1[30] & in2[30];
    assign P[53] = in1[30] ^ in2[30];
    assign G[54] = in1[29] & in2[29];
    assign P[54] = in1[29] ^ in2[29];
    assign G[55] = in1[28] & in2[28];
    assign P[55] = in1[28] ^ in2[28];
    assign G[56] = in1[27] & in2[27];
    assign P[56] = in1[27] ^ in2[27];
    assign G[57] = in1[26] & in2[26];
    assign P[57] = in1[26] ^ in2[26];
    assign G[58] = in1[25] & in2[25];
    assign P[58] = in1[25] ^ in2[25];
    assign G[59] = in1[24] & in2[24];
    assign P[59] = in1[24] ^ in2[24];
    assign G[60] = in1[23] & in2[23];
    assign P[60] = in1[23] ^ in2[23];
    assign G[61] = in1[22] & in2[22];
    assign P[61] = in1[22] ^ in2[22];
    assign G[62] = in1[21] & in2[21];
    assign P[62] = in1[21] ^ in2[21];
    assign G[63] = in1[20] & in2[20];
    assign P[63] = in1[20] ^ in2[20];
    assign G[64] = in1[19] & in2[19];
    assign P[64] = in1[19] ^ in2[19];
    assign G[65] = in1[18] & in2[18];
    assign P[65] = in1[18] ^ in2[18];
    assign G[66] = in1[17] & in2[17];
    assign P[66] = in1[17] ^ in2[17];
    assign G[67] = in1[16] & in2[16];
    assign P[67] = in1[16] ^ in2[16];
    assign G[68] = in1[15] & in2[15];
    assign P[68] = in1[15] ^ in2[15];
    assign G[69] = in1[14] & in2[14];
    assign P[69] = in1[14] ^ in2[14];
    assign G[70] = in1[13] & in2[13];
    assign P[70] = in1[13] ^ in2[13];
    assign G[71] = in1[12] & in2[12];
    assign P[71] = in1[12] ^ in2[12];
    assign G[72] = in1[11] & in2[11];
    assign P[72] = in1[11] ^ in2[11];
    assign G[73] = in1[10] & in2[10];
    assign P[73] = in1[10] ^ in2[10];
    assign G[74] = in1[9] & in2[9];
    assign P[74] = in1[9] ^ in2[9];
    assign G[75] = in1[8] & in2[8];
    assign P[75] = in1[8] ^ in2[8];
    assign G[76] = in1[7] & in2[7];
    assign P[76] = in1[7] ^ in2[7];
    assign G[77] = in1[6] & in2[6];
    assign P[77] = in1[6] ^ in2[6];
    assign G[78] = in1[5] & in2[5];
    assign P[78] = in1[5] ^ in2[5];
    assign G[79] = in1[4] & in2[4];
    assign P[79] = in1[4] ^ in2[4];
    assign G[80] = in1[3] & in2[3];
    assign P[80] = in1[3] ^ in2[3];
    assign G[81] = in1[2] & in2[2];
    assign P[81] = in1[2] ^ in2[2];
    assign G[82] = in1[1] & in2[1];
    assign P[82] = in1[1] ^ in2[1];
    assign G[83] = in1[0] & in2[0];
    assign P[83] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign cout = G[83] | (P[83] & C[83]);
    assign sum = P ^ C;
endmodule

module CLA_83(output [82:0] sum, output cout, input [82:0] in1, input [82:0] in2);

    wire[82:0] G;
    wire[82:0] C;
    wire[82:0] P;

    assign G[0] = in1[82] & in2[82];
    assign P[0] = in1[82] ^ in2[82];
    assign G[1] = in1[81] & in2[81];
    assign P[1] = in1[81] ^ in2[81];
    assign G[2] = in1[80] & in2[80];
    assign P[2] = in1[80] ^ in2[80];
    assign G[3] = in1[79] & in2[79];
    assign P[3] = in1[79] ^ in2[79];
    assign G[4] = in1[78] & in2[78];
    assign P[4] = in1[78] ^ in2[78];
    assign G[5] = in1[77] & in2[77];
    assign P[5] = in1[77] ^ in2[77];
    assign G[6] = in1[76] & in2[76];
    assign P[6] = in1[76] ^ in2[76];
    assign G[7] = in1[75] & in2[75];
    assign P[7] = in1[75] ^ in2[75];
    assign G[8] = in1[74] & in2[74];
    assign P[8] = in1[74] ^ in2[74];
    assign G[9] = in1[73] & in2[73];
    assign P[9] = in1[73] ^ in2[73];
    assign G[10] = in1[72] & in2[72];
    assign P[10] = in1[72] ^ in2[72];
    assign G[11] = in1[71] & in2[71];
    assign P[11] = in1[71] ^ in2[71];
    assign G[12] = in1[70] & in2[70];
    assign P[12] = in1[70] ^ in2[70];
    assign G[13] = in1[69] & in2[69];
    assign P[13] = in1[69] ^ in2[69];
    assign G[14] = in1[68] & in2[68];
    assign P[14] = in1[68] ^ in2[68];
    assign G[15] = in1[67] & in2[67];
    assign P[15] = in1[67] ^ in2[67];
    assign G[16] = in1[66] & in2[66];
    assign P[16] = in1[66] ^ in2[66];
    assign G[17] = in1[65] & in2[65];
    assign P[17] = in1[65] ^ in2[65];
    assign G[18] = in1[64] & in2[64];
    assign P[18] = in1[64] ^ in2[64];
    assign G[19] = in1[63] & in2[63];
    assign P[19] = in1[63] ^ in2[63];
    assign G[20] = in1[62] & in2[62];
    assign P[20] = in1[62] ^ in2[62];
    assign G[21] = in1[61] & in2[61];
    assign P[21] = in1[61] ^ in2[61];
    assign G[22] = in1[60] & in2[60];
    assign P[22] = in1[60] ^ in2[60];
    assign G[23] = in1[59] & in2[59];
    assign P[23] = in1[59] ^ in2[59];
    assign G[24] = in1[58] & in2[58];
    assign P[24] = in1[58] ^ in2[58];
    assign G[25] = in1[57] & in2[57];
    assign P[25] = in1[57] ^ in2[57];
    assign G[26] = in1[56] & in2[56];
    assign P[26] = in1[56] ^ in2[56];
    assign G[27] = in1[55] & in2[55];
    assign P[27] = in1[55] ^ in2[55];
    assign G[28] = in1[54] & in2[54];
    assign P[28] = in1[54] ^ in2[54];
    assign G[29] = in1[53] & in2[53];
    assign P[29] = in1[53] ^ in2[53];
    assign G[30] = in1[52] & in2[52];
    assign P[30] = in1[52] ^ in2[52];
    assign G[31] = in1[51] & in2[51];
    assign P[31] = in1[51] ^ in2[51];
    assign G[32] = in1[50] & in2[50];
    assign P[32] = in1[50] ^ in2[50];
    assign G[33] = in1[49] & in2[49];
    assign P[33] = in1[49] ^ in2[49];
    assign G[34] = in1[48] & in2[48];
    assign P[34] = in1[48] ^ in2[48];
    assign G[35] = in1[47] & in2[47];
    assign P[35] = in1[47] ^ in2[47];
    assign G[36] = in1[46] & in2[46];
    assign P[36] = in1[46] ^ in2[46];
    assign G[37] = in1[45] & in2[45];
    assign P[37] = in1[45] ^ in2[45];
    assign G[38] = in1[44] & in2[44];
    assign P[38] = in1[44] ^ in2[44];
    assign G[39] = in1[43] & in2[43];
    assign P[39] = in1[43] ^ in2[43];
    assign G[40] = in1[42] & in2[42];
    assign P[40] = in1[42] ^ in2[42];
    assign G[41] = in1[41] & in2[41];
    assign P[41] = in1[41] ^ in2[41];
    assign G[42] = in1[40] & in2[40];
    assign P[42] = in1[40] ^ in2[40];
    assign G[43] = in1[39] & in2[39];
    assign P[43] = in1[39] ^ in2[39];
    assign G[44] = in1[38] & in2[38];
    assign P[44] = in1[38] ^ in2[38];
    assign G[45] = in1[37] & in2[37];
    assign P[45] = in1[37] ^ in2[37];
    assign G[46] = in1[36] & in2[36];
    assign P[46] = in1[36] ^ in2[36];
    assign G[47] = in1[35] & in2[35];
    assign P[47] = in1[35] ^ in2[35];
    assign G[48] = in1[34] & in2[34];
    assign P[48] = in1[34] ^ in2[34];
    assign G[49] = in1[33] & in2[33];
    assign P[49] = in1[33] ^ in2[33];
    assign G[50] = in1[32] & in2[32];
    assign P[50] = in1[32] ^ in2[32];
    assign G[51] = in1[31] & in2[31];
    assign P[51] = in1[31] ^ in2[31];
    assign G[52] = in1[30] & in2[30];
    assign P[52] = in1[30] ^ in2[30];
    assign G[53] = in1[29] & in2[29];
    assign P[53] = in1[29] ^ in2[29];
    assign G[54] = in1[28] & in2[28];
    assign P[54] = in1[28] ^ in2[28];
    assign G[55] = in1[27] & in2[27];
    assign P[55] = in1[27] ^ in2[27];
    assign G[56] = in1[26] & in2[26];
    assign P[56] = in1[26] ^ in2[26];
    assign G[57] = in1[25] & in2[25];
    assign P[57] = in1[25] ^ in2[25];
    assign G[58] = in1[24] & in2[24];
    assign P[58] = in1[24] ^ in2[24];
    assign G[59] = in1[23] & in2[23];
    assign P[59] = in1[23] ^ in2[23];
    assign G[60] = in1[22] & in2[22];
    assign P[60] = in1[22] ^ in2[22];
    assign G[61] = in1[21] & in2[21];
    assign P[61] = in1[21] ^ in2[21];
    assign G[62] = in1[20] & in2[20];
    assign P[62] = in1[20] ^ in2[20];
    assign G[63] = in1[19] & in2[19];
    assign P[63] = in1[19] ^ in2[19];
    assign G[64] = in1[18] & in2[18];
    assign P[64] = in1[18] ^ in2[18];
    assign G[65] = in1[17] & in2[17];
    assign P[65] = in1[17] ^ in2[17];
    assign G[66] = in1[16] & in2[16];
    assign P[66] = in1[16] ^ in2[16];
    assign G[67] = in1[15] & in2[15];
    assign P[67] = in1[15] ^ in2[15];
    assign G[68] = in1[14] & in2[14];
    assign P[68] = in1[14] ^ in2[14];
    assign G[69] = in1[13] & in2[13];
    assign P[69] = in1[13] ^ in2[13];
    assign G[70] = in1[12] & in2[12];
    assign P[70] = in1[12] ^ in2[12];
    assign G[71] = in1[11] & in2[11];
    assign P[71] = in1[11] ^ in2[11];
    assign G[72] = in1[10] & in2[10];
    assign P[72] = in1[10] ^ in2[10];
    assign G[73] = in1[9] & in2[9];
    assign P[73] = in1[9] ^ in2[9];
    assign G[74] = in1[8] & in2[8];
    assign P[74] = in1[8] ^ in2[8];
    assign G[75] = in1[7] & in2[7];
    assign P[75] = in1[7] ^ in2[7];
    assign G[76] = in1[6] & in2[6];
    assign P[76] = in1[6] ^ in2[6];
    assign G[77] = in1[5] & in2[5];
    assign P[77] = in1[5] ^ in2[5];
    assign G[78] = in1[4] & in2[4];
    assign P[78] = in1[4] ^ in2[4];
    assign G[79] = in1[3] & in2[3];
    assign P[79] = in1[3] ^ in2[3];
    assign G[80] = in1[2] & in2[2];
    assign P[80] = in1[2] ^ in2[2];
    assign G[81] = in1[1] & in2[1];
    assign P[81] = in1[1] ^ in2[1];
    assign G[82] = in1[0] & in2[0];
    assign P[82] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign cout = G[82] | (P[82] & C[82]);
    assign sum = P ^ C;
endmodule

module CLA_82(output [81:0] sum, output cout, input [81:0] in1, input [81:0] in2);

    wire[81:0] G;
    wire[81:0] C;
    wire[81:0] P;

    assign G[0] = in1[81] & in2[81];
    assign P[0] = in1[81] ^ in2[81];
    assign G[1] = in1[80] & in2[80];
    assign P[1] = in1[80] ^ in2[80];
    assign G[2] = in1[79] & in2[79];
    assign P[2] = in1[79] ^ in2[79];
    assign G[3] = in1[78] & in2[78];
    assign P[3] = in1[78] ^ in2[78];
    assign G[4] = in1[77] & in2[77];
    assign P[4] = in1[77] ^ in2[77];
    assign G[5] = in1[76] & in2[76];
    assign P[5] = in1[76] ^ in2[76];
    assign G[6] = in1[75] & in2[75];
    assign P[6] = in1[75] ^ in2[75];
    assign G[7] = in1[74] & in2[74];
    assign P[7] = in1[74] ^ in2[74];
    assign G[8] = in1[73] & in2[73];
    assign P[8] = in1[73] ^ in2[73];
    assign G[9] = in1[72] & in2[72];
    assign P[9] = in1[72] ^ in2[72];
    assign G[10] = in1[71] & in2[71];
    assign P[10] = in1[71] ^ in2[71];
    assign G[11] = in1[70] & in2[70];
    assign P[11] = in1[70] ^ in2[70];
    assign G[12] = in1[69] & in2[69];
    assign P[12] = in1[69] ^ in2[69];
    assign G[13] = in1[68] & in2[68];
    assign P[13] = in1[68] ^ in2[68];
    assign G[14] = in1[67] & in2[67];
    assign P[14] = in1[67] ^ in2[67];
    assign G[15] = in1[66] & in2[66];
    assign P[15] = in1[66] ^ in2[66];
    assign G[16] = in1[65] & in2[65];
    assign P[16] = in1[65] ^ in2[65];
    assign G[17] = in1[64] & in2[64];
    assign P[17] = in1[64] ^ in2[64];
    assign G[18] = in1[63] & in2[63];
    assign P[18] = in1[63] ^ in2[63];
    assign G[19] = in1[62] & in2[62];
    assign P[19] = in1[62] ^ in2[62];
    assign G[20] = in1[61] & in2[61];
    assign P[20] = in1[61] ^ in2[61];
    assign G[21] = in1[60] & in2[60];
    assign P[21] = in1[60] ^ in2[60];
    assign G[22] = in1[59] & in2[59];
    assign P[22] = in1[59] ^ in2[59];
    assign G[23] = in1[58] & in2[58];
    assign P[23] = in1[58] ^ in2[58];
    assign G[24] = in1[57] & in2[57];
    assign P[24] = in1[57] ^ in2[57];
    assign G[25] = in1[56] & in2[56];
    assign P[25] = in1[56] ^ in2[56];
    assign G[26] = in1[55] & in2[55];
    assign P[26] = in1[55] ^ in2[55];
    assign G[27] = in1[54] & in2[54];
    assign P[27] = in1[54] ^ in2[54];
    assign G[28] = in1[53] & in2[53];
    assign P[28] = in1[53] ^ in2[53];
    assign G[29] = in1[52] & in2[52];
    assign P[29] = in1[52] ^ in2[52];
    assign G[30] = in1[51] & in2[51];
    assign P[30] = in1[51] ^ in2[51];
    assign G[31] = in1[50] & in2[50];
    assign P[31] = in1[50] ^ in2[50];
    assign G[32] = in1[49] & in2[49];
    assign P[32] = in1[49] ^ in2[49];
    assign G[33] = in1[48] & in2[48];
    assign P[33] = in1[48] ^ in2[48];
    assign G[34] = in1[47] & in2[47];
    assign P[34] = in1[47] ^ in2[47];
    assign G[35] = in1[46] & in2[46];
    assign P[35] = in1[46] ^ in2[46];
    assign G[36] = in1[45] & in2[45];
    assign P[36] = in1[45] ^ in2[45];
    assign G[37] = in1[44] & in2[44];
    assign P[37] = in1[44] ^ in2[44];
    assign G[38] = in1[43] & in2[43];
    assign P[38] = in1[43] ^ in2[43];
    assign G[39] = in1[42] & in2[42];
    assign P[39] = in1[42] ^ in2[42];
    assign G[40] = in1[41] & in2[41];
    assign P[40] = in1[41] ^ in2[41];
    assign G[41] = in1[40] & in2[40];
    assign P[41] = in1[40] ^ in2[40];
    assign G[42] = in1[39] & in2[39];
    assign P[42] = in1[39] ^ in2[39];
    assign G[43] = in1[38] & in2[38];
    assign P[43] = in1[38] ^ in2[38];
    assign G[44] = in1[37] & in2[37];
    assign P[44] = in1[37] ^ in2[37];
    assign G[45] = in1[36] & in2[36];
    assign P[45] = in1[36] ^ in2[36];
    assign G[46] = in1[35] & in2[35];
    assign P[46] = in1[35] ^ in2[35];
    assign G[47] = in1[34] & in2[34];
    assign P[47] = in1[34] ^ in2[34];
    assign G[48] = in1[33] & in2[33];
    assign P[48] = in1[33] ^ in2[33];
    assign G[49] = in1[32] & in2[32];
    assign P[49] = in1[32] ^ in2[32];
    assign G[50] = in1[31] & in2[31];
    assign P[50] = in1[31] ^ in2[31];
    assign G[51] = in1[30] & in2[30];
    assign P[51] = in1[30] ^ in2[30];
    assign G[52] = in1[29] & in2[29];
    assign P[52] = in1[29] ^ in2[29];
    assign G[53] = in1[28] & in2[28];
    assign P[53] = in1[28] ^ in2[28];
    assign G[54] = in1[27] & in2[27];
    assign P[54] = in1[27] ^ in2[27];
    assign G[55] = in1[26] & in2[26];
    assign P[55] = in1[26] ^ in2[26];
    assign G[56] = in1[25] & in2[25];
    assign P[56] = in1[25] ^ in2[25];
    assign G[57] = in1[24] & in2[24];
    assign P[57] = in1[24] ^ in2[24];
    assign G[58] = in1[23] & in2[23];
    assign P[58] = in1[23] ^ in2[23];
    assign G[59] = in1[22] & in2[22];
    assign P[59] = in1[22] ^ in2[22];
    assign G[60] = in1[21] & in2[21];
    assign P[60] = in1[21] ^ in2[21];
    assign G[61] = in1[20] & in2[20];
    assign P[61] = in1[20] ^ in2[20];
    assign G[62] = in1[19] & in2[19];
    assign P[62] = in1[19] ^ in2[19];
    assign G[63] = in1[18] & in2[18];
    assign P[63] = in1[18] ^ in2[18];
    assign G[64] = in1[17] & in2[17];
    assign P[64] = in1[17] ^ in2[17];
    assign G[65] = in1[16] & in2[16];
    assign P[65] = in1[16] ^ in2[16];
    assign G[66] = in1[15] & in2[15];
    assign P[66] = in1[15] ^ in2[15];
    assign G[67] = in1[14] & in2[14];
    assign P[67] = in1[14] ^ in2[14];
    assign G[68] = in1[13] & in2[13];
    assign P[68] = in1[13] ^ in2[13];
    assign G[69] = in1[12] & in2[12];
    assign P[69] = in1[12] ^ in2[12];
    assign G[70] = in1[11] & in2[11];
    assign P[70] = in1[11] ^ in2[11];
    assign G[71] = in1[10] & in2[10];
    assign P[71] = in1[10] ^ in2[10];
    assign G[72] = in1[9] & in2[9];
    assign P[72] = in1[9] ^ in2[9];
    assign G[73] = in1[8] & in2[8];
    assign P[73] = in1[8] ^ in2[8];
    assign G[74] = in1[7] & in2[7];
    assign P[74] = in1[7] ^ in2[7];
    assign G[75] = in1[6] & in2[6];
    assign P[75] = in1[6] ^ in2[6];
    assign G[76] = in1[5] & in2[5];
    assign P[76] = in1[5] ^ in2[5];
    assign G[77] = in1[4] & in2[4];
    assign P[77] = in1[4] ^ in2[4];
    assign G[78] = in1[3] & in2[3];
    assign P[78] = in1[3] ^ in2[3];
    assign G[79] = in1[2] & in2[2];
    assign P[79] = in1[2] ^ in2[2];
    assign G[80] = in1[1] & in2[1];
    assign P[80] = in1[1] ^ in2[1];
    assign G[81] = in1[0] & in2[0];
    assign P[81] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign cout = G[81] | (P[81] & C[81]);
    assign sum = P ^ C;
endmodule

module CLA_81(output [80:0] sum, output cout, input [80:0] in1, input [80:0] in2);

    wire[80:0] G;
    wire[80:0] C;
    wire[80:0] P;

    assign G[0] = in1[80] & in2[80];
    assign P[0] = in1[80] ^ in2[80];
    assign G[1] = in1[79] & in2[79];
    assign P[1] = in1[79] ^ in2[79];
    assign G[2] = in1[78] & in2[78];
    assign P[2] = in1[78] ^ in2[78];
    assign G[3] = in1[77] & in2[77];
    assign P[3] = in1[77] ^ in2[77];
    assign G[4] = in1[76] & in2[76];
    assign P[4] = in1[76] ^ in2[76];
    assign G[5] = in1[75] & in2[75];
    assign P[5] = in1[75] ^ in2[75];
    assign G[6] = in1[74] & in2[74];
    assign P[6] = in1[74] ^ in2[74];
    assign G[7] = in1[73] & in2[73];
    assign P[7] = in1[73] ^ in2[73];
    assign G[8] = in1[72] & in2[72];
    assign P[8] = in1[72] ^ in2[72];
    assign G[9] = in1[71] & in2[71];
    assign P[9] = in1[71] ^ in2[71];
    assign G[10] = in1[70] & in2[70];
    assign P[10] = in1[70] ^ in2[70];
    assign G[11] = in1[69] & in2[69];
    assign P[11] = in1[69] ^ in2[69];
    assign G[12] = in1[68] & in2[68];
    assign P[12] = in1[68] ^ in2[68];
    assign G[13] = in1[67] & in2[67];
    assign P[13] = in1[67] ^ in2[67];
    assign G[14] = in1[66] & in2[66];
    assign P[14] = in1[66] ^ in2[66];
    assign G[15] = in1[65] & in2[65];
    assign P[15] = in1[65] ^ in2[65];
    assign G[16] = in1[64] & in2[64];
    assign P[16] = in1[64] ^ in2[64];
    assign G[17] = in1[63] & in2[63];
    assign P[17] = in1[63] ^ in2[63];
    assign G[18] = in1[62] & in2[62];
    assign P[18] = in1[62] ^ in2[62];
    assign G[19] = in1[61] & in2[61];
    assign P[19] = in1[61] ^ in2[61];
    assign G[20] = in1[60] & in2[60];
    assign P[20] = in1[60] ^ in2[60];
    assign G[21] = in1[59] & in2[59];
    assign P[21] = in1[59] ^ in2[59];
    assign G[22] = in1[58] & in2[58];
    assign P[22] = in1[58] ^ in2[58];
    assign G[23] = in1[57] & in2[57];
    assign P[23] = in1[57] ^ in2[57];
    assign G[24] = in1[56] & in2[56];
    assign P[24] = in1[56] ^ in2[56];
    assign G[25] = in1[55] & in2[55];
    assign P[25] = in1[55] ^ in2[55];
    assign G[26] = in1[54] & in2[54];
    assign P[26] = in1[54] ^ in2[54];
    assign G[27] = in1[53] & in2[53];
    assign P[27] = in1[53] ^ in2[53];
    assign G[28] = in1[52] & in2[52];
    assign P[28] = in1[52] ^ in2[52];
    assign G[29] = in1[51] & in2[51];
    assign P[29] = in1[51] ^ in2[51];
    assign G[30] = in1[50] & in2[50];
    assign P[30] = in1[50] ^ in2[50];
    assign G[31] = in1[49] & in2[49];
    assign P[31] = in1[49] ^ in2[49];
    assign G[32] = in1[48] & in2[48];
    assign P[32] = in1[48] ^ in2[48];
    assign G[33] = in1[47] & in2[47];
    assign P[33] = in1[47] ^ in2[47];
    assign G[34] = in1[46] & in2[46];
    assign P[34] = in1[46] ^ in2[46];
    assign G[35] = in1[45] & in2[45];
    assign P[35] = in1[45] ^ in2[45];
    assign G[36] = in1[44] & in2[44];
    assign P[36] = in1[44] ^ in2[44];
    assign G[37] = in1[43] & in2[43];
    assign P[37] = in1[43] ^ in2[43];
    assign G[38] = in1[42] & in2[42];
    assign P[38] = in1[42] ^ in2[42];
    assign G[39] = in1[41] & in2[41];
    assign P[39] = in1[41] ^ in2[41];
    assign G[40] = in1[40] & in2[40];
    assign P[40] = in1[40] ^ in2[40];
    assign G[41] = in1[39] & in2[39];
    assign P[41] = in1[39] ^ in2[39];
    assign G[42] = in1[38] & in2[38];
    assign P[42] = in1[38] ^ in2[38];
    assign G[43] = in1[37] & in2[37];
    assign P[43] = in1[37] ^ in2[37];
    assign G[44] = in1[36] & in2[36];
    assign P[44] = in1[36] ^ in2[36];
    assign G[45] = in1[35] & in2[35];
    assign P[45] = in1[35] ^ in2[35];
    assign G[46] = in1[34] & in2[34];
    assign P[46] = in1[34] ^ in2[34];
    assign G[47] = in1[33] & in2[33];
    assign P[47] = in1[33] ^ in2[33];
    assign G[48] = in1[32] & in2[32];
    assign P[48] = in1[32] ^ in2[32];
    assign G[49] = in1[31] & in2[31];
    assign P[49] = in1[31] ^ in2[31];
    assign G[50] = in1[30] & in2[30];
    assign P[50] = in1[30] ^ in2[30];
    assign G[51] = in1[29] & in2[29];
    assign P[51] = in1[29] ^ in2[29];
    assign G[52] = in1[28] & in2[28];
    assign P[52] = in1[28] ^ in2[28];
    assign G[53] = in1[27] & in2[27];
    assign P[53] = in1[27] ^ in2[27];
    assign G[54] = in1[26] & in2[26];
    assign P[54] = in1[26] ^ in2[26];
    assign G[55] = in1[25] & in2[25];
    assign P[55] = in1[25] ^ in2[25];
    assign G[56] = in1[24] & in2[24];
    assign P[56] = in1[24] ^ in2[24];
    assign G[57] = in1[23] & in2[23];
    assign P[57] = in1[23] ^ in2[23];
    assign G[58] = in1[22] & in2[22];
    assign P[58] = in1[22] ^ in2[22];
    assign G[59] = in1[21] & in2[21];
    assign P[59] = in1[21] ^ in2[21];
    assign G[60] = in1[20] & in2[20];
    assign P[60] = in1[20] ^ in2[20];
    assign G[61] = in1[19] & in2[19];
    assign P[61] = in1[19] ^ in2[19];
    assign G[62] = in1[18] & in2[18];
    assign P[62] = in1[18] ^ in2[18];
    assign G[63] = in1[17] & in2[17];
    assign P[63] = in1[17] ^ in2[17];
    assign G[64] = in1[16] & in2[16];
    assign P[64] = in1[16] ^ in2[16];
    assign G[65] = in1[15] & in2[15];
    assign P[65] = in1[15] ^ in2[15];
    assign G[66] = in1[14] & in2[14];
    assign P[66] = in1[14] ^ in2[14];
    assign G[67] = in1[13] & in2[13];
    assign P[67] = in1[13] ^ in2[13];
    assign G[68] = in1[12] & in2[12];
    assign P[68] = in1[12] ^ in2[12];
    assign G[69] = in1[11] & in2[11];
    assign P[69] = in1[11] ^ in2[11];
    assign G[70] = in1[10] & in2[10];
    assign P[70] = in1[10] ^ in2[10];
    assign G[71] = in1[9] & in2[9];
    assign P[71] = in1[9] ^ in2[9];
    assign G[72] = in1[8] & in2[8];
    assign P[72] = in1[8] ^ in2[8];
    assign G[73] = in1[7] & in2[7];
    assign P[73] = in1[7] ^ in2[7];
    assign G[74] = in1[6] & in2[6];
    assign P[74] = in1[6] ^ in2[6];
    assign G[75] = in1[5] & in2[5];
    assign P[75] = in1[5] ^ in2[5];
    assign G[76] = in1[4] & in2[4];
    assign P[76] = in1[4] ^ in2[4];
    assign G[77] = in1[3] & in2[3];
    assign P[77] = in1[3] ^ in2[3];
    assign G[78] = in1[2] & in2[2];
    assign P[78] = in1[2] ^ in2[2];
    assign G[79] = in1[1] & in2[1];
    assign P[79] = in1[1] ^ in2[1];
    assign G[80] = in1[0] & in2[0];
    assign P[80] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign cout = G[80] | (P[80] & C[80]);
    assign sum = P ^ C;
endmodule

module CLA_80(output [79:0] sum, output cout, input [79:0] in1, input [79:0] in2);

    wire[79:0] G;
    wire[79:0] C;
    wire[79:0] P;

    assign G[0] = in1[79] & in2[79];
    assign P[0] = in1[79] ^ in2[79];
    assign G[1] = in1[78] & in2[78];
    assign P[1] = in1[78] ^ in2[78];
    assign G[2] = in1[77] & in2[77];
    assign P[2] = in1[77] ^ in2[77];
    assign G[3] = in1[76] & in2[76];
    assign P[3] = in1[76] ^ in2[76];
    assign G[4] = in1[75] & in2[75];
    assign P[4] = in1[75] ^ in2[75];
    assign G[5] = in1[74] & in2[74];
    assign P[5] = in1[74] ^ in2[74];
    assign G[6] = in1[73] & in2[73];
    assign P[6] = in1[73] ^ in2[73];
    assign G[7] = in1[72] & in2[72];
    assign P[7] = in1[72] ^ in2[72];
    assign G[8] = in1[71] & in2[71];
    assign P[8] = in1[71] ^ in2[71];
    assign G[9] = in1[70] & in2[70];
    assign P[9] = in1[70] ^ in2[70];
    assign G[10] = in1[69] & in2[69];
    assign P[10] = in1[69] ^ in2[69];
    assign G[11] = in1[68] & in2[68];
    assign P[11] = in1[68] ^ in2[68];
    assign G[12] = in1[67] & in2[67];
    assign P[12] = in1[67] ^ in2[67];
    assign G[13] = in1[66] & in2[66];
    assign P[13] = in1[66] ^ in2[66];
    assign G[14] = in1[65] & in2[65];
    assign P[14] = in1[65] ^ in2[65];
    assign G[15] = in1[64] & in2[64];
    assign P[15] = in1[64] ^ in2[64];
    assign G[16] = in1[63] & in2[63];
    assign P[16] = in1[63] ^ in2[63];
    assign G[17] = in1[62] & in2[62];
    assign P[17] = in1[62] ^ in2[62];
    assign G[18] = in1[61] & in2[61];
    assign P[18] = in1[61] ^ in2[61];
    assign G[19] = in1[60] & in2[60];
    assign P[19] = in1[60] ^ in2[60];
    assign G[20] = in1[59] & in2[59];
    assign P[20] = in1[59] ^ in2[59];
    assign G[21] = in1[58] & in2[58];
    assign P[21] = in1[58] ^ in2[58];
    assign G[22] = in1[57] & in2[57];
    assign P[22] = in1[57] ^ in2[57];
    assign G[23] = in1[56] & in2[56];
    assign P[23] = in1[56] ^ in2[56];
    assign G[24] = in1[55] & in2[55];
    assign P[24] = in1[55] ^ in2[55];
    assign G[25] = in1[54] & in2[54];
    assign P[25] = in1[54] ^ in2[54];
    assign G[26] = in1[53] & in2[53];
    assign P[26] = in1[53] ^ in2[53];
    assign G[27] = in1[52] & in2[52];
    assign P[27] = in1[52] ^ in2[52];
    assign G[28] = in1[51] & in2[51];
    assign P[28] = in1[51] ^ in2[51];
    assign G[29] = in1[50] & in2[50];
    assign P[29] = in1[50] ^ in2[50];
    assign G[30] = in1[49] & in2[49];
    assign P[30] = in1[49] ^ in2[49];
    assign G[31] = in1[48] & in2[48];
    assign P[31] = in1[48] ^ in2[48];
    assign G[32] = in1[47] & in2[47];
    assign P[32] = in1[47] ^ in2[47];
    assign G[33] = in1[46] & in2[46];
    assign P[33] = in1[46] ^ in2[46];
    assign G[34] = in1[45] & in2[45];
    assign P[34] = in1[45] ^ in2[45];
    assign G[35] = in1[44] & in2[44];
    assign P[35] = in1[44] ^ in2[44];
    assign G[36] = in1[43] & in2[43];
    assign P[36] = in1[43] ^ in2[43];
    assign G[37] = in1[42] & in2[42];
    assign P[37] = in1[42] ^ in2[42];
    assign G[38] = in1[41] & in2[41];
    assign P[38] = in1[41] ^ in2[41];
    assign G[39] = in1[40] & in2[40];
    assign P[39] = in1[40] ^ in2[40];
    assign G[40] = in1[39] & in2[39];
    assign P[40] = in1[39] ^ in2[39];
    assign G[41] = in1[38] & in2[38];
    assign P[41] = in1[38] ^ in2[38];
    assign G[42] = in1[37] & in2[37];
    assign P[42] = in1[37] ^ in2[37];
    assign G[43] = in1[36] & in2[36];
    assign P[43] = in1[36] ^ in2[36];
    assign G[44] = in1[35] & in2[35];
    assign P[44] = in1[35] ^ in2[35];
    assign G[45] = in1[34] & in2[34];
    assign P[45] = in1[34] ^ in2[34];
    assign G[46] = in1[33] & in2[33];
    assign P[46] = in1[33] ^ in2[33];
    assign G[47] = in1[32] & in2[32];
    assign P[47] = in1[32] ^ in2[32];
    assign G[48] = in1[31] & in2[31];
    assign P[48] = in1[31] ^ in2[31];
    assign G[49] = in1[30] & in2[30];
    assign P[49] = in1[30] ^ in2[30];
    assign G[50] = in1[29] & in2[29];
    assign P[50] = in1[29] ^ in2[29];
    assign G[51] = in1[28] & in2[28];
    assign P[51] = in1[28] ^ in2[28];
    assign G[52] = in1[27] & in2[27];
    assign P[52] = in1[27] ^ in2[27];
    assign G[53] = in1[26] & in2[26];
    assign P[53] = in1[26] ^ in2[26];
    assign G[54] = in1[25] & in2[25];
    assign P[54] = in1[25] ^ in2[25];
    assign G[55] = in1[24] & in2[24];
    assign P[55] = in1[24] ^ in2[24];
    assign G[56] = in1[23] & in2[23];
    assign P[56] = in1[23] ^ in2[23];
    assign G[57] = in1[22] & in2[22];
    assign P[57] = in1[22] ^ in2[22];
    assign G[58] = in1[21] & in2[21];
    assign P[58] = in1[21] ^ in2[21];
    assign G[59] = in1[20] & in2[20];
    assign P[59] = in1[20] ^ in2[20];
    assign G[60] = in1[19] & in2[19];
    assign P[60] = in1[19] ^ in2[19];
    assign G[61] = in1[18] & in2[18];
    assign P[61] = in1[18] ^ in2[18];
    assign G[62] = in1[17] & in2[17];
    assign P[62] = in1[17] ^ in2[17];
    assign G[63] = in1[16] & in2[16];
    assign P[63] = in1[16] ^ in2[16];
    assign G[64] = in1[15] & in2[15];
    assign P[64] = in1[15] ^ in2[15];
    assign G[65] = in1[14] & in2[14];
    assign P[65] = in1[14] ^ in2[14];
    assign G[66] = in1[13] & in2[13];
    assign P[66] = in1[13] ^ in2[13];
    assign G[67] = in1[12] & in2[12];
    assign P[67] = in1[12] ^ in2[12];
    assign G[68] = in1[11] & in2[11];
    assign P[68] = in1[11] ^ in2[11];
    assign G[69] = in1[10] & in2[10];
    assign P[69] = in1[10] ^ in2[10];
    assign G[70] = in1[9] & in2[9];
    assign P[70] = in1[9] ^ in2[9];
    assign G[71] = in1[8] & in2[8];
    assign P[71] = in1[8] ^ in2[8];
    assign G[72] = in1[7] & in2[7];
    assign P[72] = in1[7] ^ in2[7];
    assign G[73] = in1[6] & in2[6];
    assign P[73] = in1[6] ^ in2[6];
    assign G[74] = in1[5] & in2[5];
    assign P[74] = in1[5] ^ in2[5];
    assign G[75] = in1[4] & in2[4];
    assign P[75] = in1[4] ^ in2[4];
    assign G[76] = in1[3] & in2[3];
    assign P[76] = in1[3] ^ in2[3];
    assign G[77] = in1[2] & in2[2];
    assign P[77] = in1[2] ^ in2[2];
    assign G[78] = in1[1] & in2[1];
    assign P[78] = in1[1] ^ in2[1];
    assign G[79] = in1[0] & in2[0];
    assign P[79] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign cout = G[79] | (P[79] & C[79]);
    assign sum = P ^ C;
endmodule

module CLA_79(output [78:0] sum, output cout, input [78:0] in1, input [78:0] in2);

    wire[78:0] G;
    wire[78:0] C;
    wire[78:0] P;

    assign G[0] = in1[78] & in2[78];
    assign P[0] = in1[78] ^ in2[78];
    assign G[1] = in1[77] & in2[77];
    assign P[1] = in1[77] ^ in2[77];
    assign G[2] = in1[76] & in2[76];
    assign P[2] = in1[76] ^ in2[76];
    assign G[3] = in1[75] & in2[75];
    assign P[3] = in1[75] ^ in2[75];
    assign G[4] = in1[74] & in2[74];
    assign P[4] = in1[74] ^ in2[74];
    assign G[5] = in1[73] & in2[73];
    assign P[5] = in1[73] ^ in2[73];
    assign G[6] = in1[72] & in2[72];
    assign P[6] = in1[72] ^ in2[72];
    assign G[7] = in1[71] & in2[71];
    assign P[7] = in1[71] ^ in2[71];
    assign G[8] = in1[70] & in2[70];
    assign P[8] = in1[70] ^ in2[70];
    assign G[9] = in1[69] & in2[69];
    assign P[9] = in1[69] ^ in2[69];
    assign G[10] = in1[68] & in2[68];
    assign P[10] = in1[68] ^ in2[68];
    assign G[11] = in1[67] & in2[67];
    assign P[11] = in1[67] ^ in2[67];
    assign G[12] = in1[66] & in2[66];
    assign P[12] = in1[66] ^ in2[66];
    assign G[13] = in1[65] & in2[65];
    assign P[13] = in1[65] ^ in2[65];
    assign G[14] = in1[64] & in2[64];
    assign P[14] = in1[64] ^ in2[64];
    assign G[15] = in1[63] & in2[63];
    assign P[15] = in1[63] ^ in2[63];
    assign G[16] = in1[62] & in2[62];
    assign P[16] = in1[62] ^ in2[62];
    assign G[17] = in1[61] & in2[61];
    assign P[17] = in1[61] ^ in2[61];
    assign G[18] = in1[60] & in2[60];
    assign P[18] = in1[60] ^ in2[60];
    assign G[19] = in1[59] & in2[59];
    assign P[19] = in1[59] ^ in2[59];
    assign G[20] = in1[58] & in2[58];
    assign P[20] = in1[58] ^ in2[58];
    assign G[21] = in1[57] & in2[57];
    assign P[21] = in1[57] ^ in2[57];
    assign G[22] = in1[56] & in2[56];
    assign P[22] = in1[56] ^ in2[56];
    assign G[23] = in1[55] & in2[55];
    assign P[23] = in1[55] ^ in2[55];
    assign G[24] = in1[54] & in2[54];
    assign P[24] = in1[54] ^ in2[54];
    assign G[25] = in1[53] & in2[53];
    assign P[25] = in1[53] ^ in2[53];
    assign G[26] = in1[52] & in2[52];
    assign P[26] = in1[52] ^ in2[52];
    assign G[27] = in1[51] & in2[51];
    assign P[27] = in1[51] ^ in2[51];
    assign G[28] = in1[50] & in2[50];
    assign P[28] = in1[50] ^ in2[50];
    assign G[29] = in1[49] & in2[49];
    assign P[29] = in1[49] ^ in2[49];
    assign G[30] = in1[48] & in2[48];
    assign P[30] = in1[48] ^ in2[48];
    assign G[31] = in1[47] & in2[47];
    assign P[31] = in1[47] ^ in2[47];
    assign G[32] = in1[46] & in2[46];
    assign P[32] = in1[46] ^ in2[46];
    assign G[33] = in1[45] & in2[45];
    assign P[33] = in1[45] ^ in2[45];
    assign G[34] = in1[44] & in2[44];
    assign P[34] = in1[44] ^ in2[44];
    assign G[35] = in1[43] & in2[43];
    assign P[35] = in1[43] ^ in2[43];
    assign G[36] = in1[42] & in2[42];
    assign P[36] = in1[42] ^ in2[42];
    assign G[37] = in1[41] & in2[41];
    assign P[37] = in1[41] ^ in2[41];
    assign G[38] = in1[40] & in2[40];
    assign P[38] = in1[40] ^ in2[40];
    assign G[39] = in1[39] & in2[39];
    assign P[39] = in1[39] ^ in2[39];
    assign G[40] = in1[38] & in2[38];
    assign P[40] = in1[38] ^ in2[38];
    assign G[41] = in1[37] & in2[37];
    assign P[41] = in1[37] ^ in2[37];
    assign G[42] = in1[36] & in2[36];
    assign P[42] = in1[36] ^ in2[36];
    assign G[43] = in1[35] & in2[35];
    assign P[43] = in1[35] ^ in2[35];
    assign G[44] = in1[34] & in2[34];
    assign P[44] = in1[34] ^ in2[34];
    assign G[45] = in1[33] & in2[33];
    assign P[45] = in1[33] ^ in2[33];
    assign G[46] = in1[32] & in2[32];
    assign P[46] = in1[32] ^ in2[32];
    assign G[47] = in1[31] & in2[31];
    assign P[47] = in1[31] ^ in2[31];
    assign G[48] = in1[30] & in2[30];
    assign P[48] = in1[30] ^ in2[30];
    assign G[49] = in1[29] & in2[29];
    assign P[49] = in1[29] ^ in2[29];
    assign G[50] = in1[28] & in2[28];
    assign P[50] = in1[28] ^ in2[28];
    assign G[51] = in1[27] & in2[27];
    assign P[51] = in1[27] ^ in2[27];
    assign G[52] = in1[26] & in2[26];
    assign P[52] = in1[26] ^ in2[26];
    assign G[53] = in1[25] & in2[25];
    assign P[53] = in1[25] ^ in2[25];
    assign G[54] = in1[24] & in2[24];
    assign P[54] = in1[24] ^ in2[24];
    assign G[55] = in1[23] & in2[23];
    assign P[55] = in1[23] ^ in2[23];
    assign G[56] = in1[22] & in2[22];
    assign P[56] = in1[22] ^ in2[22];
    assign G[57] = in1[21] & in2[21];
    assign P[57] = in1[21] ^ in2[21];
    assign G[58] = in1[20] & in2[20];
    assign P[58] = in1[20] ^ in2[20];
    assign G[59] = in1[19] & in2[19];
    assign P[59] = in1[19] ^ in2[19];
    assign G[60] = in1[18] & in2[18];
    assign P[60] = in1[18] ^ in2[18];
    assign G[61] = in1[17] & in2[17];
    assign P[61] = in1[17] ^ in2[17];
    assign G[62] = in1[16] & in2[16];
    assign P[62] = in1[16] ^ in2[16];
    assign G[63] = in1[15] & in2[15];
    assign P[63] = in1[15] ^ in2[15];
    assign G[64] = in1[14] & in2[14];
    assign P[64] = in1[14] ^ in2[14];
    assign G[65] = in1[13] & in2[13];
    assign P[65] = in1[13] ^ in2[13];
    assign G[66] = in1[12] & in2[12];
    assign P[66] = in1[12] ^ in2[12];
    assign G[67] = in1[11] & in2[11];
    assign P[67] = in1[11] ^ in2[11];
    assign G[68] = in1[10] & in2[10];
    assign P[68] = in1[10] ^ in2[10];
    assign G[69] = in1[9] & in2[9];
    assign P[69] = in1[9] ^ in2[9];
    assign G[70] = in1[8] & in2[8];
    assign P[70] = in1[8] ^ in2[8];
    assign G[71] = in1[7] & in2[7];
    assign P[71] = in1[7] ^ in2[7];
    assign G[72] = in1[6] & in2[6];
    assign P[72] = in1[6] ^ in2[6];
    assign G[73] = in1[5] & in2[5];
    assign P[73] = in1[5] ^ in2[5];
    assign G[74] = in1[4] & in2[4];
    assign P[74] = in1[4] ^ in2[4];
    assign G[75] = in1[3] & in2[3];
    assign P[75] = in1[3] ^ in2[3];
    assign G[76] = in1[2] & in2[2];
    assign P[76] = in1[2] ^ in2[2];
    assign G[77] = in1[1] & in2[1];
    assign P[77] = in1[1] ^ in2[1];
    assign G[78] = in1[0] & in2[0];
    assign P[78] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign cout = G[78] | (P[78] & C[78]);
    assign sum = P ^ C;
endmodule

module CLA_78(output [77:0] sum, output cout, input [77:0] in1, input [77:0] in2);

    wire[77:0] G;
    wire[77:0] C;
    wire[77:0] P;

    assign G[0] = in1[77] & in2[77];
    assign P[0] = in1[77] ^ in2[77];
    assign G[1] = in1[76] & in2[76];
    assign P[1] = in1[76] ^ in2[76];
    assign G[2] = in1[75] & in2[75];
    assign P[2] = in1[75] ^ in2[75];
    assign G[3] = in1[74] & in2[74];
    assign P[3] = in1[74] ^ in2[74];
    assign G[4] = in1[73] & in2[73];
    assign P[4] = in1[73] ^ in2[73];
    assign G[5] = in1[72] & in2[72];
    assign P[5] = in1[72] ^ in2[72];
    assign G[6] = in1[71] & in2[71];
    assign P[6] = in1[71] ^ in2[71];
    assign G[7] = in1[70] & in2[70];
    assign P[7] = in1[70] ^ in2[70];
    assign G[8] = in1[69] & in2[69];
    assign P[8] = in1[69] ^ in2[69];
    assign G[9] = in1[68] & in2[68];
    assign P[9] = in1[68] ^ in2[68];
    assign G[10] = in1[67] & in2[67];
    assign P[10] = in1[67] ^ in2[67];
    assign G[11] = in1[66] & in2[66];
    assign P[11] = in1[66] ^ in2[66];
    assign G[12] = in1[65] & in2[65];
    assign P[12] = in1[65] ^ in2[65];
    assign G[13] = in1[64] & in2[64];
    assign P[13] = in1[64] ^ in2[64];
    assign G[14] = in1[63] & in2[63];
    assign P[14] = in1[63] ^ in2[63];
    assign G[15] = in1[62] & in2[62];
    assign P[15] = in1[62] ^ in2[62];
    assign G[16] = in1[61] & in2[61];
    assign P[16] = in1[61] ^ in2[61];
    assign G[17] = in1[60] & in2[60];
    assign P[17] = in1[60] ^ in2[60];
    assign G[18] = in1[59] & in2[59];
    assign P[18] = in1[59] ^ in2[59];
    assign G[19] = in1[58] & in2[58];
    assign P[19] = in1[58] ^ in2[58];
    assign G[20] = in1[57] & in2[57];
    assign P[20] = in1[57] ^ in2[57];
    assign G[21] = in1[56] & in2[56];
    assign P[21] = in1[56] ^ in2[56];
    assign G[22] = in1[55] & in2[55];
    assign P[22] = in1[55] ^ in2[55];
    assign G[23] = in1[54] & in2[54];
    assign P[23] = in1[54] ^ in2[54];
    assign G[24] = in1[53] & in2[53];
    assign P[24] = in1[53] ^ in2[53];
    assign G[25] = in1[52] & in2[52];
    assign P[25] = in1[52] ^ in2[52];
    assign G[26] = in1[51] & in2[51];
    assign P[26] = in1[51] ^ in2[51];
    assign G[27] = in1[50] & in2[50];
    assign P[27] = in1[50] ^ in2[50];
    assign G[28] = in1[49] & in2[49];
    assign P[28] = in1[49] ^ in2[49];
    assign G[29] = in1[48] & in2[48];
    assign P[29] = in1[48] ^ in2[48];
    assign G[30] = in1[47] & in2[47];
    assign P[30] = in1[47] ^ in2[47];
    assign G[31] = in1[46] & in2[46];
    assign P[31] = in1[46] ^ in2[46];
    assign G[32] = in1[45] & in2[45];
    assign P[32] = in1[45] ^ in2[45];
    assign G[33] = in1[44] & in2[44];
    assign P[33] = in1[44] ^ in2[44];
    assign G[34] = in1[43] & in2[43];
    assign P[34] = in1[43] ^ in2[43];
    assign G[35] = in1[42] & in2[42];
    assign P[35] = in1[42] ^ in2[42];
    assign G[36] = in1[41] & in2[41];
    assign P[36] = in1[41] ^ in2[41];
    assign G[37] = in1[40] & in2[40];
    assign P[37] = in1[40] ^ in2[40];
    assign G[38] = in1[39] & in2[39];
    assign P[38] = in1[39] ^ in2[39];
    assign G[39] = in1[38] & in2[38];
    assign P[39] = in1[38] ^ in2[38];
    assign G[40] = in1[37] & in2[37];
    assign P[40] = in1[37] ^ in2[37];
    assign G[41] = in1[36] & in2[36];
    assign P[41] = in1[36] ^ in2[36];
    assign G[42] = in1[35] & in2[35];
    assign P[42] = in1[35] ^ in2[35];
    assign G[43] = in1[34] & in2[34];
    assign P[43] = in1[34] ^ in2[34];
    assign G[44] = in1[33] & in2[33];
    assign P[44] = in1[33] ^ in2[33];
    assign G[45] = in1[32] & in2[32];
    assign P[45] = in1[32] ^ in2[32];
    assign G[46] = in1[31] & in2[31];
    assign P[46] = in1[31] ^ in2[31];
    assign G[47] = in1[30] & in2[30];
    assign P[47] = in1[30] ^ in2[30];
    assign G[48] = in1[29] & in2[29];
    assign P[48] = in1[29] ^ in2[29];
    assign G[49] = in1[28] & in2[28];
    assign P[49] = in1[28] ^ in2[28];
    assign G[50] = in1[27] & in2[27];
    assign P[50] = in1[27] ^ in2[27];
    assign G[51] = in1[26] & in2[26];
    assign P[51] = in1[26] ^ in2[26];
    assign G[52] = in1[25] & in2[25];
    assign P[52] = in1[25] ^ in2[25];
    assign G[53] = in1[24] & in2[24];
    assign P[53] = in1[24] ^ in2[24];
    assign G[54] = in1[23] & in2[23];
    assign P[54] = in1[23] ^ in2[23];
    assign G[55] = in1[22] & in2[22];
    assign P[55] = in1[22] ^ in2[22];
    assign G[56] = in1[21] & in2[21];
    assign P[56] = in1[21] ^ in2[21];
    assign G[57] = in1[20] & in2[20];
    assign P[57] = in1[20] ^ in2[20];
    assign G[58] = in1[19] & in2[19];
    assign P[58] = in1[19] ^ in2[19];
    assign G[59] = in1[18] & in2[18];
    assign P[59] = in1[18] ^ in2[18];
    assign G[60] = in1[17] & in2[17];
    assign P[60] = in1[17] ^ in2[17];
    assign G[61] = in1[16] & in2[16];
    assign P[61] = in1[16] ^ in2[16];
    assign G[62] = in1[15] & in2[15];
    assign P[62] = in1[15] ^ in2[15];
    assign G[63] = in1[14] & in2[14];
    assign P[63] = in1[14] ^ in2[14];
    assign G[64] = in1[13] & in2[13];
    assign P[64] = in1[13] ^ in2[13];
    assign G[65] = in1[12] & in2[12];
    assign P[65] = in1[12] ^ in2[12];
    assign G[66] = in1[11] & in2[11];
    assign P[66] = in1[11] ^ in2[11];
    assign G[67] = in1[10] & in2[10];
    assign P[67] = in1[10] ^ in2[10];
    assign G[68] = in1[9] & in2[9];
    assign P[68] = in1[9] ^ in2[9];
    assign G[69] = in1[8] & in2[8];
    assign P[69] = in1[8] ^ in2[8];
    assign G[70] = in1[7] & in2[7];
    assign P[70] = in1[7] ^ in2[7];
    assign G[71] = in1[6] & in2[6];
    assign P[71] = in1[6] ^ in2[6];
    assign G[72] = in1[5] & in2[5];
    assign P[72] = in1[5] ^ in2[5];
    assign G[73] = in1[4] & in2[4];
    assign P[73] = in1[4] ^ in2[4];
    assign G[74] = in1[3] & in2[3];
    assign P[74] = in1[3] ^ in2[3];
    assign G[75] = in1[2] & in2[2];
    assign P[75] = in1[2] ^ in2[2];
    assign G[76] = in1[1] & in2[1];
    assign P[76] = in1[1] ^ in2[1];
    assign G[77] = in1[0] & in2[0];
    assign P[77] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign cout = G[77] | (P[77] & C[77]);
    assign sum = P ^ C;
endmodule

module CLA_77(output [76:0] sum, output cout, input [76:0] in1, input [76:0] in2);

    wire[76:0] G;
    wire[76:0] C;
    wire[76:0] P;

    assign G[0] = in1[76] & in2[76];
    assign P[0] = in1[76] ^ in2[76];
    assign G[1] = in1[75] & in2[75];
    assign P[1] = in1[75] ^ in2[75];
    assign G[2] = in1[74] & in2[74];
    assign P[2] = in1[74] ^ in2[74];
    assign G[3] = in1[73] & in2[73];
    assign P[3] = in1[73] ^ in2[73];
    assign G[4] = in1[72] & in2[72];
    assign P[4] = in1[72] ^ in2[72];
    assign G[5] = in1[71] & in2[71];
    assign P[5] = in1[71] ^ in2[71];
    assign G[6] = in1[70] & in2[70];
    assign P[6] = in1[70] ^ in2[70];
    assign G[7] = in1[69] & in2[69];
    assign P[7] = in1[69] ^ in2[69];
    assign G[8] = in1[68] & in2[68];
    assign P[8] = in1[68] ^ in2[68];
    assign G[9] = in1[67] & in2[67];
    assign P[9] = in1[67] ^ in2[67];
    assign G[10] = in1[66] & in2[66];
    assign P[10] = in1[66] ^ in2[66];
    assign G[11] = in1[65] & in2[65];
    assign P[11] = in1[65] ^ in2[65];
    assign G[12] = in1[64] & in2[64];
    assign P[12] = in1[64] ^ in2[64];
    assign G[13] = in1[63] & in2[63];
    assign P[13] = in1[63] ^ in2[63];
    assign G[14] = in1[62] & in2[62];
    assign P[14] = in1[62] ^ in2[62];
    assign G[15] = in1[61] & in2[61];
    assign P[15] = in1[61] ^ in2[61];
    assign G[16] = in1[60] & in2[60];
    assign P[16] = in1[60] ^ in2[60];
    assign G[17] = in1[59] & in2[59];
    assign P[17] = in1[59] ^ in2[59];
    assign G[18] = in1[58] & in2[58];
    assign P[18] = in1[58] ^ in2[58];
    assign G[19] = in1[57] & in2[57];
    assign P[19] = in1[57] ^ in2[57];
    assign G[20] = in1[56] & in2[56];
    assign P[20] = in1[56] ^ in2[56];
    assign G[21] = in1[55] & in2[55];
    assign P[21] = in1[55] ^ in2[55];
    assign G[22] = in1[54] & in2[54];
    assign P[22] = in1[54] ^ in2[54];
    assign G[23] = in1[53] & in2[53];
    assign P[23] = in1[53] ^ in2[53];
    assign G[24] = in1[52] & in2[52];
    assign P[24] = in1[52] ^ in2[52];
    assign G[25] = in1[51] & in2[51];
    assign P[25] = in1[51] ^ in2[51];
    assign G[26] = in1[50] & in2[50];
    assign P[26] = in1[50] ^ in2[50];
    assign G[27] = in1[49] & in2[49];
    assign P[27] = in1[49] ^ in2[49];
    assign G[28] = in1[48] & in2[48];
    assign P[28] = in1[48] ^ in2[48];
    assign G[29] = in1[47] & in2[47];
    assign P[29] = in1[47] ^ in2[47];
    assign G[30] = in1[46] & in2[46];
    assign P[30] = in1[46] ^ in2[46];
    assign G[31] = in1[45] & in2[45];
    assign P[31] = in1[45] ^ in2[45];
    assign G[32] = in1[44] & in2[44];
    assign P[32] = in1[44] ^ in2[44];
    assign G[33] = in1[43] & in2[43];
    assign P[33] = in1[43] ^ in2[43];
    assign G[34] = in1[42] & in2[42];
    assign P[34] = in1[42] ^ in2[42];
    assign G[35] = in1[41] & in2[41];
    assign P[35] = in1[41] ^ in2[41];
    assign G[36] = in1[40] & in2[40];
    assign P[36] = in1[40] ^ in2[40];
    assign G[37] = in1[39] & in2[39];
    assign P[37] = in1[39] ^ in2[39];
    assign G[38] = in1[38] & in2[38];
    assign P[38] = in1[38] ^ in2[38];
    assign G[39] = in1[37] & in2[37];
    assign P[39] = in1[37] ^ in2[37];
    assign G[40] = in1[36] & in2[36];
    assign P[40] = in1[36] ^ in2[36];
    assign G[41] = in1[35] & in2[35];
    assign P[41] = in1[35] ^ in2[35];
    assign G[42] = in1[34] & in2[34];
    assign P[42] = in1[34] ^ in2[34];
    assign G[43] = in1[33] & in2[33];
    assign P[43] = in1[33] ^ in2[33];
    assign G[44] = in1[32] & in2[32];
    assign P[44] = in1[32] ^ in2[32];
    assign G[45] = in1[31] & in2[31];
    assign P[45] = in1[31] ^ in2[31];
    assign G[46] = in1[30] & in2[30];
    assign P[46] = in1[30] ^ in2[30];
    assign G[47] = in1[29] & in2[29];
    assign P[47] = in1[29] ^ in2[29];
    assign G[48] = in1[28] & in2[28];
    assign P[48] = in1[28] ^ in2[28];
    assign G[49] = in1[27] & in2[27];
    assign P[49] = in1[27] ^ in2[27];
    assign G[50] = in1[26] & in2[26];
    assign P[50] = in1[26] ^ in2[26];
    assign G[51] = in1[25] & in2[25];
    assign P[51] = in1[25] ^ in2[25];
    assign G[52] = in1[24] & in2[24];
    assign P[52] = in1[24] ^ in2[24];
    assign G[53] = in1[23] & in2[23];
    assign P[53] = in1[23] ^ in2[23];
    assign G[54] = in1[22] & in2[22];
    assign P[54] = in1[22] ^ in2[22];
    assign G[55] = in1[21] & in2[21];
    assign P[55] = in1[21] ^ in2[21];
    assign G[56] = in1[20] & in2[20];
    assign P[56] = in1[20] ^ in2[20];
    assign G[57] = in1[19] & in2[19];
    assign P[57] = in1[19] ^ in2[19];
    assign G[58] = in1[18] & in2[18];
    assign P[58] = in1[18] ^ in2[18];
    assign G[59] = in1[17] & in2[17];
    assign P[59] = in1[17] ^ in2[17];
    assign G[60] = in1[16] & in2[16];
    assign P[60] = in1[16] ^ in2[16];
    assign G[61] = in1[15] & in2[15];
    assign P[61] = in1[15] ^ in2[15];
    assign G[62] = in1[14] & in2[14];
    assign P[62] = in1[14] ^ in2[14];
    assign G[63] = in1[13] & in2[13];
    assign P[63] = in1[13] ^ in2[13];
    assign G[64] = in1[12] & in2[12];
    assign P[64] = in1[12] ^ in2[12];
    assign G[65] = in1[11] & in2[11];
    assign P[65] = in1[11] ^ in2[11];
    assign G[66] = in1[10] & in2[10];
    assign P[66] = in1[10] ^ in2[10];
    assign G[67] = in1[9] & in2[9];
    assign P[67] = in1[9] ^ in2[9];
    assign G[68] = in1[8] & in2[8];
    assign P[68] = in1[8] ^ in2[8];
    assign G[69] = in1[7] & in2[7];
    assign P[69] = in1[7] ^ in2[7];
    assign G[70] = in1[6] & in2[6];
    assign P[70] = in1[6] ^ in2[6];
    assign G[71] = in1[5] & in2[5];
    assign P[71] = in1[5] ^ in2[5];
    assign G[72] = in1[4] & in2[4];
    assign P[72] = in1[4] ^ in2[4];
    assign G[73] = in1[3] & in2[3];
    assign P[73] = in1[3] ^ in2[3];
    assign G[74] = in1[2] & in2[2];
    assign P[74] = in1[2] ^ in2[2];
    assign G[75] = in1[1] & in2[1];
    assign P[75] = in1[1] ^ in2[1];
    assign G[76] = in1[0] & in2[0];
    assign P[76] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign cout = G[76] | (P[76] & C[76]);
    assign sum = P ^ C;
endmodule

module CLA_76(output [75:0] sum, output cout, input [75:0] in1, input [75:0] in2);

    wire[75:0] G;
    wire[75:0] C;
    wire[75:0] P;

    assign G[0] = in1[75] & in2[75];
    assign P[0] = in1[75] ^ in2[75];
    assign G[1] = in1[74] & in2[74];
    assign P[1] = in1[74] ^ in2[74];
    assign G[2] = in1[73] & in2[73];
    assign P[2] = in1[73] ^ in2[73];
    assign G[3] = in1[72] & in2[72];
    assign P[3] = in1[72] ^ in2[72];
    assign G[4] = in1[71] & in2[71];
    assign P[4] = in1[71] ^ in2[71];
    assign G[5] = in1[70] & in2[70];
    assign P[5] = in1[70] ^ in2[70];
    assign G[6] = in1[69] & in2[69];
    assign P[6] = in1[69] ^ in2[69];
    assign G[7] = in1[68] & in2[68];
    assign P[7] = in1[68] ^ in2[68];
    assign G[8] = in1[67] & in2[67];
    assign P[8] = in1[67] ^ in2[67];
    assign G[9] = in1[66] & in2[66];
    assign P[9] = in1[66] ^ in2[66];
    assign G[10] = in1[65] & in2[65];
    assign P[10] = in1[65] ^ in2[65];
    assign G[11] = in1[64] & in2[64];
    assign P[11] = in1[64] ^ in2[64];
    assign G[12] = in1[63] & in2[63];
    assign P[12] = in1[63] ^ in2[63];
    assign G[13] = in1[62] & in2[62];
    assign P[13] = in1[62] ^ in2[62];
    assign G[14] = in1[61] & in2[61];
    assign P[14] = in1[61] ^ in2[61];
    assign G[15] = in1[60] & in2[60];
    assign P[15] = in1[60] ^ in2[60];
    assign G[16] = in1[59] & in2[59];
    assign P[16] = in1[59] ^ in2[59];
    assign G[17] = in1[58] & in2[58];
    assign P[17] = in1[58] ^ in2[58];
    assign G[18] = in1[57] & in2[57];
    assign P[18] = in1[57] ^ in2[57];
    assign G[19] = in1[56] & in2[56];
    assign P[19] = in1[56] ^ in2[56];
    assign G[20] = in1[55] & in2[55];
    assign P[20] = in1[55] ^ in2[55];
    assign G[21] = in1[54] & in2[54];
    assign P[21] = in1[54] ^ in2[54];
    assign G[22] = in1[53] & in2[53];
    assign P[22] = in1[53] ^ in2[53];
    assign G[23] = in1[52] & in2[52];
    assign P[23] = in1[52] ^ in2[52];
    assign G[24] = in1[51] & in2[51];
    assign P[24] = in1[51] ^ in2[51];
    assign G[25] = in1[50] & in2[50];
    assign P[25] = in1[50] ^ in2[50];
    assign G[26] = in1[49] & in2[49];
    assign P[26] = in1[49] ^ in2[49];
    assign G[27] = in1[48] & in2[48];
    assign P[27] = in1[48] ^ in2[48];
    assign G[28] = in1[47] & in2[47];
    assign P[28] = in1[47] ^ in2[47];
    assign G[29] = in1[46] & in2[46];
    assign P[29] = in1[46] ^ in2[46];
    assign G[30] = in1[45] & in2[45];
    assign P[30] = in1[45] ^ in2[45];
    assign G[31] = in1[44] & in2[44];
    assign P[31] = in1[44] ^ in2[44];
    assign G[32] = in1[43] & in2[43];
    assign P[32] = in1[43] ^ in2[43];
    assign G[33] = in1[42] & in2[42];
    assign P[33] = in1[42] ^ in2[42];
    assign G[34] = in1[41] & in2[41];
    assign P[34] = in1[41] ^ in2[41];
    assign G[35] = in1[40] & in2[40];
    assign P[35] = in1[40] ^ in2[40];
    assign G[36] = in1[39] & in2[39];
    assign P[36] = in1[39] ^ in2[39];
    assign G[37] = in1[38] & in2[38];
    assign P[37] = in1[38] ^ in2[38];
    assign G[38] = in1[37] & in2[37];
    assign P[38] = in1[37] ^ in2[37];
    assign G[39] = in1[36] & in2[36];
    assign P[39] = in1[36] ^ in2[36];
    assign G[40] = in1[35] & in2[35];
    assign P[40] = in1[35] ^ in2[35];
    assign G[41] = in1[34] & in2[34];
    assign P[41] = in1[34] ^ in2[34];
    assign G[42] = in1[33] & in2[33];
    assign P[42] = in1[33] ^ in2[33];
    assign G[43] = in1[32] & in2[32];
    assign P[43] = in1[32] ^ in2[32];
    assign G[44] = in1[31] & in2[31];
    assign P[44] = in1[31] ^ in2[31];
    assign G[45] = in1[30] & in2[30];
    assign P[45] = in1[30] ^ in2[30];
    assign G[46] = in1[29] & in2[29];
    assign P[46] = in1[29] ^ in2[29];
    assign G[47] = in1[28] & in2[28];
    assign P[47] = in1[28] ^ in2[28];
    assign G[48] = in1[27] & in2[27];
    assign P[48] = in1[27] ^ in2[27];
    assign G[49] = in1[26] & in2[26];
    assign P[49] = in1[26] ^ in2[26];
    assign G[50] = in1[25] & in2[25];
    assign P[50] = in1[25] ^ in2[25];
    assign G[51] = in1[24] & in2[24];
    assign P[51] = in1[24] ^ in2[24];
    assign G[52] = in1[23] & in2[23];
    assign P[52] = in1[23] ^ in2[23];
    assign G[53] = in1[22] & in2[22];
    assign P[53] = in1[22] ^ in2[22];
    assign G[54] = in1[21] & in2[21];
    assign P[54] = in1[21] ^ in2[21];
    assign G[55] = in1[20] & in2[20];
    assign P[55] = in1[20] ^ in2[20];
    assign G[56] = in1[19] & in2[19];
    assign P[56] = in1[19] ^ in2[19];
    assign G[57] = in1[18] & in2[18];
    assign P[57] = in1[18] ^ in2[18];
    assign G[58] = in1[17] & in2[17];
    assign P[58] = in1[17] ^ in2[17];
    assign G[59] = in1[16] & in2[16];
    assign P[59] = in1[16] ^ in2[16];
    assign G[60] = in1[15] & in2[15];
    assign P[60] = in1[15] ^ in2[15];
    assign G[61] = in1[14] & in2[14];
    assign P[61] = in1[14] ^ in2[14];
    assign G[62] = in1[13] & in2[13];
    assign P[62] = in1[13] ^ in2[13];
    assign G[63] = in1[12] & in2[12];
    assign P[63] = in1[12] ^ in2[12];
    assign G[64] = in1[11] & in2[11];
    assign P[64] = in1[11] ^ in2[11];
    assign G[65] = in1[10] & in2[10];
    assign P[65] = in1[10] ^ in2[10];
    assign G[66] = in1[9] & in2[9];
    assign P[66] = in1[9] ^ in2[9];
    assign G[67] = in1[8] & in2[8];
    assign P[67] = in1[8] ^ in2[8];
    assign G[68] = in1[7] & in2[7];
    assign P[68] = in1[7] ^ in2[7];
    assign G[69] = in1[6] & in2[6];
    assign P[69] = in1[6] ^ in2[6];
    assign G[70] = in1[5] & in2[5];
    assign P[70] = in1[5] ^ in2[5];
    assign G[71] = in1[4] & in2[4];
    assign P[71] = in1[4] ^ in2[4];
    assign G[72] = in1[3] & in2[3];
    assign P[72] = in1[3] ^ in2[3];
    assign G[73] = in1[2] & in2[2];
    assign P[73] = in1[2] ^ in2[2];
    assign G[74] = in1[1] & in2[1];
    assign P[74] = in1[1] ^ in2[1];
    assign G[75] = in1[0] & in2[0];
    assign P[75] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign cout = G[75] | (P[75] & C[75]);
    assign sum = P ^ C;
endmodule

module CLA_75(output [74:0] sum, output cout, input [74:0] in1, input [74:0] in2);

    wire[74:0] G;
    wire[74:0] C;
    wire[74:0] P;

    assign G[0] = in1[74] & in2[74];
    assign P[0] = in1[74] ^ in2[74];
    assign G[1] = in1[73] & in2[73];
    assign P[1] = in1[73] ^ in2[73];
    assign G[2] = in1[72] & in2[72];
    assign P[2] = in1[72] ^ in2[72];
    assign G[3] = in1[71] & in2[71];
    assign P[3] = in1[71] ^ in2[71];
    assign G[4] = in1[70] & in2[70];
    assign P[4] = in1[70] ^ in2[70];
    assign G[5] = in1[69] & in2[69];
    assign P[5] = in1[69] ^ in2[69];
    assign G[6] = in1[68] & in2[68];
    assign P[6] = in1[68] ^ in2[68];
    assign G[7] = in1[67] & in2[67];
    assign P[7] = in1[67] ^ in2[67];
    assign G[8] = in1[66] & in2[66];
    assign P[8] = in1[66] ^ in2[66];
    assign G[9] = in1[65] & in2[65];
    assign P[9] = in1[65] ^ in2[65];
    assign G[10] = in1[64] & in2[64];
    assign P[10] = in1[64] ^ in2[64];
    assign G[11] = in1[63] & in2[63];
    assign P[11] = in1[63] ^ in2[63];
    assign G[12] = in1[62] & in2[62];
    assign P[12] = in1[62] ^ in2[62];
    assign G[13] = in1[61] & in2[61];
    assign P[13] = in1[61] ^ in2[61];
    assign G[14] = in1[60] & in2[60];
    assign P[14] = in1[60] ^ in2[60];
    assign G[15] = in1[59] & in2[59];
    assign P[15] = in1[59] ^ in2[59];
    assign G[16] = in1[58] & in2[58];
    assign P[16] = in1[58] ^ in2[58];
    assign G[17] = in1[57] & in2[57];
    assign P[17] = in1[57] ^ in2[57];
    assign G[18] = in1[56] & in2[56];
    assign P[18] = in1[56] ^ in2[56];
    assign G[19] = in1[55] & in2[55];
    assign P[19] = in1[55] ^ in2[55];
    assign G[20] = in1[54] & in2[54];
    assign P[20] = in1[54] ^ in2[54];
    assign G[21] = in1[53] & in2[53];
    assign P[21] = in1[53] ^ in2[53];
    assign G[22] = in1[52] & in2[52];
    assign P[22] = in1[52] ^ in2[52];
    assign G[23] = in1[51] & in2[51];
    assign P[23] = in1[51] ^ in2[51];
    assign G[24] = in1[50] & in2[50];
    assign P[24] = in1[50] ^ in2[50];
    assign G[25] = in1[49] & in2[49];
    assign P[25] = in1[49] ^ in2[49];
    assign G[26] = in1[48] & in2[48];
    assign P[26] = in1[48] ^ in2[48];
    assign G[27] = in1[47] & in2[47];
    assign P[27] = in1[47] ^ in2[47];
    assign G[28] = in1[46] & in2[46];
    assign P[28] = in1[46] ^ in2[46];
    assign G[29] = in1[45] & in2[45];
    assign P[29] = in1[45] ^ in2[45];
    assign G[30] = in1[44] & in2[44];
    assign P[30] = in1[44] ^ in2[44];
    assign G[31] = in1[43] & in2[43];
    assign P[31] = in1[43] ^ in2[43];
    assign G[32] = in1[42] & in2[42];
    assign P[32] = in1[42] ^ in2[42];
    assign G[33] = in1[41] & in2[41];
    assign P[33] = in1[41] ^ in2[41];
    assign G[34] = in1[40] & in2[40];
    assign P[34] = in1[40] ^ in2[40];
    assign G[35] = in1[39] & in2[39];
    assign P[35] = in1[39] ^ in2[39];
    assign G[36] = in1[38] & in2[38];
    assign P[36] = in1[38] ^ in2[38];
    assign G[37] = in1[37] & in2[37];
    assign P[37] = in1[37] ^ in2[37];
    assign G[38] = in1[36] & in2[36];
    assign P[38] = in1[36] ^ in2[36];
    assign G[39] = in1[35] & in2[35];
    assign P[39] = in1[35] ^ in2[35];
    assign G[40] = in1[34] & in2[34];
    assign P[40] = in1[34] ^ in2[34];
    assign G[41] = in1[33] & in2[33];
    assign P[41] = in1[33] ^ in2[33];
    assign G[42] = in1[32] & in2[32];
    assign P[42] = in1[32] ^ in2[32];
    assign G[43] = in1[31] & in2[31];
    assign P[43] = in1[31] ^ in2[31];
    assign G[44] = in1[30] & in2[30];
    assign P[44] = in1[30] ^ in2[30];
    assign G[45] = in1[29] & in2[29];
    assign P[45] = in1[29] ^ in2[29];
    assign G[46] = in1[28] & in2[28];
    assign P[46] = in1[28] ^ in2[28];
    assign G[47] = in1[27] & in2[27];
    assign P[47] = in1[27] ^ in2[27];
    assign G[48] = in1[26] & in2[26];
    assign P[48] = in1[26] ^ in2[26];
    assign G[49] = in1[25] & in2[25];
    assign P[49] = in1[25] ^ in2[25];
    assign G[50] = in1[24] & in2[24];
    assign P[50] = in1[24] ^ in2[24];
    assign G[51] = in1[23] & in2[23];
    assign P[51] = in1[23] ^ in2[23];
    assign G[52] = in1[22] & in2[22];
    assign P[52] = in1[22] ^ in2[22];
    assign G[53] = in1[21] & in2[21];
    assign P[53] = in1[21] ^ in2[21];
    assign G[54] = in1[20] & in2[20];
    assign P[54] = in1[20] ^ in2[20];
    assign G[55] = in1[19] & in2[19];
    assign P[55] = in1[19] ^ in2[19];
    assign G[56] = in1[18] & in2[18];
    assign P[56] = in1[18] ^ in2[18];
    assign G[57] = in1[17] & in2[17];
    assign P[57] = in1[17] ^ in2[17];
    assign G[58] = in1[16] & in2[16];
    assign P[58] = in1[16] ^ in2[16];
    assign G[59] = in1[15] & in2[15];
    assign P[59] = in1[15] ^ in2[15];
    assign G[60] = in1[14] & in2[14];
    assign P[60] = in1[14] ^ in2[14];
    assign G[61] = in1[13] & in2[13];
    assign P[61] = in1[13] ^ in2[13];
    assign G[62] = in1[12] & in2[12];
    assign P[62] = in1[12] ^ in2[12];
    assign G[63] = in1[11] & in2[11];
    assign P[63] = in1[11] ^ in2[11];
    assign G[64] = in1[10] & in2[10];
    assign P[64] = in1[10] ^ in2[10];
    assign G[65] = in1[9] & in2[9];
    assign P[65] = in1[9] ^ in2[9];
    assign G[66] = in1[8] & in2[8];
    assign P[66] = in1[8] ^ in2[8];
    assign G[67] = in1[7] & in2[7];
    assign P[67] = in1[7] ^ in2[7];
    assign G[68] = in1[6] & in2[6];
    assign P[68] = in1[6] ^ in2[6];
    assign G[69] = in1[5] & in2[5];
    assign P[69] = in1[5] ^ in2[5];
    assign G[70] = in1[4] & in2[4];
    assign P[70] = in1[4] ^ in2[4];
    assign G[71] = in1[3] & in2[3];
    assign P[71] = in1[3] ^ in2[3];
    assign G[72] = in1[2] & in2[2];
    assign P[72] = in1[2] ^ in2[2];
    assign G[73] = in1[1] & in2[1];
    assign P[73] = in1[1] ^ in2[1];
    assign G[74] = in1[0] & in2[0];
    assign P[74] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign cout = G[74] | (P[74] & C[74]);
    assign sum = P ^ C;
endmodule

module CLA_74(output [73:0] sum, output cout, input [73:0] in1, input [73:0] in2);

    wire[73:0] G;
    wire[73:0] C;
    wire[73:0] P;

    assign G[0] = in1[73] & in2[73];
    assign P[0] = in1[73] ^ in2[73];
    assign G[1] = in1[72] & in2[72];
    assign P[1] = in1[72] ^ in2[72];
    assign G[2] = in1[71] & in2[71];
    assign P[2] = in1[71] ^ in2[71];
    assign G[3] = in1[70] & in2[70];
    assign P[3] = in1[70] ^ in2[70];
    assign G[4] = in1[69] & in2[69];
    assign P[4] = in1[69] ^ in2[69];
    assign G[5] = in1[68] & in2[68];
    assign P[5] = in1[68] ^ in2[68];
    assign G[6] = in1[67] & in2[67];
    assign P[6] = in1[67] ^ in2[67];
    assign G[7] = in1[66] & in2[66];
    assign P[7] = in1[66] ^ in2[66];
    assign G[8] = in1[65] & in2[65];
    assign P[8] = in1[65] ^ in2[65];
    assign G[9] = in1[64] & in2[64];
    assign P[9] = in1[64] ^ in2[64];
    assign G[10] = in1[63] & in2[63];
    assign P[10] = in1[63] ^ in2[63];
    assign G[11] = in1[62] & in2[62];
    assign P[11] = in1[62] ^ in2[62];
    assign G[12] = in1[61] & in2[61];
    assign P[12] = in1[61] ^ in2[61];
    assign G[13] = in1[60] & in2[60];
    assign P[13] = in1[60] ^ in2[60];
    assign G[14] = in1[59] & in2[59];
    assign P[14] = in1[59] ^ in2[59];
    assign G[15] = in1[58] & in2[58];
    assign P[15] = in1[58] ^ in2[58];
    assign G[16] = in1[57] & in2[57];
    assign P[16] = in1[57] ^ in2[57];
    assign G[17] = in1[56] & in2[56];
    assign P[17] = in1[56] ^ in2[56];
    assign G[18] = in1[55] & in2[55];
    assign P[18] = in1[55] ^ in2[55];
    assign G[19] = in1[54] & in2[54];
    assign P[19] = in1[54] ^ in2[54];
    assign G[20] = in1[53] & in2[53];
    assign P[20] = in1[53] ^ in2[53];
    assign G[21] = in1[52] & in2[52];
    assign P[21] = in1[52] ^ in2[52];
    assign G[22] = in1[51] & in2[51];
    assign P[22] = in1[51] ^ in2[51];
    assign G[23] = in1[50] & in2[50];
    assign P[23] = in1[50] ^ in2[50];
    assign G[24] = in1[49] & in2[49];
    assign P[24] = in1[49] ^ in2[49];
    assign G[25] = in1[48] & in2[48];
    assign P[25] = in1[48] ^ in2[48];
    assign G[26] = in1[47] & in2[47];
    assign P[26] = in1[47] ^ in2[47];
    assign G[27] = in1[46] & in2[46];
    assign P[27] = in1[46] ^ in2[46];
    assign G[28] = in1[45] & in2[45];
    assign P[28] = in1[45] ^ in2[45];
    assign G[29] = in1[44] & in2[44];
    assign P[29] = in1[44] ^ in2[44];
    assign G[30] = in1[43] & in2[43];
    assign P[30] = in1[43] ^ in2[43];
    assign G[31] = in1[42] & in2[42];
    assign P[31] = in1[42] ^ in2[42];
    assign G[32] = in1[41] & in2[41];
    assign P[32] = in1[41] ^ in2[41];
    assign G[33] = in1[40] & in2[40];
    assign P[33] = in1[40] ^ in2[40];
    assign G[34] = in1[39] & in2[39];
    assign P[34] = in1[39] ^ in2[39];
    assign G[35] = in1[38] & in2[38];
    assign P[35] = in1[38] ^ in2[38];
    assign G[36] = in1[37] & in2[37];
    assign P[36] = in1[37] ^ in2[37];
    assign G[37] = in1[36] & in2[36];
    assign P[37] = in1[36] ^ in2[36];
    assign G[38] = in1[35] & in2[35];
    assign P[38] = in1[35] ^ in2[35];
    assign G[39] = in1[34] & in2[34];
    assign P[39] = in1[34] ^ in2[34];
    assign G[40] = in1[33] & in2[33];
    assign P[40] = in1[33] ^ in2[33];
    assign G[41] = in1[32] & in2[32];
    assign P[41] = in1[32] ^ in2[32];
    assign G[42] = in1[31] & in2[31];
    assign P[42] = in1[31] ^ in2[31];
    assign G[43] = in1[30] & in2[30];
    assign P[43] = in1[30] ^ in2[30];
    assign G[44] = in1[29] & in2[29];
    assign P[44] = in1[29] ^ in2[29];
    assign G[45] = in1[28] & in2[28];
    assign P[45] = in1[28] ^ in2[28];
    assign G[46] = in1[27] & in2[27];
    assign P[46] = in1[27] ^ in2[27];
    assign G[47] = in1[26] & in2[26];
    assign P[47] = in1[26] ^ in2[26];
    assign G[48] = in1[25] & in2[25];
    assign P[48] = in1[25] ^ in2[25];
    assign G[49] = in1[24] & in2[24];
    assign P[49] = in1[24] ^ in2[24];
    assign G[50] = in1[23] & in2[23];
    assign P[50] = in1[23] ^ in2[23];
    assign G[51] = in1[22] & in2[22];
    assign P[51] = in1[22] ^ in2[22];
    assign G[52] = in1[21] & in2[21];
    assign P[52] = in1[21] ^ in2[21];
    assign G[53] = in1[20] & in2[20];
    assign P[53] = in1[20] ^ in2[20];
    assign G[54] = in1[19] & in2[19];
    assign P[54] = in1[19] ^ in2[19];
    assign G[55] = in1[18] & in2[18];
    assign P[55] = in1[18] ^ in2[18];
    assign G[56] = in1[17] & in2[17];
    assign P[56] = in1[17] ^ in2[17];
    assign G[57] = in1[16] & in2[16];
    assign P[57] = in1[16] ^ in2[16];
    assign G[58] = in1[15] & in2[15];
    assign P[58] = in1[15] ^ in2[15];
    assign G[59] = in1[14] & in2[14];
    assign P[59] = in1[14] ^ in2[14];
    assign G[60] = in1[13] & in2[13];
    assign P[60] = in1[13] ^ in2[13];
    assign G[61] = in1[12] & in2[12];
    assign P[61] = in1[12] ^ in2[12];
    assign G[62] = in1[11] & in2[11];
    assign P[62] = in1[11] ^ in2[11];
    assign G[63] = in1[10] & in2[10];
    assign P[63] = in1[10] ^ in2[10];
    assign G[64] = in1[9] & in2[9];
    assign P[64] = in1[9] ^ in2[9];
    assign G[65] = in1[8] & in2[8];
    assign P[65] = in1[8] ^ in2[8];
    assign G[66] = in1[7] & in2[7];
    assign P[66] = in1[7] ^ in2[7];
    assign G[67] = in1[6] & in2[6];
    assign P[67] = in1[6] ^ in2[6];
    assign G[68] = in1[5] & in2[5];
    assign P[68] = in1[5] ^ in2[5];
    assign G[69] = in1[4] & in2[4];
    assign P[69] = in1[4] ^ in2[4];
    assign G[70] = in1[3] & in2[3];
    assign P[70] = in1[3] ^ in2[3];
    assign G[71] = in1[2] & in2[2];
    assign P[71] = in1[2] ^ in2[2];
    assign G[72] = in1[1] & in2[1];
    assign P[72] = in1[1] ^ in2[1];
    assign G[73] = in1[0] & in2[0];
    assign P[73] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign cout = G[73] | (P[73] & C[73]);
    assign sum = P ^ C;
endmodule

module CLA_73(output [72:0] sum, output cout, input [72:0] in1, input [72:0] in2);

    wire[72:0] G;
    wire[72:0] C;
    wire[72:0] P;

    assign G[0] = in1[72] & in2[72];
    assign P[0] = in1[72] ^ in2[72];
    assign G[1] = in1[71] & in2[71];
    assign P[1] = in1[71] ^ in2[71];
    assign G[2] = in1[70] & in2[70];
    assign P[2] = in1[70] ^ in2[70];
    assign G[3] = in1[69] & in2[69];
    assign P[3] = in1[69] ^ in2[69];
    assign G[4] = in1[68] & in2[68];
    assign P[4] = in1[68] ^ in2[68];
    assign G[5] = in1[67] & in2[67];
    assign P[5] = in1[67] ^ in2[67];
    assign G[6] = in1[66] & in2[66];
    assign P[6] = in1[66] ^ in2[66];
    assign G[7] = in1[65] & in2[65];
    assign P[7] = in1[65] ^ in2[65];
    assign G[8] = in1[64] & in2[64];
    assign P[8] = in1[64] ^ in2[64];
    assign G[9] = in1[63] & in2[63];
    assign P[9] = in1[63] ^ in2[63];
    assign G[10] = in1[62] & in2[62];
    assign P[10] = in1[62] ^ in2[62];
    assign G[11] = in1[61] & in2[61];
    assign P[11] = in1[61] ^ in2[61];
    assign G[12] = in1[60] & in2[60];
    assign P[12] = in1[60] ^ in2[60];
    assign G[13] = in1[59] & in2[59];
    assign P[13] = in1[59] ^ in2[59];
    assign G[14] = in1[58] & in2[58];
    assign P[14] = in1[58] ^ in2[58];
    assign G[15] = in1[57] & in2[57];
    assign P[15] = in1[57] ^ in2[57];
    assign G[16] = in1[56] & in2[56];
    assign P[16] = in1[56] ^ in2[56];
    assign G[17] = in1[55] & in2[55];
    assign P[17] = in1[55] ^ in2[55];
    assign G[18] = in1[54] & in2[54];
    assign P[18] = in1[54] ^ in2[54];
    assign G[19] = in1[53] & in2[53];
    assign P[19] = in1[53] ^ in2[53];
    assign G[20] = in1[52] & in2[52];
    assign P[20] = in1[52] ^ in2[52];
    assign G[21] = in1[51] & in2[51];
    assign P[21] = in1[51] ^ in2[51];
    assign G[22] = in1[50] & in2[50];
    assign P[22] = in1[50] ^ in2[50];
    assign G[23] = in1[49] & in2[49];
    assign P[23] = in1[49] ^ in2[49];
    assign G[24] = in1[48] & in2[48];
    assign P[24] = in1[48] ^ in2[48];
    assign G[25] = in1[47] & in2[47];
    assign P[25] = in1[47] ^ in2[47];
    assign G[26] = in1[46] & in2[46];
    assign P[26] = in1[46] ^ in2[46];
    assign G[27] = in1[45] & in2[45];
    assign P[27] = in1[45] ^ in2[45];
    assign G[28] = in1[44] & in2[44];
    assign P[28] = in1[44] ^ in2[44];
    assign G[29] = in1[43] & in2[43];
    assign P[29] = in1[43] ^ in2[43];
    assign G[30] = in1[42] & in2[42];
    assign P[30] = in1[42] ^ in2[42];
    assign G[31] = in1[41] & in2[41];
    assign P[31] = in1[41] ^ in2[41];
    assign G[32] = in1[40] & in2[40];
    assign P[32] = in1[40] ^ in2[40];
    assign G[33] = in1[39] & in2[39];
    assign P[33] = in1[39] ^ in2[39];
    assign G[34] = in1[38] & in2[38];
    assign P[34] = in1[38] ^ in2[38];
    assign G[35] = in1[37] & in2[37];
    assign P[35] = in1[37] ^ in2[37];
    assign G[36] = in1[36] & in2[36];
    assign P[36] = in1[36] ^ in2[36];
    assign G[37] = in1[35] & in2[35];
    assign P[37] = in1[35] ^ in2[35];
    assign G[38] = in1[34] & in2[34];
    assign P[38] = in1[34] ^ in2[34];
    assign G[39] = in1[33] & in2[33];
    assign P[39] = in1[33] ^ in2[33];
    assign G[40] = in1[32] & in2[32];
    assign P[40] = in1[32] ^ in2[32];
    assign G[41] = in1[31] & in2[31];
    assign P[41] = in1[31] ^ in2[31];
    assign G[42] = in1[30] & in2[30];
    assign P[42] = in1[30] ^ in2[30];
    assign G[43] = in1[29] & in2[29];
    assign P[43] = in1[29] ^ in2[29];
    assign G[44] = in1[28] & in2[28];
    assign P[44] = in1[28] ^ in2[28];
    assign G[45] = in1[27] & in2[27];
    assign P[45] = in1[27] ^ in2[27];
    assign G[46] = in1[26] & in2[26];
    assign P[46] = in1[26] ^ in2[26];
    assign G[47] = in1[25] & in2[25];
    assign P[47] = in1[25] ^ in2[25];
    assign G[48] = in1[24] & in2[24];
    assign P[48] = in1[24] ^ in2[24];
    assign G[49] = in1[23] & in2[23];
    assign P[49] = in1[23] ^ in2[23];
    assign G[50] = in1[22] & in2[22];
    assign P[50] = in1[22] ^ in2[22];
    assign G[51] = in1[21] & in2[21];
    assign P[51] = in1[21] ^ in2[21];
    assign G[52] = in1[20] & in2[20];
    assign P[52] = in1[20] ^ in2[20];
    assign G[53] = in1[19] & in2[19];
    assign P[53] = in1[19] ^ in2[19];
    assign G[54] = in1[18] & in2[18];
    assign P[54] = in1[18] ^ in2[18];
    assign G[55] = in1[17] & in2[17];
    assign P[55] = in1[17] ^ in2[17];
    assign G[56] = in1[16] & in2[16];
    assign P[56] = in1[16] ^ in2[16];
    assign G[57] = in1[15] & in2[15];
    assign P[57] = in1[15] ^ in2[15];
    assign G[58] = in1[14] & in2[14];
    assign P[58] = in1[14] ^ in2[14];
    assign G[59] = in1[13] & in2[13];
    assign P[59] = in1[13] ^ in2[13];
    assign G[60] = in1[12] & in2[12];
    assign P[60] = in1[12] ^ in2[12];
    assign G[61] = in1[11] & in2[11];
    assign P[61] = in1[11] ^ in2[11];
    assign G[62] = in1[10] & in2[10];
    assign P[62] = in1[10] ^ in2[10];
    assign G[63] = in1[9] & in2[9];
    assign P[63] = in1[9] ^ in2[9];
    assign G[64] = in1[8] & in2[8];
    assign P[64] = in1[8] ^ in2[8];
    assign G[65] = in1[7] & in2[7];
    assign P[65] = in1[7] ^ in2[7];
    assign G[66] = in1[6] & in2[6];
    assign P[66] = in1[6] ^ in2[6];
    assign G[67] = in1[5] & in2[5];
    assign P[67] = in1[5] ^ in2[5];
    assign G[68] = in1[4] & in2[4];
    assign P[68] = in1[4] ^ in2[4];
    assign G[69] = in1[3] & in2[3];
    assign P[69] = in1[3] ^ in2[3];
    assign G[70] = in1[2] & in2[2];
    assign P[70] = in1[2] ^ in2[2];
    assign G[71] = in1[1] & in2[1];
    assign P[71] = in1[1] ^ in2[1];
    assign G[72] = in1[0] & in2[0];
    assign P[72] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign cout = G[72] | (P[72] & C[72]);
    assign sum = P ^ C;
endmodule

module CLA_72(output [71:0] sum, output cout, input [71:0] in1, input [71:0] in2);

    wire[71:0] G;
    wire[71:0] C;
    wire[71:0] P;

    assign G[0] = in1[71] & in2[71];
    assign P[0] = in1[71] ^ in2[71];
    assign G[1] = in1[70] & in2[70];
    assign P[1] = in1[70] ^ in2[70];
    assign G[2] = in1[69] & in2[69];
    assign P[2] = in1[69] ^ in2[69];
    assign G[3] = in1[68] & in2[68];
    assign P[3] = in1[68] ^ in2[68];
    assign G[4] = in1[67] & in2[67];
    assign P[4] = in1[67] ^ in2[67];
    assign G[5] = in1[66] & in2[66];
    assign P[5] = in1[66] ^ in2[66];
    assign G[6] = in1[65] & in2[65];
    assign P[6] = in1[65] ^ in2[65];
    assign G[7] = in1[64] & in2[64];
    assign P[7] = in1[64] ^ in2[64];
    assign G[8] = in1[63] & in2[63];
    assign P[8] = in1[63] ^ in2[63];
    assign G[9] = in1[62] & in2[62];
    assign P[9] = in1[62] ^ in2[62];
    assign G[10] = in1[61] & in2[61];
    assign P[10] = in1[61] ^ in2[61];
    assign G[11] = in1[60] & in2[60];
    assign P[11] = in1[60] ^ in2[60];
    assign G[12] = in1[59] & in2[59];
    assign P[12] = in1[59] ^ in2[59];
    assign G[13] = in1[58] & in2[58];
    assign P[13] = in1[58] ^ in2[58];
    assign G[14] = in1[57] & in2[57];
    assign P[14] = in1[57] ^ in2[57];
    assign G[15] = in1[56] & in2[56];
    assign P[15] = in1[56] ^ in2[56];
    assign G[16] = in1[55] & in2[55];
    assign P[16] = in1[55] ^ in2[55];
    assign G[17] = in1[54] & in2[54];
    assign P[17] = in1[54] ^ in2[54];
    assign G[18] = in1[53] & in2[53];
    assign P[18] = in1[53] ^ in2[53];
    assign G[19] = in1[52] & in2[52];
    assign P[19] = in1[52] ^ in2[52];
    assign G[20] = in1[51] & in2[51];
    assign P[20] = in1[51] ^ in2[51];
    assign G[21] = in1[50] & in2[50];
    assign P[21] = in1[50] ^ in2[50];
    assign G[22] = in1[49] & in2[49];
    assign P[22] = in1[49] ^ in2[49];
    assign G[23] = in1[48] & in2[48];
    assign P[23] = in1[48] ^ in2[48];
    assign G[24] = in1[47] & in2[47];
    assign P[24] = in1[47] ^ in2[47];
    assign G[25] = in1[46] & in2[46];
    assign P[25] = in1[46] ^ in2[46];
    assign G[26] = in1[45] & in2[45];
    assign P[26] = in1[45] ^ in2[45];
    assign G[27] = in1[44] & in2[44];
    assign P[27] = in1[44] ^ in2[44];
    assign G[28] = in1[43] & in2[43];
    assign P[28] = in1[43] ^ in2[43];
    assign G[29] = in1[42] & in2[42];
    assign P[29] = in1[42] ^ in2[42];
    assign G[30] = in1[41] & in2[41];
    assign P[30] = in1[41] ^ in2[41];
    assign G[31] = in1[40] & in2[40];
    assign P[31] = in1[40] ^ in2[40];
    assign G[32] = in1[39] & in2[39];
    assign P[32] = in1[39] ^ in2[39];
    assign G[33] = in1[38] & in2[38];
    assign P[33] = in1[38] ^ in2[38];
    assign G[34] = in1[37] & in2[37];
    assign P[34] = in1[37] ^ in2[37];
    assign G[35] = in1[36] & in2[36];
    assign P[35] = in1[36] ^ in2[36];
    assign G[36] = in1[35] & in2[35];
    assign P[36] = in1[35] ^ in2[35];
    assign G[37] = in1[34] & in2[34];
    assign P[37] = in1[34] ^ in2[34];
    assign G[38] = in1[33] & in2[33];
    assign P[38] = in1[33] ^ in2[33];
    assign G[39] = in1[32] & in2[32];
    assign P[39] = in1[32] ^ in2[32];
    assign G[40] = in1[31] & in2[31];
    assign P[40] = in1[31] ^ in2[31];
    assign G[41] = in1[30] & in2[30];
    assign P[41] = in1[30] ^ in2[30];
    assign G[42] = in1[29] & in2[29];
    assign P[42] = in1[29] ^ in2[29];
    assign G[43] = in1[28] & in2[28];
    assign P[43] = in1[28] ^ in2[28];
    assign G[44] = in1[27] & in2[27];
    assign P[44] = in1[27] ^ in2[27];
    assign G[45] = in1[26] & in2[26];
    assign P[45] = in1[26] ^ in2[26];
    assign G[46] = in1[25] & in2[25];
    assign P[46] = in1[25] ^ in2[25];
    assign G[47] = in1[24] & in2[24];
    assign P[47] = in1[24] ^ in2[24];
    assign G[48] = in1[23] & in2[23];
    assign P[48] = in1[23] ^ in2[23];
    assign G[49] = in1[22] & in2[22];
    assign P[49] = in1[22] ^ in2[22];
    assign G[50] = in1[21] & in2[21];
    assign P[50] = in1[21] ^ in2[21];
    assign G[51] = in1[20] & in2[20];
    assign P[51] = in1[20] ^ in2[20];
    assign G[52] = in1[19] & in2[19];
    assign P[52] = in1[19] ^ in2[19];
    assign G[53] = in1[18] & in2[18];
    assign P[53] = in1[18] ^ in2[18];
    assign G[54] = in1[17] & in2[17];
    assign P[54] = in1[17] ^ in2[17];
    assign G[55] = in1[16] & in2[16];
    assign P[55] = in1[16] ^ in2[16];
    assign G[56] = in1[15] & in2[15];
    assign P[56] = in1[15] ^ in2[15];
    assign G[57] = in1[14] & in2[14];
    assign P[57] = in1[14] ^ in2[14];
    assign G[58] = in1[13] & in2[13];
    assign P[58] = in1[13] ^ in2[13];
    assign G[59] = in1[12] & in2[12];
    assign P[59] = in1[12] ^ in2[12];
    assign G[60] = in1[11] & in2[11];
    assign P[60] = in1[11] ^ in2[11];
    assign G[61] = in1[10] & in2[10];
    assign P[61] = in1[10] ^ in2[10];
    assign G[62] = in1[9] & in2[9];
    assign P[62] = in1[9] ^ in2[9];
    assign G[63] = in1[8] & in2[8];
    assign P[63] = in1[8] ^ in2[8];
    assign G[64] = in1[7] & in2[7];
    assign P[64] = in1[7] ^ in2[7];
    assign G[65] = in1[6] & in2[6];
    assign P[65] = in1[6] ^ in2[6];
    assign G[66] = in1[5] & in2[5];
    assign P[66] = in1[5] ^ in2[5];
    assign G[67] = in1[4] & in2[4];
    assign P[67] = in1[4] ^ in2[4];
    assign G[68] = in1[3] & in2[3];
    assign P[68] = in1[3] ^ in2[3];
    assign G[69] = in1[2] & in2[2];
    assign P[69] = in1[2] ^ in2[2];
    assign G[70] = in1[1] & in2[1];
    assign P[70] = in1[1] ^ in2[1];
    assign G[71] = in1[0] & in2[0];
    assign P[71] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign cout = G[71] | (P[71] & C[71]);
    assign sum = P ^ C;
endmodule

module CLA_71(output [70:0] sum, output cout, input [70:0] in1, input [70:0] in2);

    wire[70:0] G;
    wire[70:0] C;
    wire[70:0] P;

    assign G[0] = in1[70] & in2[70];
    assign P[0] = in1[70] ^ in2[70];
    assign G[1] = in1[69] & in2[69];
    assign P[1] = in1[69] ^ in2[69];
    assign G[2] = in1[68] & in2[68];
    assign P[2] = in1[68] ^ in2[68];
    assign G[3] = in1[67] & in2[67];
    assign P[3] = in1[67] ^ in2[67];
    assign G[4] = in1[66] & in2[66];
    assign P[4] = in1[66] ^ in2[66];
    assign G[5] = in1[65] & in2[65];
    assign P[5] = in1[65] ^ in2[65];
    assign G[6] = in1[64] & in2[64];
    assign P[6] = in1[64] ^ in2[64];
    assign G[7] = in1[63] & in2[63];
    assign P[7] = in1[63] ^ in2[63];
    assign G[8] = in1[62] & in2[62];
    assign P[8] = in1[62] ^ in2[62];
    assign G[9] = in1[61] & in2[61];
    assign P[9] = in1[61] ^ in2[61];
    assign G[10] = in1[60] & in2[60];
    assign P[10] = in1[60] ^ in2[60];
    assign G[11] = in1[59] & in2[59];
    assign P[11] = in1[59] ^ in2[59];
    assign G[12] = in1[58] & in2[58];
    assign P[12] = in1[58] ^ in2[58];
    assign G[13] = in1[57] & in2[57];
    assign P[13] = in1[57] ^ in2[57];
    assign G[14] = in1[56] & in2[56];
    assign P[14] = in1[56] ^ in2[56];
    assign G[15] = in1[55] & in2[55];
    assign P[15] = in1[55] ^ in2[55];
    assign G[16] = in1[54] & in2[54];
    assign P[16] = in1[54] ^ in2[54];
    assign G[17] = in1[53] & in2[53];
    assign P[17] = in1[53] ^ in2[53];
    assign G[18] = in1[52] & in2[52];
    assign P[18] = in1[52] ^ in2[52];
    assign G[19] = in1[51] & in2[51];
    assign P[19] = in1[51] ^ in2[51];
    assign G[20] = in1[50] & in2[50];
    assign P[20] = in1[50] ^ in2[50];
    assign G[21] = in1[49] & in2[49];
    assign P[21] = in1[49] ^ in2[49];
    assign G[22] = in1[48] & in2[48];
    assign P[22] = in1[48] ^ in2[48];
    assign G[23] = in1[47] & in2[47];
    assign P[23] = in1[47] ^ in2[47];
    assign G[24] = in1[46] & in2[46];
    assign P[24] = in1[46] ^ in2[46];
    assign G[25] = in1[45] & in2[45];
    assign P[25] = in1[45] ^ in2[45];
    assign G[26] = in1[44] & in2[44];
    assign P[26] = in1[44] ^ in2[44];
    assign G[27] = in1[43] & in2[43];
    assign P[27] = in1[43] ^ in2[43];
    assign G[28] = in1[42] & in2[42];
    assign P[28] = in1[42] ^ in2[42];
    assign G[29] = in1[41] & in2[41];
    assign P[29] = in1[41] ^ in2[41];
    assign G[30] = in1[40] & in2[40];
    assign P[30] = in1[40] ^ in2[40];
    assign G[31] = in1[39] & in2[39];
    assign P[31] = in1[39] ^ in2[39];
    assign G[32] = in1[38] & in2[38];
    assign P[32] = in1[38] ^ in2[38];
    assign G[33] = in1[37] & in2[37];
    assign P[33] = in1[37] ^ in2[37];
    assign G[34] = in1[36] & in2[36];
    assign P[34] = in1[36] ^ in2[36];
    assign G[35] = in1[35] & in2[35];
    assign P[35] = in1[35] ^ in2[35];
    assign G[36] = in1[34] & in2[34];
    assign P[36] = in1[34] ^ in2[34];
    assign G[37] = in1[33] & in2[33];
    assign P[37] = in1[33] ^ in2[33];
    assign G[38] = in1[32] & in2[32];
    assign P[38] = in1[32] ^ in2[32];
    assign G[39] = in1[31] & in2[31];
    assign P[39] = in1[31] ^ in2[31];
    assign G[40] = in1[30] & in2[30];
    assign P[40] = in1[30] ^ in2[30];
    assign G[41] = in1[29] & in2[29];
    assign P[41] = in1[29] ^ in2[29];
    assign G[42] = in1[28] & in2[28];
    assign P[42] = in1[28] ^ in2[28];
    assign G[43] = in1[27] & in2[27];
    assign P[43] = in1[27] ^ in2[27];
    assign G[44] = in1[26] & in2[26];
    assign P[44] = in1[26] ^ in2[26];
    assign G[45] = in1[25] & in2[25];
    assign P[45] = in1[25] ^ in2[25];
    assign G[46] = in1[24] & in2[24];
    assign P[46] = in1[24] ^ in2[24];
    assign G[47] = in1[23] & in2[23];
    assign P[47] = in1[23] ^ in2[23];
    assign G[48] = in1[22] & in2[22];
    assign P[48] = in1[22] ^ in2[22];
    assign G[49] = in1[21] & in2[21];
    assign P[49] = in1[21] ^ in2[21];
    assign G[50] = in1[20] & in2[20];
    assign P[50] = in1[20] ^ in2[20];
    assign G[51] = in1[19] & in2[19];
    assign P[51] = in1[19] ^ in2[19];
    assign G[52] = in1[18] & in2[18];
    assign P[52] = in1[18] ^ in2[18];
    assign G[53] = in1[17] & in2[17];
    assign P[53] = in1[17] ^ in2[17];
    assign G[54] = in1[16] & in2[16];
    assign P[54] = in1[16] ^ in2[16];
    assign G[55] = in1[15] & in2[15];
    assign P[55] = in1[15] ^ in2[15];
    assign G[56] = in1[14] & in2[14];
    assign P[56] = in1[14] ^ in2[14];
    assign G[57] = in1[13] & in2[13];
    assign P[57] = in1[13] ^ in2[13];
    assign G[58] = in1[12] & in2[12];
    assign P[58] = in1[12] ^ in2[12];
    assign G[59] = in1[11] & in2[11];
    assign P[59] = in1[11] ^ in2[11];
    assign G[60] = in1[10] & in2[10];
    assign P[60] = in1[10] ^ in2[10];
    assign G[61] = in1[9] & in2[9];
    assign P[61] = in1[9] ^ in2[9];
    assign G[62] = in1[8] & in2[8];
    assign P[62] = in1[8] ^ in2[8];
    assign G[63] = in1[7] & in2[7];
    assign P[63] = in1[7] ^ in2[7];
    assign G[64] = in1[6] & in2[6];
    assign P[64] = in1[6] ^ in2[6];
    assign G[65] = in1[5] & in2[5];
    assign P[65] = in1[5] ^ in2[5];
    assign G[66] = in1[4] & in2[4];
    assign P[66] = in1[4] ^ in2[4];
    assign G[67] = in1[3] & in2[3];
    assign P[67] = in1[3] ^ in2[3];
    assign G[68] = in1[2] & in2[2];
    assign P[68] = in1[2] ^ in2[2];
    assign G[69] = in1[1] & in2[1];
    assign P[69] = in1[1] ^ in2[1];
    assign G[70] = in1[0] & in2[0];
    assign P[70] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign cout = G[70] | (P[70] & C[70]);
    assign sum = P ^ C;
endmodule

module CLA_70(output [69:0] sum, output cout, input [69:0] in1, input [69:0] in2);

    wire[69:0] G;
    wire[69:0] C;
    wire[69:0] P;

    assign G[0] = in1[69] & in2[69];
    assign P[0] = in1[69] ^ in2[69];
    assign G[1] = in1[68] & in2[68];
    assign P[1] = in1[68] ^ in2[68];
    assign G[2] = in1[67] & in2[67];
    assign P[2] = in1[67] ^ in2[67];
    assign G[3] = in1[66] & in2[66];
    assign P[3] = in1[66] ^ in2[66];
    assign G[4] = in1[65] & in2[65];
    assign P[4] = in1[65] ^ in2[65];
    assign G[5] = in1[64] & in2[64];
    assign P[5] = in1[64] ^ in2[64];
    assign G[6] = in1[63] & in2[63];
    assign P[6] = in1[63] ^ in2[63];
    assign G[7] = in1[62] & in2[62];
    assign P[7] = in1[62] ^ in2[62];
    assign G[8] = in1[61] & in2[61];
    assign P[8] = in1[61] ^ in2[61];
    assign G[9] = in1[60] & in2[60];
    assign P[9] = in1[60] ^ in2[60];
    assign G[10] = in1[59] & in2[59];
    assign P[10] = in1[59] ^ in2[59];
    assign G[11] = in1[58] & in2[58];
    assign P[11] = in1[58] ^ in2[58];
    assign G[12] = in1[57] & in2[57];
    assign P[12] = in1[57] ^ in2[57];
    assign G[13] = in1[56] & in2[56];
    assign P[13] = in1[56] ^ in2[56];
    assign G[14] = in1[55] & in2[55];
    assign P[14] = in1[55] ^ in2[55];
    assign G[15] = in1[54] & in2[54];
    assign P[15] = in1[54] ^ in2[54];
    assign G[16] = in1[53] & in2[53];
    assign P[16] = in1[53] ^ in2[53];
    assign G[17] = in1[52] & in2[52];
    assign P[17] = in1[52] ^ in2[52];
    assign G[18] = in1[51] & in2[51];
    assign P[18] = in1[51] ^ in2[51];
    assign G[19] = in1[50] & in2[50];
    assign P[19] = in1[50] ^ in2[50];
    assign G[20] = in1[49] & in2[49];
    assign P[20] = in1[49] ^ in2[49];
    assign G[21] = in1[48] & in2[48];
    assign P[21] = in1[48] ^ in2[48];
    assign G[22] = in1[47] & in2[47];
    assign P[22] = in1[47] ^ in2[47];
    assign G[23] = in1[46] & in2[46];
    assign P[23] = in1[46] ^ in2[46];
    assign G[24] = in1[45] & in2[45];
    assign P[24] = in1[45] ^ in2[45];
    assign G[25] = in1[44] & in2[44];
    assign P[25] = in1[44] ^ in2[44];
    assign G[26] = in1[43] & in2[43];
    assign P[26] = in1[43] ^ in2[43];
    assign G[27] = in1[42] & in2[42];
    assign P[27] = in1[42] ^ in2[42];
    assign G[28] = in1[41] & in2[41];
    assign P[28] = in1[41] ^ in2[41];
    assign G[29] = in1[40] & in2[40];
    assign P[29] = in1[40] ^ in2[40];
    assign G[30] = in1[39] & in2[39];
    assign P[30] = in1[39] ^ in2[39];
    assign G[31] = in1[38] & in2[38];
    assign P[31] = in1[38] ^ in2[38];
    assign G[32] = in1[37] & in2[37];
    assign P[32] = in1[37] ^ in2[37];
    assign G[33] = in1[36] & in2[36];
    assign P[33] = in1[36] ^ in2[36];
    assign G[34] = in1[35] & in2[35];
    assign P[34] = in1[35] ^ in2[35];
    assign G[35] = in1[34] & in2[34];
    assign P[35] = in1[34] ^ in2[34];
    assign G[36] = in1[33] & in2[33];
    assign P[36] = in1[33] ^ in2[33];
    assign G[37] = in1[32] & in2[32];
    assign P[37] = in1[32] ^ in2[32];
    assign G[38] = in1[31] & in2[31];
    assign P[38] = in1[31] ^ in2[31];
    assign G[39] = in1[30] & in2[30];
    assign P[39] = in1[30] ^ in2[30];
    assign G[40] = in1[29] & in2[29];
    assign P[40] = in1[29] ^ in2[29];
    assign G[41] = in1[28] & in2[28];
    assign P[41] = in1[28] ^ in2[28];
    assign G[42] = in1[27] & in2[27];
    assign P[42] = in1[27] ^ in2[27];
    assign G[43] = in1[26] & in2[26];
    assign P[43] = in1[26] ^ in2[26];
    assign G[44] = in1[25] & in2[25];
    assign P[44] = in1[25] ^ in2[25];
    assign G[45] = in1[24] & in2[24];
    assign P[45] = in1[24] ^ in2[24];
    assign G[46] = in1[23] & in2[23];
    assign P[46] = in1[23] ^ in2[23];
    assign G[47] = in1[22] & in2[22];
    assign P[47] = in1[22] ^ in2[22];
    assign G[48] = in1[21] & in2[21];
    assign P[48] = in1[21] ^ in2[21];
    assign G[49] = in1[20] & in2[20];
    assign P[49] = in1[20] ^ in2[20];
    assign G[50] = in1[19] & in2[19];
    assign P[50] = in1[19] ^ in2[19];
    assign G[51] = in1[18] & in2[18];
    assign P[51] = in1[18] ^ in2[18];
    assign G[52] = in1[17] & in2[17];
    assign P[52] = in1[17] ^ in2[17];
    assign G[53] = in1[16] & in2[16];
    assign P[53] = in1[16] ^ in2[16];
    assign G[54] = in1[15] & in2[15];
    assign P[54] = in1[15] ^ in2[15];
    assign G[55] = in1[14] & in2[14];
    assign P[55] = in1[14] ^ in2[14];
    assign G[56] = in1[13] & in2[13];
    assign P[56] = in1[13] ^ in2[13];
    assign G[57] = in1[12] & in2[12];
    assign P[57] = in1[12] ^ in2[12];
    assign G[58] = in1[11] & in2[11];
    assign P[58] = in1[11] ^ in2[11];
    assign G[59] = in1[10] & in2[10];
    assign P[59] = in1[10] ^ in2[10];
    assign G[60] = in1[9] & in2[9];
    assign P[60] = in1[9] ^ in2[9];
    assign G[61] = in1[8] & in2[8];
    assign P[61] = in1[8] ^ in2[8];
    assign G[62] = in1[7] & in2[7];
    assign P[62] = in1[7] ^ in2[7];
    assign G[63] = in1[6] & in2[6];
    assign P[63] = in1[6] ^ in2[6];
    assign G[64] = in1[5] & in2[5];
    assign P[64] = in1[5] ^ in2[5];
    assign G[65] = in1[4] & in2[4];
    assign P[65] = in1[4] ^ in2[4];
    assign G[66] = in1[3] & in2[3];
    assign P[66] = in1[3] ^ in2[3];
    assign G[67] = in1[2] & in2[2];
    assign P[67] = in1[2] ^ in2[2];
    assign G[68] = in1[1] & in2[1];
    assign P[68] = in1[1] ^ in2[1];
    assign G[69] = in1[0] & in2[0];
    assign P[69] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign cout = G[69] | (P[69] & C[69]);
    assign sum = P ^ C;
endmodule

module CLA_69(output [68:0] sum, output cout, input [68:0] in1, input [68:0] in2);

    wire[68:0] G;
    wire[68:0] C;
    wire[68:0] P;

    assign G[0] = in1[68] & in2[68];
    assign P[0] = in1[68] ^ in2[68];
    assign G[1] = in1[67] & in2[67];
    assign P[1] = in1[67] ^ in2[67];
    assign G[2] = in1[66] & in2[66];
    assign P[2] = in1[66] ^ in2[66];
    assign G[3] = in1[65] & in2[65];
    assign P[3] = in1[65] ^ in2[65];
    assign G[4] = in1[64] & in2[64];
    assign P[4] = in1[64] ^ in2[64];
    assign G[5] = in1[63] & in2[63];
    assign P[5] = in1[63] ^ in2[63];
    assign G[6] = in1[62] & in2[62];
    assign P[6] = in1[62] ^ in2[62];
    assign G[7] = in1[61] & in2[61];
    assign P[7] = in1[61] ^ in2[61];
    assign G[8] = in1[60] & in2[60];
    assign P[8] = in1[60] ^ in2[60];
    assign G[9] = in1[59] & in2[59];
    assign P[9] = in1[59] ^ in2[59];
    assign G[10] = in1[58] & in2[58];
    assign P[10] = in1[58] ^ in2[58];
    assign G[11] = in1[57] & in2[57];
    assign P[11] = in1[57] ^ in2[57];
    assign G[12] = in1[56] & in2[56];
    assign P[12] = in1[56] ^ in2[56];
    assign G[13] = in1[55] & in2[55];
    assign P[13] = in1[55] ^ in2[55];
    assign G[14] = in1[54] & in2[54];
    assign P[14] = in1[54] ^ in2[54];
    assign G[15] = in1[53] & in2[53];
    assign P[15] = in1[53] ^ in2[53];
    assign G[16] = in1[52] & in2[52];
    assign P[16] = in1[52] ^ in2[52];
    assign G[17] = in1[51] & in2[51];
    assign P[17] = in1[51] ^ in2[51];
    assign G[18] = in1[50] & in2[50];
    assign P[18] = in1[50] ^ in2[50];
    assign G[19] = in1[49] & in2[49];
    assign P[19] = in1[49] ^ in2[49];
    assign G[20] = in1[48] & in2[48];
    assign P[20] = in1[48] ^ in2[48];
    assign G[21] = in1[47] & in2[47];
    assign P[21] = in1[47] ^ in2[47];
    assign G[22] = in1[46] & in2[46];
    assign P[22] = in1[46] ^ in2[46];
    assign G[23] = in1[45] & in2[45];
    assign P[23] = in1[45] ^ in2[45];
    assign G[24] = in1[44] & in2[44];
    assign P[24] = in1[44] ^ in2[44];
    assign G[25] = in1[43] & in2[43];
    assign P[25] = in1[43] ^ in2[43];
    assign G[26] = in1[42] & in2[42];
    assign P[26] = in1[42] ^ in2[42];
    assign G[27] = in1[41] & in2[41];
    assign P[27] = in1[41] ^ in2[41];
    assign G[28] = in1[40] & in2[40];
    assign P[28] = in1[40] ^ in2[40];
    assign G[29] = in1[39] & in2[39];
    assign P[29] = in1[39] ^ in2[39];
    assign G[30] = in1[38] & in2[38];
    assign P[30] = in1[38] ^ in2[38];
    assign G[31] = in1[37] & in2[37];
    assign P[31] = in1[37] ^ in2[37];
    assign G[32] = in1[36] & in2[36];
    assign P[32] = in1[36] ^ in2[36];
    assign G[33] = in1[35] & in2[35];
    assign P[33] = in1[35] ^ in2[35];
    assign G[34] = in1[34] & in2[34];
    assign P[34] = in1[34] ^ in2[34];
    assign G[35] = in1[33] & in2[33];
    assign P[35] = in1[33] ^ in2[33];
    assign G[36] = in1[32] & in2[32];
    assign P[36] = in1[32] ^ in2[32];
    assign G[37] = in1[31] & in2[31];
    assign P[37] = in1[31] ^ in2[31];
    assign G[38] = in1[30] & in2[30];
    assign P[38] = in1[30] ^ in2[30];
    assign G[39] = in1[29] & in2[29];
    assign P[39] = in1[29] ^ in2[29];
    assign G[40] = in1[28] & in2[28];
    assign P[40] = in1[28] ^ in2[28];
    assign G[41] = in1[27] & in2[27];
    assign P[41] = in1[27] ^ in2[27];
    assign G[42] = in1[26] & in2[26];
    assign P[42] = in1[26] ^ in2[26];
    assign G[43] = in1[25] & in2[25];
    assign P[43] = in1[25] ^ in2[25];
    assign G[44] = in1[24] & in2[24];
    assign P[44] = in1[24] ^ in2[24];
    assign G[45] = in1[23] & in2[23];
    assign P[45] = in1[23] ^ in2[23];
    assign G[46] = in1[22] & in2[22];
    assign P[46] = in1[22] ^ in2[22];
    assign G[47] = in1[21] & in2[21];
    assign P[47] = in1[21] ^ in2[21];
    assign G[48] = in1[20] & in2[20];
    assign P[48] = in1[20] ^ in2[20];
    assign G[49] = in1[19] & in2[19];
    assign P[49] = in1[19] ^ in2[19];
    assign G[50] = in1[18] & in2[18];
    assign P[50] = in1[18] ^ in2[18];
    assign G[51] = in1[17] & in2[17];
    assign P[51] = in1[17] ^ in2[17];
    assign G[52] = in1[16] & in2[16];
    assign P[52] = in1[16] ^ in2[16];
    assign G[53] = in1[15] & in2[15];
    assign P[53] = in1[15] ^ in2[15];
    assign G[54] = in1[14] & in2[14];
    assign P[54] = in1[14] ^ in2[14];
    assign G[55] = in1[13] & in2[13];
    assign P[55] = in1[13] ^ in2[13];
    assign G[56] = in1[12] & in2[12];
    assign P[56] = in1[12] ^ in2[12];
    assign G[57] = in1[11] & in2[11];
    assign P[57] = in1[11] ^ in2[11];
    assign G[58] = in1[10] & in2[10];
    assign P[58] = in1[10] ^ in2[10];
    assign G[59] = in1[9] & in2[9];
    assign P[59] = in1[9] ^ in2[9];
    assign G[60] = in1[8] & in2[8];
    assign P[60] = in1[8] ^ in2[8];
    assign G[61] = in1[7] & in2[7];
    assign P[61] = in1[7] ^ in2[7];
    assign G[62] = in1[6] & in2[6];
    assign P[62] = in1[6] ^ in2[6];
    assign G[63] = in1[5] & in2[5];
    assign P[63] = in1[5] ^ in2[5];
    assign G[64] = in1[4] & in2[4];
    assign P[64] = in1[4] ^ in2[4];
    assign G[65] = in1[3] & in2[3];
    assign P[65] = in1[3] ^ in2[3];
    assign G[66] = in1[2] & in2[2];
    assign P[66] = in1[2] ^ in2[2];
    assign G[67] = in1[1] & in2[1];
    assign P[67] = in1[1] ^ in2[1];
    assign G[68] = in1[0] & in2[0];
    assign P[68] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign cout = G[68] | (P[68] & C[68]);
    assign sum = P ^ C;
endmodule

module CLA_68(output [67:0] sum, output cout, input [67:0] in1, input [67:0] in2);

    wire[67:0] G;
    wire[67:0] C;
    wire[67:0] P;

    assign G[0] = in1[67] & in2[67];
    assign P[0] = in1[67] ^ in2[67];
    assign G[1] = in1[66] & in2[66];
    assign P[1] = in1[66] ^ in2[66];
    assign G[2] = in1[65] & in2[65];
    assign P[2] = in1[65] ^ in2[65];
    assign G[3] = in1[64] & in2[64];
    assign P[3] = in1[64] ^ in2[64];
    assign G[4] = in1[63] & in2[63];
    assign P[4] = in1[63] ^ in2[63];
    assign G[5] = in1[62] & in2[62];
    assign P[5] = in1[62] ^ in2[62];
    assign G[6] = in1[61] & in2[61];
    assign P[6] = in1[61] ^ in2[61];
    assign G[7] = in1[60] & in2[60];
    assign P[7] = in1[60] ^ in2[60];
    assign G[8] = in1[59] & in2[59];
    assign P[8] = in1[59] ^ in2[59];
    assign G[9] = in1[58] & in2[58];
    assign P[9] = in1[58] ^ in2[58];
    assign G[10] = in1[57] & in2[57];
    assign P[10] = in1[57] ^ in2[57];
    assign G[11] = in1[56] & in2[56];
    assign P[11] = in1[56] ^ in2[56];
    assign G[12] = in1[55] & in2[55];
    assign P[12] = in1[55] ^ in2[55];
    assign G[13] = in1[54] & in2[54];
    assign P[13] = in1[54] ^ in2[54];
    assign G[14] = in1[53] & in2[53];
    assign P[14] = in1[53] ^ in2[53];
    assign G[15] = in1[52] & in2[52];
    assign P[15] = in1[52] ^ in2[52];
    assign G[16] = in1[51] & in2[51];
    assign P[16] = in1[51] ^ in2[51];
    assign G[17] = in1[50] & in2[50];
    assign P[17] = in1[50] ^ in2[50];
    assign G[18] = in1[49] & in2[49];
    assign P[18] = in1[49] ^ in2[49];
    assign G[19] = in1[48] & in2[48];
    assign P[19] = in1[48] ^ in2[48];
    assign G[20] = in1[47] & in2[47];
    assign P[20] = in1[47] ^ in2[47];
    assign G[21] = in1[46] & in2[46];
    assign P[21] = in1[46] ^ in2[46];
    assign G[22] = in1[45] & in2[45];
    assign P[22] = in1[45] ^ in2[45];
    assign G[23] = in1[44] & in2[44];
    assign P[23] = in1[44] ^ in2[44];
    assign G[24] = in1[43] & in2[43];
    assign P[24] = in1[43] ^ in2[43];
    assign G[25] = in1[42] & in2[42];
    assign P[25] = in1[42] ^ in2[42];
    assign G[26] = in1[41] & in2[41];
    assign P[26] = in1[41] ^ in2[41];
    assign G[27] = in1[40] & in2[40];
    assign P[27] = in1[40] ^ in2[40];
    assign G[28] = in1[39] & in2[39];
    assign P[28] = in1[39] ^ in2[39];
    assign G[29] = in1[38] & in2[38];
    assign P[29] = in1[38] ^ in2[38];
    assign G[30] = in1[37] & in2[37];
    assign P[30] = in1[37] ^ in2[37];
    assign G[31] = in1[36] & in2[36];
    assign P[31] = in1[36] ^ in2[36];
    assign G[32] = in1[35] & in2[35];
    assign P[32] = in1[35] ^ in2[35];
    assign G[33] = in1[34] & in2[34];
    assign P[33] = in1[34] ^ in2[34];
    assign G[34] = in1[33] & in2[33];
    assign P[34] = in1[33] ^ in2[33];
    assign G[35] = in1[32] & in2[32];
    assign P[35] = in1[32] ^ in2[32];
    assign G[36] = in1[31] & in2[31];
    assign P[36] = in1[31] ^ in2[31];
    assign G[37] = in1[30] & in2[30];
    assign P[37] = in1[30] ^ in2[30];
    assign G[38] = in1[29] & in2[29];
    assign P[38] = in1[29] ^ in2[29];
    assign G[39] = in1[28] & in2[28];
    assign P[39] = in1[28] ^ in2[28];
    assign G[40] = in1[27] & in2[27];
    assign P[40] = in1[27] ^ in2[27];
    assign G[41] = in1[26] & in2[26];
    assign P[41] = in1[26] ^ in2[26];
    assign G[42] = in1[25] & in2[25];
    assign P[42] = in1[25] ^ in2[25];
    assign G[43] = in1[24] & in2[24];
    assign P[43] = in1[24] ^ in2[24];
    assign G[44] = in1[23] & in2[23];
    assign P[44] = in1[23] ^ in2[23];
    assign G[45] = in1[22] & in2[22];
    assign P[45] = in1[22] ^ in2[22];
    assign G[46] = in1[21] & in2[21];
    assign P[46] = in1[21] ^ in2[21];
    assign G[47] = in1[20] & in2[20];
    assign P[47] = in1[20] ^ in2[20];
    assign G[48] = in1[19] & in2[19];
    assign P[48] = in1[19] ^ in2[19];
    assign G[49] = in1[18] & in2[18];
    assign P[49] = in1[18] ^ in2[18];
    assign G[50] = in1[17] & in2[17];
    assign P[50] = in1[17] ^ in2[17];
    assign G[51] = in1[16] & in2[16];
    assign P[51] = in1[16] ^ in2[16];
    assign G[52] = in1[15] & in2[15];
    assign P[52] = in1[15] ^ in2[15];
    assign G[53] = in1[14] & in2[14];
    assign P[53] = in1[14] ^ in2[14];
    assign G[54] = in1[13] & in2[13];
    assign P[54] = in1[13] ^ in2[13];
    assign G[55] = in1[12] & in2[12];
    assign P[55] = in1[12] ^ in2[12];
    assign G[56] = in1[11] & in2[11];
    assign P[56] = in1[11] ^ in2[11];
    assign G[57] = in1[10] & in2[10];
    assign P[57] = in1[10] ^ in2[10];
    assign G[58] = in1[9] & in2[9];
    assign P[58] = in1[9] ^ in2[9];
    assign G[59] = in1[8] & in2[8];
    assign P[59] = in1[8] ^ in2[8];
    assign G[60] = in1[7] & in2[7];
    assign P[60] = in1[7] ^ in2[7];
    assign G[61] = in1[6] & in2[6];
    assign P[61] = in1[6] ^ in2[6];
    assign G[62] = in1[5] & in2[5];
    assign P[62] = in1[5] ^ in2[5];
    assign G[63] = in1[4] & in2[4];
    assign P[63] = in1[4] ^ in2[4];
    assign G[64] = in1[3] & in2[3];
    assign P[64] = in1[3] ^ in2[3];
    assign G[65] = in1[2] & in2[2];
    assign P[65] = in1[2] ^ in2[2];
    assign G[66] = in1[1] & in2[1];
    assign P[66] = in1[1] ^ in2[1];
    assign G[67] = in1[0] & in2[0];
    assign P[67] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign cout = G[67] | (P[67] & C[67]);
    assign sum = P ^ C;
endmodule

module CLA_67(output [66:0] sum, output cout, input [66:0] in1, input [66:0] in2);

    wire[66:0] G;
    wire[66:0] C;
    wire[66:0] P;

    assign G[0] = in1[66] & in2[66];
    assign P[0] = in1[66] ^ in2[66];
    assign G[1] = in1[65] & in2[65];
    assign P[1] = in1[65] ^ in2[65];
    assign G[2] = in1[64] & in2[64];
    assign P[2] = in1[64] ^ in2[64];
    assign G[3] = in1[63] & in2[63];
    assign P[3] = in1[63] ^ in2[63];
    assign G[4] = in1[62] & in2[62];
    assign P[4] = in1[62] ^ in2[62];
    assign G[5] = in1[61] & in2[61];
    assign P[5] = in1[61] ^ in2[61];
    assign G[6] = in1[60] & in2[60];
    assign P[6] = in1[60] ^ in2[60];
    assign G[7] = in1[59] & in2[59];
    assign P[7] = in1[59] ^ in2[59];
    assign G[8] = in1[58] & in2[58];
    assign P[8] = in1[58] ^ in2[58];
    assign G[9] = in1[57] & in2[57];
    assign P[9] = in1[57] ^ in2[57];
    assign G[10] = in1[56] & in2[56];
    assign P[10] = in1[56] ^ in2[56];
    assign G[11] = in1[55] & in2[55];
    assign P[11] = in1[55] ^ in2[55];
    assign G[12] = in1[54] & in2[54];
    assign P[12] = in1[54] ^ in2[54];
    assign G[13] = in1[53] & in2[53];
    assign P[13] = in1[53] ^ in2[53];
    assign G[14] = in1[52] & in2[52];
    assign P[14] = in1[52] ^ in2[52];
    assign G[15] = in1[51] & in2[51];
    assign P[15] = in1[51] ^ in2[51];
    assign G[16] = in1[50] & in2[50];
    assign P[16] = in1[50] ^ in2[50];
    assign G[17] = in1[49] & in2[49];
    assign P[17] = in1[49] ^ in2[49];
    assign G[18] = in1[48] & in2[48];
    assign P[18] = in1[48] ^ in2[48];
    assign G[19] = in1[47] & in2[47];
    assign P[19] = in1[47] ^ in2[47];
    assign G[20] = in1[46] & in2[46];
    assign P[20] = in1[46] ^ in2[46];
    assign G[21] = in1[45] & in2[45];
    assign P[21] = in1[45] ^ in2[45];
    assign G[22] = in1[44] & in2[44];
    assign P[22] = in1[44] ^ in2[44];
    assign G[23] = in1[43] & in2[43];
    assign P[23] = in1[43] ^ in2[43];
    assign G[24] = in1[42] & in2[42];
    assign P[24] = in1[42] ^ in2[42];
    assign G[25] = in1[41] & in2[41];
    assign P[25] = in1[41] ^ in2[41];
    assign G[26] = in1[40] & in2[40];
    assign P[26] = in1[40] ^ in2[40];
    assign G[27] = in1[39] & in2[39];
    assign P[27] = in1[39] ^ in2[39];
    assign G[28] = in1[38] & in2[38];
    assign P[28] = in1[38] ^ in2[38];
    assign G[29] = in1[37] & in2[37];
    assign P[29] = in1[37] ^ in2[37];
    assign G[30] = in1[36] & in2[36];
    assign P[30] = in1[36] ^ in2[36];
    assign G[31] = in1[35] & in2[35];
    assign P[31] = in1[35] ^ in2[35];
    assign G[32] = in1[34] & in2[34];
    assign P[32] = in1[34] ^ in2[34];
    assign G[33] = in1[33] & in2[33];
    assign P[33] = in1[33] ^ in2[33];
    assign G[34] = in1[32] & in2[32];
    assign P[34] = in1[32] ^ in2[32];
    assign G[35] = in1[31] & in2[31];
    assign P[35] = in1[31] ^ in2[31];
    assign G[36] = in1[30] & in2[30];
    assign P[36] = in1[30] ^ in2[30];
    assign G[37] = in1[29] & in2[29];
    assign P[37] = in1[29] ^ in2[29];
    assign G[38] = in1[28] & in2[28];
    assign P[38] = in1[28] ^ in2[28];
    assign G[39] = in1[27] & in2[27];
    assign P[39] = in1[27] ^ in2[27];
    assign G[40] = in1[26] & in2[26];
    assign P[40] = in1[26] ^ in2[26];
    assign G[41] = in1[25] & in2[25];
    assign P[41] = in1[25] ^ in2[25];
    assign G[42] = in1[24] & in2[24];
    assign P[42] = in1[24] ^ in2[24];
    assign G[43] = in1[23] & in2[23];
    assign P[43] = in1[23] ^ in2[23];
    assign G[44] = in1[22] & in2[22];
    assign P[44] = in1[22] ^ in2[22];
    assign G[45] = in1[21] & in2[21];
    assign P[45] = in1[21] ^ in2[21];
    assign G[46] = in1[20] & in2[20];
    assign P[46] = in1[20] ^ in2[20];
    assign G[47] = in1[19] & in2[19];
    assign P[47] = in1[19] ^ in2[19];
    assign G[48] = in1[18] & in2[18];
    assign P[48] = in1[18] ^ in2[18];
    assign G[49] = in1[17] & in2[17];
    assign P[49] = in1[17] ^ in2[17];
    assign G[50] = in1[16] & in2[16];
    assign P[50] = in1[16] ^ in2[16];
    assign G[51] = in1[15] & in2[15];
    assign P[51] = in1[15] ^ in2[15];
    assign G[52] = in1[14] & in2[14];
    assign P[52] = in1[14] ^ in2[14];
    assign G[53] = in1[13] & in2[13];
    assign P[53] = in1[13] ^ in2[13];
    assign G[54] = in1[12] & in2[12];
    assign P[54] = in1[12] ^ in2[12];
    assign G[55] = in1[11] & in2[11];
    assign P[55] = in1[11] ^ in2[11];
    assign G[56] = in1[10] & in2[10];
    assign P[56] = in1[10] ^ in2[10];
    assign G[57] = in1[9] & in2[9];
    assign P[57] = in1[9] ^ in2[9];
    assign G[58] = in1[8] & in2[8];
    assign P[58] = in1[8] ^ in2[8];
    assign G[59] = in1[7] & in2[7];
    assign P[59] = in1[7] ^ in2[7];
    assign G[60] = in1[6] & in2[6];
    assign P[60] = in1[6] ^ in2[6];
    assign G[61] = in1[5] & in2[5];
    assign P[61] = in1[5] ^ in2[5];
    assign G[62] = in1[4] & in2[4];
    assign P[62] = in1[4] ^ in2[4];
    assign G[63] = in1[3] & in2[3];
    assign P[63] = in1[3] ^ in2[3];
    assign G[64] = in1[2] & in2[2];
    assign P[64] = in1[2] ^ in2[2];
    assign G[65] = in1[1] & in2[1];
    assign P[65] = in1[1] ^ in2[1];
    assign G[66] = in1[0] & in2[0];
    assign P[66] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign cout = G[66] | (P[66] & C[66]);
    assign sum = P ^ C;
endmodule

module CLA_66(output [65:0] sum, output cout, input [65:0] in1, input [65:0] in2);

    wire[65:0] G;
    wire[65:0] C;
    wire[65:0] P;

    assign G[0] = in1[65] & in2[65];
    assign P[0] = in1[65] ^ in2[65];
    assign G[1] = in1[64] & in2[64];
    assign P[1] = in1[64] ^ in2[64];
    assign G[2] = in1[63] & in2[63];
    assign P[2] = in1[63] ^ in2[63];
    assign G[3] = in1[62] & in2[62];
    assign P[3] = in1[62] ^ in2[62];
    assign G[4] = in1[61] & in2[61];
    assign P[4] = in1[61] ^ in2[61];
    assign G[5] = in1[60] & in2[60];
    assign P[5] = in1[60] ^ in2[60];
    assign G[6] = in1[59] & in2[59];
    assign P[6] = in1[59] ^ in2[59];
    assign G[7] = in1[58] & in2[58];
    assign P[7] = in1[58] ^ in2[58];
    assign G[8] = in1[57] & in2[57];
    assign P[8] = in1[57] ^ in2[57];
    assign G[9] = in1[56] & in2[56];
    assign P[9] = in1[56] ^ in2[56];
    assign G[10] = in1[55] & in2[55];
    assign P[10] = in1[55] ^ in2[55];
    assign G[11] = in1[54] & in2[54];
    assign P[11] = in1[54] ^ in2[54];
    assign G[12] = in1[53] & in2[53];
    assign P[12] = in1[53] ^ in2[53];
    assign G[13] = in1[52] & in2[52];
    assign P[13] = in1[52] ^ in2[52];
    assign G[14] = in1[51] & in2[51];
    assign P[14] = in1[51] ^ in2[51];
    assign G[15] = in1[50] & in2[50];
    assign P[15] = in1[50] ^ in2[50];
    assign G[16] = in1[49] & in2[49];
    assign P[16] = in1[49] ^ in2[49];
    assign G[17] = in1[48] & in2[48];
    assign P[17] = in1[48] ^ in2[48];
    assign G[18] = in1[47] & in2[47];
    assign P[18] = in1[47] ^ in2[47];
    assign G[19] = in1[46] & in2[46];
    assign P[19] = in1[46] ^ in2[46];
    assign G[20] = in1[45] & in2[45];
    assign P[20] = in1[45] ^ in2[45];
    assign G[21] = in1[44] & in2[44];
    assign P[21] = in1[44] ^ in2[44];
    assign G[22] = in1[43] & in2[43];
    assign P[22] = in1[43] ^ in2[43];
    assign G[23] = in1[42] & in2[42];
    assign P[23] = in1[42] ^ in2[42];
    assign G[24] = in1[41] & in2[41];
    assign P[24] = in1[41] ^ in2[41];
    assign G[25] = in1[40] & in2[40];
    assign P[25] = in1[40] ^ in2[40];
    assign G[26] = in1[39] & in2[39];
    assign P[26] = in1[39] ^ in2[39];
    assign G[27] = in1[38] & in2[38];
    assign P[27] = in1[38] ^ in2[38];
    assign G[28] = in1[37] & in2[37];
    assign P[28] = in1[37] ^ in2[37];
    assign G[29] = in1[36] & in2[36];
    assign P[29] = in1[36] ^ in2[36];
    assign G[30] = in1[35] & in2[35];
    assign P[30] = in1[35] ^ in2[35];
    assign G[31] = in1[34] & in2[34];
    assign P[31] = in1[34] ^ in2[34];
    assign G[32] = in1[33] & in2[33];
    assign P[32] = in1[33] ^ in2[33];
    assign G[33] = in1[32] & in2[32];
    assign P[33] = in1[32] ^ in2[32];
    assign G[34] = in1[31] & in2[31];
    assign P[34] = in1[31] ^ in2[31];
    assign G[35] = in1[30] & in2[30];
    assign P[35] = in1[30] ^ in2[30];
    assign G[36] = in1[29] & in2[29];
    assign P[36] = in1[29] ^ in2[29];
    assign G[37] = in1[28] & in2[28];
    assign P[37] = in1[28] ^ in2[28];
    assign G[38] = in1[27] & in2[27];
    assign P[38] = in1[27] ^ in2[27];
    assign G[39] = in1[26] & in2[26];
    assign P[39] = in1[26] ^ in2[26];
    assign G[40] = in1[25] & in2[25];
    assign P[40] = in1[25] ^ in2[25];
    assign G[41] = in1[24] & in2[24];
    assign P[41] = in1[24] ^ in2[24];
    assign G[42] = in1[23] & in2[23];
    assign P[42] = in1[23] ^ in2[23];
    assign G[43] = in1[22] & in2[22];
    assign P[43] = in1[22] ^ in2[22];
    assign G[44] = in1[21] & in2[21];
    assign P[44] = in1[21] ^ in2[21];
    assign G[45] = in1[20] & in2[20];
    assign P[45] = in1[20] ^ in2[20];
    assign G[46] = in1[19] & in2[19];
    assign P[46] = in1[19] ^ in2[19];
    assign G[47] = in1[18] & in2[18];
    assign P[47] = in1[18] ^ in2[18];
    assign G[48] = in1[17] & in2[17];
    assign P[48] = in1[17] ^ in2[17];
    assign G[49] = in1[16] & in2[16];
    assign P[49] = in1[16] ^ in2[16];
    assign G[50] = in1[15] & in2[15];
    assign P[50] = in1[15] ^ in2[15];
    assign G[51] = in1[14] & in2[14];
    assign P[51] = in1[14] ^ in2[14];
    assign G[52] = in1[13] & in2[13];
    assign P[52] = in1[13] ^ in2[13];
    assign G[53] = in1[12] & in2[12];
    assign P[53] = in1[12] ^ in2[12];
    assign G[54] = in1[11] & in2[11];
    assign P[54] = in1[11] ^ in2[11];
    assign G[55] = in1[10] & in2[10];
    assign P[55] = in1[10] ^ in2[10];
    assign G[56] = in1[9] & in2[9];
    assign P[56] = in1[9] ^ in2[9];
    assign G[57] = in1[8] & in2[8];
    assign P[57] = in1[8] ^ in2[8];
    assign G[58] = in1[7] & in2[7];
    assign P[58] = in1[7] ^ in2[7];
    assign G[59] = in1[6] & in2[6];
    assign P[59] = in1[6] ^ in2[6];
    assign G[60] = in1[5] & in2[5];
    assign P[60] = in1[5] ^ in2[5];
    assign G[61] = in1[4] & in2[4];
    assign P[61] = in1[4] ^ in2[4];
    assign G[62] = in1[3] & in2[3];
    assign P[62] = in1[3] ^ in2[3];
    assign G[63] = in1[2] & in2[2];
    assign P[63] = in1[2] ^ in2[2];
    assign G[64] = in1[1] & in2[1];
    assign P[64] = in1[1] ^ in2[1];
    assign G[65] = in1[0] & in2[0];
    assign P[65] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign cout = G[65] | (P[65] & C[65]);
    assign sum = P ^ C;
endmodule

module CLA_65(output [64:0] sum, output cout, input [64:0] in1, input [64:0] in2);

    wire[64:0] G;
    wire[64:0] C;
    wire[64:0] P;

    assign G[0] = in1[64] & in2[64];
    assign P[0] = in1[64] ^ in2[64];
    assign G[1] = in1[63] & in2[63];
    assign P[1] = in1[63] ^ in2[63];
    assign G[2] = in1[62] & in2[62];
    assign P[2] = in1[62] ^ in2[62];
    assign G[3] = in1[61] & in2[61];
    assign P[3] = in1[61] ^ in2[61];
    assign G[4] = in1[60] & in2[60];
    assign P[4] = in1[60] ^ in2[60];
    assign G[5] = in1[59] & in2[59];
    assign P[5] = in1[59] ^ in2[59];
    assign G[6] = in1[58] & in2[58];
    assign P[6] = in1[58] ^ in2[58];
    assign G[7] = in1[57] & in2[57];
    assign P[7] = in1[57] ^ in2[57];
    assign G[8] = in1[56] & in2[56];
    assign P[8] = in1[56] ^ in2[56];
    assign G[9] = in1[55] & in2[55];
    assign P[9] = in1[55] ^ in2[55];
    assign G[10] = in1[54] & in2[54];
    assign P[10] = in1[54] ^ in2[54];
    assign G[11] = in1[53] & in2[53];
    assign P[11] = in1[53] ^ in2[53];
    assign G[12] = in1[52] & in2[52];
    assign P[12] = in1[52] ^ in2[52];
    assign G[13] = in1[51] & in2[51];
    assign P[13] = in1[51] ^ in2[51];
    assign G[14] = in1[50] & in2[50];
    assign P[14] = in1[50] ^ in2[50];
    assign G[15] = in1[49] & in2[49];
    assign P[15] = in1[49] ^ in2[49];
    assign G[16] = in1[48] & in2[48];
    assign P[16] = in1[48] ^ in2[48];
    assign G[17] = in1[47] & in2[47];
    assign P[17] = in1[47] ^ in2[47];
    assign G[18] = in1[46] & in2[46];
    assign P[18] = in1[46] ^ in2[46];
    assign G[19] = in1[45] & in2[45];
    assign P[19] = in1[45] ^ in2[45];
    assign G[20] = in1[44] & in2[44];
    assign P[20] = in1[44] ^ in2[44];
    assign G[21] = in1[43] & in2[43];
    assign P[21] = in1[43] ^ in2[43];
    assign G[22] = in1[42] & in2[42];
    assign P[22] = in1[42] ^ in2[42];
    assign G[23] = in1[41] & in2[41];
    assign P[23] = in1[41] ^ in2[41];
    assign G[24] = in1[40] & in2[40];
    assign P[24] = in1[40] ^ in2[40];
    assign G[25] = in1[39] & in2[39];
    assign P[25] = in1[39] ^ in2[39];
    assign G[26] = in1[38] & in2[38];
    assign P[26] = in1[38] ^ in2[38];
    assign G[27] = in1[37] & in2[37];
    assign P[27] = in1[37] ^ in2[37];
    assign G[28] = in1[36] & in2[36];
    assign P[28] = in1[36] ^ in2[36];
    assign G[29] = in1[35] & in2[35];
    assign P[29] = in1[35] ^ in2[35];
    assign G[30] = in1[34] & in2[34];
    assign P[30] = in1[34] ^ in2[34];
    assign G[31] = in1[33] & in2[33];
    assign P[31] = in1[33] ^ in2[33];
    assign G[32] = in1[32] & in2[32];
    assign P[32] = in1[32] ^ in2[32];
    assign G[33] = in1[31] & in2[31];
    assign P[33] = in1[31] ^ in2[31];
    assign G[34] = in1[30] & in2[30];
    assign P[34] = in1[30] ^ in2[30];
    assign G[35] = in1[29] & in2[29];
    assign P[35] = in1[29] ^ in2[29];
    assign G[36] = in1[28] & in2[28];
    assign P[36] = in1[28] ^ in2[28];
    assign G[37] = in1[27] & in2[27];
    assign P[37] = in1[27] ^ in2[27];
    assign G[38] = in1[26] & in2[26];
    assign P[38] = in1[26] ^ in2[26];
    assign G[39] = in1[25] & in2[25];
    assign P[39] = in1[25] ^ in2[25];
    assign G[40] = in1[24] & in2[24];
    assign P[40] = in1[24] ^ in2[24];
    assign G[41] = in1[23] & in2[23];
    assign P[41] = in1[23] ^ in2[23];
    assign G[42] = in1[22] & in2[22];
    assign P[42] = in1[22] ^ in2[22];
    assign G[43] = in1[21] & in2[21];
    assign P[43] = in1[21] ^ in2[21];
    assign G[44] = in1[20] & in2[20];
    assign P[44] = in1[20] ^ in2[20];
    assign G[45] = in1[19] & in2[19];
    assign P[45] = in1[19] ^ in2[19];
    assign G[46] = in1[18] & in2[18];
    assign P[46] = in1[18] ^ in2[18];
    assign G[47] = in1[17] & in2[17];
    assign P[47] = in1[17] ^ in2[17];
    assign G[48] = in1[16] & in2[16];
    assign P[48] = in1[16] ^ in2[16];
    assign G[49] = in1[15] & in2[15];
    assign P[49] = in1[15] ^ in2[15];
    assign G[50] = in1[14] & in2[14];
    assign P[50] = in1[14] ^ in2[14];
    assign G[51] = in1[13] & in2[13];
    assign P[51] = in1[13] ^ in2[13];
    assign G[52] = in1[12] & in2[12];
    assign P[52] = in1[12] ^ in2[12];
    assign G[53] = in1[11] & in2[11];
    assign P[53] = in1[11] ^ in2[11];
    assign G[54] = in1[10] & in2[10];
    assign P[54] = in1[10] ^ in2[10];
    assign G[55] = in1[9] & in2[9];
    assign P[55] = in1[9] ^ in2[9];
    assign G[56] = in1[8] & in2[8];
    assign P[56] = in1[8] ^ in2[8];
    assign G[57] = in1[7] & in2[7];
    assign P[57] = in1[7] ^ in2[7];
    assign G[58] = in1[6] & in2[6];
    assign P[58] = in1[6] ^ in2[6];
    assign G[59] = in1[5] & in2[5];
    assign P[59] = in1[5] ^ in2[5];
    assign G[60] = in1[4] & in2[4];
    assign P[60] = in1[4] ^ in2[4];
    assign G[61] = in1[3] & in2[3];
    assign P[61] = in1[3] ^ in2[3];
    assign G[62] = in1[2] & in2[2];
    assign P[62] = in1[2] ^ in2[2];
    assign G[63] = in1[1] & in2[1];
    assign P[63] = in1[1] ^ in2[1];
    assign G[64] = in1[0] & in2[0];
    assign P[64] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign cout = G[64] | (P[64] & C[64]);
    assign sum = P ^ C;
endmodule

module CLA_64(output [63:0] sum, output cout, input [63:0] in1, input [63:0] in2);

    wire[63:0] G;
    wire[63:0] C;
    wire[63:0] P;

    assign G[0] = in1[63] & in2[63];
    assign P[0] = in1[63] ^ in2[63];
    assign G[1] = in1[62] & in2[62];
    assign P[1] = in1[62] ^ in2[62];
    assign G[2] = in1[61] & in2[61];
    assign P[2] = in1[61] ^ in2[61];
    assign G[3] = in1[60] & in2[60];
    assign P[3] = in1[60] ^ in2[60];
    assign G[4] = in1[59] & in2[59];
    assign P[4] = in1[59] ^ in2[59];
    assign G[5] = in1[58] & in2[58];
    assign P[5] = in1[58] ^ in2[58];
    assign G[6] = in1[57] & in2[57];
    assign P[6] = in1[57] ^ in2[57];
    assign G[7] = in1[56] & in2[56];
    assign P[7] = in1[56] ^ in2[56];
    assign G[8] = in1[55] & in2[55];
    assign P[8] = in1[55] ^ in2[55];
    assign G[9] = in1[54] & in2[54];
    assign P[9] = in1[54] ^ in2[54];
    assign G[10] = in1[53] & in2[53];
    assign P[10] = in1[53] ^ in2[53];
    assign G[11] = in1[52] & in2[52];
    assign P[11] = in1[52] ^ in2[52];
    assign G[12] = in1[51] & in2[51];
    assign P[12] = in1[51] ^ in2[51];
    assign G[13] = in1[50] & in2[50];
    assign P[13] = in1[50] ^ in2[50];
    assign G[14] = in1[49] & in2[49];
    assign P[14] = in1[49] ^ in2[49];
    assign G[15] = in1[48] & in2[48];
    assign P[15] = in1[48] ^ in2[48];
    assign G[16] = in1[47] & in2[47];
    assign P[16] = in1[47] ^ in2[47];
    assign G[17] = in1[46] & in2[46];
    assign P[17] = in1[46] ^ in2[46];
    assign G[18] = in1[45] & in2[45];
    assign P[18] = in1[45] ^ in2[45];
    assign G[19] = in1[44] & in2[44];
    assign P[19] = in1[44] ^ in2[44];
    assign G[20] = in1[43] & in2[43];
    assign P[20] = in1[43] ^ in2[43];
    assign G[21] = in1[42] & in2[42];
    assign P[21] = in1[42] ^ in2[42];
    assign G[22] = in1[41] & in2[41];
    assign P[22] = in1[41] ^ in2[41];
    assign G[23] = in1[40] & in2[40];
    assign P[23] = in1[40] ^ in2[40];
    assign G[24] = in1[39] & in2[39];
    assign P[24] = in1[39] ^ in2[39];
    assign G[25] = in1[38] & in2[38];
    assign P[25] = in1[38] ^ in2[38];
    assign G[26] = in1[37] & in2[37];
    assign P[26] = in1[37] ^ in2[37];
    assign G[27] = in1[36] & in2[36];
    assign P[27] = in1[36] ^ in2[36];
    assign G[28] = in1[35] & in2[35];
    assign P[28] = in1[35] ^ in2[35];
    assign G[29] = in1[34] & in2[34];
    assign P[29] = in1[34] ^ in2[34];
    assign G[30] = in1[33] & in2[33];
    assign P[30] = in1[33] ^ in2[33];
    assign G[31] = in1[32] & in2[32];
    assign P[31] = in1[32] ^ in2[32];
    assign G[32] = in1[31] & in2[31];
    assign P[32] = in1[31] ^ in2[31];
    assign G[33] = in1[30] & in2[30];
    assign P[33] = in1[30] ^ in2[30];
    assign G[34] = in1[29] & in2[29];
    assign P[34] = in1[29] ^ in2[29];
    assign G[35] = in1[28] & in2[28];
    assign P[35] = in1[28] ^ in2[28];
    assign G[36] = in1[27] & in2[27];
    assign P[36] = in1[27] ^ in2[27];
    assign G[37] = in1[26] & in2[26];
    assign P[37] = in1[26] ^ in2[26];
    assign G[38] = in1[25] & in2[25];
    assign P[38] = in1[25] ^ in2[25];
    assign G[39] = in1[24] & in2[24];
    assign P[39] = in1[24] ^ in2[24];
    assign G[40] = in1[23] & in2[23];
    assign P[40] = in1[23] ^ in2[23];
    assign G[41] = in1[22] & in2[22];
    assign P[41] = in1[22] ^ in2[22];
    assign G[42] = in1[21] & in2[21];
    assign P[42] = in1[21] ^ in2[21];
    assign G[43] = in1[20] & in2[20];
    assign P[43] = in1[20] ^ in2[20];
    assign G[44] = in1[19] & in2[19];
    assign P[44] = in1[19] ^ in2[19];
    assign G[45] = in1[18] & in2[18];
    assign P[45] = in1[18] ^ in2[18];
    assign G[46] = in1[17] & in2[17];
    assign P[46] = in1[17] ^ in2[17];
    assign G[47] = in1[16] & in2[16];
    assign P[47] = in1[16] ^ in2[16];
    assign G[48] = in1[15] & in2[15];
    assign P[48] = in1[15] ^ in2[15];
    assign G[49] = in1[14] & in2[14];
    assign P[49] = in1[14] ^ in2[14];
    assign G[50] = in1[13] & in2[13];
    assign P[50] = in1[13] ^ in2[13];
    assign G[51] = in1[12] & in2[12];
    assign P[51] = in1[12] ^ in2[12];
    assign G[52] = in1[11] & in2[11];
    assign P[52] = in1[11] ^ in2[11];
    assign G[53] = in1[10] & in2[10];
    assign P[53] = in1[10] ^ in2[10];
    assign G[54] = in1[9] & in2[9];
    assign P[54] = in1[9] ^ in2[9];
    assign G[55] = in1[8] & in2[8];
    assign P[55] = in1[8] ^ in2[8];
    assign G[56] = in1[7] & in2[7];
    assign P[56] = in1[7] ^ in2[7];
    assign G[57] = in1[6] & in2[6];
    assign P[57] = in1[6] ^ in2[6];
    assign G[58] = in1[5] & in2[5];
    assign P[58] = in1[5] ^ in2[5];
    assign G[59] = in1[4] & in2[4];
    assign P[59] = in1[4] ^ in2[4];
    assign G[60] = in1[3] & in2[3];
    assign P[60] = in1[3] ^ in2[3];
    assign G[61] = in1[2] & in2[2];
    assign P[61] = in1[2] ^ in2[2];
    assign G[62] = in1[1] & in2[1];
    assign P[62] = in1[1] ^ in2[1];
    assign G[63] = in1[0] & in2[0];
    assign P[63] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign cout = G[63] | (P[63] & C[63]);
    assign sum = P ^ C;
endmodule

module CLA_63(output [62:0] sum, output cout, input [62:0] in1, input [62:0] in2);

    wire[62:0] G;
    wire[62:0] C;
    wire[62:0] P;

    assign G[0] = in1[62] & in2[62];
    assign P[0] = in1[62] ^ in2[62];
    assign G[1] = in1[61] & in2[61];
    assign P[1] = in1[61] ^ in2[61];
    assign G[2] = in1[60] & in2[60];
    assign P[2] = in1[60] ^ in2[60];
    assign G[3] = in1[59] & in2[59];
    assign P[3] = in1[59] ^ in2[59];
    assign G[4] = in1[58] & in2[58];
    assign P[4] = in1[58] ^ in2[58];
    assign G[5] = in1[57] & in2[57];
    assign P[5] = in1[57] ^ in2[57];
    assign G[6] = in1[56] & in2[56];
    assign P[6] = in1[56] ^ in2[56];
    assign G[7] = in1[55] & in2[55];
    assign P[7] = in1[55] ^ in2[55];
    assign G[8] = in1[54] & in2[54];
    assign P[8] = in1[54] ^ in2[54];
    assign G[9] = in1[53] & in2[53];
    assign P[9] = in1[53] ^ in2[53];
    assign G[10] = in1[52] & in2[52];
    assign P[10] = in1[52] ^ in2[52];
    assign G[11] = in1[51] & in2[51];
    assign P[11] = in1[51] ^ in2[51];
    assign G[12] = in1[50] & in2[50];
    assign P[12] = in1[50] ^ in2[50];
    assign G[13] = in1[49] & in2[49];
    assign P[13] = in1[49] ^ in2[49];
    assign G[14] = in1[48] & in2[48];
    assign P[14] = in1[48] ^ in2[48];
    assign G[15] = in1[47] & in2[47];
    assign P[15] = in1[47] ^ in2[47];
    assign G[16] = in1[46] & in2[46];
    assign P[16] = in1[46] ^ in2[46];
    assign G[17] = in1[45] & in2[45];
    assign P[17] = in1[45] ^ in2[45];
    assign G[18] = in1[44] & in2[44];
    assign P[18] = in1[44] ^ in2[44];
    assign G[19] = in1[43] & in2[43];
    assign P[19] = in1[43] ^ in2[43];
    assign G[20] = in1[42] & in2[42];
    assign P[20] = in1[42] ^ in2[42];
    assign G[21] = in1[41] & in2[41];
    assign P[21] = in1[41] ^ in2[41];
    assign G[22] = in1[40] & in2[40];
    assign P[22] = in1[40] ^ in2[40];
    assign G[23] = in1[39] & in2[39];
    assign P[23] = in1[39] ^ in2[39];
    assign G[24] = in1[38] & in2[38];
    assign P[24] = in1[38] ^ in2[38];
    assign G[25] = in1[37] & in2[37];
    assign P[25] = in1[37] ^ in2[37];
    assign G[26] = in1[36] & in2[36];
    assign P[26] = in1[36] ^ in2[36];
    assign G[27] = in1[35] & in2[35];
    assign P[27] = in1[35] ^ in2[35];
    assign G[28] = in1[34] & in2[34];
    assign P[28] = in1[34] ^ in2[34];
    assign G[29] = in1[33] & in2[33];
    assign P[29] = in1[33] ^ in2[33];
    assign G[30] = in1[32] & in2[32];
    assign P[30] = in1[32] ^ in2[32];
    assign G[31] = in1[31] & in2[31];
    assign P[31] = in1[31] ^ in2[31];
    assign G[32] = in1[30] & in2[30];
    assign P[32] = in1[30] ^ in2[30];
    assign G[33] = in1[29] & in2[29];
    assign P[33] = in1[29] ^ in2[29];
    assign G[34] = in1[28] & in2[28];
    assign P[34] = in1[28] ^ in2[28];
    assign G[35] = in1[27] & in2[27];
    assign P[35] = in1[27] ^ in2[27];
    assign G[36] = in1[26] & in2[26];
    assign P[36] = in1[26] ^ in2[26];
    assign G[37] = in1[25] & in2[25];
    assign P[37] = in1[25] ^ in2[25];
    assign G[38] = in1[24] & in2[24];
    assign P[38] = in1[24] ^ in2[24];
    assign G[39] = in1[23] & in2[23];
    assign P[39] = in1[23] ^ in2[23];
    assign G[40] = in1[22] & in2[22];
    assign P[40] = in1[22] ^ in2[22];
    assign G[41] = in1[21] & in2[21];
    assign P[41] = in1[21] ^ in2[21];
    assign G[42] = in1[20] & in2[20];
    assign P[42] = in1[20] ^ in2[20];
    assign G[43] = in1[19] & in2[19];
    assign P[43] = in1[19] ^ in2[19];
    assign G[44] = in1[18] & in2[18];
    assign P[44] = in1[18] ^ in2[18];
    assign G[45] = in1[17] & in2[17];
    assign P[45] = in1[17] ^ in2[17];
    assign G[46] = in1[16] & in2[16];
    assign P[46] = in1[16] ^ in2[16];
    assign G[47] = in1[15] & in2[15];
    assign P[47] = in1[15] ^ in2[15];
    assign G[48] = in1[14] & in2[14];
    assign P[48] = in1[14] ^ in2[14];
    assign G[49] = in1[13] & in2[13];
    assign P[49] = in1[13] ^ in2[13];
    assign G[50] = in1[12] & in2[12];
    assign P[50] = in1[12] ^ in2[12];
    assign G[51] = in1[11] & in2[11];
    assign P[51] = in1[11] ^ in2[11];
    assign G[52] = in1[10] & in2[10];
    assign P[52] = in1[10] ^ in2[10];
    assign G[53] = in1[9] & in2[9];
    assign P[53] = in1[9] ^ in2[9];
    assign G[54] = in1[8] & in2[8];
    assign P[54] = in1[8] ^ in2[8];
    assign G[55] = in1[7] & in2[7];
    assign P[55] = in1[7] ^ in2[7];
    assign G[56] = in1[6] & in2[6];
    assign P[56] = in1[6] ^ in2[6];
    assign G[57] = in1[5] & in2[5];
    assign P[57] = in1[5] ^ in2[5];
    assign G[58] = in1[4] & in2[4];
    assign P[58] = in1[4] ^ in2[4];
    assign G[59] = in1[3] & in2[3];
    assign P[59] = in1[3] ^ in2[3];
    assign G[60] = in1[2] & in2[2];
    assign P[60] = in1[2] ^ in2[2];
    assign G[61] = in1[1] & in2[1];
    assign P[61] = in1[1] ^ in2[1];
    assign G[62] = in1[0] & in2[0];
    assign P[62] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign cout = G[62] | (P[62] & C[62]);
    assign sum = P ^ C;
endmodule

module CLA_62(output [61:0] sum, output cout, input [61:0] in1, input [61:0] in2);

    wire[61:0] G;
    wire[61:0] C;
    wire[61:0] P;

    assign G[0] = in1[61] & in2[61];
    assign P[0] = in1[61] ^ in2[61];
    assign G[1] = in1[60] & in2[60];
    assign P[1] = in1[60] ^ in2[60];
    assign G[2] = in1[59] & in2[59];
    assign P[2] = in1[59] ^ in2[59];
    assign G[3] = in1[58] & in2[58];
    assign P[3] = in1[58] ^ in2[58];
    assign G[4] = in1[57] & in2[57];
    assign P[4] = in1[57] ^ in2[57];
    assign G[5] = in1[56] & in2[56];
    assign P[5] = in1[56] ^ in2[56];
    assign G[6] = in1[55] & in2[55];
    assign P[6] = in1[55] ^ in2[55];
    assign G[7] = in1[54] & in2[54];
    assign P[7] = in1[54] ^ in2[54];
    assign G[8] = in1[53] & in2[53];
    assign P[8] = in1[53] ^ in2[53];
    assign G[9] = in1[52] & in2[52];
    assign P[9] = in1[52] ^ in2[52];
    assign G[10] = in1[51] & in2[51];
    assign P[10] = in1[51] ^ in2[51];
    assign G[11] = in1[50] & in2[50];
    assign P[11] = in1[50] ^ in2[50];
    assign G[12] = in1[49] & in2[49];
    assign P[12] = in1[49] ^ in2[49];
    assign G[13] = in1[48] & in2[48];
    assign P[13] = in1[48] ^ in2[48];
    assign G[14] = in1[47] & in2[47];
    assign P[14] = in1[47] ^ in2[47];
    assign G[15] = in1[46] & in2[46];
    assign P[15] = in1[46] ^ in2[46];
    assign G[16] = in1[45] & in2[45];
    assign P[16] = in1[45] ^ in2[45];
    assign G[17] = in1[44] & in2[44];
    assign P[17] = in1[44] ^ in2[44];
    assign G[18] = in1[43] & in2[43];
    assign P[18] = in1[43] ^ in2[43];
    assign G[19] = in1[42] & in2[42];
    assign P[19] = in1[42] ^ in2[42];
    assign G[20] = in1[41] & in2[41];
    assign P[20] = in1[41] ^ in2[41];
    assign G[21] = in1[40] & in2[40];
    assign P[21] = in1[40] ^ in2[40];
    assign G[22] = in1[39] & in2[39];
    assign P[22] = in1[39] ^ in2[39];
    assign G[23] = in1[38] & in2[38];
    assign P[23] = in1[38] ^ in2[38];
    assign G[24] = in1[37] & in2[37];
    assign P[24] = in1[37] ^ in2[37];
    assign G[25] = in1[36] & in2[36];
    assign P[25] = in1[36] ^ in2[36];
    assign G[26] = in1[35] & in2[35];
    assign P[26] = in1[35] ^ in2[35];
    assign G[27] = in1[34] & in2[34];
    assign P[27] = in1[34] ^ in2[34];
    assign G[28] = in1[33] & in2[33];
    assign P[28] = in1[33] ^ in2[33];
    assign G[29] = in1[32] & in2[32];
    assign P[29] = in1[32] ^ in2[32];
    assign G[30] = in1[31] & in2[31];
    assign P[30] = in1[31] ^ in2[31];
    assign G[31] = in1[30] & in2[30];
    assign P[31] = in1[30] ^ in2[30];
    assign G[32] = in1[29] & in2[29];
    assign P[32] = in1[29] ^ in2[29];
    assign G[33] = in1[28] & in2[28];
    assign P[33] = in1[28] ^ in2[28];
    assign G[34] = in1[27] & in2[27];
    assign P[34] = in1[27] ^ in2[27];
    assign G[35] = in1[26] & in2[26];
    assign P[35] = in1[26] ^ in2[26];
    assign G[36] = in1[25] & in2[25];
    assign P[36] = in1[25] ^ in2[25];
    assign G[37] = in1[24] & in2[24];
    assign P[37] = in1[24] ^ in2[24];
    assign G[38] = in1[23] & in2[23];
    assign P[38] = in1[23] ^ in2[23];
    assign G[39] = in1[22] & in2[22];
    assign P[39] = in1[22] ^ in2[22];
    assign G[40] = in1[21] & in2[21];
    assign P[40] = in1[21] ^ in2[21];
    assign G[41] = in1[20] & in2[20];
    assign P[41] = in1[20] ^ in2[20];
    assign G[42] = in1[19] & in2[19];
    assign P[42] = in1[19] ^ in2[19];
    assign G[43] = in1[18] & in2[18];
    assign P[43] = in1[18] ^ in2[18];
    assign G[44] = in1[17] & in2[17];
    assign P[44] = in1[17] ^ in2[17];
    assign G[45] = in1[16] & in2[16];
    assign P[45] = in1[16] ^ in2[16];
    assign G[46] = in1[15] & in2[15];
    assign P[46] = in1[15] ^ in2[15];
    assign G[47] = in1[14] & in2[14];
    assign P[47] = in1[14] ^ in2[14];
    assign G[48] = in1[13] & in2[13];
    assign P[48] = in1[13] ^ in2[13];
    assign G[49] = in1[12] & in2[12];
    assign P[49] = in1[12] ^ in2[12];
    assign G[50] = in1[11] & in2[11];
    assign P[50] = in1[11] ^ in2[11];
    assign G[51] = in1[10] & in2[10];
    assign P[51] = in1[10] ^ in2[10];
    assign G[52] = in1[9] & in2[9];
    assign P[52] = in1[9] ^ in2[9];
    assign G[53] = in1[8] & in2[8];
    assign P[53] = in1[8] ^ in2[8];
    assign G[54] = in1[7] & in2[7];
    assign P[54] = in1[7] ^ in2[7];
    assign G[55] = in1[6] & in2[6];
    assign P[55] = in1[6] ^ in2[6];
    assign G[56] = in1[5] & in2[5];
    assign P[56] = in1[5] ^ in2[5];
    assign G[57] = in1[4] & in2[4];
    assign P[57] = in1[4] ^ in2[4];
    assign G[58] = in1[3] & in2[3];
    assign P[58] = in1[3] ^ in2[3];
    assign G[59] = in1[2] & in2[2];
    assign P[59] = in1[2] ^ in2[2];
    assign G[60] = in1[1] & in2[1];
    assign P[60] = in1[1] ^ in2[1];
    assign G[61] = in1[0] & in2[0];
    assign P[61] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign cout = G[61] | (P[61] & C[61]);
    assign sum = P ^ C;
endmodule

module CLA_61(output [60:0] sum, output cout, input [60:0] in1, input [60:0] in2);

    wire[60:0] G;
    wire[60:0] C;
    wire[60:0] P;

    assign G[0] = in1[60] & in2[60];
    assign P[0] = in1[60] ^ in2[60];
    assign G[1] = in1[59] & in2[59];
    assign P[1] = in1[59] ^ in2[59];
    assign G[2] = in1[58] & in2[58];
    assign P[2] = in1[58] ^ in2[58];
    assign G[3] = in1[57] & in2[57];
    assign P[3] = in1[57] ^ in2[57];
    assign G[4] = in1[56] & in2[56];
    assign P[4] = in1[56] ^ in2[56];
    assign G[5] = in1[55] & in2[55];
    assign P[5] = in1[55] ^ in2[55];
    assign G[6] = in1[54] & in2[54];
    assign P[6] = in1[54] ^ in2[54];
    assign G[7] = in1[53] & in2[53];
    assign P[7] = in1[53] ^ in2[53];
    assign G[8] = in1[52] & in2[52];
    assign P[8] = in1[52] ^ in2[52];
    assign G[9] = in1[51] & in2[51];
    assign P[9] = in1[51] ^ in2[51];
    assign G[10] = in1[50] & in2[50];
    assign P[10] = in1[50] ^ in2[50];
    assign G[11] = in1[49] & in2[49];
    assign P[11] = in1[49] ^ in2[49];
    assign G[12] = in1[48] & in2[48];
    assign P[12] = in1[48] ^ in2[48];
    assign G[13] = in1[47] & in2[47];
    assign P[13] = in1[47] ^ in2[47];
    assign G[14] = in1[46] & in2[46];
    assign P[14] = in1[46] ^ in2[46];
    assign G[15] = in1[45] & in2[45];
    assign P[15] = in1[45] ^ in2[45];
    assign G[16] = in1[44] & in2[44];
    assign P[16] = in1[44] ^ in2[44];
    assign G[17] = in1[43] & in2[43];
    assign P[17] = in1[43] ^ in2[43];
    assign G[18] = in1[42] & in2[42];
    assign P[18] = in1[42] ^ in2[42];
    assign G[19] = in1[41] & in2[41];
    assign P[19] = in1[41] ^ in2[41];
    assign G[20] = in1[40] & in2[40];
    assign P[20] = in1[40] ^ in2[40];
    assign G[21] = in1[39] & in2[39];
    assign P[21] = in1[39] ^ in2[39];
    assign G[22] = in1[38] & in2[38];
    assign P[22] = in1[38] ^ in2[38];
    assign G[23] = in1[37] & in2[37];
    assign P[23] = in1[37] ^ in2[37];
    assign G[24] = in1[36] & in2[36];
    assign P[24] = in1[36] ^ in2[36];
    assign G[25] = in1[35] & in2[35];
    assign P[25] = in1[35] ^ in2[35];
    assign G[26] = in1[34] & in2[34];
    assign P[26] = in1[34] ^ in2[34];
    assign G[27] = in1[33] & in2[33];
    assign P[27] = in1[33] ^ in2[33];
    assign G[28] = in1[32] & in2[32];
    assign P[28] = in1[32] ^ in2[32];
    assign G[29] = in1[31] & in2[31];
    assign P[29] = in1[31] ^ in2[31];
    assign G[30] = in1[30] & in2[30];
    assign P[30] = in1[30] ^ in2[30];
    assign G[31] = in1[29] & in2[29];
    assign P[31] = in1[29] ^ in2[29];
    assign G[32] = in1[28] & in2[28];
    assign P[32] = in1[28] ^ in2[28];
    assign G[33] = in1[27] & in2[27];
    assign P[33] = in1[27] ^ in2[27];
    assign G[34] = in1[26] & in2[26];
    assign P[34] = in1[26] ^ in2[26];
    assign G[35] = in1[25] & in2[25];
    assign P[35] = in1[25] ^ in2[25];
    assign G[36] = in1[24] & in2[24];
    assign P[36] = in1[24] ^ in2[24];
    assign G[37] = in1[23] & in2[23];
    assign P[37] = in1[23] ^ in2[23];
    assign G[38] = in1[22] & in2[22];
    assign P[38] = in1[22] ^ in2[22];
    assign G[39] = in1[21] & in2[21];
    assign P[39] = in1[21] ^ in2[21];
    assign G[40] = in1[20] & in2[20];
    assign P[40] = in1[20] ^ in2[20];
    assign G[41] = in1[19] & in2[19];
    assign P[41] = in1[19] ^ in2[19];
    assign G[42] = in1[18] & in2[18];
    assign P[42] = in1[18] ^ in2[18];
    assign G[43] = in1[17] & in2[17];
    assign P[43] = in1[17] ^ in2[17];
    assign G[44] = in1[16] & in2[16];
    assign P[44] = in1[16] ^ in2[16];
    assign G[45] = in1[15] & in2[15];
    assign P[45] = in1[15] ^ in2[15];
    assign G[46] = in1[14] & in2[14];
    assign P[46] = in1[14] ^ in2[14];
    assign G[47] = in1[13] & in2[13];
    assign P[47] = in1[13] ^ in2[13];
    assign G[48] = in1[12] & in2[12];
    assign P[48] = in1[12] ^ in2[12];
    assign G[49] = in1[11] & in2[11];
    assign P[49] = in1[11] ^ in2[11];
    assign G[50] = in1[10] & in2[10];
    assign P[50] = in1[10] ^ in2[10];
    assign G[51] = in1[9] & in2[9];
    assign P[51] = in1[9] ^ in2[9];
    assign G[52] = in1[8] & in2[8];
    assign P[52] = in1[8] ^ in2[8];
    assign G[53] = in1[7] & in2[7];
    assign P[53] = in1[7] ^ in2[7];
    assign G[54] = in1[6] & in2[6];
    assign P[54] = in1[6] ^ in2[6];
    assign G[55] = in1[5] & in2[5];
    assign P[55] = in1[5] ^ in2[5];
    assign G[56] = in1[4] & in2[4];
    assign P[56] = in1[4] ^ in2[4];
    assign G[57] = in1[3] & in2[3];
    assign P[57] = in1[3] ^ in2[3];
    assign G[58] = in1[2] & in2[2];
    assign P[58] = in1[2] ^ in2[2];
    assign G[59] = in1[1] & in2[1];
    assign P[59] = in1[1] ^ in2[1];
    assign G[60] = in1[0] & in2[0];
    assign P[60] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign cout = G[60] | (P[60] & C[60]);
    assign sum = P ^ C;
endmodule

module CLA_60(output [59:0] sum, output cout, input [59:0] in1, input [59:0] in2);

    wire[59:0] G;
    wire[59:0] C;
    wire[59:0] P;

    assign G[0] = in1[59] & in2[59];
    assign P[0] = in1[59] ^ in2[59];
    assign G[1] = in1[58] & in2[58];
    assign P[1] = in1[58] ^ in2[58];
    assign G[2] = in1[57] & in2[57];
    assign P[2] = in1[57] ^ in2[57];
    assign G[3] = in1[56] & in2[56];
    assign P[3] = in1[56] ^ in2[56];
    assign G[4] = in1[55] & in2[55];
    assign P[4] = in1[55] ^ in2[55];
    assign G[5] = in1[54] & in2[54];
    assign P[5] = in1[54] ^ in2[54];
    assign G[6] = in1[53] & in2[53];
    assign P[6] = in1[53] ^ in2[53];
    assign G[7] = in1[52] & in2[52];
    assign P[7] = in1[52] ^ in2[52];
    assign G[8] = in1[51] & in2[51];
    assign P[8] = in1[51] ^ in2[51];
    assign G[9] = in1[50] & in2[50];
    assign P[9] = in1[50] ^ in2[50];
    assign G[10] = in1[49] & in2[49];
    assign P[10] = in1[49] ^ in2[49];
    assign G[11] = in1[48] & in2[48];
    assign P[11] = in1[48] ^ in2[48];
    assign G[12] = in1[47] & in2[47];
    assign P[12] = in1[47] ^ in2[47];
    assign G[13] = in1[46] & in2[46];
    assign P[13] = in1[46] ^ in2[46];
    assign G[14] = in1[45] & in2[45];
    assign P[14] = in1[45] ^ in2[45];
    assign G[15] = in1[44] & in2[44];
    assign P[15] = in1[44] ^ in2[44];
    assign G[16] = in1[43] & in2[43];
    assign P[16] = in1[43] ^ in2[43];
    assign G[17] = in1[42] & in2[42];
    assign P[17] = in1[42] ^ in2[42];
    assign G[18] = in1[41] & in2[41];
    assign P[18] = in1[41] ^ in2[41];
    assign G[19] = in1[40] & in2[40];
    assign P[19] = in1[40] ^ in2[40];
    assign G[20] = in1[39] & in2[39];
    assign P[20] = in1[39] ^ in2[39];
    assign G[21] = in1[38] & in2[38];
    assign P[21] = in1[38] ^ in2[38];
    assign G[22] = in1[37] & in2[37];
    assign P[22] = in1[37] ^ in2[37];
    assign G[23] = in1[36] & in2[36];
    assign P[23] = in1[36] ^ in2[36];
    assign G[24] = in1[35] & in2[35];
    assign P[24] = in1[35] ^ in2[35];
    assign G[25] = in1[34] & in2[34];
    assign P[25] = in1[34] ^ in2[34];
    assign G[26] = in1[33] & in2[33];
    assign P[26] = in1[33] ^ in2[33];
    assign G[27] = in1[32] & in2[32];
    assign P[27] = in1[32] ^ in2[32];
    assign G[28] = in1[31] & in2[31];
    assign P[28] = in1[31] ^ in2[31];
    assign G[29] = in1[30] & in2[30];
    assign P[29] = in1[30] ^ in2[30];
    assign G[30] = in1[29] & in2[29];
    assign P[30] = in1[29] ^ in2[29];
    assign G[31] = in1[28] & in2[28];
    assign P[31] = in1[28] ^ in2[28];
    assign G[32] = in1[27] & in2[27];
    assign P[32] = in1[27] ^ in2[27];
    assign G[33] = in1[26] & in2[26];
    assign P[33] = in1[26] ^ in2[26];
    assign G[34] = in1[25] & in2[25];
    assign P[34] = in1[25] ^ in2[25];
    assign G[35] = in1[24] & in2[24];
    assign P[35] = in1[24] ^ in2[24];
    assign G[36] = in1[23] & in2[23];
    assign P[36] = in1[23] ^ in2[23];
    assign G[37] = in1[22] & in2[22];
    assign P[37] = in1[22] ^ in2[22];
    assign G[38] = in1[21] & in2[21];
    assign P[38] = in1[21] ^ in2[21];
    assign G[39] = in1[20] & in2[20];
    assign P[39] = in1[20] ^ in2[20];
    assign G[40] = in1[19] & in2[19];
    assign P[40] = in1[19] ^ in2[19];
    assign G[41] = in1[18] & in2[18];
    assign P[41] = in1[18] ^ in2[18];
    assign G[42] = in1[17] & in2[17];
    assign P[42] = in1[17] ^ in2[17];
    assign G[43] = in1[16] & in2[16];
    assign P[43] = in1[16] ^ in2[16];
    assign G[44] = in1[15] & in2[15];
    assign P[44] = in1[15] ^ in2[15];
    assign G[45] = in1[14] & in2[14];
    assign P[45] = in1[14] ^ in2[14];
    assign G[46] = in1[13] & in2[13];
    assign P[46] = in1[13] ^ in2[13];
    assign G[47] = in1[12] & in2[12];
    assign P[47] = in1[12] ^ in2[12];
    assign G[48] = in1[11] & in2[11];
    assign P[48] = in1[11] ^ in2[11];
    assign G[49] = in1[10] & in2[10];
    assign P[49] = in1[10] ^ in2[10];
    assign G[50] = in1[9] & in2[9];
    assign P[50] = in1[9] ^ in2[9];
    assign G[51] = in1[8] & in2[8];
    assign P[51] = in1[8] ^ in2[8];
    assign G[52] = in1[7] & in2[7];
    assign P[52] = in1[7] ^ in2[7];
    assign G[53] = in1[6] & in2[6];
    assign P[53] = in1[6] ^ in2[6];
    assign G[54] = in1[5] & in2[5];
    assign P[54] = in1[5] ^ in2[5];
    assign G[55] = in1[4] & in2[4];
    assign P[55] = in1[4] ^ in2[4];
    assign G[56] = in1[3] & in2[3];
    assign P[56] = in1[3] ^ in2[3];
    assign G[57] = in1[2] & in2[2];
    assign P[57] = in1[2] ^ in2[2];
    assign G[58] = in1[1] & in2[1];
    assign P[58] = in1[1] ^ in2[1];
    assign G[59] = in1[0] & in2[0];
    assign P[59] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign cout = G[59] | (P[59] & C[59]);
    assign sum = P ^ C;
endmodule

module CLA_59(output [58:0] sum, output cout, input [58:0] in1, input [58:0] in2);

    wire[58:0] G;
    wire[58:0] C;
    wire[58:0] P;

    assign G[0] = in1[58] & in2[58];
    assign P[0] = in1[58] ^ in2[58];
    assign G[1] = in1[57] & in2[57];
    assign P[1] = in1[57] ^ in2[57];
    assign G[2] = in1[56] & in2[56];
    assign P[2] = in1[56] ^ in2[56];
    assign G[3] = in1[55] & in2[55];
    assign P[3] = in1[55] ^ in2[55];
    assign G[4] = in1[54] & in2[54];
    assign P[4] = in1[54] ^ in2[54];
    assign G[5] = in1[53] & in2[53];
    assign P[5] = in1[53] ^ in2[53];
    assign G[6] = in1[52] & in2[52];
    assign P[6] = in1[52] ^ in2[52];
    assign G[7] = in1[51] & in2[51];
    assign P[7] = in1[51] ^ in2[51];
    assign G[8] = in1[50] & in2[50];
    assign P[8] = in1[50] ^ in2[50];
    assign G[9] = in1[49] & in2[49];
    assign P[9] = in1[49] ^ in2[49];
    assign G[10] = in1[48] & in2[48];
    assign P[10] = in1[48] ^ in2[48];
    assign G[11] = in1[47] & in2[47];
    assign P[11] = in1[47] ^ in2[47];
    assign G[12] = in1[46] & in2[46];
    assign P[12] = in1[46] ^ in2[46];
    assign G[13] = in1[45] & in2[45];
    assign P[13] = in1[45] ^ in2[45];
    assign G[14] = in1[44] & in2[44];
    assign P[14] = in1[44] ^ in2[44];
    assign G[15] = in1[43] & in2[43];
    assign P[15] = in1[43] ^ in2[43];
    assign G[16] = in1[42] & in2[42];
    assign P[16] = in1[42] ^ in2[42];
    assign G[17] = in1[41] & in2[41];
    assign P[17] = in1[41] ^ in2[41];
    assign G[18] = in1[40] & in2[40];
    assign P[18] = in1[40] ^ in2[40];
    assign G[19] = in1[39] & in2[39];
    assign P[19] = in1[39] ^ in2[39];
    assign G[20] = in1[38] & in2[38];
    assign P[20] = in1[38] ^ in2[38];
    assign G[21] = in1[37] & in2[37];
    assign P[21] = in1[37] ^ in2[37];
    assign G[22] = in1[36] & in2[36];
    assign P[22] = in1[36] ^ in2[36];
    assign G[23] = in1[35] & in2[35];
    assign P[23] = in1[35] ^ in2[35];
    assign G[24] = in1[34] & in2[34];
    assign P[24] = in1[34] ^ in2[34];
    assign G[25] = in1[33] & in2[33];
    assign P[25] = in1[33] ^ in2[33];
    assign G[26] = in1[32] & in2[32];
    assign P[26] = in1[32] ^ in2[32];
    assign G[27] = in1[31] & in2[31];
    assign P[27] = in1[31] ^ in2[31];
    assign G[28] = in1[30] & in2[30];
    assign P[28] = in1[30] ^ in2[30];
    assign G[29] = in1[29] & in2[29];
    assign P[29] = in1[29] ^ in2[29];
    assign G[30] = in1[28] & in2[28];
    assign P[30] = in1[28] ^ in2[28];
    assign G[31] = in1[27] & in2[27];
    assign P[31] = in1[27] ^ in2[27];
    assign G[32] = in1[26] & in2[26];
    assign P[32] = in1[26] ^ in2[26];
    assign G[33] = in1[25] & in2[25];
    assign P[33] = in1[25] ^ in2[25];
    assign G[34] = in1[24] & in2[24];
    assign P[34] = in1[24] ^ in2[24];
    assign G[35] = in1[23] & in2[23];
    assign P[35] = in1[23] ^ in2[23];
    assign G[36] = in1[22] & in2[22];
    assign P[36] = in1[22] ^ in2[22];
    assign G[37] = in1[21] & in2[21];
    assign P[37] = in1[21] ^ in2[21];
    assign G[38] = in1[20] & in2[20];
    assign P[38] = in1[20] ^ in2[20];
    assign G[39] = in1[19] & in2[19];
    assign P[39] = in1[19] ^ in2[19];
    assign G[40] = in1[18] & in2[18];
    assign P[40] = in1[18] ^ in2[18];
    assign G[41] = in1[17] & in2[17];
    assign P[41] = in1[17] ^ in2[17];
    assign G[42] = in1[16] & in2[16];
    assign P[42] = in1[16] ^ in2[16];
    assign G[43] = in1[15] & in2[15];
    assign P[43] = in1[15] ^ in2[15];
    assign G[44] = in1[14] & in2[14];
    assign P[44] = in1[14] ^ in2[14];
    assign G[45] = in1[13] & in2[13];
    assign P[45] = in1[13] ^ in2[13];
    assign G[46] = in1[12] & in2[12];
    assign P[46] = in1[12] ^ in2[12];
    assign G[47] = in1[11] & in2[11];
    assign P[47] = in1[11] ^ in2[11];
    assign G[48] = in1[10] & in2[10];
    assign P[48] = in1[10] ^ in2[10];
    assign G[49] = in1[9] & in2[9];
    assign P[49] = in1[9] ^ in2[9];
    assign G[50] = in1[8] & in2[8];
    assign P[50] = in1[8] ^ in2[8];
    assign G[51] = in1[7] & in2[7];
    assign P[51] = in1[7] ^ in2[7];
    assign G[52] = in1[6] & in2[6];
    assign P[52] = in1[6] ^ in2[6];
    assign G[53] = in1[5] & in2[5];
    assign P[53] = in1[5] ^ in2[5];
    assign G[54] = in1[4] & in2[4];
    assign P[54] = in1[4] ^ in2[4];
    assign G[55] = in1[3] & in2[3];
    assign P[55] = in1[3] ^ in2[3];
    assign G[56] = in1[2] & in2[2];
    assign P[56] = in1[2] ^ in2[2];
    assign G[57] = in1[1] & in2[1];
    assign P[57] = in1[1] ^ in2[1];
    assign G[58] = in1[0] & in2[0];
    assign P[58] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign cout = G[58] | (P[58] & C[58]);
    assign sum = P ^ C;
endmodule

module CLA_58(output [57:0] sum, output cout, input [57:0] in1, input [57:0] in2);

    wire[57:0] G;
    wire[57:0] C;
    wire[57:0] P;

    assign G[0] = in1[57] & in2[57];
    assign P[0] = in1[57] ^ in2[57];
    assign G[1] = in1[56] & in2[56];
    assign P[1] = in1[56] ^ in2[56];
    assign G[2] = in1[55] & in2[55];
    assign P[2] = in1[55] ^ in2[55];
    assign G[3] = in1[54] & in2[54];
    assign P[3] = in1[54] ^ in2[54];
    assign G[4] = in1[53] & in2[53];
    assign P[4] = in1[53] ^ in2[53];
    assign G[5] = in1[52] & in2[52];
    assign P[5] = in1[52] ^ in2[52];
    assign G[6] = in1[51] & in2[51];
    assign P[6] = in1[51] ^ in2[51];
    assign G[7] = in1[50] & in2[50];
    assign P[7] = in1[50] ^ in2[50];
    assign G[8] = in1[49] & in2[49];
    assign P[8] = in1[49] ^ in2[49];
    assign G[9] = in1[48] & in2[48];
    assign P[9] = in1[48] ^ in2[48];
    assign G[10] = in1[47] & in2[47];
    assign P[10] = in1[47] ^ in2[47];
    assign G[11] = in1[46] & in2[46];
    assign P[11] = in1[46] ^ in2[46];
    assign G[12] = in1[45] & in2[45];
    assign P[12] = in1[45] ^ in2[45];
    assign G[13] = in1[44] & in2[44];
    assign P[13] = in1[44] ^ in2[44];
    assign G[14] = in1[43] & in2[43];
    assign P[14] = in1[43] ^ in2[43];
    assign G[15] = in1[42] & in2[42];
    assign P[15] = in1[42] ^ in2[42];
    assign G[16] = in1[41] & in2[41];
    assign P[16] = in1[41] ^ in2[41];
    assign G[17] = in1[40] & in2[40];
    assign P[17] = in1[40] ^ in2[40];
    assign G[18] = in1[39] & in2[39];
    assign P[18] = in1[39] ^ in2[39];
    assign G[19] = in1[38] & in2[38];
    assign P[19] = in1[38] ^ in2[38];
    assign G[20] = in1[37] & in2[37];
    assign P[20] = in1[37] ^ in2[37];
    assign G[21] = in1[36] & in2[36];
    assign P[21] = in1[36] ^ in2[36];
    assign G[22] = in1[35] & in2[35];
    assign P[22] = in1[35] ^ in2[35];
    assign G[23] = in1[34] & in2[34];
    assign P[23] = in1[34] ^ in2[34];
    assign G[24] = in1[33] & in2[33];
    assign P[24] = in1[33] ^ in2[33];
    assign G[25] = in1[32] & in2[32];
    assign P[25] = in1[32] ^ in2[32];
    assign G[26] = in1[31] & in2[31];
    assign P[26] = in1[31] ^ in2[31];
    assign G[27] = in1[30] & in2[30];
    assign P[27] = in1[30] ^ in2[30];
    assign G[28] = in1[29] & in2[29];
    assign P[28] = in1[29] ^ in2[29];
    assign G[29] = in1[28] & in2[28];
    assign P[29] = in1[28] ^ in2[28];
    assign G[30] = in1[27] & in2[27];
    assign P[30] = in1[27] ^ in2[27];
    assign G[31] = in1[26] & in2[26];
    assign P[31] = in1[26] ^ in2[26];
    assign G[32] = in1[25] & in2[25];
    assign P[32] = in1[25] ^ in2[25];
    assign G[33] = in1[24] & in2[24];
    assign P[33] = in1[24] ^ in2[24];
    assign G[34] = in1[23] & in2[23];
    assign P[34] = in1[23] ^ in2[23];
    assign G[35] = in1[22] & in2[22];
    assign P[35] = in1[22] ^ in2[22];
    assign G[36] = in1[21] & in2[21];
    assign P[36] = in1[21] ^ in2[21];
    assign G[37] = in1[20] & in2[20];
    assign P[37] = in1[20] ^ in2[20];
    assign G[38] = in1[19] & in2[19];
    assign P[38] = in1[19] ^ in2[19];
    assign G[39] = in1[18] & in2[18];
    assign P[39] = in1[18] ^ in2[18];
    assign G[40] = in1[17] & in2[17];
    assign P[40] = in1[17] ^ in2[17];
    assign G[41] = in1[16] & in2[16];
    assign P[41] = in1[16] ^ in2[16];
    assign G[42] = in1[15] & in2[15];
    assign P[42] = in1[15] ^ in2[15];
    assign G[43] = in1[14] & in2[14];
    assign P[43] = in1[14] ^ in2[14];
    assign G[44] = in1[13] & in2[13];
    assign P[44] = in1[13] ^ in2[13];
    assign G[45] = in1[12] & in2[12];
    assign P[45] = in1[12] ^ in2[12];
    assign G[46] = in1[11] & in2[11];
    assign P[46] = in1[11] ^ in2[11];
    assign G[47] = in1[10] & in2[10];
    assign P[47] = in1[10] ^ in2[10];
    assign G[48] = in1[9] & in2[9];
    assign P[48] = in1[9] ^ in2[9];
    assign G[49] = in1[8] & in2[8];
    assign P[49] = in1[8] ^ in2[8];
    assign G[50] = in1[7] & in2[7];
    assign P[50] = in1[7] ^ in2[7];
    assign G[51] = in1[6] & in2[6];
    assign P[51] = in1[6] ^ in2[6];
    assign G[52] = in1[5] & in2[5];
    assign P[52] = in1[5] ^ in2[5];
    assign G[53] = in1[4] & in2[4];
    assign P[53] = in1[4] ^ in2[4];
    assign G[54] = in1[3] & in2[3];
    assign P[54] = in1[3] ^ in2[3];
    assign G[55] = in1[2] & in2[2];
    assign P[55] = in1[2] ^ in2[2];
    assign G[56] = in1[1] & in2[1];
    assign P[56] = in1[1] ^ in2[1];
    assign G[57] = in1[0] & in2[0];
    assign P[57] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign cout = G[57] | (P[57] & C[57]);
    assign sum = P ^ C;
endmodule

module CLA_57(output [56:0] sum, output cout, input [56:0] in1, input [56:0] in2);

    wire[56:0] G;
    wire[56:0] C;
    wire[56:0] P;

    assign G[0] = in1[56] & in2[56];
    assign P[0] = in1[56] ^ in2[56];
    assign G[1] = in1[55] & in2[55];
    assign P[1] = in1[55] ^ in2[55];
    assign G[2] = in1[54] & in2[54];
    assign P[2] = in1[54] ^ in2[54];
    assign G[3] = in1[53] & in2[53];
    assign P[3] = in1[53] ^ in2[53];
    assign G[4] = in1[52] & in2[52];
    assign P[4] = in1[52] ^ in2[52];
    assign G[5] = in1[51] & in2[51];
    assign P[5] = in1[51] ^ in2[51];
    assign G[6] = in1[50] & in2[50];
    assign P[6] = in1[50] ^ in2[50];
    assign G[7] = in1[49] & in2[49];
    assign P[7] = in1[49] ^ in2[49];
    assign G[8] = in1[48] & in2[48];
    assign P[8] = in1[48] ^ in2[48];
    assign G[9] = in1[47] & in2[47];
    assign P[9] = in1[47] ^ in2[47];
    assign G[10] = in1[46] & in2[46];
    assign P[10] = in1[46] ^ in2[46];
    assign G[11] = in1[45] & in2[45];
    assign P[11] = in1[45] ^ in2[45];
    assign G[12] = in1[44] & in2[44];
    assign P[12] = in1[44] ^ in2[44];
    assign G[13] = in1[43] & in2[43];
    assign P[13] = in1[43] ^ in2[43];
    assign G[14] = in1[42] & in2[42];
    assign P[14] = in1[42] ^ in2[42];
    assign G[15] = in1[41] & in2[41];
    assign P[15] = in1[41] ^ in2[41];
    assign G[16] = in1[40] & in2[40];
    assign P[16] = in1[40] ^ in2[40];
    assign G[17] = in1[39] & in2[39];
    assign P[17] = in1[39] ^ in2[39];
    assign G[18] = in1[38] & in2[38];
    assign P[18] = in1[38] ^ in2[38];
    assign G[19] = in1[37] & in2[37];
    assign P[19] = in1[37] ^ in2[37];
    assign G[20] = in1[36] & in2[36];
    assign P[20] = in1[36] ^ in2[36];
    assign G[21] = in1[35] & in2[35];
    assign P[21] = in1[35] ^ in2[35];
    assign G[22] = in1[34] & in2[34];
    assign P[22] = in1[34] ^ in2[34];
    assign G[23] = in1[33] & in2[33];
    assign P[23] = in1[33] ^ in2[33];
    assign G[24] = in1[32] & in2[32];
    assign P[24] = in1[32] ^ in2[32];
    assign G[25] = in1[31] & in2[31];
    assign P[25] = in1[31] ^ in2[31];
    assign G[26] = in1[30] & in2[30];
    assign P[26] = in1[30] ^ in2[30];
    assign G[27] = in1[29] & in2[29];
    assign P[27] = in1[29] ^ in2[29];
    assign G[28] = in1[28] & in2[28];
    assign P[28] = in1[28] ^ in2[28];
    assign G[29] = in1[27] & in2[27];
    assign P[29] = in1[27] ^ in2[27];
    assign G[30] = in1[26] & in2[26];
    assign P[30] = in1[26] ^ in2[26];
    assign G[31] = in1[25] & in2[25];
    assign P[31] = in1[25] ^ in2[25];
    assign G[32] = in1[24] & in2[24];
    assign P[32] = in1[24] ^ in2[24];
    assign G[33] = in1[23] & in2[23];
    assign P[33] = in1[23] ^ in2[23];
    assign G[34] = in1[22] & in2[22];
    assign P[34] = in1[22] ^ in2[22];
    assign G[35] = in1[21] & in2[21];
    assign P[35] = in1[21] ^ in2[21];
    assign G[36] = in1[20] & in2[20];
    assign P[36] = in1[20] ^ in2[20];
    assign G[37] = in1[19] & in2[19];
    assign P[37] = in1[19] ^ in2[19];
    assign G[38] = in1[18] & in2[18];
    assign P[38] = in1[18] ^ in2[18];
    assign G[39] = in1[17] & in2[17];
    assign P[39] = in1[17] ^ in2[17];
    assign G[40] = in1[16] & in2[16];
    assign P[40] = in1[16] ^ in2[16];
    assign G[41] = in1[15] & in2[15];
    assign P[41] = in1[15] ^ in2[15];
    assign G[42] = in1[14] & in2[14];
    assign P[42] = in1[14] ^ in2[14];
    assign G[43] = in1[13] & in2[13];
    assign P[43] = in1[13] ^ in2[13];
    assign G[44] = in1[12] & in2[12];
    assign P[44] = in1[12] ^ in2[12];
    assign G[45] = in1[11] & in2[11];
    assign P[45] = in1[11] ^ in2[11];
    assign G[46] = in1[10] & in2[10];
    assign P[46] = in1[10] ^ in2[10];
    assign G[47] = in1[9] & in2[9];
    assign P[47] = in1[9] ^ in2[9];
    assign G[48] = in1[8] & in2[8];
    assign P[48] = in1[8] ^ in2[8];
    assign G[49] = in1[7] & in2[7];
    assign P[49] = in1[7] ^ in2[7];
    assign G[50] = in1[6] & in2[6];
    assign P[50] = in1[6] ^ in2[6];
    assign G[51] = in1[5] & in2[5];
    assign P[51] = in1[5] ^ in2[5];
    assign G[52] = in1[4] & in2[4];
    assign P[52] = in1[4] ^ in2[4];
    assign G[53] = in1[3] & in2[3];
    assign P[53] = in1[3] ^ in2[3];
    assign G[54] = in1[2] & in2[2];
    assign P[54] = in1[2] ^ in2[2];
    assign G[55] = in1[1] & in2[1];
    assign P[55] = in1[1] ^ in2[1];
    assign G[56] = in1[0] & in2[0];
    assign P[56] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign cout = G[56] | (P[56] & C[56]);
    assign sum = P ^ C;
endmodule

module CLA_56(output [55:0] sum, output cout, input [55:0] in1, input [55:0] in2);

    wire[55:0] G;
    wire[55:0] C;
    wire[55:0] P;

    assign G[0] = in1[55] & in2[55];
    assign P[0] = in1[55] ^ in2[55];
    assign G[1] = in1[54] & in2[54];
    assign P[1] = in1[54] ^ in2[54];
    assign G[2] = in1[53] & in2[53];
    assign P[2] = in1[53] ^ in2[53];
    assign G[3] = in1[52] & in2[52];
    assign P[3] = in1[52] ^ in2[52];
    assign G[4] = in1[51] & in2[51];
    assign P[4] = in1[51] ^ in2[51];
    assign G[5] = in1[50] & in2[50];
    assign P[5] = in1[50] ^ in2[50];
    assign G[6] = in1[49] & in2[49];
    assign P[6] = in1[49] ^ in2[49];
    assign G[7] = in1[48] & in2[48];
    assign P[7] = in1[48] ^ in2[48];
    assign G[8] = in1[47] & in2[47];
    assign P[8] = in1[47] ^ in2[47];
    assign G[9] = in1[46] & in2[46];
    assign P[9] = in1[46] ^ in2[46];
    assign G[10] = in1[45] & in2[45];
    assign P[10] = in1[45] ^ in2[45];
    assign G[11] = in1[44] & in2[44];
    assign P[11] = in1[44] ^ in2[44];
    assign G[12] = in1[43] & in2[43];
    assign P[12] = in1[43] ^ in2[43];
    assign G[13] = in1[42] & in2[42];
    assign P[13] = in1[42] ^ in2[42];
    assign G[14] = in1[41] & in2[41];
    assign P[14] = in1[41] ^ in2[41];
    assign G[15] = in1[40] & in2[40];
    assign P[15] = in1[40] ^ in2[40];
    assign G[16] = in1[39] & in2[39];
    assign P[16] = in1[39] ^ in2[39];
    assign G[17] = in1[38] & in2[38];
    assign P[17] = in1[38] ^ in2[38];
    assign G[18] = in1[37] & in2[37];
    assign P[18] = in1[37] ^ in2[37];
    assign G[19] = in1[36] & in2[36];
    assign P[19] = in1[36] ^ in2[36];
    assign G[20] = in1[35] & in2[35];
    assign P[20] = in1[35] ^ in2[35];
    assign G[21] = in1[34] & in2[34];
    assign P[21] = in1[34] ^ in2[34];
    assign G[22] = in1[33] & in2[33];
    assign P[22] = in1[33] ^ in2[33];
    assign G[23] = in1[32] & in2[32];
    assign P[23] = in1[32] ^ in2[32];
    assign G[24] = in1[31] & in2[31];
    assign P[24] = in1[31] ^ in2[31];
    assign G[25] = in1[30] & in2[30];
    assign P[25] = in1[30] ^ in2[30];
    assign G[26] = in1[29] & in2[29];
    assign P[26] = in1[29] ^ in2[29];
    assign G[27] = in1[28] & in2[28];
    assign P[27] = in1[28] ^ in2[28];
    assign G[28] = in1[27] & in2[27];
    assign P[28] = in1[27] ^ in2[27];
    assign G[29] = in1[26] & in2[26];
    assign P[29] = in1[26] ^ in2[26];
    assign G[30] = in1[25] & in2[25];
    assign P[30] = in1[25] ^ in2[25];
    assign G[31] = in1[24] & in2[24];
    assign P[31] = in1[24] ^ in2[24];
    assign G[32] = in1[23] & in2[23];
    assign P[32] = in1[23] ^ in2[23];
    assign G[33] = in1[22] & in2[22];
    assign P[33] = in1[22] ^ in2[22];
    assign G[34] = in1[21] & in2[21];
    assign P[34] = in1[21] ^ in2[21];
    assign G[35] = in1[20] & in2[20];
    assign P[35] = in1[20] ^ in2[20];
    assign G[36] = in1[19] & in2[19];
    assign P[36] = in1[19] ^ in2[19];
    assign G[37] = in1[18] & in2[18];
    assign P[37] = in1[18] ^ in2[18];
    assign G[38] = in1[17] & in2[17];
    assign P[38] = in1[17] ^ in2[17];
    assign G[39] = in1[16] & in2[16];
    assign P[39] = in1[16] ^ in2[16];
    assign G[40] = in1[15] & in2[15];
    assign P[40] = in1[15] ^ in2[15];
    assign G[41] = in1[14] & in2[14];
    assign P[41] = in1[14] ^ in2[14];
    assign G[42] = in1[13] & in2[13];
    assign P[42] = in1[13] ^ in2[13];
    assign G[43] = in1[12] & in2[12];
    assign P[43] = in1[12] ^ in2[12];
    assign G[44] = in1[11] & in2[11];
    assign P[44] = in1[11] ^ in2[11];
    assign G[45] = in1[10] & in2[10];
    assign P[45] = in1[10] ^ in2[10];
    assign G[46] = in1[9] & in2[9];
    assign P[46] = in1[9] ^ in2[9];
    assign G[47] = in1[8] & in2[8];
    assign P[47] = in1[8] ^ in2[8];
    assign G[48] = in1[7] & in2[7];
    assign P[48] = in1[7] ^ in2[7];
    assign G[49] = in1[6] & in2[6];
    assign P[49] = in1[6] ^ in2[6];
    assign G[50] = in1[5] & in2[5];
    assign P[50] = in1[5] ^ in2[5];
    assign G[51] = in1[4] & in2[4];
    assign P[51] = in1[4] ^ in2[4];
    assign G[52] = in1[3] & in2[3];
    assign P[52] = in1[3] ^ in2[3];
    assign G[53] = in1[2] & in2[2];
    assign P[53] = in1[2] ^ in2[2];
    assign G[54] = in1[1] & in2[1];
    assign P[54] = in1[1] ^ in2[1];
    assign G[55] = in1[0] & in2[0];
    assign P[55] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign cout = G[55] | (P[55] & C[55]);
    assign sum = P ^ C;
endmodule

module CLA_55(output [54:0] sum, output cout, input [54:0] in1, input [54:0] in2);

    wire[54:0] G;
    wire[54:0] C;
    wire[54:0] P;

    assign G[0] = in1[54] & in2[54];
    assign P[0] = in1[54] ^ in2[54];
    assign G[1] = in1[53] & in2[53];
    assign P[1] = in1[53] ^ in2[53];
    assign G[2] = in1[52] & in2[52];
    assign P[2] = in1[52] ^ in2[52];
    assign G[3] = in1[51] & in2[51];
    assign P[3] = in1[51] ^ in2[51];
    assign G[4] = in1[50] & in2[50];
    assign P[4] = in1[50] ^ in2[50];
    assign G[5] = in1[49] & in2[49];
    assign P[5] = in1[49] ^ in2[49];
    assign G[6] = in1[48] & in2[48];
    assign P[6] = in1[48] ^ in2[48];
    assign G[7] = in1[47] & in2[47];
    assign P[7] = in1[47] ^ in2[47];
    assign G[8] = in1[46] & in2[46];
    assign P[8] = in1[46] ^ in2[46];
    assign G[9] = in1[45] & in2[45];
    assign P[9] = in1[45] ^ in2[45];
    assign G[10] = in1[44] & in2[44];
    assign P[10] = in1[44] ^ in2[44];
    assign G[11] = in1[43] & in2[43];
    assign P[11] = in1[43] ^ in2[43];
    assign G[12] = in1[42] & in2[42];
    assign P[12] = in1[42] ^ in2[42];
    assign G[13] = in1[41] & in2[41];
    assign P[13] = in1[41] ^ in2[41];
    assign G[14] = in1[40] & in2[40];
    assign P[14] = in1[40] ^ in2[40];
    assign G[15] = in1[39] & in2[39];
    assign P[15] = in1[39] ^ in2[39];
    assign G[16] = in1[38] & in2[38];
    assign P[16] = in1[38] ^ in2[38];
    assign G[17] = in1[37] & in2[37];
    assign P[17] = in1[37] ^ in2[37];
    assign G[18] = in1[36] & in2[36];
    assign P[18] = in1[36] ^ in2[36];
    assign G[19] = in1[35] & in2[35];
    assign P[19] = in1[35] ^ in2[35];
    assign G[20] = in1[34] & in2[34];
    assign P[20] = in1[34] ^ in2[34];
    assign G[21] = in1[33] & in2[33];
    assign P[21] = in1[33] ^ in2[33];
    assign G[22] = in1[32] & in2[32];
    assign P[22] = in1[32] ^ in2[32];
    assign G[23] = in1[31] & in2[31];
    assign P[23] = in1[31] ^ in2[31];
    assign G[24] = in1[30] & in2[30];
    assign P[24] = in1[30] ^ in2[30];
    assign G[25] = in1[29] & in2[29];
    assign P[25] = in1[29] ^ in2[29];
    assign G[26] = in1[28] & in2[28];
    assign P[26] = in1[28] ^ in2[28];
    assign G[27] = in1[27] & in2[27];
    assign P[27] = in1[27] ^ in2[27];
    assign G[28] = in1[26] & in2[26];
    assign P[28] = in1[26] ^ in2[26];
    assign G[29] = in1[25] & in2[25];
    assign P[29] = in1[25] ^ in2[25];
    assign G[30] = in1[24] & in2[24];
    assign P[30] = in1[24] ^ in2[24];
    assign G[31] = in1[23] & in2[23];
    assign P[31] = in1[23] ^ in2[23];
    assign G[32] = in1[22] & in2[22];
    assign P[32] = in1[22] ^ in2[22];
    assign G[33] = in1[21] & in2[21];
    assign P[33] = in1[21] ^ in2[21];
    assign G[34] = in1[20] & in2[20];
    assign P[34] = in1[20] ^ in2[20];
    assign G[35] = in1[19] & in2[19];
    assign P[35] = in1[19] ^ in2[19];
    assign G[36] = in1[18] & in2[18];
    assign P[36] = in1[18] ^ in2[18];
    assign G[37] = in1[17] & in2[17];
    assign P[37] = in1[17] ^ in2[17];
    assign G[38] = in1[16] & in2[16];
    assign P[38] = in1[16] ^ in2[16];
    assign G[39] = in1[15] & in2[15];
    assign P[39] = in1[15] ^ in2[15];
    assign G[40] = in1[14] & in2[14];
    assign P[40] = in1[14] ^ in2[14];
    assign G[41] = in1[13] & in2[13];
    assign P[41] = in1[13] ^ in2[13];
    assign G[42] = in1[12] & in2[12];
    assign P[42] = in1[12] ^ in2[12];
    assign G[43] = in1[11] & in2[11];
    assign P[43] = in1[11] ^ in2[11];
    assign G[44] = in1[10] & in2[10];
    assign P[44] = in1[10] ^ in2[10];
    assign G[45] = in1[9] & in2[9];
    assign P[45] = in1[9] ^ in2[9];
    assign G[46] = in1[8] & in2[8];
    assign P[46] = in1[8] ^ in2[8];
    assign G[47] = in1[7] & in2[7];
    assign P[47] = in1[7] ^ in2[7];
    assign G[48] = in1[6] & in2[6];
    assign P[48] = in1[6] ^ in2[6];
    assign G[49] = in1[5] & in2[5];
    assign P[49] = in1[5] ^ in2[5];
    assign G[50] = in1[4] & in2[4];
    assign P[50] = in1[4] ^ in2[4];
    assign G[51] = in1[3] & in2[3];
    assign P[51] = in1[3] ^ in2[3];
    assign G[52] = in1[2] & in2[2];
    assign P[52] = in1[2] ^ in2[2];
    assign G[53] = in1[1] & in2[1];
    assign P[53] = in1[1] ^ in2[1];
    assign G[54] = in1[0] & in2[0];
    assign P[54] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign cout = G[54] | (P[54] & C[54]);
    assign sum = P ^ C;
endmodule

module CLA_54(output [53:0] sum, output cout, input [53:0] in1, input [53:0] in2);

    wire[53:0] G;
    wire[53:0] C;
    wire[53:0] P;

    assign G[0] = in1[53] & in2[53];
    assign P[0] = in1[53] ^ in2[53];
    assign G[1] = in1[52] & in2[52];
    assign P[1] = in1[52] ^ in2[52];
    assign G[2] = in1[51] & in2[51];
    assign P[2] = in1[51] ^ in2[51];
    assign G[3] = in1[50] & in2[50];
    assign P[3] = in1[50] ^ in2[50];
    assign G[4] = in1[49] & in2[49];
    assign P[4] = in1[49] ^ in2[49];
    assign G[5] = in1[48] & in2[48];
    assign P[5] = in1[48] ^ in2[48];
    assign G[6] = in1[47] & in2[47];
    assign P[6] = in1[47] ^ in2[47];
    assign G[7] = in1[46] & in2[46];
    assign P[7] = in1[46] ^ in2[46];
    assign G[8] = in1[45] & in2[45];
    assign P[8] = in1[45] ^ in2[45];
    assign G[9] = in1[44] & in2[44];
    assign P[9] = in1[44] ^ in2[44];
    assign G[10] = in1[43] & in2[43];
    assign P[10] = in1[43] ^ in2[43];
    assign G[11] = in1[42] & in2[42];
    assign P[11] = in1[42] ^ in2[42];
    assign G[12] = in1[41] & in2[41];
    assign P[12] = in1[41] ^ in2[41];
    assign G[13] = in1[40] & in2[40];
    assign P[13] = in1[40] ^ in2[40];
    assign G[14] = in1[39] & in2[39];
    assign P[14] = in1[39] ^ in2[39];
    assign G[15] = in1[38] & in2[38];
    assign P[15] = in1[38] ^ in2[38];
    assign G[16] = in1[37] & in2[37];
    assign P[16] = in1[37] ^ in2[37];
    assign G[17] = in1[36] & in2[36];
    assign P[17] = in1[36] ^ in2[36];
    assign G[18] = in1[35] & in2[35];
    assign P[18] = in1[35] ^ in2[35];
    assign G[19] = in1[34] & in2[34];
    assign P[19] = in1[34] ^ in2[34];
    assign G[20] = in1[33] & in2[33];
    assign P[20] = in1[33] ^ in2[33];
    assign G[21] = in1[32] & in2[32];
    assign P[21] = in1[32] ^ in2[32];
    assign G[22] = in1[31] & in2[31];
    assign P[22] = in1[31] ^ in2[31];
    assign G[23] = in1[30] & in2[30];
    assign P[23] = in1[30] ^ in2[30];
    assign G[24] = in1[29] & in2[29];
    assign P[24] = in1[29] ^ in2[29];
    assign G[25] = in1[28] & in2[28];
    assign P[25] = in1[28] ^ in2[28];
    assign G[26] = in1[27] & in2[27];
    assign P[26] = in1[27] ^ in2[27];
    assign G[27] = in1[26] & in2[26];
    assign P[27] = in1[26] ^ in2[26];
    assign G[28] = in1[25] & in2[25];
    assign P[28] = in1[25] ^ in2[25];
    assign G[29] = in1[24] & in2[24];
    assign P[29] = in1[24] ^ in2[24];
    assign G[30] = in1[23] & in2[23];
    assign P[30] = in1[23] ^ in2[23];
    assign G[31] = in1[22] & in2[22];
    assign P[31] = in1[22] ^ in2[22];
    assign G[32] = in1[21] & in2[21];
    assign P[32] = in1[21] ^ in2[21];
    assign G[33] = in1[20] & in2[20];
    assign P[33] = in1[20] ^ in2[20];
    assign G[34] = in1[19] & in2[19];
    assign P[34] = in1[19] ^ in2[19];
    assign G[35] = in1[18] & in2[18];
    assign P[35] = in1[18] ^ in2[18];
    assign G[36] = in1[17] & in2[17];
    assign P[36] = in1[17] ^ in2[17];
    assign G[37] = in1[16] & in2[16];
    assign P[37] = in1[16] ^ in2[16];
    assign G[38] = in1[15] & in2[15];
    assign P[38] = in1[15] ^ in2[15];
    assign G[39] = in1[14] & in2[14];
    assign P[39] = in1[14] ^ in2[14];
    assign G[40] = in1[13] & in2[13];
    assign P[40] = in1[13] ^ in2[13];
    assign G[41] = in1[12] & in2[12];
    assign P[41] = in1[12] ^ in2[12];
    assign G[42] = in1[11] & in2[11];
    assign P[42] = in1[11] ^ in2[11];
    assign G[43] = in1[10] & in2[10];
    assign P[43] = in1[10] ^ in2[10];
    assign G[44] = in1[9] & in2[9];
    assign P[44] = in1[9] ^ in2[9];
    assign G[45] = in1[8] & in2[8];
    assign P[45] = in1[8] ^ in2[8];
    assign G[46] = in1[7] & in2[7];
    assign P[46] = in1[7] ^ in2[7];
    assign G[47] = in1[6] & in2[6];
    assign P[47] = in1[6] ^ in2[6];
    assign G[48] = in1[5] & in2[5];
    assign P[48] = in1[5] ^ in2[5];
    assign G[49] = in1[4] & in2[4];
    assign P[49] = in1[4] ^ in2[4];
    assign G[50] = in1[3] & in2[3];
    assign P[50] = in1[3] ^ in2[3];
    assign G[51] = in1[2] & in2[2];
    assign P[51] = in1[2] ^ in2[2];
    assign G[52] = in1[1] & in2[1];
    assign P[52] = in1[1] ^ in2[1];
    assign G[53] = in1[0] & in2[0];
    assign P[53] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign cout = G[53] | (P[53] & C[53]);
    assign sum = P ^ C;
endmodule

module CLA_53(output [52:0] sum, output cout, input [52:0] in1, input [52:0] in2);

    wire[52:0] G;
    wire[52:0] C;
    wire[52:0] P;

    assign G[0] = in1[52] & in2[52];
    assign P[0] = in1[52] ^ in2[52];
    assign G[1] = in1[51] & in2[51];
    assign P[1] = in1[51] ^ in2[51];
    assign G[2] = in1[50] & in2[50];
    assign P[2] = in1[50] ^ in2[50];
    assign G[3] = in1[49] & in2[49];
    assign P[3] = in1[49] ^ in2[49];
    assign G[4] = in1[48] & in2[48];
    assign P[4] = in1[48] ^ in2[48];
    assign G[5] = in1[47] & in2[47];
    assign P[5] = in1[47] ^ in2[47];
    assign G[6] = in1[46] & in2[46];
    assign P[6] = in1[46] ^ in2[46];
    assign G[7] = in1[45] & in2[45];
    assign P[7] = in1[45] ^ in2[45];
    assign G[8] = in1[44] & in2[44];
    assign P[8] = in1[44] ^ in2[44];
    assign G[9] = in1[43] & in2[43];
    assign P[9] = in1[43] ^ in2[43];
    assign G[10] = in1[42] & in2[42];
    assign P[10] = in1[42] ^ in2[42];
    assign G[11] = in1[41] & in2[41];
    assign P[11] = in1[41] ^ in2[41];
    assign G[12] = in1[40] & in2[40];
    assign P[12] = in1[40] ^ in2[40];
    assign G[13] = in1[39] & in2[39];
    assign P[13] = in1[39] ^ in2[39];
    assign G[14] = in1[38] & in2[38];
    assign P[14] = in1[38] ^ in2[38];
    assign G[15] = in1[37] & in2[37];
    assign P[15] = in1[37] ^ in2[37];
    assign G[16] = in1[36] & in2[36];
    assign P[16] = in1[36] ^ in2[36];
    assign G[17] = in1[35] & in2[35];
    assign P[17] = in1[35] ^ in2[35];
    assign G[18] = in1[34] & in2[34];
    assign P[18] = in1[34] ^ in2[34];
    assign G[19] = in1[33] & in2[33];
    assign P[19] = in1[33] ^ in2[33];
    assign G[20] = in1[32] & in2[32];
    assign P[20] = in1[32] ^ in2[32];
    assign G[21] = in1[31] & in2[31];
    assign P[21] = in1[31] ^ in2[31];
    assign G[22] = in1[30] & in2[30];
    assign P[22] = in1[30] ^ in2[30];
    assign G[23] = in1[29] & in2[29];
    assign P[23] = in1[29] ^ in2[29];
    assign G[24] = in1[28] & in2[28];
    assign P[24] = in1[28] ^ in2[28];
    assign G[25] = in1[27] & in2[27];
    assign P[25] = in1[27] ^ in2[27];
    assign G[26] = in1[26] & in2[26];
    assign P[26] = in1[26] ^ in2[26];
    assign G[27] = in1[25] & in2[25];
    assign P[27] = in1[25] ^ in2[25];
    assign G[28] = in1[24] & in2[24];
    assign P[28] = in1[24] ^ in2[24];
    assign G[29] = in1[23] & in2[23];
    assign P[29] = in1[23] ^ in2[23];
    assign G[30] = in1[22] & in2[22];
    assign P[30] = in1[22] ^ in2[22];
    assign G[31] = in1[21] & in2[21];
    assign P[31] = in1[21] ^ in2[21];
    assign G[32] = in1[20] & in2[20];
    assign P[32] = in1[20] ^ in2[20];
    assign G[33] = in1[19] & in2[19];
    assign P[33] = in1[19] ^ in2[19];
    assign G[34] = in1[18] & in2[18];
    assign P[34] = in1[18] ^ in2[18];
    assign G[35] = in1[17] & in2[17];
    assign P[35] = in1[17] ^ in2[17];
    assign G[36] = in1[16] & in2[16];
    assign P[36] = in1[16] ^ in2[16];
    assign G[37] = in1[15] & in2[15];
    assign P[37] = in1[15] ^ in2[15];
    assign G[38] = in1[14] & in2[14];
    assign P[38] = in1[14] ^ in2[14];
    assign G[39] = in1[13] & in2[13];
    assign P[39] = in1[13] ^ in2[13];
    assign G[40] = in1[12] & in2[12];
    assign P[40] = in1[12] ^ in2[12];
    assign G[41] = in1[11] & in2[11];
    assign P[41] = in1[11] ^ in2[11];
    assign G[42] = in1[10] & in2[10];
    assign P[42] = in1[10] ^ in2[10];
    assign G[43] = in1[9] & in2[9];
    assign P[43] = in1[9] ^ in2[9];
    assign G[44] = in1[8] & in2[8];
    assign P[44] = in1[8] ^ in2[8];
    assign G[45] = in1[7] & in2[7];
    assign P[45] = in1[7] ^ in2[7];
    assign G[46] = in1[6] & in2[6];
    assign P[46] = in1[6] ^ in2[6];
    assign G[47] = in1[5] & in2[5];
    assign P[47] = in1[5] ^ in2[5];
    assign G[48] = in1[4] & in2[4];
    assign P[48] = in1[4] ^ in2[4];
    assign G[49] = in1[3] & in2[3];
    assign P[49] = in1[3] ^ in2[3];
    assign G[50] = in1[2] & in2[2];
    assign P[50] = in1[2] ^ in2[2];
    assign G[51] = in1[1] & in2[1];
    assign P[51] = in1[1] ^ in2[1];
    assign G[52] = in1[0] & in2[0];
    assign P[52] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign cout = G[52] | (P[52] & C[52]);
    assign sum = P ^ C;
endmodule

module CLA_52(output [51:0] sum, output cout, input [51:0] in1, input [51:0] in2);

    wire[51:0] G;
    wire[51:0] C;
    wire[51:0] P;

    assign G[0] = in1[51] & in2[51];
    assign P[0] = in1[51] ^ in2[51];
    assign G[1] = in1[50] & in2[50];
    assign P[1] = in1[50] ^ in2[50];
    assign G[2] = in1[49] & in2[49];
    assign P[2] = in1[49] ^ in2[49];
    assign G[3] = in1[48] & in2[48];
    assign P[3] = in1[48] ^ in2[48];
    assign G[4] = in1[47] & in2[47];
    assign P[4] = in1[47] ^ in2[47];
    assign G[5] = in1[46] & in2[46];
    assign P[5] = in1[46] ^ in2[46];
    assign G[6] = in1[45] & in2[45];
    assign P[6] = in1[45] ^ in2[45];
    assign G[7] = in1[44] & in2[44];
    assign P[7] = in1[44] ^ in2[44];
    assign G[8] = in1[43] & in2[43];
    assign P[8] = in1[43] ^ in2[43];
    assign G[9] = in1[42] & in2[42];
    assign P[9] = in1[42] ^ in2[42];
    assign G[10] = in1[41] & in2[41];
    assign P[10] = in1[41] ^ in2[41];
    assign G[11] = in1[40] & in2[40];
    assign P[11] = in1[40] ^ in2[40];
    assign G[12] = in1[39] & in2[39];
    assign P[12] = in1[39] ^ in2[39];
    assign G[13] = in1[38] & in2[38];
    assign P[13] = in1[38] ^ in2[38];
    assign G[14] = in1[37] & in2[37];
    assign P[14] = in1[37] ^ in2[37];
    assign G[15] = in1[36] & in2[36];
    assign P[15] = in1[36] ^ in2[36];
    assign G[16] = in1[35] & in2[35];
    assign P[16] = in1[35] ^ in2[35];
    assign G[17] = in1[34] & in2[34];
    assign P[17] = in1[34] ^ in2[34];
    assign G[18] = in1[33] & in2[33];
    assign P[18] = in1[33] ^ in2[33];
    assign G[19] = in1[32] & in2[32];
    assign P[19] = in1[32] ^ in2[32];
    assign G[20] = in1[31] & in2[31];
    assign P[20] = in1[31] ^ in2[31];
    assign G[21] = in1[30] & in2[30];
    assign P[21] = in1[30] ^ in2[30];
    assign G[22] = in1[29] & in2[29];
    assign P[22] = in1[29] ^ in2[29];
    assign G[23] = in1[28] & in2[28];
    assign P[23] = in1[28] ^ in2[28];
    assign G[24] = in1[27] & in2[27];
    assign P[24] = in1[27] ^ in2[27];
    assign G[25] = in1[26] & in2[26];
    assign P[25] = in1[26] ^ in2[26];
    assign G[26] = in1[25] & in2[25];
    assign P[26] = in1[25] ^ in2[25];
    assign G[27] = in1[24] & in2[24];
    assign P[27] = in1[24] ^ in2[24];
    assign G[28] = in1[23] & in2[23];
    assign P[28] = in1[23] ^ in2[23];
    assign G[29] = in1[22] & in2[22];
    assign P[29] = in1[22] ^ in2[22];
    assign G[30] = in1[21] & in2[21];
    assign P[30] = in1[21] ^ in2[21];
    assign G[31] = in1[20] & in2[20];
    assign P[31] = in1[20] ^ in2[20];
    assign G[32] = in1[19] & in2[19];
    assign P[32] = in1[19] ^ in2[19];
    assign G[33] = in1[18] & in2[18];
    assign P[33] = in1[18] ^ in2[18];
    assign G[34] = in1[17] & in2[17];
    assign P[34] = in1[17] ^ in2[17];
    assign G[35] = in1[16] & in2[16];
    assign P[35] = in1[16] ^ in2[16];
    assign G[36] = in1[15] & in2[15];
    assign P[36] = in1[15] ^ in2[15];
    assign G[37] = in1[14] & in2[14];
    assign P[37] = in1[14] ^ in2[14];
    assign G[38] = in1[13] & in2[13];
    assign P[38] = in1[13] ^ in2[13];
    assign G[39] = in1[12] & in2[12];
    assign P[39] = in1[12] ^ in2[12];
    assign G[40] = in1[11] & in2[11];
    assign P[40] = in1[11] ^ in2[11];
    assign G[41] = in1[10] & in2[10];
    assign P[41] = in1[10] ^ in2[10];
    assign G[42] = in1[9] & in2[9];
    assign P[42] = in1[9] ^ in2[9];
    assign G[43] = in1[8] & in2[8];
    assign P[43] = in1[8] ^ in2[8];
    assign G[44] = in1[7] & in2[7];
    assign P[44] = in1[7] ^ in2[7];
    assign G[45] = in1[6] & in2[6];
    assign P[45] = in1[6] ^ in2[6];
    assign G[46] = in1[5] & in2[5];
    assign P[46] = in1[5] ^ in2[5];
    assign G[47] = in1[4] & in2[4];
    assign P[47] = in1[4] ^ in2[4];
    assign G[48] = in1[3] & in2[3];
    assign P[48] = in1[3] ^ in2[3];
    assign G[49] = in1[2] & in2[2];
    assign P[49] = in1[2] ^ in2[2];
    assign G[50] = in1[1] & in2[1];
    assign P[50] = in1[1] ^ in2[1];
    assign G[51] = in1[0] & in2[0];
    assign P[51] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign cout = G[51] | (P[51] & C[51]);
    assign sum = P ^ C;
endmodule

module CLA_51(output [50:0] sum, output cout, input [50:0] in1, input [50:0] in2);

    wire[50:0] G;
    wire[50:0] C;
    wire[50:0] P;

    assign G[0] = in1[50] & in2[50];
    assign P[0] = in1[50] ^ in2[50];
    assign G[1] = in1[49] & in2[49];
    assign P[1] = in1[49] ^ in2[49];
    assign G[2] = in1[48] & in2[48];
    assign P[2] = in1[48] ^ in2[48];
    assign G[3] = in1[47] & in2[47];
    assign P[3] = in1[47] ^ in2[47];
    assign G[4] = in1[46] & in2[46];
    assign P[4] = in1[46] ^ in2[46];
    assign G[5] = in1[45] & in2[45];
    assign P[5] = in1[45] ^ in2[45];
    assign G[6] = in1[44] & in2[44];
    assign P[6] = in1[44] ^ in2[44];
    assign G[7] = in1[43] & in2[43];
    assign P[7] = in1[43] ^ in2[43];
    assign G[8] = in1[42] & in2[42];
    assign P[8] = in1[42] ^ in2[42];
    assign G[9] = in1[41] & in2[41];
    assign P[9] = in1[41] ^ in2[41];
    assign G[10] = in1[40] & in2[40];
    assign P[10] = in1[40] ^ in2[40];
    assign G[11] = in1[39] & in2[39];
    assign P[11] = in1[39] ^ in2[39];
    assign G[12] = in1[38] & in2[38];
    assign P[12] = in1[38] ^ in2[38];
    assign G[13] = in1[37] & in2[37];
    assign P[13] = in1[37] ^ in2[37];
    assign G[14] = in1[36] & in2[36];
    assign P[14] = in1[36] ^ in2[36];
    assign G[15] = in1[35] & in2[35];
    assign P[15] = in1[35] ^ in2[35];
    assign G[16] = in1[34] & in2[34];
    assign P[16] = in1[34] ^ in2[34];
    assign G[17] = in1[33] & in2[33];
    assign P[17] = in1[33] ^ in2[33];
    assign G[18] = in1[32] & in2[32];
    assign P[18] = in1[32] ^ in2[32];
    assign G[19] = in1[31] & in2[31];
    assign P[19] = in1[31] ^ in2[31];
    assign G[20] = in1[30] & in2[30];
    assign P[20] = in1[30] ^ in2[30];
    assign G[21] = in1[29] & in2[29];
    assign P[21] = in1[29] ^ in2[29];
    assign G[22] = in1[28] & in2[28];
    assign P[22] = in1[28] ^ in2[28];
    assign G[23] = in1[27] & in2[27];
    assign P[23] = in1[27] ^ in2[27];
    assign G[24] = in1[26] & in2[26];
    assign P[24] = in1[26] ^ in2[26];
    assign G[25] = in1[25] & in2[25];
    assign P[25] = in1[25] ^ in2[25];
    assign G[26] = in1[24] & in2[24];
    assign P[26] = in1[24] ^ in2[24];
    assign G[27] = in1[23] & in2[23];
    assign P[27] = in1[23] ^ in2[23];
    assign G[28] = in1[22] & in2[22];
    assign P[28] = in1[22] ^ in2[22];
    assign G[29] = in1[21] & in2[21];
    assign P[29] = in1[21] ^ in2[21];
    assign G[30] = in1[20] & in2[20];
    assign P[30] = in1[20] ^ in2[20];
    assign G[31] = in1[19] & in2[19];
    assign P[31] = in1[19] ^ in2[19];
    assign G[32] = in1[18] & in2[18];
    assign P[32] = in1[18] ^ in2[18];
    assign G[33] = in1[17] & in2[17];
    assign P[33] = in1[17] ^ in2[17];
    assign G[34] = in1[16] & in2[16];
    assign P[34] = in1[16] ^ in2[16];
    assign G[35] = in1[15] & in2[15];
    assign P[35] = in1[15] ^ in2[15];
    assign G[36] = in1[14] & in2[14];
    assign P[36] = in1[14] ^ in2[14];
    assign G[37] = in1[13] & in2[13];
    assign P[37] = in1[13] ^ in2[13];
    assign G[38] = in1[12] & in2[12];
    assign P[38] = in1[12] ^ in2[12];
    assign G[39] = in1[11] & in2[11];
    assign P[39] = in1[11] ^ in2[11];
    assign G[40] = in1[10] & in2[10];
    assign P[40] = in1[10] ^ in2[10];
    assign G[41] = in1[9] & in2[9];
    assign P[41] = in1[9] ^ in2[9];
    assign G[42] = in1[8] & in2[8];
    assign P[42] = in1[8] ^ in2[8];
    assign G[43] = in1[7] & in2[7];
    assign P[43] = in1[7] ^ in2[7];
    assign G[44] = in1[6] & in2[6];
    assign P[44] = in1[6] ^ in2[6];
    assign G[45] = in1[5] & in2[5];
    assign P[45] = in1[5] ^ in2[5];
    assign G[46] = in1[4] & in2[4];
    assign P[46] = in1[4] ^ in2[4];
    assign G[47] = in1[3] & in2[3];
    assign P[47] = in1[3] ^ in2[3];
    assign G[48] = in1[2] & in2[2];
    assign P[48] = in1[2] ^ in2[2];
    assign G[49] = in1[1] & in2[1];
    assign P[49] = in1[1] ^ in2[1];
    assign G[50] = in1[0] & in2[0];
    assign P[50] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign cout = G[50] | (P[50] & C[50]);
    assign sum = P ^ C;
endmodule

module CLA_50(output [49:0] sum, output cout, input [49:0] in1, input [49:0] in2);

    wire[49:0] G;
    wire[49:0] C;
    wire[49:0] P;

    assign G[0] = in1[49] & in2[49];
    assign P[0] = in1[49] ^ in2[49];
    assign G[1] = in1[48] & in2[48];
    assign P[1] = in1[48] ^ in2[48];
    assign G[2] = in1[47] & in2[47];
    assign P[2] = in1[47] ^ in2[47];
    assign G[3] = in1[46] & in2[46];
    assign P[3] = in1[46] ^ in2[46];
    assign G[4] = in1[45] & in2[45];
    assign P[4] = in1[45] ^ in2[45];
    assign G[5] = in1[44] & in2[44];
    assign P[5] = in1[44] ^ in2[44];
    assign G[6] = in1[43] & in2[43];
    assign P[6] = in1[43] ^ in2[43];
    assign G[7] = in1[42] & in2[42];
    assign P[7] = in1[42] ^ in2[42];
    assign G[8] = in1[41] & in2[41];
    assign P[8] = in1[41] ^ in2[41];
    assign G[9] = in1[40] & in2[40];
    assign P[9] = in1[40] ^ in2[40];
    assign G[10] = in1[39] & in2[39];
    assign P[10] = in1[39] ^ in2[39];
    assign G[11] = in1[38] & in2[38];
    assign P[11] = in1[38] ^ in2[38];
    assign G[12] = in1[37] & in2[37];
    assign P[12] = in1[37] ^ in2[37];
    assign G[13] = in1[36] & in2[36];
    assign P[13] = in1[36] ^ in2[36];
    assign G[14] = in1[35] & in2[35];
    assign P[14] = in1[35] ^ in2[35];
    assign G[15] = in1[34] & in2[34];
    assign P[15] = in1[34] ^ in2[34];
    assign G[16] = in1[33] & in2[33];
    assign P[16] = in1[33] ^ in2[33];
    assign G[17] = in1[32] & in2[32];
    assign P[17] = in1[32] ^ in2[32];
    assign G[18] = in1[31] & in2[31];
    assign P[18] = in1[31] ^ in2[31];
    assign G[19] = in1[30] & in2[30];
    assign P[19] = in1[30] ^ in2[30];
    assign G[20] = in1[29] & in2[29];
    assign P[20] = in1[29] ^ in2[29];
    assign G[21] = in1[28] & in2[28];
    assign P[21] = in1[28] ^ in2[28];
    assign G[22] = in1[27] & in2[27];
    assign P[22] = in1[27] ^ in2[27];
    assign G[23] = in1[26] & in2[26];
    assign P[23] = in1[26] ^ in2[26];
    assign G[24] = in1[25] & in2[25];
    assign P[24] = in1[25] ^ in2[25];
    assign G[25] = in1[24] & in2[24];
    assign P[25] = in1[24] ^ in2[24];
    assign G[26] = in1[23] & in2[23];
    assign P[26] = in1[23] ^ in2[23];
    assign G[27] = in1[22] & in2[22];
    assign P[27] = in1[22] ^ in2[22];
    assign G[28] = in1[21] & in2[21];
    assign P[28] = in1[21] ^ in2[21];
    assign G[29] = in1[20] & in2[20];
    assign P[29] = in1[20] ^ in2[20];
    assign G[30] = in1[19] & in2[19];
    assign P[30] = in1[19] ^ in2[19];
    assign G[31] = in1[18] & in2[18];
    assign P[31] = in1[18] ^ in2[18];
    assign G[32] = in1[17] & in2[17];
    assign P[32] = in1[17] ^ in2[17];
    assign G[33] = in1[16] & in2[16];
    assign P[33] = in1[16] ^ in2[16];
    assign G[34] = in1[15] & in2[15];
    assign P[34] = in1[15] ^ in2[15];
    assign G[35] = in1[14] & in2[14];
    assign P[35] = in1[14] ^ in2[14];
    assign G[36] = in1[13] & in2[13];
    assign P[36] = in1[13] ^ in2[13];
    assign G[37] = in1[12] & in2[12];
    assign P[37] = in1[12] ^ in2[12];
    assign G[38] = in1[11] & in2[11];
    assign P[38] = in1[11] ^ in2[11];
    assign G[39] = in1[10] & in2[10];
    assign P[39] = in1[10] ^ in2[10];
    assign G[40] = in1[9] & in2[9];
    assign P[40] = in1[9] ^ in2[9];
    assign G[41] = in1[8] & in2[8];
    assign P[41] = in1[8] ^ in2[8];
    assign G[42] = in1[7] & in2[7];
    assign P[42] = in1[7] ^ in2[7];
    assign G[43] = in1[6] & in2[6];
    assign P[43] = in1[6] ^ in2[6];
    assign G[44] = in1[5] & in2[5];
    assign P[44] = in1[5] ^ in2[5];
    assign G[45] = in1[4] & in2[4];
    assign P[45] = in1[4] ^ in2[4];
    assign G[46] = in1[3] & in2[3];
    assign P[46] = in1[3] ^ in2[3];
    assign G[47] = in1[2] & in2[2];
    assign P[47] = in1[2] ^ in2[2];
    assign G[48] = in1[1] & in2[1];
    assign P[48] = in1[1] ^ in2[1];
    assign G[49] = in1[0] & in2[0];
    assign P[49] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign cout = G[49] | (P[49] & C[49]);
    assign sum = P ^ C;
endmodule

module CLA_49(output [48:0] sum, output cout, input [48:0] in1, input [48:0] in2);

    wire[48:0] G;
    wire[48:0] C;
    wire[48:0] P;

    assign G[0] = in1[48] & in2[48];
    assign P[0] = in1[48] ^ in2[48];
    assign G[1] = in1[47] & in2[47];
    assign P[1] = in1[47] ^ in2[47];
    assign G[2] = in1[46] & in2[46];
    assign P[2] = in1[46] ^ in2[46];
    assign G[3] = in1[45] & in2[45];
    assign P[3] = in1[45] ^ in2[45];
    assign G[4] = in1[44] & in2[44];
    assign P[4] = in1[44] ^ in2[44];
    assign G[5] = in1[43] & in2[43];
    assign P[5] = in1[43] ^ in2[43];
    assign G[6] = in1[42] & in2[42];
    assign P[6] = in1[42] ^ in2[42];
    assign G[7] = in1[41] & in2[41];
    assign P[7] = in1[41] ^ in2[41];
    assign G[8] = in1[40] & in2[40];
    assign P[8] = in1[40] ^ in2[40];
    assign G[9] = in1[39] & in2[39];
    assign P[9] = in1[39] ^ in2[39];
    assign G[10] = in1[38] & in2[38];
    assign P[10] = in1[38] ^ in2[38];
    assign G[11] = in1[37] & in2[37];
    assign P[11] = in1[37] ^ in2[37];
    assign G[12] = in1[36] & in2[36];
    assign P[12] = in1[36] ^ in2[36];
    assign G[13] = in1[35] & in2[35];
    assign P[13] = in1[35] ^ in2[35];
    assign G[14] = in1[34] & in2[34];
    assign P[14] = in1[34] ^ in2[34];
    assign G[15] = in1[33] & in2[33];
    assign P[15] = in1[33] ^ in2[33];
    assign G[16] = in1[32] & in2[32];
    assign P[16] = in1[32] ^ in2[32];
    assign G[17] = in1[31] & in2[31];
    assign P[17] = in1[31] ^ in2[31];
    assign G[18] = in1[30] & in2[30];
    assign P[18] = in1[30] ^ in2[30];
    assign G[19] = in1[29] & in2[29];
    assign P[19] = in1[29] ^ in2[29];
    assign G[20] = in1[28] & in2[28];
    assign P[20] = in1[28] ^ in2[28];
    assign G[21] = in1[27] & in2[27];
    assign P[21] = in1[27] ^ in2[27];
    assign G[22] = in1[26] & in2[26];
    assign P[22] = in1[26] ^ in2[26];
    assign G[23] = in1[25] & in2[25];
    assign P[23] = in1[25] ^ in2[25];
    assign G[24] = in1[24] & in2[24];
    assign P[24] = in1[24] ^ in2[24];
    assign G[25] = in1[23] & in2[23];
    assign P[25] = in1[23] ^ in2[23];
    assign G[26] = in1[22] & in2[22];
    assign P[26] = in1[22] ^ in2[22];
    assign G[27] = in1[21] & in2[21];
    assign P[27] = in1[21] ^ in2[21];
    assign G[28] = in1[20] & in2[20];
    assign P[28] = in1[20] ^ in2[20];
    assign G[29] = in1[19] & in2[19];
    assign P[29] = in1[19] ^ in2[19];
    assign G[30] = in1[18] & in2[18];
    assign P[30] = in1[18] ^ in2[18];
    assign G[31] = in1[17] & in2[17];
    assign P[31] = in1[17] ^ in2[17];
    assign G[32] = in1[16] & in2[16];
    assign P[32] = in1[16] ^ in2[16];
    assign G[33] = in1[15] & in2[15];
    assign P[33] = in1[15] ^ in2[15];
    assign G[34] = in1[14] & in2[14];
    assign P[34] = in1[14] ^ in2[14];
    assign G[35] = in1[13] & in2[13];
    assign P[35] = in1[13] ^ in2[13];
    assign G[36] = in1[12] & in2[12];
    assign P[36] = in1[12] ^ in2[12];
    assign G[37] = in1[11] & in2[11];
    assign P[37] = in1[11] ^ in2[11];
    assign G[38] = in1[10] & in2[10];
    assign P[38] = in1[10] ^ in2[10];
    assign G[39] = in1[9] & in2[9];
    assign P[39] = in1[9] ^ in2[9];
    assign G[40] = in1[8] & in2[8];
    assign P[40] = in1[8] ^ in2[8];
    assign G[41] = in1[7] & in2[7];
    assign P[41] = in1[7] ^ in2[7];
    assign G[42] = in1[6] & in2[6];
    assign P[42] = in1[6] ^ in2[6];
    assign G[43] = in1[5] & in2[5];
    assign P[43] = in1[5] ^ in2[5];
    assign G[44] = in1[4] & in2[4];
    assign P[44] = in1[4] ^ in2[4];
    assign G[45] = in1[3] & in2[3];
    assign P[45] = in1[3] ^ in2[3];
    assign G[46] = in1[2] & in2[2];
    assign P[46] = in1[2] ^ in2[2];
    assign G[47] = in1[1] & in2[1];
    assign P[47] = in1[1] ^ in2[1];
    assign G[48] = in1[0] & in2[0];
    assign P[48] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign cout = G[48] | (P[48] & C[48]);
    assign sum = P ^ C;
endmodule

module CLA_48(output [47:0] sum, output cout, input [47:0] in1, input [47:0] in2);

    wire[47:0] G;
    wire[47:0] C;
    wire[47:0] P;

    assign G[0] = in1[47] & in2[47];
    assign P[0] = in1[47] ^ in2[47];
    assign G[1] = in1[46] & in2[46];
    assign P[1] = in1[46] ^ in2[46];
    assign G[2] = in1[45] & in2[45];
    assign P[2] = in1[45] ^ in2[45];
    assign G[3] = in1[44] & in2[44];
    assign P[3] = in1[44] ^ in2[44];
    assign G[4] = in1[43] & in2[43];
    assign P[4] = in1[43] ^ in2[43];
    assign G[5] = in1[42] & in2[42];
    assign P[5] = in1[42] ^ in2[42];
    assign G[6] = in1[41] & in2[41];
    assign P[6] = in1[41] ^ in2[41];
    assign G[7] = in1[40] & in2[40];
    assign P[7] = in1[40] ^ in2[40];
    assign G[8] = in1[39] & in2[39];
    assign P[8] = in1[39] ^ in2[39];
    assign G[9] = in1[38] & in2[38];
    assign P[9] = in1[38] ^ in2[38];
    assign G[10] = in1[37] & in2[37];
    assign P[10] = in1[37] ^ in2[37];
    assign G[11] = in1[36] & in2[36];
    assign P[11] = in1[36] ^ in2[36];
    assign G[12] = in1[35] & in2[35];
    assign P[12] = in1[35] ^ in2[35];
    assign G[13] = in1[34] & in2[34];
    assign P[13] = in1[34] ^ in2[34];
    assign G[14] = in1[33] & in2[33];
    assign P[14] = in1[33] ^ in2[33];
    assign G[15] = in1[32] & in2[32];
    assign P[15] = in1[32] ^ in2[32];
    assign G[16] = in1[31] & in2[31];
    assign P[16] = in1[31] ^ in2[31];
    assign G[17] = in1[30] & in2[30];
    assign P[17] = in1[30] ^ in2[30];
    assign G[18] = in1[29] & in2[29];
    assign P[18] = in1[29] ^ in2[29];
    assign G[19] = in1[28] & in2[28];
    assign P[19] = in1[28] ^ in2[28];
    assign G[20] = in1[27] & in2[27];
    assign P[20] = in1[27] ^ in2[27];
    assign G[21] = in1[26] & in2[26];
    assign P[21] = in1[26] ^ in2[26];
    assign G[22] = in1[25] & in2[25];
    assign P[22] = in1[25] ^ in2[25];
    assign G[23] = in1[24] & in2[24];
    assign P[23] = in1[24] ^ in2[24];
    assign G[24] = in1[23] & in2[23];
    assign P[24] = in1[23] ^ in2[23];
    assign G[25] = in1[22] & in2[22];
    assign P[25] = in1[22] ^ in2[22];
    assign G[26] = in1[21] & in2[21];
    assign P[26] = in1[21] ^ in2[21];
    assign G[27] = in1[20] & in2[20];
    assign P[27] = in1[20] ^ in2[20];
    assign G[28] = in1[19] & in2[19];
    assign P[28] = in1[19] ^ in2[19];
    assign G[29] = in1[18] & in2[18];
    assign P[29] = in1[18] ^ in2[18];
    assign G[30] = in1[17] & in2[17];
    assign P[30] = in1[17] ^ in2[17];
    assign G[31] = in1[16] & in2[16];
    assign P[31] = in1[16] ^ in2[16];
    assign G[32] = in1[15] & in2[15];
    assign P[32] = in1[15] ^ in2[15];
    assign G[33] = in1[14] & in2[14];
    assign P[33] = in1[14] ^ in2[14];
    assign G[34] = in1[13] & in2[13];
    assign P[34] = in1[13] ^ in2[13];
    assign G[35] = in1[12] & in2[12];
    assign P[35] = in1[12] ^ in2[12];
    assign G[36] = in1[11] & in2[11];
    assign P[36] = in1[11] ^ in2[11];
    assign G[37] = in1[10] & in2[10];
    assign P[37] = in1[10] ^ in2[10];
    assign G[38] = in1[9] & in2[9];
    assign P[38] = in1[9] ^ in2[9];
    assign G[39] = in1[8] & in2[8];
    assign P[39] = in1[8] ^ in2[8];
    assign G[40] = in1[7] & in2[7];
    assign P[40] = in1[7] ^ in2[7];
    assign G[41] = in1[6] & in2[6];
    assign P[41] = in1[6] ^ in2[6];
    assign G[42] = in1[5] & in2[5];
    assign P[42] = in1[5] ^ in2[5];
    assign G[43] = in1[4] & in2[4];
    assign P[43] = in1[4] ^ in2[4];
    assign G[44] = in1[3] & in2[3];
    assign P[44] = in1[3] ^ in2[3];
    assign G[45] = in1[2] & in2[2];
    assign P[45] = in1[2] ^ in2[2];
    assign G[46] = in1[1] & in2[1];
    assign P[46] = in1[1] ^ in2[1];
    assign G[47] = in1[0] & in2[0];
    assign P[47] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign cout = G[47] | (P[47] & C[47]);
    assign sum = P ^ C;
endmodule

module CLA_47(output [46:0] sum, output cout, input [46:0] in1, input [46:0] in2);

    wire[46:0] G;
    wire[46:0] C;
    wire[46:0] P;

    assign G[0] = in1[46] & in2[46];
    assign P[0] = in1[46] ^ in2[46];
    assign G[1] = in1[45] & in2[45];
    assign P[1] = in1[45] ^ in2[45];
    assign G[2] = in1[44] & in2[44];
    assign P[2] = in1[44] ^ in2[44];
    assign G[3] = in1[43] & in2[43];
    assign P[3] = in1[43] ^ in2[43];
    assign G[4] = in1[42] & in2[42];
    assign P[4] = in1[42] ^ in2[42];
    assign G[5] = in1[41] & in2[41];
    assign P[5] = in1[41] ^ in2[41];
    assign G[6] = in1[40] & in2[40];
    assign P[6] = in1[40] ^ in2[40];
    assign G[7] = in1[39] & in2[39];
    assign P[7] = in1[39] ^ in2[39];
    assign G[8] = in1[38] & in2[38];
    assign P[8] = in1[38] ^ in2[38];
    assign G[9] = in1[37] & in2[37];
    assign P[9] = in1[37] ^ in2[37];
    assign G[10] = in1[36] & in2[36];
    assign P[10] = in1[36] ^ in2[36];
    assign G[11] = in1[35] & in2[35];
    assign P[11] = in1[35] ^ in2[35];
    assign G[12] = in1[34] & in2[34];
    assign P[12] = in1[34] ^ in2[34];
    assign G[13] = in1[33] & in2[33];
    assign P[13] = in1[33] ^ in2[33];
    assign G[14] = in1[32] & in2[32];
    assign P[14] = in1[32] ^ in2[32];
    assign G[15] = in1[31] & in2[31];
    assign P[15] = in1[31] ^ in2[31];
    assign G[16] = in1[30] & in2[30];
    assign P[16] = in1[30] ^ in2[30];
    assign G[17] = in1[29] & in2[29];
    assign P[17] = in1[29] ^ in2[29];
    assign G[18] = in1[28] & in2[28];
    assign P[18] = in1[28] ^ in2[28];
    assign G[19] = in1[27] & in2[27];
    assign P[19] = in1[27] ^ in2[27];
    assign G[20] = in1[26] & in2[26];
    assign P[20] = in1[26] ^ in2[26];
    assign G[21] = in1[25] & in2[25];
    assign P[21] = in1[25] ^ in2[25];
    assign G[22] = in1[24] & in2[24];
    assign P[22] = in1[24] ^ in2[24];
    assign G[23] = in1[23] & in2[23];
    assign P[23] = in1[23] ^ in2[23];
    assign G[24] = in1[22] & in2[22];
    assign P[24] = in1[22] ^ in2[22];
    assign G[25] = in1[21] & in2[21];
    assign P[25] = in1[21] ^ in2[21];
    assign G[26] = in1[20] & in2[20];
    assign P[26] = in1[20] ^ in2[20];
    assign G[27] = in1[19] & in2[19];
    assign P[27] = in1[19] ^ in2[19];
    assign G[28] = in1[18] & in2[18];
    assign P[28] = in1[18] ^ in2[18];
    assign G[29] = in1[17] & in2[17];
    assign P[29] = in1[17] ^ in2[17];
    assign G[30] = in1[16] & in2[16];
    assign P[30] = in1[16] ^ in2[16];
    assign G[31] = in1[15] & in2[15];
    assign P[31] = in1[15] ^ in2[15];
    assign G[32] = in1[14] & in2[14];
    assign P[32] = in1[14] ^ in2[14];
    assign G[33] = in1[13] & in2[13];
    assign P[33] = in1[13] ^ in2[13];
    assign G[34] = in1[12] & in2[12];
    assign P[34] = in1[12] ^ in2[12];
    assign G[35] = in1[11] & in2[11];
    assign P[35] = in1[11] ^ in2[11];
    assign G[36] = in1[10] & in2[10];
    assign P[36] = in1[10] ^ in2[10];
    assign G[37] = in1[9] & in2[9];
    assign P[37] = in1[9] ^ in2[9];
    assign G[38] = in1[8] & in2[8];
    assign P[38] = in1[8] ^ in2[8];
    assign G[39] = in1[7] & in2[7];
    assign P[39] = in1[7] ^ in2[7];
    assign G[40] = in1[6] & in2[6];
    assign P[40] = in1[6] ^ in2[6];
    assign G[41] = in1[5] & in2[5];
    assign P[41] = in1[5] ^ in2[5];
    assign G[42] = in1[4] & in2[4];
    assign P[42] = in1[4] ^ in2[4];
    assign G[43] = in1[3] & in2[3];
    assign P[43] = in1[3] ^ in2[3];
    assign G[44] = in1[2] & in2[2];
    assign P[44] = in1[2] ^ in2[2];
    assign G[45] = in1[1] & in2[1];
    assign P[45] = in1[1] ^ in2[1];
    assign G[46] = in1[0] & in2[0];
    assign P[46] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign cout = G[46] | (P[46] & C[46]);
    assign sum = P ^ C;
endmodule

module CLA_46(output [45:0] sum, output cout, input [45:0] in1, input [45:0] in2);

    wire[45:0] G;
    wire[45:0] C;
    wire[45:0] P;

    assign G[0] = in1[45] & in2[45];
    assign P[0] = in1[45] ^ in2[45];
    assign G[1] = in1[44] & in2[44];
    assign P[1] = in1[44] ^ in2[44];
    assign G[2] = in1[43] & in2[43];
    assign P[2] = in1[43] ^ in2[43];
    assign G[3] = in1[42] & in2[42];
    assign P[3] = in1[42] ^ in2[42];
    assign G[4] = in1[41] & in2[41];
    assign P[4] = in1[41] ^ in2[41];
    assign G[5] = in1[40] & in2[40];
    assign P[5] = in1[40] ^ in2[40];
    assign G[6] = in1[39] & in2[39];
    assign P[6] = in1[39] ^ in2[39];
    assign G[7] = in1[38] & in2[38];
    assign P[7] = in1[38] ^ in2[38];
    assign G[8] = in1[37] & in2[37];
    assign P[8] = in1[37] ^ in2[37];
    assign G[9] = in1[36] & in2[36];
    assign P[9] = in1[36] ^ in2[36];
    assign G[10] = in1[35] & in2[35];
    assign P[10] = in1[35] ^ in2[35];
    assign G[11] = in1[34] & in2[34];
    assign P[11] = in1[34] ^ in2[34];
    assign G[12] = in1[33] & in2[33];
    assign P[12] = in1[33] ^ in2[33];
    assign G[13] = in1[32] & in2[32];
    assign P[13] = in1[32] ^ in2[32];
    assign G[14] = in1[31] & in2[31];
    assign P[14] = in1[31] ^ in2[31];
    assign G[15] = in1[30] & in2[30];
    assign P[15] = in1[30] ^ in2[30];
    assign G[16] = in1[29] & in2[29];
    assign P[16] = in1[29] ^ in2[29];
    assign G[17] = in1[28] & in2[28];
    assign P[17] = in1[28] ^ in2[28];
    assign G[18] = in1[27] & in2[27];
    assign P[18] = in1[27] ^ in2[27];
    assign G[19] = in1[26] & in2[26];
    assign P[19] = in1[26] ^ in2[26];
    assign G[20] = in1[25] & in2[25];
    assign P[20] = in1[25] ^ in2[25];
    assign G[21] = in1[24] & in2[24];
    assign P[21] = in1[24] ^ in2[24];
    assign G[22] = in1[23] & in2[23];
    assign P[22] = in1[23] ^ in2[23];
    assign G[23] = in1[22] & in2[22];
    assign P[23] = in1[22] ^ in2[22];
    assign G[24] = in1[21] & in2[21];
    assign P[24] = in1[21] ^ in2[21];
    assign G[25] = in1[20] & in2[20];
    assign P[25] = in1[20] ^ in2[20];
    assign G[26] = in1[19] & in2[19];
    assign P[26] = in1[19] ^ in2[19];
    assign G[27] = in1[18] & in2[18];
    assign P[27] = in1[18] ^ in2[18];
    assign G[28] = in1[17] & in2[17];
    assign P[28] = in1[17] ^ in2[17];
    assign G[29] = in1[16] & in2[16];
    assign P[29] = in1[16] ^ in2[16];
    assign G[30] = in1[15] & in2[15];
    assign P[30] = in1[15] ^ in2[15];
    assign G[31] = in1[14] & in2[14];
    assign P[31] = in1[14] ^ in2[14];
    assign G[32] = in1[13] & in2[13];
    assign P[32] = in1[13] ^ in2[13];
    assign G[33] = in1[12] & in2[12];
    assign P[33] = in1[12] ^ in2[12];
    assign G[34] = in1[11] & in2[11];
    assign P[34] = in1[11] ^ in2[11];
    assign G[35] = in1[10] & in2[10];
    assign P[35] = in1[10] ^ in2[10];
    assign G[36] = in1[9] & in2[9];
    assign P[36] = in1[9] ^ in2[9];
    assign G[37] = in1[8] & in2[8];
    assign P[37] = in1[8] ^ in2[8];
    assign G[38] = in1[7] & in2[7];
    assign P[38] = in1[7] ^ in2[7];
    assign G[39] = in1[6] & in2[6];
    assign P[39] = in1[6] ^ in2[6];
    assign G[40] = in1[5] & in2[5];
    assign P[40] = in1[5] ^ in2[5];
    assign G[41] = in1[4] & in2[4];
    assign P[41] = in1[4] ^ in2[4];
    assign G[42] = in1[3] & in2[3];
    assign P[42] = in1[3] ^ in2[3];
    assign G[43] = in1[2] & in2[2];
    assign P[43] = in1[2] ^ in2[2];
    assign G[44] = in1[1] & in2[1];
    assign P[44] = in1[1] ^ in2[1];
    assign G[45] = in1[0] & in2[0];
    assign P[45] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign cout = G[45] | (P[45] & C[45]);
    assign sum = P ^ C;
endmodule

module CLA_45(output [44:0] sum, output cout, input [44:0] in1, input [44:0] in2);

    wire[44:0] G;
    wire[44:0] C;
    wire[44:0] P;

    assign G[0] = in1[44] & in2[44];
    assign P[0] = in1[44] ^ in2[44];
    assign G[1] = in1[43] & in2[43];
    assign P[1] = in1[43] ^ in2[43];
    assign G[2] = in1[42] & in2[42];
    assign P[2] = in1[42] ^ in2[42];
    assign G[3] = in1[41] & in2[41];
    assign P[3] = in1[41] ^ in2[41];
    assign G[4] = in1[40] & in2[40];
    assign P[4] = in1[40] ^ in2[40];
    assign G[5] = in1[39] & in2[39];
    assign P[5] = in1[39] ^ in2[39];
    assign G[6] = in1[38] & in2[38];
    assign P[6] = in1[38] ^ in2[38];
    assign G[7] = in1[37] & in2[37];
    assign P[7] = in1[37] ^ in2[37];
    assign G[8] = in1[36] & in2[36];
    assign P[8] = in1[36] ^ in2[36];
    assign G[9] = in1[35] & in2[35];
    assign P[9] = in1[35] ^ in2[35];
    assign G[10] = in1[34] & in2[34];
    assign P[10] = in1[34] ^ in2[34];
    assign G[11] = in1[33] & in2[33];
    assign P[11] = in1[33] ^ in2[33];
    assign G[12] = in1[32] & in2[32];
    assign P[12] = in1[32] ^ in2[32];
    assign G[13] = in1[31] & in2[31];
    assign P[13] = in1[31] ^ in2[31];
    assign G[14] = in1[30] & in2[30];
    assign P[14] = in1[30] ^ in2[30];
    assign G[15] = in1[29] & in2[29];
    assign P[15] = in1[29] ^ in2[29];
    assign G[16] = in1[28] & in2[28];
    assign P[16] = in1[28] ^ in2[28];
    assign G[17] = in1[27] & in2[27];
    assign P[17] = in1[27] ^ in2[27];
    assign G[18] = in1[26] & in2[26];
    assign P[18] = in1[26] ^ in2[26];
    assign G[19] = in1[25] & in2[25];
    assign P[19] = in1[25] ^ in2[25];
    assign G[20] = in1[24] & in2[24];
    assign P[20] = in1[24] ^ in2[24];
    assign G[21] = in1[23] & in2[23];
    assign P[21] = in1[23] ^ in2[23];
    assign G[22] = in1[22] & in2[22];
    assign P[22] = in1[22] ^ in2[22];
    assign G[23] = in1[21] & in2[21];
    assign P[23] = in1[21] ^ in2[21];
    assign G[24] = in1[20] & in2[20];
    assign P[24] = in1[20] ^ in2[20];
    assign G[25] = in1[19] & in2[19];
    assign P[25] = in1[19] ^ in2[19];
    assign G[26] = in1[18] & in2[18];
    assign P[26] = in1[18] ^ in2[18];
    assign G[27] = in1[17] & in2[17];
    assign P[27] = in1[17] ^ in2[17];
    assign G[28] = in1[16] & in2[16];
    assign P[28] = in1[16] ^ in2[16];
    assign G[29] = in1[15] & in2[15];
    assign P[29] = in1[15] ^ in2[15];
    assign G[30] = in1[14] & in2[14];
    assign P[30] = in1[14] ^ in2[14];
    assign G[31] = in1[13] & in2[13];
    assign P[31] = in1[13] ^ in2[13];
    assign G[32] = in1[12] & in2[12];
    assign P[32] = in1[12] ^ in2[12];
    assign G[33] = in1[11] & in2[11];
    assign P[33] = in1[11] ^ in2[11];
    assign G[34] = in1[10] & in2[10];
    assign P[34] = in1[10] ^ in2[10];
    assign G[35] = in1[9] & in2[9];
    assign P[35] = in1[9] ^ in2[9];
    assign G[36] = in1[8] & in2[8];
    assign P[36] = in1[8] ^ in2[8];
    assign G[37] = in1[7] & in2[7];
    assign P[37] = in1[7] ^ in2[7];
    assign G[38] = in1[6] & in2[6];
    assign P[38] = in1[6] ^ in2[6];
    assign G[39] = in1[5] & in2[5];
    assign P[39] = in1[5] ^ in2[5];
    assign G[40] = in1[4] & in2[4];
    assign P[40] = in1[4] ^ in2[4];
    assign G[41] = in1[3] & in2[3];
    assign P[41] = in1[3] ^ in2[3];
    assign G[42] = in1[2] & in2[2];
    assign P[42] = in1[2] ^ in2[2];
    assign G[43] = in1[1] & in2[1];
    assign P[43] = in1[1] ^ in2[1];
    assign G[44] = in1[0] & in2[0];
    assign P[44] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign cout = G[44] | (P[44] & C[44]);
    assign sum = P ^ C;
endmodule

module CLA_44(output [43:0] sum, output cout, input [43:0] in1, input [43:0] in2);

    wire[43:0] G;
    wire[43:0] C;
    wire[43:0] P;

    assign G[0] = in1[43] & in2[43];
    assign P[0] = in1[43] ^ in2[43];
    assign G[1] = in1[42] & in2[42];
    assign P[1] = in1[42] ^ in2[42];
    assign G[2] = in1[41] & in2[41];
    assign P[2] = in1[41] ^ in2[41];
    assign G[3] = in1[40] & in2[40];
    assign P[3] = in1[40] ^ in2[40];
    assign G[4] = in1[39] & in2[39];
    assign P[4] = in1[39] ^ in2[39];
    assign G[5] = in1[38] & in2[38];
    assign P[5] = in1[38] ^ in2[38];
    assign G[6] = in1[37] & in2[37];
    assign P[6] = in1[37] ^ in2[37];
    assign G[7] = in1[36] & in2[36];
    assign P[7] = in1[36] ^ in2[36];
    assign G[8] = in1[35] & in2[35];
    assign P[8] = in1[35] ^ in2[35];
    assign G[9] = in1[34] & in2[34];
    assign P[9] = in1[34] ^ in2[34];
    assign G[10] = in1[33] & in2[33];
    assign P[10] = in1[33] ^ in2[33];
    assign G[11] = in1[32] & in2[32];
    assign P[11] = in1[32] ^ in2[32];
    assign G[12] = in1[31] & in2[31];
    assign P[12] = in1[31] ^ in2[31];
    assign G[13] = in1[30] & in2[30];
    assign P[13] = in1[30] ^ in2[30];
    assign G[14] = in1[29] & in2[29];
    assign P[14] = in1[29] ^ in2[29];
    assign G[15] = in1[28] & in2[28];
    assign P[15] = in1[28] ^ in2[28];
    assign G[16] = in1[27] & in2[27];
    assign P[16] = in1[27] ^ in2[27];
    assign G[17] = in1[26] & in2[26];
    assign P[17] = in1[26] ^ in2[26];
    assign G[18] = in1[25] & in2[25];
    assign P[18] = in1[25] ^ in2[25];
    assign G[19] = in1[24] & in2[24];
    assign P[19] = in1[24] ^ in2[24];
    assign G[20] = in1[23] & in2[23];
    assign P[20] = in1[23] ^ in2[23];
    assign G[21] = in1[22] & in2[22];
    assign P[21] = in1[22] ^ in2[22];
    assign G[22] = in1[21] & in2[21];
    assign P[22] = in1[21] ^ in2[21];
    assign G[23] = in1[20] & in2[20];
    assign P[23] = in1[20] ^ in2[20];
    assign G[24] = in1[19] & in2[19];
    assign P[24] = in1[19] ^ in2[19];
    assign G[25] = in1[18] & in2[18];
    assign P[25] = in1[18] ^ in2[18];
    assign G[26] = in1[17] & in2[17];
    assign P[26] = in1[17] ^ in2[17];
    assign G[27] = in1[16] & in2[16];
    assign P[27] = in1[16] ^ in2[16];
    assign G[28] = in1[15] & in2[15];
    assign P[28] = in1[15] ^ in2[15];
    assign G[29] = in1[14] & in2[14];
    assign P[29] = in1[14] ^ in2[14];
    assign G[30] = in1[13] & in2[13];
    assign P[30] = in1[13] ^ in2[13];
    assign G[31] = in1[12] & in2[12];
    assign P[31] = in1[12] ^ in2[12];
    assign G[32] = in1[11] & in2[11];
    assign P[32] = in1[11] ^ in2[11];
    assign G[33] = in1[10] & in2[10];
    assign P[33] = in1[10] ^ in2[10];
    assign G[34] = in1[9] & in2[9];
    assign P[34] = in1[9] ^ in2[9];
    assign G[35] = in1[8] & in2[8];
    assign P[35] = in1[8] ^ in2[8];
    assign G[36] = in1[7] & in2[7];
    assign P[36] = in1[7] ^ in2[7];
    assign G[37] = in1[6] & in2[6];
    assign P[37] = in1[6] ^ in2[6];
    assign G[38] = in1[5] & in2[5];
    assign P[38] = in1[5] ^ in2[5];
    assign G[39] = in1[4] & in2[4];
    assign P[39] = in1[4] ^ in2[4];
    assign G[40] = in1[3] & in2[3];
    assign P[40] = in1[3] ^ in2[3];
    assign G[41] = in1[2] & in2[2];
    assign P[41] = in1[2] ^ in2[2];
    assign G[42] = in1[1] & in2[1];
    assign P[42] = in1[1] ^ in2[1];
    assign G[43] = in1[0] & in2[0];
    assign P[43] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign cout = G[43] | (P[43] & C[43]);
    assign sum = P ^ C;
endmodule

module CLA_43(output [42:0] sum, output cout, input [42:0] in1, input [42:0] in2);

    wire[42:0] G;
    wire[42:0] C;
    wire[42:0] P;

    assign G[0] = in1[42] & in2[42];
    assign P[0] = in1[42] ^ in2[42];
    assign G[1] = in1[41] & in2[41];
    assign P[1] = in1[41] ^ in2[41];
    assign G[2] = in1[40] & in2[40];
    assign P[2] = in1[40] ^ in2[40];
    assign G[3] = in1[39] & in2[39];
    assign P[3] = in1[39] ^ in2[39];
    assign G[4] = in1[38] & in2[38];
    assign P[4] = in1[38] ^ in2[38];
    assign G[5] = in1[37] & in2[37];
    assign P[5] = in1[37] ^ in2[37];
    assign G[6] = in1[36] & in2[36];
    assign P[6] = in1[36] ^ in2[36];
    assign G[7] = in1[35] & in2[35];
    assign P[7] = in1[35] ^ in2[35];
    assign G[8] = in1[34] & in2[34];
    assign P[8] = in1[34] ^ in2[34];
    assign G[9] = in1[33] & in2[33];
    assign P[9] = in1[33] ^ in2[33];
    assign G[10] = in1[32] & in2[32];
    assign P[10] = in1[32] ^ in2[32];
    assign G[11] = in1[31] & in2[31];
    assign P[11] = in1[31] ^ in2[31];
    assign G[12] = in1[30] & in2[30];
    assign P[12] = in1[30] ^ in2[30];
    assign G[13] = in1[29] & in2[29];
    assign P[13] = in1[29] ^ in2[29];
    assign G[14] = in1[28] & in2[28];
    assign P[14] = in1[28] ^ in2[28];
    assign G[15] = in1[27] & in2[27];
    assign P[15] = in1[27] ^ in2[27];
    assign G[16] = in1[26] & in2[26];
    assign P[16] = in1[26] ^ in2[26];
    assign G[17] = in1[25] & in2[25];
    assign P[17] = in1[25] ^ in2[25];
    assign G[18] = in1[24] & in2[24];
    assign P[18] = in1[24] ^ in2[24];
    assign G[19] = in1[23] & in2[23];
    assign P[19] = in1[23] ^ in2[23];
    assign G[20] = in1[22] & in2[22];
    assign P[20] = in1[22] ^ in2[22];
    assign G[21] = in1[21] & in2[21];
    assign P[21] = in1[21] ^ in2[21];
    assign G[22] = in1[20] & in2[20];
    assign P[22] = in1[20] ^ in2[20];
    assign G[23] = in1[19] & in2[19];
    assign P[23] = in1[19] ^ in2[19];
    assign G[24] = in1[18] & in2[18];
    assign P[24] = in1[18] ^ in2[18];
    assign G[25] = in1[17] & in2[17];
    assign P[25] = in1[17] ^ in2[17];
    assign G[26] = in1[16] & in2[16];
    assign P[26] = in1[16] ^ in2[16];
    assign G[27] = in1[15] & in2[15];
    assign P[27] = in1[15] ^ in2[15];
    assign G[28] = in1[14] & in2[14];
    assign P[28] = in1[14] ^ in2[14];
    assign G[29] = in1[13] & in2[13];
    assign P[29] = in1[13] ^ in2[13];
    assign G[30] = in1[12] & in2[12];
    assign P[30] = in1[12] ^ in2[12];
    assign G[31] = in1[11] & in2[11];
    assign P[31] = in1[11] ^ in2[11];
    assign G[32] = in1[10] & in2[10];
    assign P[32] = in1[10] ^ in2[10];
    assign G[33] = in1[9] & in2[9];
    assign P[33] = in1[9] ^ in2[9];
    assign G[34] = in1[8] & in2[8];
    assign P[34] = in1[8] ^ in2[8];
    assign G[35] = in1[7] & in2[7];
    assign P[35] = in1[7] ^ in2[7];
    assign G[36] = in1[6] & in2[6];
    assign P[36] = in1[6] ^ in2[6];
    assign G[37] = in1[5] & in2[5];
    assign P[37] = in1[5] ^ in2[5];
    assign G[38] = in1[4] & in2[4];
    assign P[38] = in1[4] ^ in2[4];
    assign G[39] = in1[3] & in2[3];
    assign P[39] = in1[3] ^ in2[3];
    assign G[40] = in1[2] & in2[2];
    assign P[40] = in1[2] ^ in2[2];
    assign G[41] = in1[1] & in2[1];
    assign P[41] = in1[1] ^ in2[1];
    assign G[42] = in1[0] & in2[0];
    assign P[42] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign cout = G[42] | (P[42] & C[42]);
    assign sum = P ^ C;
endmodule

module CLA_42(output [41:0] sum, output cout, input [41:0] in1, input [41:0] in2);

    wire[41:0] G;
    wire[41:0] C;
    wire[41:0] P;

    assign G[0] = in1[41] & in2[41];
    assign P[0] = in1[41] ^ in2[41];
    assign G[1] = in1[40] & in2[40];
    assign P[1] = in1[40] ^ in2[40];
    assign G[2] = in1[39] & in2[39];
    assign P[2] = in1[39] ^ in2[39];
    assign G[3] = in1[38] & in2[38];
    assign P[3] = in1[38] ^ in2[38];
    assign G[4] = in1[37] & in2[37];
    assign P[4] = in1[37] ^ in2[37];
    assign G[5] = in1[36] & in2[36];
    assign P[5] = in1[36] ^ in2[36];
    assign G[6] = in1[35] & in2[35];
    assign P[6] = in1[35] ^ in2[35];
    assign G[7] = in1[34] & in2[34];
    assign P[7] = in1[34] ^ in2[34];
    assign G[8] = in1[33] & in2[33];
    assign P[8] = in1[33] ^ in2[33];
    assign G[9] = in1[32] & in2[32];
    assign P[9] = in1[32] ^ in2[32];
    assign G[10] = in1[31] & in2[31];
    assign P[10] = in1[31] ^ in2[31];
    assign G[11] = in1[30] & in2[30];
    assign P[11] = in1[30] ^ in2[30];
    assign G[12] = in1[29] & in2[29];
    assign P[12] = in1[29] ^ in2[29];
    assign G[13] = in1[28] & in2[28];
    assign P[13] = in1[28] ^ in2[28];
    assign G[14] = in1[27] & in2[27];
    assign P[14] = in1[27] ^ in2[27];
    assign G[15] = in1[26] & in2[26];
    assign P[15] = in1[26] ^ in2[26];
    assign G[16] = in1[25] & in2[25];
    assign P[16] = in1[25] ^ in2[25];
    assign G[17] = in1[24] & in2[24];
    assign P[17] = in1[24] ^ in2[24];
    assign G[18] = in1[23] & in2[23];
    assign P[18] = in1[23] ^ in2[23];
    assign G[19] = in1[22] & in2[22];
    assign P[19] = in1[22] ^ in2[22];
    assign G[20] = in1[21] & in2[21];
    assign P[20] = in1[21] ^ in2[21];
    assign G[21] = in1[20] & in2[20];
    assign P[21] = in1[20] ^ in2[20];
    assign G[22] = in1[19] & in2[19];
    assign P[22] = in1[19] ^ in2[19];
    assign G[23] = in1[18] & in2[18];
    assign P[23] = in1[18] ^ in2[18];
    assign G[24] = in1[17] & in2[17];
    assign P[24] = in1[17] ^ in2[17];
    assign G[25] = in1[16] & in2[16];
    assign P[25] = in1[16] ^ in2[16];
    assign G[26] = in1[15] & in2[15];
    assign P[26] = in1[15] ^ in2[15];
    assign G[27] = in1[14] & in2[14];
    assign P[27] = in1[14] ^ in2[14];
    assign G[28] = in1[13] & in2[13];
    assign P[28] = in1[13] ^ in2[13];
    assign G[29] = in1[12] & in2[12];
    assign P[29] = in1[12] ^ in2[12];
    assign G[30] = in1[11] & in2[11];
    assign P[30] = in1[11] ^ in2[11];
    assign G[31] = in1[10] & in2[10];
    assign P[31] = in1[10] ^ in2[10];
    assign G[32] = in1[9] & in2[9];
    assign P[32] = in1[9] ^ in2[9];
    assign G[33] = in1[8] & in2[8];
    assign P[33] = in1[8] ^ in2[8];
    assign G[34] = in1[7] & in2[7];
    assign P[34] = in1[7] ^ in2[7];
    assign G[35] = in1[6] & in2[6];
    assign P[35] = in1[6] ^ in2[6];
    assign G[36] = in1[5] & in2[5];
    assign P[36] = in1[5] ^ in2[5];
    assign G[37] = in1[4] & in2[4];
    assign P[37] = in1[4] ^ in2[4];
    assign G[38] = in1[3] & in2[3];
    assign P[38] = in1[3] ^ in2[3];
    assign G[39] = in1[2] & in2[2];
    assign P[39] = in1[2] ^ in2[2];
    assign G[40] = in1[1] & in2[1];
    assign P[40] = in1[1] ^ in2[1];
    assign G[41] = in1[0] & in2[0];
    assign P[41] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign cout = G[41] | (P[41] & C[41]);
    assign sum = P ^ C;
endmodule

module CLA_41(output [40:0] sum, output cout, input [40:0] in1, input [40:0] in2);

    wire[40:0] G;
    wire[40:0] C;
    wire[40:0] P;

    assign G[0] = in1[40] & in2[40];
    assign P[0] = in1[40] ^ in2[40];
    assign G[1] = in1[39] & in2[39];
    assign P[1] = in1[39] ^ in2[39];
    assign G[2] = in1[38] & in2[38];
    assign P[2] = in1[38] ^ in2[38];
    assign G[3] = in1[37] & in2[37];
    assign P[3] = in1[37] ^ in2[37];
    assign G[4] = in1[36] & in2[36];
    assign P[4] = in1[36] ^ in2[36];
    assign G[5] = in1[35] & in2[35];
    assign P[5] = in1[35] ^ in2[35];
    assign G[6] = in1[34] & in2[34];
    assign P[6] = in1[34] ^ in2[34];
    assign G[7] = in1[33] & in2[33];
    assign P[7] = in1[33] ^ in2[33];
    assign G[8] = in1[32] & in2[32];
    assign P[8] = in1[32] ^ in2[32];
    assign G[9] = in1[31] & in2[31];
    assign P[9] = in1[31] ^ in2[31];
    assign G[10] = in1[30] & in2[30];
    assign P[10] = in1[30] ^ in2[30];
    assign G[11] = in1[29] & in2[29];
    assign P[11] = in1[29] ^ in2[29];
    assign G[12] = in1[28] & in2[28];
    assign P[12] = in1[28] ^ in2[28];
    assign G[13] = in1[27] & in2[27];
    assign P[13] = in1[27] ^ in2[27];
    assign G[14] = in1[26] & in2[26];
    assign P[14] = in1[26] ^ in2[26];
    assign G[15] = in1[25] & in2[25];
    assign P[15] = in1[25] ^ in2[25];
    assign G[16] = in1[24] & in2[24];
    assign P[16] = in1[24] ^ in2[24];
    assign G[17] = in1[23] & in2[23];
    assign P[17] = in1[23] ^ in2[23];
    assign G[18] = in1[22] & in2[22];
    assign P[18] = in1[22] ^ in2[22];
    assign G[19] = in1[21] & in2[21];
    assign P[19] = in1[21] ^ in2[21];
    assign G[20] = in1[20] & in2[20];
    assign P[20] = in1[20] ^ in2[20];
    assign G[21] = in1[19] & in2[19];
    assign P[21] = in1[19] ^ in2[19];
    assign G[22] = in1[18] & in2[18];
    assign P[22] = in1[18] ^ in2[18];
    assign G[23] = in1[17] & in2[17];
    assign P[23] = in1[17] ^ in2[17];
    assign G[24] = in1[16] & in2[16];
    assign P[24] = in1[16] ^ in2[16];
    assign G[25] = in1[15] & in2[15];
    assign P[25] = in1[15] ^ in2[15];
    assign G[26] = in1[14] & in2[14];
    assign P[26] = in1[14] ^ in2[14];
    assign G[27] = in1[13] & in2[13];
    assign P[27] = in1[13] ^ in2[13];
    assign G[28] = in1[12] & in2[12];
    assign P[28] = in1[12] ^ in2[12];
    assign G[29] = in1[11] & in2[11];
    assign P[29] = in1[11] ^ in2[11];
    assign G[30] = in1[10] & in2[10];
    assign P[30] = in1[10] ^ in2[10];
    assign G[31] = in1[9] & in2[9];
    assign P[31] = in1[9] ^ in2[9];
    assign G[32] = in1[8] & in2[8];
    assign P[32] = in1[8] ^ in2[8];
    assign G[33] = in1[7] & in2[7];
    assign P[33] = in1[7] ^ in2[7];
    assign G[34] = in1[6] & in2[6];
    assign P[34] = in1[6] ^ in2[6];
    assign G[35] = in1[5] & in2[5];
    assign P[35] = in1[5] ^ in2[5];
    assign G[36] = in1[4] & in2[4];
    assign P[36] = in1[4] ^ in2[4];
    assign G[37] = in1[3] & in2[3];
    assign P[37] = in1[3] ^ in2[3];
    assign G[38] = in1[2] & in2[2];
    assign P[38] = in1[2] ^ in2[2];
    assign G[39] = in1[1] & in2[1];
    assign P[39] = in1[1] ^ in2[1];
    assign G[40] = in1[0] & in2[0];
    assign P[40] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign cout = G[40] | (P[40] & C[40]);
    assign sum = P ^ C;
endmodule

module CLA_40(output [39:0] sum, output cout, input [39:0] in1, input [39:0] in2);

    wire[39:0] G;
    wire[39:0] C;
    wire[39:0] P;

    assign G[0] = in1[39] & in2[39];
    assign P[0] = in1[39] ^ in2[39];
    assign G[1] = in1[38] & in2[38];
    assign P[1] = in1[38] ^ in2[38];
    assign G[2] = in1[37] & in2[37];
    assign P[2] = in1[37] ^ in2[37];
    assign G[3] = in1[36] & in2[36];
    assign P[3] = in1[36] ^ in2[36];
    assign G[4] = in1[35] & in2[35];
    assign P[4] = in1[35] ^ in2[35];
    assign G[5] = in1[34] & in2[34];
    assign P[5] = in1[34] ^ in2[34];
    assign G[6] = in1[33] & in2[33];
    assign P[6] = in1[33] ^ in2[33];
    assign G[7] = in1[32] & in2[32];
    assign P[7] = in1[32] ^ in2[32];
    assign G[8] = in1[31] & in2[31];
    assign P[8] = in1[31] ^ in2[31];
    assign G[9] = in1[30] & in2[30];
    assign P[9] = in1[30] ^ in2[30];
    assign G[10] = in1[29] & in2[29];
    assign P[10] = in1[29] ^ in2[29];
    assign G[11] = in1[28] & in2[28];
    assign P[11] = in1[28] ^ in2[28];
    assign G[12] = in1[27] & in2[27];
    assign P[12] = in1[27] ^ in2[27];
    assign G[13] = in1[26] & in2[26];
    assign P[13] = in1[26] ^ in2[26];
    assign G[14] = in1[25] & in2[25];
    assign P[14] = in1[25] ^ in2[25];
    assign G[15] = in1[24] & in2[24];
    assign P[15] = in1[24] ^ in2[24];
    assign G[16] = in1[23] & in2[23];
    assign P[16] = in1[23] ^ in2[23];
    assign G[17] = in1[22] & in2[22];
    assign P[17] = in1[22] ^ in2[22];
    assign G[18] = in1[21] & in2[21];
    assign P[18] = in1[21] ^ in2[21];
    assign G[19] = in1[20] & in2[20];
    assign P[19] = in1[20] ^ in2[20];
    assign G[20] = in1[19] & in2[19];
    assign P[20] = in1[19] ^ in2[19];
    assign G[21] = in1[18] & in2[18];
    assign P[21] = in1[18] ^ in2[18];
    assign G[22] = in1[17] & in2[17];
    assign P[22] = in1[17] ^ in2[17];
    assign G[23] = in1[16] & in2[16];
    assign P[23] = in1[16] ^ in2[16];
    assign G[24] = in1[15] & in2[15];
    assign P[24] = in1[15] ^ in2[15];
    assign G[25] = in1[14] & in2[14];
    assign P[25] = in1[14] ^ in2[14];
    assign G[26] = in1[13] & in2[13];
    assign P[26] = in1[13] ^ in2[13];
    assign G[27] = in1[12] & in2[12];
    assign P[27] = in1[12] ^ in2[12];
    assign G[28] = in1[11] & in2[11];
    assign P[28] = in1[11] ^ in2[11];
    assign G[29] = in1[10] & in2[10];
    assign P[29] = in1[10] ^ in2[10];
    assign G[30] = in1[9] & in2[9];
    assign P[30] = in1[9] ^ in2[9];
    assign G[31] = in1[8] & in2[8];
    assign P[31] = in1[8] ^ in2[8];
    assign G[32] = in1[7] & in2[7];
    assign P[32] = in1[7] ^ in2[7];
    assign G[33] = in1[6] & in2[6];
    assign P[33] = in1[6] ^ in2[6];
    assign G[34] = in1[5] & in2[5];
    assign P[34] = in1[5] ^ in2[5];
    assign G[35] = in1[4] & in2[4];
    assign P[35] = in1[4] ^ in2[4];
    assign G[36] = in1[3] & in2[3];
    assign P[36] = in1[3] ^ in2[3];
    assign G[37] = in1[2] & in2[2];
    assign P[37] = in1[2] ^ in2[2];
    assign G[38] = in1[1] & in2[1];
    assign P[38] = in1[1] ^ in2[1];
    assign G[39] = in1[0] & in2[0];
    assign P[39] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign cout = G[39] | (P[39] & C[39]);
    assign sum = P ^ C;
endmodule

module CLA_39(output [38:0] sum, output cout, input [38:0] in1, input [38:0] in2);

    wire[38:0] G;
    wire[38:0] C;
    wire[38:0] P;

    assign G[0] = in1[38] & in2[38];
    assign P[0] = in1[38] ^ in2[38];
    assign G[1] = in1[37] & in2[37];
    assign P[1] = in1[37] ^ in2[37];
    assign G[2] = in1[36] & in2[36];
    assign P[2] = in1[36] ^ in2[36];
    assign G[3] = in1[35] & in2[35];
    assign P[3] = in1[35] ^ in2[35];
    assign G[4] = in1[34] & in2[34];
    assign P[4] = in1[34] ^ in2[34];
    assign G[5] = in1[33] & in2[33];
    assign P[5] = in1[33] ^ in2[33];
    assign G[6] = in1[32] & in2[32];
    assign P[6] = in1[32] ^ in2[32];
    assign G[7] = in1[31] & in2[31];
    assign P[7] = in1[31] ^ in2[31];
    assign G[8] = in1[30] & in2[30];
    assign P[8] = in1[30] ^ in2[30];
    assign G[9] = in1[29] & in2[29];
    assign P[9] = in1[29] ^ in2[29];
    assign G[10] = in1[28] & in2[28];
    assign P[10] = in1[28] ^ in2[28];
    assign G[11] = in1[27] & in2[27];
    assign P[11] = in1[27] ^ in2[27];
    assign G[12] = in1[26] & in2[26];
    assign P[12] = in1[26] ^ in2[26];
    assign G[13] = in1[25] & in2[25];
    assign P[13] = in1[25] ^ in2[25];
    assign G[14] = in1[24] & in2[24];
    assign P[14] = in1[24] ^ in2[24];
    assign G[15] = in1[23] & in2[23];
    assign P[15] = in1[23] ^ in2[23];
    assign G[16] = in1[22] & in2[22];
    assign P[16] = in1[22] ^ in2[22];
    assign G[17] = in1[21] & in2[21];
    assign P[17] = in1[21] ^ in2[21];
    assign G[18] = in1[20] & in2[20];
    assign P[18] = in1[20] ^ in2[20];
    assign G[19] = in1[19] & in2[19];
    assign P[19] = in1[19] ^ in2[19];
    assign G[20] = in1[18] & in2[18];
    assign P[20] = in1[18] ^ in2[18];
    assign G[21] = in1[17] & in2[17];
    assign P[21] = in1[17] ^ in2[17];
    assign G[22] = in1[16] & in2[16];
    assign P[22] = in1[16] ^ in2[16];
    assign G[23] = in1[15] & in2[15];
    assign P[23] = in1[15] ^ in2[15];
    assign G[24] = in1[14] & in2[14];
    assign P[24] = in1[14] ^ in2[14];
    assign G[25] = in1[13] & in2[13];
    assign P[25] = in1[13] ^ in2[13];
    assign G[26] = in1[12] & in2[12];
    assign P[26] = in1[12] ^ in2[12];
    assign G[27] = in1[11] & in2[11];
    assign P[27] = in1[11] ^ in2[11];
    assign G[28] = in1[10] & in2[10];
    assign P[28] = in1[10] ^ in2[10];
    assign G[29] = in1[9] & in2[9];
    assign P[29] = in1[9] ^ in2[9];
    assign G[30] = in1[8] & in2[8];
    assign P[30] = in1[8] ^ in2[8];
    assign G[31] = in1[7] & in2[7];
    assign P[31] = in1[7] ^ in2[7];
    assign G[32] = in1[6] & in2[6];
    assign P[32] = in1[6] ^ in2[6];
    assign G[33] = in1[5] & in2[5];
    assign P[33] = in1[5] ^ in2[5];
    assign G[34] = in1[4] & in2[4];
    assign P[34] = in1[4] ^ in2[4];
    assign G[35] = in1[3] & in2[3];
    assign P[35] = in1[3] ^ in2[3];
    assign G[36] = in1[2] & in2[2];
    assign P[36] = in1[2] ^ in2[2];
    assign G[37] = in1[1] & in2[1];
    assign P[37] = in1[1] ^ in2[1];
    assign G[38] = in1[0] & in2[0];
    assign P[38] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign cout = G[38] | (P[38] & C[38]);
    assign sum = P ^ C;
endmodule

module CLA_38(output [37:0] sum, output cout, input [37:0] in1, input [37:0] in2);

    wire[37:0] G;
    wire[37:0] C;
    wire[37:0] P;

    assign G[0] = in1[37] & in2[37];
    assign P[0] = in1[37] ^ in2[37];
    assign G[1] = in1[36] & in2[36];
    assign P[1] = in1[36] ^ in2[36];
    assign G[2] = in1[35] & in2[35];
    assign P[2] = in1[35] ^ in2[35];
    assign G[3] = in1[34] & in2[34];
    assign P[3] = in1[34] ^ in2[34];
    assign G[4] = in1[33] & in2[33];
    assign P[4] = in1[33] ^ in2[33];
    assign G[5] = in1[32] & in2[32];
    assign P[5] = in1[32] ^ in2[32];
    assign G[6] = in1[31] & in2[31];
    assign P[6] = in1[31] ^ in2[31];
    assign G[7] = in1[30] & in2[30];
    assign P[7] = in1[30] ^ in2[30];
    assign G[8] = in1[29] & in2[29];
    assign P[8] = in1[29] ^ in2[29];
    assign G[9] = in1[28] & in2[28];
    assign P[9] = in1[28] ^ in2[28];
    assign G[10] = in1[27] & in2[27];
    assign P[10] = in1[27] ^ in2[27];
    assign G[11] = in1[26] & in2[26];
    assign P[11] = in1[26] ^ in2[26];
    assign G[12] = in1[25] & in2[25];
    assign P[12] = in1[25] ^ in2[25];
    assign G[13] = in1[24] & in2[24];
    assign P[13] = in1[24] ^ in2[24];
    assign G[14] = in1[23] & in2[23];
    assign P[14] = in1[23] ^ in2[23];
    assign G[15] = in1[22] & in2[22];
    assign P[15] = in1[22] ^ in2[22];
    assign G[16] = in1[21] & in2[21];
    assign P[16] = in1[21] ^ in2[21];
    assign G[17] = in1[20] & in2[20];
    assign P[17] = in1[20] ^ in2[20];
    assign G[18] = in1[19] & in2[19];
    assign P[18] = in1[19] ^ in2[19];
    assign G[19] = in1[18] & in2[18];
    assign P[19] = in1[18] ^ in2[18];
    assign G[20] = in1[17] & in2[17];
    assign P[20] = in1[17] ^ in2[17];
    assign G[21] = in1[16] & in2[16];
    assign P[21] = in1[16] ^ in2[16];
    assign G[22] = in1[15] & in2[15];
    assign P[22] = in1[15] ^ in2[15];
    assign G[23] = in1[14] & in2[14];
    assign P[23] = in1[14] ^ in2[14];
    assign G[24] = in1[13] & in2[13];
    assign P[24] = in1[13] ^ in2[13];
    assign G[25] = in1[12] & in2[12];
    assign P[25] = in1[12] ^ in2[12];
    assign G[26] = in1[11] & in2[11];
    assign P[26] = in1[11] ^ in2[11];
    assign G[27] = in1[10] & in2[10];
    assign P[27] = in1[10] ^ in2[10];
    assign G[28] = in1[9] & in2[9];
    assign P[28] = in1[9] ^ in2[9];
    assign G[29] = in1[8] & in2[8];
    assign P[29] = in1[8] ^ in2[8];
    assign G[30] = in1[7] & in2[7];
    assign P[30] = in1[7] ^ in2[7];
    assign G[31] = in1[6] & in2[6];
    assign P[31] = in1[6] ^ in2[6];
    assign G[32] = in1[5] & in2[5];
    assign P[32] = in1[5] ^ in2[5];
    assign G[33] = in1[4] & in2[4];
    assign P[33] = in1[4] ^ in2[4];
    assign G[34] = in1[3] & in2[3];
    assign P[34] = in1[3] ^ in2[3];
    assign G[35] = in1[2] & in2[2];
    assign P[35] = in1[2] ^ in2[2];
    assign G[36] = in1[1] & in2[1];
    assign P[36] = in1[1] ^ in2[1];
    assign G[37] = in1[0] & in2[0];
    assign P[37] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign cout = G[37] | (P[37] & C[37]);
    assign sum = P ^ C;
endmodule

module CLA_37(output [36:0] sum, output cout, input [36:0] in1, input [36:0] in2);

    wire[36:0] G;
    wire[36:0] C;
    wire[36:0] P;

    assign G[0] = in1[36] & in2[36];
    assign P[0] = in1[36] ^ in2[36];
    assign G[1] = in1[35] & in2[35];
    assign P[1] = in1[35] ^ in2[35];
    assign G[2] = in1[34] & in2[34];
    assign P[2] = in1[34] ^ in2[34];
    assign G[3] = in1[33] & in2[33];
    assign P[3] = in1[33] ^ in2[33];
    assign G[4] = in1[32] & in2[32];
    assign P[4] = in1[32] ^ in2[32];
    assign G[5] = in1[31] & in2[31];
    assign P[5] = in1[31] ^ in2[31];
    assign G[6] = in1[30] & in2[30];
    assign P[6] = in1[30] ^ in2[30];
    assign G[7] = in1[29] & in2[29];
    assign P[7] = in1[29] ^ in2[29];
    assign G[8] = in1[28] & in2[28];
    assign P[8] = in1[28] ^ in2[28];
    assign G[9] = in1[27] & in2[27];
    assign P[9] = in1[27] ^ in2[27];
    assign G[10] = in1[26] & in2[26];
    assign P[10] = in1[26] ^ in2[26];
    assign G[11] = in1[25] & in2[25];
    assign P[11] = in1[25] ^ in2[25];
    assign G[12] = in1[24] & in2[24];
    assign P[12] = in1[24] ^ in2[24];
    assign G[13] = in1[23] & in2[23];
    assign P[13] = in1[23] ^ in2[23];
    assign G[14] = in1[22] & in2[22];
    assign P[14] = in1[22] ^ in2[22];
    assign G[15] = in1[21] & in2[21];
    assign P[15] = in1[21] ^ in2[21];
    assign G[16] = in1[20] & in2[20];
    assign P[16] = in1[20] ^ in2[20];
    assign G[17] = in1[19] & in2[19];
    assign P[17] = in1[19] ^ in2[19];
    assign G[18] = in1[18] & in2[18];
    assign P[18] = in1[18] ^ in2[18];
    assign G[19] = in1[17] & in2[17];
    assign P[19] = in1[17] ^ in2[17];
    assign G[20] = in1[16] & in2[16];
    assign P[20] = in1[16] ^ in2[16];
    assign G[21] = in1[15] & in2[15];
    assign P[21] = in1[15] ^ in2[15];
    assign G[22] = in1[14] & in2[14];
    assign P[22] = in1[14] ^ in2[14];
    assign G[23] = in1[13] & in2[13];
    assign P[23] = in1[13] ^ in2[13];
    assign G[24] = in1[12] & in2[12];
    assign P[24] = in1[12] ^ in2[12];
    assign G[25] = in1[11] & in2[11];
    assign P[25] = in1[11] ^ in2[11];
    assign G[26] = in1[10] & in2[10];
    assign P[26] = in1[10] ^ in2[10];
    assign G[27] = in1[9] & in2[9];
    assign P[27] = in1[9] ^ in2[9];
    assign G[28] = in1[8] & in2[8];
    assign P[28] = in1[8] ^ in2[8];
    assign G[29] = in1[7] & in2[7];
    assign P[29] = in1[7] ^ in2[7];
    assign G[30] = in1[6] & in2[6];
    assign P[30] = in1[6] ^ in2[6];
    assign G[31] = in1[5] & in2[5];
    assign P[31] = in1[5] ^ in2[5];
    assign G[32] = in1[4] & in2[4];
    assign P[32] = in1[4] ^ in2[4];
    assign G[33] = in1[3] & in2[3];
    assign P[33] = in1[3] ^ in2[3];
    assign G[34] = in1[2] & in2[2];
    assign P[34] = in1[2] ^ in2[2];
    assign G[35] = in1[1] & in2[1];
    assign P[35] = in1[1] ^ in2[1];
    assign G[36] = in1[0] & in2[0];
    assign P[36] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign cout = G[36] | (P[36] & C[36]);
    assign sum = P ^ C;
endmodule

module CLA_36(output [35:0] sum, output cout, input [35:0] in1, input [35:0] in2);

    wire[35:0] G;
    wire[35:0] C;
    wire[35:0] P;

    assign G[0] = in1[35] & in2[35];
    assign P[0] = in1[35] ^ in2[35];
    assign G[1] = in1[34] & in2[34];
    assign P[1] = in1[34] ^ in2[34];
    assign G[2] = in1[33] & in2[33];
    assign P[2] = in1[33] ^ in2[33];
    assign G[3] = in1[32] & in2[32];
    assign P[3] = in1[32] ^ in2[32];
    assign G[4] = in1[31] & in2[31];
    assign P[4] = in1[31] ^ in2[31];
    assign G[5] = in1[30] & in2[30];
    assign P[5] = in1[30] ^ in2[30];
    assign G[6] = in1[29] & in2[29];
    assign P[6] = in1[29] ^ in2[29];
    assign G[7] = in1[28] & in2[28];
    assign P[7] = in1[28] ^ in2[28];
    assign G[8] = in1[27] & in2[27];
    assign P[8] = in1[27] ^ in2[27];
    assign G[9] = in1[26] & in2[26];
    assign P[9] = in1[26] ^ in2[26];
    assign G[10] = in1[25] & in2[25];
    assign P[10] = in1[25] ^ in2[25];
    assign G[11] = in1[24] & in2[24];
    assign P[11] = in1[24] ^ in2[24];
    assign G[12] = in1[23] & in2[23];
    assign P[12] = in1[23] ^ in2[23];
    assign G[13] = in1[22] & in2[22];
    assign P[13] = in1[22] ^ in2[22];
    assign G[14] = in1[21] & in2[21];
    assign P[14] = in1[21] ^ in2[21];
    assign G[15] = in1[20] & in2[20];
    assign P[15] = in1[20] ^ in2[20];
    assign G[16] = in1[19] & in2[19];
    assign P[16] = in1[19] ^ in2[19];
    assign G[17] = in1[18] & in2[18];
    assign P[17] = in1[18] ^ in2[18];
    assign G[18] = in1[17] & in2[17];
    assign P[18] = in1[17] ^ in2[17];
    assign G[19] = in1[16] & in2[16];
    assign P[19] = in1[16] ^ in2[16];
    assign G[20] = in1[15] & in2[15];
    assign P[20] = in1[15] ^ in2[15];
    assign G[21] = in1[14] & in2[14];
    assign P[21] = in1[14] ^ in2[14];
    assign G[22] = in1[13] & in2[13];
    assign P[22] = in1[13] ^ in2[13];
    assign G[23] = in1[12] & in2[12];
    assign P[23] = in1[12] ^ in2[12];
    assign G[24] = in1[11] & in2[11];
    assign P[24] = in1[11] ^ in2[11];
    assign G[25] = in1[10] & in2[10];
    assign P[25] = in1[10] ^ in2[10];
    assign G[26] = in1[9] & in2[9];
    assign P[26] = in1[9] ^ in2[9];
    assign G[27] = in1[8] & in2[8];
    assign P[27] = in1[8] ^ in2[8];
    assign G[28] = in1[7] & in2[7];
    assign P[28] = in1[7] ^ in2[7];
    assign G[29] = in1[6] & in2[6];
    assign P[29] = in1[6] ^ in2[6];
    assign G[30] = in1[5] & in2[5];
    assign P[30] = in1[5] ^ in2[5];
    assign G[31] = in1[4] & in2[4];
    assign P[31] = in1[4] ^ in2[4];
    assign G[32] = in1[3] & in2[3];
    assign P[32] = in1[3] ^ in2[3];
    assign G[33] = in1[2] & in2[2];
    assign P[33] = in1[2] ^ in2[2];
    assign G[34] = in1[1] & in2[1];
    assign P[34] = in1[1] ^ in2[1];
    assign G[35] = in1[0] & in2[0];
    assign P[35] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign cout = G[35] | (P[35] & C[35]);
    assign sum = P ^ C;
endmodule

module CLA_35(output [34:0] sum, output cout, input [34:0] in1, input [34:0] in2);

    wire[34:0] G;
    wire[34:0] C;
    wire[34:0] P;

    assign G[0] = in1[34] & in2[34];
    assign P[0] = in1[34] ^ in2[34];
    assign G[1] = in1[33] & in2[33];
    assign P[1] = in1[33] ^ in2[33];
    assign G[2] = in1[32] & in2[32];
    assign P[2] = in1[32] ^ in2[32];
    assign G[3] = in1[31] & in2[31];
    assign P[3] = in1[31] ^ in2[31];
    assign G[4] = in1[30] & in2[30];
    assign P[4] = in1[30] ^ in2[30];
    assign G[5] = in1[29] & in2[29];
    assign P[5] = in1[29] ^ in2[29];
    assign G[6] = in1[28] & in2[28];
    assign P[6] = in1[28] ^ in2[28];
    assign G[7] = in1[27] & in2[27];
    assign P[7] = in1[27] ^ in2[27];
    assign G[8] = in1[26] & in2[26];
    assign P[8] = in1[26] ^ in2[26];
    assign G[9] = in1[25] & in2[25];
    assign P[9] = in1[25] ^ in2[25];
    assign G[10] = in1[24] & in2[24];
    assign P[10] = in1[24] ^ in2[24];
    assign G[11] = in1[23] & in2[23];
    assign P[11] = in1[23] ^ in2[23];
    assign G[12] = in1[22] & in2[22];
    assign P[12] = in1[22] ^ in2[22];
    assign G[13] = in1[21] & in2[21];
    assign P[13] = in1[21] ^ in2[21];
    assign G[14] = in1[20] & in2[20];
    assign P[14] = in1[20] ^ in2[20];
    assign G[15] = in1[19] & in2[19];
    assign P[15] = in1[19] ^ in2[19];
    assign G[16] = in1[18] & in2[18];
    assign P[16] = in1[18] ^ in2[18];
    assign G[17] = in1[17] & in2[17];
    assign P[17] = in1[17] ^ in2[17];
    assign G[18] = in1[16] & in2[16];
    assign P[18] = in1[16] ^ in2[16];
    assign G[19] = in1[15] & in2[15];
    assign P[19] = in1[15] ^ in2[15];
    assign G[20] = in1[14] & in2[14];
    assign P[20] = in1[14] ^ in2[14];
    assign G[21] = in1[13] & in2[13];
    assign P[21] = in1[13] ^ in2[13];
    assign G[22] = in1[12] & in2[12];
    assign P[22] = in1[12] ^ in2[12];
    assign G[23] = in1[11] & in2[11];
    assign P[23] = in1[11] ^ in2[11];
    assign G[24] = in1[10] & in2[10];
    assign P[24] = in1[10] ^ in2[10];
    assign G[25] = in1[9] & in2[9];
    assign P[25] = in1[9] ^ in2[9];
    assign G[26] = in1[8] & in2[8];
    assign P[26] = in1[8] ^ in2[8];
    assign G[27] = in1[7] & in2[7];
    assign P[27] = in1[7] ^ in2[7];
    assign G[28] = in1[6] & in2[6];
    assign P[28] = in1[6] ^ in2[6];
    assign G[29] = in1[5] & in2[5];
    assign P[29] = in1[5] ^ in2[5];
    assign G[30] = in1[4] & in2[4];
    assign P[30] = in1[4] ^ in2[4];
    assign G[31] = in1[3] & in2[3];
    assign P[31] = in1[3] ^ in2[3];
    assign G[32] = in1[2] & in2[2];
    assign P[32] = in1[2] ^ in2[2];
    assign G[33] = in1[1] & in2[1];
    assign P[33] = in1[1] ^ in2[1];
    assign G[34] = in1[0] & in2[0];
    assign P[34] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign cout = G[34] | (P[34] & C[34]);
    assign sum = P ^ C;
endmodule

module CLA_34(output [33:0] sum, output cout, input [33:0] in1, input [33:0] in2);

    wire[33:0] G;
    wire[33:0] C;
    wire[33:0] P;

    assign G[0] = in1[33] & in2[33];
    assign P[0] = in1[33] ^ in2[33];
    assign G[1] = in1[32] & in2[32];
    assign P[1] = in1[32] ^ in2[32];
    assign G[2] = in1[31] & in2[31];
    assign P[2] = in1[31] ^ in2[31];
    assign G[3] = in1[30] & in2[30];
    assign P[3] = in1[30] ^ in2[30];
    assign G[4] = in1[29] & in2[29];
    assign P[4] = in1[29] ^ in2[29];
    assign G[5] = in1[28] & in2[28];
    assign P[5] = in1[28] ^ in2[28];
    assign G[6] = in1[27] & in2[27];
    assign P[6] = in1[27] ^ in2[27];
    assign G[7] = in1[26] & in2[26];
    assign P[7] = in1[26] ^ in2[26];
    assign G[8] = in1[25] & in2[25];
    assign P[8] = in1[25] ^ in2[25];
    assign G[9] = in1[24] & in2[24];
    assign P[9] = in1[24] ^ in2[24];
    assign G[10] = in1[23] & in2[23];
    assign P[10] = in1[23] ^ in2[23];
    assign G[11] = in1[22] & in2[22];
    assign P[11] = in1[22] ^ in2[22];
    assign G[12] = in1[21] & in2[21];
    assign P[12] = in1[21] ^ in2[21];
    assign G[13] = in1[20] & in2[20];
    assign P[13] = in1[20] ^ in2[20];
    assign G[14] = in1[19] & in2[19];
    assign P[14] = in1[19] ^ in2[19];
    assign G[15] = in1[18] & in2[18];
    assign P[15] = in1[18] ^ in2[18];
    assign G[16] = in1[17] & in2[17];
    assign P[16] = in1[17] ^ in2[17];
    assign G[17] = in1[16] & in2[16];
    assign P[17] = in1[16] ^ in2[16];
    assign G[18] = in1[15] & in2[15];
    assign P[18] = in1[15] ^ in2[15];
    assign G[19] = in1[14] & in2[14];
    assign P[19] = in1[14] ^ in2[14];
    assign G[20] = in1[13] & in2[13];
    assign P[20] = in1[13] ^ in2[13];
    assign G[21] = in1[12] & in2[12];
    assign P[21] = in1[12] ^ in2[12];
    assign G[22] = in1[11] & in2[11];
    assign P[22] = in1[11] ^ in2[11];
    assign G[23] = in1[10] & in2[10];
    assign P[23] = in1[10] ^ in2[10];
    assign G[24] = in1[9] & in2[9];
    assign P[24] = in1[9] ^ in2[9];
    assign G[25] = in1[8] & in2[8];
    assign P[25] = in1[8] ^ in2[8];
    assign G[26] = in1[7] & in2[7];
    assign P[26] = in1[7] ^ in2[7];
    assign G[27] = in1[6] & in2[6];
    assign P[27] = in1[6] ^ in2[6];
    assign G[28] = in1[5] & in2[5];
    assign P[28] = in1[5] ^ in2[5];
    assign G[29] = in1[4] & in2[4];
    assign P[29] = in1[4] ^ in2[4];
    assign G[30] = in1[3] & in2[3];
    assign P[30] = in1[3] ^ in2[3];
    assign G[31] = in1[2] & in2[2];
    assign P[31] = in1[2] ^ in2[2];
    assign G[32] = in1[1] & in2[1];
    assign P[32] = in1[1] ^ in2[1];
    assign G[33] = in1[0] & in2[0];
    assign P[33] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign cout = G[33] | (P[33] & C[33]);
    assign sum = P ^ C;
endmodule

module CLA_33(output [32:0] sum, output cout, input [32:0] in1, input [32:0] in2);

    wire[32:0] G;
    wire[32:0] C;
    wire[32:0] P;

    assign G[0] = in1[32] & in2[32];
    assign P[0] = in1[32] ^ in2[32];
    assign G[1] = in1[31] & in2[31];
    assign P[1] = in1[31] ^ in2[31];
    assign G[2] = in1[30] & in2[30];
    assign P[2] = in1[30] ^ in2[30];
    assign G[3] = in1[29] & in2[29];
    assign P[3] = in1[29] ^ in2[29];
    assign G[4] = in1[28] & in2[28];
    assign P[4] = in1[28] ^ in2[28];
    assign G[5] = in1[27] & in2[27];
    assign P[5] = in1[27] ^ in2[27];
    assign G[6] = in1[26] & in2[26];
    assign P[6] = in1[26] ^ in2[26];
    assign G[7] = in1[25] & in2[25];
    assign P[7] = in1[25] ^ in2[25];
    assign G[8] = in1[24] & in2[24];
    assign P[8] = in1[24] ^ in2[24];
    assign G[9] = in1[23] & in2[23];
    assign P[9] = in1[23] ^ in2[23];
    assign G[10] = in1[22] & in2[22];
    assign P[10] = in1[22] ^ in2[22];
    assign G[11] = in1[21] & in2[21];
    assign P[11] = in1[21] ^ in2[21];
    assign G[12] = in1[20] & in2[20];
    assign P[12] = in1[20] ^ in2[20];
    assign G[13] = in1[19] & in2[19];
    assign P[13] = in1[19] ^ in2[19];
    assign G[14] = in1[18] & in2[18];
    assign P[14] = in1[18] ^ in2[18];
    assign G[15] = in1[17] & in2[17];
    assign P[15] = in1[17] ^ in2[17];
    assign G[16] = in1[16] & in2[16];
    assign P[16] = in1[16] ^ in2[16];
    assign G[17] = in1[15] & in2[15];
    assign P[17] = in1[15] ^ in2[15];
    assign G[18] = in1[14] & in2[14];
    assign P[18] = in1[14] ^ in2[14];
    assign G[19] = in1[13] & in2[13];
    assign P[19] = in1[13] ^ in2[13];
    assign G[20] = in1[12] & in2[12];
    assign P[20] = in1[12] ^ in2[12];
    assign G[21] = in1[11] & in2[11];
    assign P[21] = in1[11] ^ in2[11];
    assign G[22] = in1[10] & in2[10];
    assign P[22] = in1[10] ^ in2[10];
    assign G[23] = in1[9] & in2[9];
    assign P[23] = in1[9] ^ in2[9];
    assign G[24] = in1[8] & in2[8];
    assign P[24] = in1[8] ^ in2[8];
    assign G[25] = in1[7] & in2[7];
    assign P[25] = in1[7] ^ in2[7];
    assign G[26] = in1[6] & in2[6];
    assign P[26] = in1[6] ^ in2[6];
    assign G[27] = in1[5] & in2[5];
    assign P[27] = in1[5] ^ in2[5];
    assign G[28] = in1[4] & in2[4];
    assign P[28] = in1[4] ^ in2[4];
    assign G[29] = in1[3] & in2[3];
    assign P[29] = in1[3] ^ in2[3];
    assign G[30] = in1[2] & in2[2];
    assign P[30] = in1[2] ^ in2[2];
    assign G[31] = in1[1] & in2[1];
    assign P[31] = in1[1] ^ in2[1];
    assign G[32] = in1[0] & in2[0];
    assign P[32] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign cout = G[32] | (P[32] & C[32]);
    assign sum = P ^ C;
endmodule

module CLA_32(output [31:0] sum, output cout, input [31:0] in1, input [31:0] in2);

    wire[31:0] G;
    wire[31:0] C;
    wire[31:0] P;

    assign G[0] = in1[31] & in2[31];
    assign P[0] = in1[31] ^ in2[31];
    assign G[1] = in1[30] & in2[30];
    assign P[1] = in1[30] ^ in2[30];
    assign G[2] = in1[29] & in2[29];
    assign P[2] = in1[29] ^ in2[29];
    assign G[3] = in1[28] & in2[28];
    assign P[3] = in1[28] ^ in2[28];
    assign G[4] = in1[27] & in2[27];
    assign P[4] = in1[27] ^ in2[27];
    assign G[5] = in1[26] & in2[26];
    assign P[5] = in1[26] ^ in2[26];
    assign G[6] = in1[25] & in2[25];
    assign P[6] = in1[25] ^ in2[25];
    assign G[7] = in1[24] & in2[24];
    assign P[7] = in1[24] ^ in2[24];
    assign G[8] = in1[23] & in2[23];
    assign P[8] = in1[23] ^ in2[23];
    assign G[9] = in1[22] & in2[22];
    assign P[9] = in1[22] ^ in2[22];
    assign G[10] = in1[21] & in2[21];
    assign P[10] = in1[21] ^ in2[21];
    assign G[11] = in1[20] & in2[20];
    assign P[11] = in1[20] ^ in2[20];
    assign G[12] = in1[19] & in2[19];
    assign P[12] = in1[19] ^ in2[19];
    assign G[13] = in1[18] & in2[18];
    assign P[13] = in1[18] ^ in2[18];
    assign G[14] = in1[17] & in2[17];
    assign P[14] = in1[17] ^ in2[17];
    assign G[15] = in1[16] & in2[16];
    assign P[15] = in1[16] ^ in2[16];
    assign G[16] = in1[15] & in2[15];
    assign P[16] = in1[15] ^ in2[15];
    assign G[17] = in1[14] & in2[14];
    assign P[17] = in1[14] ^ in2[14];
    assign G[18] = in1[13] & in2[13];
    assign P[18] = in1[13] ^ in2[13];
    assign G[19] = in1[12] & in2[12];
    assign P[19] = in1[12] ^ in2[12];
    assign G[20] = in1[11] & in2[11];
    assign P[20] = in1[11] ^ in2[11];
    assign G[21] = in1[10] & in2[10];
    assign P[21] = in1[10] ^ in2[10];
    assign G[22] = in1[9] & in2[9];
    assign P[22] = in1[9] ^ in2[9];
    assign G[23] = in1[8] & in2[8];
    assign P[23] = in1[8] ^ in2[8];
    assign G[24] = in1[7] & in2[7];
    assign P[24] = in1[7] ^ in2[7];
    assign G[25] = in1[6] & in2[6];
    assign P[25] = in1[6] ^ in2[6];
    assign G[26] = in1[5] & in2[5];
    assign P[26] = in1[5] ^ in2[5];
    assign G[27] = in1[4] & in2[4];
    assign P[27] = in1[4] ^ in2[4];
    assign G[28] = in1[3] & in2[3];
    assign P[28] = in1[3] ^ in2[3];
    assign G[29] = in1[2] & in2[2];
    assign P[29] = in1[2] ^ in2[2];
    assign G[30] = in1[1] & in2[1];
    assign P[30] = in1[1] ^ in2[1];
    assign G[31] = in1[0] & in2[0];
    assign P[31] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign cout = G[31] | (P[31] & C[31]);
    assign sum = P ^ C;
endmodule

module CLA_31(output [30:0] sum, output cout, input [30:0] in1, input [30:0] in2);

    wire[30:0] G;
    wire[30:0] C;
    wire[30:0] P;

    assign G[0] = in1[30] & in2[30];
    assign P[0] = in1[30] ^ in2[30];
    assign G[1] = in1[29] & in2[29];
    assign P[1] = in1[29] ^ in2[29];
    assign G[2] = in1[28] & in2[28];
    assign P[2] = in1[28] ^ in2[28];
    assign G[3] = in1[27] & in2[27];
    assign P[3] = in1[27] ^ in2[27];
    assign G[4] = in1[26] & in2[26];
    assign P[4] = in1[26] ^ in2[26];
    assign G[5] = in1[25] & in2[25];
    assign P[5] = in1[25] ^ in2[25];
    assign G[6] = in1[24] & in2[24];
    assign P[6] = in1[24] ^ in2[24];
    assign G[7] = in1[23] & in2[23];
    assign P[7] = in1[23] ^ in2[23];
    assign G[8] = in1[22] & in2[22];
    assign P[8] = in1[22] ^ in2[22];
    assign G[9] = in1[21] & in2[21];
    assign P[9] = in1[21] ^ in2[21];
    assign G[10] = in1[20] & in2[20];
    assign P[10] = in1[20] ^ in2[20];
    assign G[11] = in1[19] & in2[19];
    assign P[11] = in1[19] ^ in2[19];
    assign G[12] = in1[18] & in2[18];
    assign P[12] = in1[18] ^ in2[18];
    assign G[13] = in1[17] & in2[17];
    assign P[13] = in1[17] ^ in2[17];
    assign G[14] = in1[16] & in2[16];
    assign P[14] = in1[16] ^ in2[16];
    assign G[15] = in1[15] & in2[15];
    assign P[15] = in1[15] ^ in2[15];
    assign G[16] = in1[14] & in2[14];
    assign P[16] = in1[14] ^ in2[14];
    assign G[17] = in1[13] & in2[13];
    assign P[17] = in1[13] ^ in2[13];
    assign G[18] = in1[12] & in2[12];
    assign P[18] = in1[12] ^ in2[12];
    assign G[19] = in1[11] & in2[11];
    assign P[19] = in1[11] ^ in2[11];
    assign G[20] = in1[10] & in2[10];
    assign P[20] = in1[10] ^ in2[10];
    assign G[21] = in1[9] & in2[9];
    assign P[21] = in1[9] ^ in2[9];
    assign G[22] = in1[8] & in2[8];
    assign P[22] = in1[8] ^ in2[8];
    assign G[23] = in1[7] & in2[7];
    assign P[23] = in1[7] ^ in2[7];
    assign G[24] = in1[6] & in2[6];
    assign P[24] = in1[6] ^ in2[6];
    assign G[25] = in1[5] & in2[5];
    assign P[25] = in1[5] ^ in2[5];
    assign G[26] = in1[4] & in2[4];
    assign P[26] = in1[4] ^ in2[4];
    assign G[27] = in1[3] & in2[3];
    assign P[27] = in1[3] ^ in2[3];
    assign G[28] = in1[2] & in2[2];
    assign P[28] = in1[2] ^ in2[2];
    assign G[29] = in1[1] & in2[1];
    assign P[29] = in1[1] ^ in2[1];
    assign G[30] = in1[0] & in2[0];
    assign P[30] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign cout = G[30] | (P[30] & C[30]);
    assign sum = P ^ C;
endmodule

module CLA_30(output [29:0] sum, output cout, input [29:0] in1, input [29:0] in2);

    wire[29:0] G;
    wire[29:0] C;
    wire[29:0] P;

    assign G[0] = in1[29] & in2[29];
    assign P[0] = in1[29] ^ in2[29];
    assign G[1] = in1[28] & in2[28];
    assign P[1] = in1[28] ^ in2[28];
    assign G[2] = in1[27] & in2[27];
    assign P[2] = in1[27] ^ in2[27];
    assign G[3] = in1[26] & in2[26];
    assign P[3] = in1[26] ^ in2[26];
    assign G[4] = in1[25] & in2[25];
    assign P[4] = in1[25] ^ in2[25];
    assign G[5] = in1[24] & in2[24];
    assign P[5] = in1[24] ^ in2[24];
    assign G[6] = in1[23] & in2[23];
    assign P[6] = in1[23] ^ in2[23];
    assign G[7] = in1[22] & in2[22];
    assign P[7] = in1[22] ^ in2[22];
    assign G[8] = in1[21] & in2[21];
    assign P[8] = in1[21] ^ in2[21];
    assign G[9] = in1[20] & in2[20];
    assign P[9] = in1[20] ^ in2[20];
    assign G[10] = in1[19] & in2[19];
    assign P[10] = in1[19] ^ in2[19];
    assign G[11] = in1[18] & in2[18];
    assign P[11] = in1[18] ^ in2[18];
    assign G[12] = in1[17] & in2[17];
    assign P[12] = in1[17] ^ in2[17];
    assign G[13] = in1[16] & in2[16];
    assign P[13] = in1[16] ^ in2[16];
    assign G[14] = in1[15] & in2[15];
    assign P[14] = in1[15] ^ in2[15];
    assign G[15] = in1[14] & in2[14];
    assign P[15] = in1[14] ^ in2[14];
    assign G[16] = in1[13] & in2[13];
    assign P[16] = in1[13] ^ in2[13];
    assign G[17] = in1[12] & in2[12];
    assign P[17] = in1[12] ^ in2[12];
    assign G[18] = in1[11] & in2[11];
    assign P[18] = in1[11] ^ in2[11];
    assign G[19] = in1[10] & in2[10];
    assign P[19] = in1[10] ^ in2[10];
    assign G[20] = in1[9] & in2[9];
    assign P[20] = in1[9] ^ in2[9];
    assign G[21] = in1[8] & in2[8];
    assign P[21] = in1[8] ^ in2[8];
    assign G[22] = in1[7] & in2[7];
    assign P[22] = in1[7] ^ in2[7];
    assign G[23] = in1[6] & in2[6];
    assign P[23] = in1[6] ^ in2[6];
    assign G[24] = in1[5] & in2[5];
    assign P[24] = in1[5] ^ in2[5];
    assign G[25] = in1[4] & in2[4];
    assign P[25] = in1[4] ^ in2[4];
    assign G[26] = in1[3] & in2[3];
    assign P[26] = in1[3] ^ in2[3];
    assign G[27] = in1[2] & in2[2];
    assign P[27] = in1[2] ^ in2[2];
    assign G[28] = in1[1] & in2[1];
    assign P[28] = in1[1] ^ in2[1];
    assign G[29] = in1[0] & in2[0];
    assign P[29] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign cout = G[29] | (P[29] & C[29]);
    assign sum = P ^ C;
endmodule

module CLA_29(output [28:0] sum, output cout, input [28:0] in1, input [28:0] in2);

    wire[28:0] G;
    wire[28:0] C;
    wire[28:0] P;

    assign G[0] = in1[28] & in2[28];
    assign P[0] = in1[28] ^ in2[28];
    assign G[1] = in1[27] & in2[27];
    assign P[1] = in1[27] ^ in2[27];
    assign G[2] = in1[26] & in2[26];
    assign P[2] = in1[26] ^ in2[26];
    assign G[3] = in1[25] & in2[25];
    assign P[3] = in1[25] ^ in2[25];
    assign G[4] = in1[24] & in2[24];
    assign P[4] = in1[24] ^ in2[24];
    assign G[5] = in1[23] & in2[23];
    assign P[5] = in1[23] ^ in2[23];
    assign G[6] = in1[22] & in2[22];
    assign P[6] = in1[22] ^ in2[22];
    assign G[7] = in1[21] & in2[21];
    assign P[7] = in1[21] ^ in2[21];
    assign G[8] = in1[20] & in2[20];
    assign P[8] = in1[20] ^ in2[20];
    assign G[9] = in1[19] & in2[19];
    assign P[9] = in1[19] ^ in2[19];
    assign G[10] = in1[18] & in2[18];
    assign P[10] = in1[18] ^ in2[18];
    assign G[11] = in1[17] & in2[17];
    assign P[11] = in1[17] ^ in2[17];
    assign G[12] = in1[16] & in2[16];
    assign P[12] = in1[16] ^ in2[16];
    assign G[13] = in1[15] & in2[15];
    assign P[13] = in1[15] ^ in2[15];
    assign G[14] = in1[14] & in2[14];
    assign P[14] = in1[14] ^ in2[14];
    assign G[15] = in1[13] & in2[13];
    assign P[15] = in1[13] ^ in2[13];
    assign G[16] = in1[12] & in2[12];
    assign P[16] = in1[12] ^ in2[12];
    assign G[17] = in1[11] & in2[11];
    assign P[17] = in1[11] ^ in2[11];
    assign G[18] = in1[10] & in2[10];
    assign P[18] = in1[10] ^ in2[10];
    assign G[19] = in1[9] & in2[9];
    assign P[19] = in1[9] ^ in2[9];
    assign G[20] = in1[8] & in2[8];
    assign P[20] = in1[8] ^ in2[8];
    assign G[21] = in1[7] & in2[7];
    assign P[21] = in1[7] ^ in2[7];
    assign G[22] = in1[6] & in2[6];
    assign P[22] = in1[6] ^ in2[6];
    assign G[23] = in1[5] & in2[5];
    assign P[23] = in1[5] ^ in2[5];
    assign G[24] = in1[4] & in2[4];
    assign P[24] = in1[4] ^ in2[4];
    assign G[25] = in1[3] & in2[3];
    assign P[25] = in1[3] ^ in2[3];
    assign G[26] = in1[2] & in2[2];
    assign P[26] = in1[2] ^ in2[2];
    assign G[27] = in1[1] & in2[1];
    assign P[27] = in1[1] ^ in2[1];
    assign G[28] = in1[0] & in2[0];
    assign P[28] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign cout = G[28] | (P[28] & C[28]);
    assign sum = P ^ C;
endmodule

module CLA_28(output [27:0] sum, output cout, input [27:0] in1, input [27:0] in2);

    wire[27:0] G;
    wire[27:0] C;
    wire[27:0] P;

    assign G[0] = in1[27] & in2[27];
    assign P[0] = in1[27] ^ in2[27];
    assign G[1] = in1[26] & in2[26];
    assign P[1] = in1[26] ^ in2[26];
    assign G[2] = in1[25] & in2[25];
    assign P[2] = in1[25] ^ in2[25];
    assign G[3] = in1[24] & in2[24];
    assign P[3] = in1[24] ^ in2[24];
    assign G[4] = in1[23] & in2[23];
    assign P[4] = in1[23] ^ in2[23];
    assign G[5] = in1[22] & in2[22];
    assign P[5] = in1[22] ^ in2[22];
    assign G[6] = in1[21] & in2[21];
    assign P[6] = in1[21] ^ in2[21];
    assign G[7] = in1[20] & in2[20];
    assign P[7] = in1[20] ^ in2[20];
    assign G[8] = in1[19] & in2[19];
    assign P[8] = in1[19] ^ in2[19];
    assign G[9] = in1[18] & in2[18];
    assign P[9] = in1[18] ^ in2[18];
    assign G[10] = in1[17] & in2[17];
    assign P[10] = in1[17] ^ in2[17];
    assign G[11] = in1[16] & in2[16];
    assign P[11] = in1[16] ^ in2[16];
    assign G[12] = in1[15] & in2[15];
    assign P[12] = in1[15] ^ in2[15];
    assign G[13] = in1[14] & in2[14];
    assign P[13] = in1[14] ^ in2[14];
    assign G[14] = in1[13] & in2[13];
    assign P[14] = in1[13] ^ in2[13];
    assign G[15] = in1[12] & in2[12];
    assign P[15] = in1[12] ^ in2[12];
    assign G[16] = in1[11] & in2[11];
    assign P[16] = in1[11] ^ in2[11];
    assign G[17] = in1[10] & in2[10];
    assign P[17] = in1[10] ^ in2[10];
    assign G[18] = in1[9] & in2[9];
    assign P[18] = in1[9] ^ in2[9];
    assign G[19] = in1[8] & in2[8];
    assign P[19] = in1[8] ^ in2[8];
    assign G[20] = in1[7] & in2[7];
    assign P[20] = in1[7] ^ in2[7];
    assign G[21] = in1[6] & in2[6];
    assign P[21] = in1[6] ^ in2[6];
    assign G[22] = in1[5] & in2[5];
    assign P[22] = in1[5] ^ in2[5];
    assign G[23] = in1[4] & in2[4];
    assign P[23] = in1[4] ^ in2[4];
    assign G[24] = in1[3] & in2[3];
    assign P[24] = in1[3] ^ in2[3];
    assign G[25] = in1[2] & in2[2];
    assign P[25] = in1[2] ^ in2[2];
    assign G[26] = in1[1] & in2[1];
    assign P[26] = in1[1] ^ in2[1];
    assign G[27] = in1[0] & in2[0];
    assign P[27] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign cout = G[27] | (P[27] & C[27]);
    assign sum = P ^ C;
endmodule

module CLA_27(output [26:0] sum, output cout, input [26:0] in1, input [26:0] in2);

    wire[26:0] G;
    wire[26:0] C;
    wire[26:0] P;

    assign G[0] = in1[26] & in2[26];
    assign P[0] = in1[26] ^ in2[26];
    assign G[1] = in1[25] & in2[25];
    assign P[1] = in1[25] ^ in2[25];
    assign G[2] = in1[24] & in2[24];
    assign P[2] = in1[24] ^ in2[24];
    assign G[3] = in1[23] & in2[23];
    assign P[3] = in1[23] ^ in2[23];
    assign G[4] = in1[22] & in2[22];
    assign P[4] = in1[22] ^ in2[22];
    assign G[5] = in1[21] & in2[21];
    assign P[5] = in1[21] ^ in2[21];
    assign G[6] = in1[20] & in2[20];
    assign P[6] = in1[20] ^ in2[20];
    assign G[7] = in1[19] & in2[19];
    assign P[7] = in1[19] ^ in2[19];
    assign G[8] = in1[18] & in2[18];
    assign P[8] = in1[18] ^ in2[18];
    assign G[9] = in1[17] & in2[17];
    assign P[9] = in1[17] ^ in2[17];
    assign G[10] = in1[16] & in2[16];
    assign P[10] = in1[16] ^ in2[16];
    assign G[11] = in1[15] & in2[15];
    assign P[11] = in1[15] ^ in2[15];
    assign G[12] = in1[14] & in2[14];
    assign P[12] = in1[14] ^ in2[14];
    assign G[13] = in1[13] & in2[13];
    assign P[13] = in1[13] ^ in2[13];
    assign G[14] = in1[12] & in2[12];
    assign P[14] = in1[12] ^ in2[12];
    assign G[15] = in1[11] & in2[11];
    assign P[15] = in1[11] ^ in2[11];
    assign G[16] = in1[10] & in2[10];
    assign P[16] = in1[10] ^ in2[10];
    assign G[17] = in1[9] & in2[9];
    assign P[17] = in1[9] ^ in2[9];
    assign G[18] = in1[8] & in2[8];
    assign P[18] = in1[8] ^ in2[8];
    assign G[19] = in1[7] & in2[7];
    assign P[19] = in1[7] ^ in2[7];
    assign G[20] = in1[6] & in2[6];
    assign P[20] = in1[6] ^ in2[6];
    assign G[21] = in1[5] & in2[5];
    assign P[21] = in1[5] ^ in2[5];
    assign G[22] = in1[4] & in2[4];
    assign P[22] = in1[4] ^ in2[4];
    assign G[23] = in1[3] & in2[3];
    assign P[23] = in1[3] ^ in2[3];
    assign G[24] = in1[2] & in2[2];
    assign P[24] = in1[2] ^ in2[2];
    assign G[25] = in1[1] & in2[1];
    assign P[25] = in1[1] ^ in2[1];
    assign G[26] = in1[0] & in2[0];
    assign P[26] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign cout = G[26] | (P[26] & C[26]);
    assign sum = P ^ C;
endmodule

module CLA_26(output [25:0] sum, output cout, input [25:0] in1, input [25:0] in2);

    wire[25:0] G;
    wire[25:0] C;
    wire[25:0] P;

    assign G[0] = in1[25] & in2[25];
    assign P[0] = in1[25] ^ in2[25];
    assign G[1] = in1[24] & in2[24];
    assign P[1] = in1[24] ^ in2[24];
    assign G[2] = in1[23] & in2[23];
    assign P[2] = in1[23] ^ in2[23];
    assign G[3] = in1[22] & in2[22];
    assign P[3] = in1[22] ^ in2[22];
    assign G[4] = in1[21] & in2[21];
    assign P[4] = in1[21] ^ in2[21];
    assign G[5] = in1[20] & in2[20];
    assign P[5] = in1[20] ^ in2[20];
    assign G[6] = in1[19] & in2[19];
    assign P[6] = in1[19] ^ in2[19];
    assign G[7] = in1[18] & in2[18];
    assign P[7] = in1[18] ^ in2[18];
    assign G[8] = in1[17] & in2[17];
    assign P[8] = in1[17] ^ in2[17];
    assign G[9] = in1[16] & in2[16];
    assign P[9] = in1[16] ^ in2[16];
    assign G[10] = in1[15] & in2[15];
    assign P[10] = in1[15] ^ in2[15];
    assign G[11] = in1[14] & in2[14];
    assign P[11] = in1[14] ^ in2[14];
    assign G[12] = in1[13] & in2[13];
    assign P[12] = in1[13] ^ in2[13];
    assign G[13] = in1[12] & in2[12];
    assign P[13] = in1[12] ^ in2[12];
    assign G[14] = in1[11] & in2[11];
    assign P[14] = in1[11] ^ in2[11];
    assign G[15] = in1[10] & in2[10];
    assign P[15] = in1[10] ^ in2[10];
    assign G[16] = in1[9] & in2[9];
    assign P[16] = in1[9] ^ in2[9];
    assign G[17] = in1[8] & in2[8];
    assign P[17] = in1[8] ^ in2[8];
    assign G[18] = in1[7] & in2[7];
    assign P[18] = in1[7] ^ in2[7];
    assign G[19] = in1[6] & in2[6];
    assign P[19] = in1[6] ^ in2[6];
    assign G[20] = in1[5] & in2[5];
    assign P[20] = in1[5] ^ in2[5];
    assign G[21] = in1[4] & in2[4];
    assign P[21] = in1[4] ^ in2[4];
    assign G[22] = in1[3] & in2[3];
    assign P[22] = in1[3] ^ in2[3];
    assign G[23] = in1[2] & in2[2];
    assign P[23] = in1[2] ^ in2[2];
    assign G[24] = in1[1] & in2[1];
    assign P[24] = in1[1] ^ in2[1];
    assign G[25] = in1[0] & in2[0];
    assign P[25] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign cout = G[25] | (P[25] & C[25]);
    assign sum = P ^ C;
endmodule

module CLA_25(output [24:0] sum, output cout, input [24:0] in1, input [24:0] in2);

    wire[24:0] G;
    wire[24:0] C;
    wire[24:0] P;

    assign G[0] = in1[24] & in2[24];
    assign P[0] = in1[24] ^ in2[24];
    assign G[1] = in1[23] & in2[23];
    assign P[1] = in1[23] ^ in2[23];
    assign G[2] = in1[22] & in2[22];
    assign P[2] = in1[22] ^ in2[22];
    assign G[3] = in1[21] & in2[21];
    assign P[3] = in1[21] ^ in2[21];
    assign G[4] = in1[20] & in2[20];
    assign P[4] = in1[20] ^ in2[20];
    assign G[5] = in1[19] & in2[19];
    assign P[5] = in1[19] ^ in2[19];
    assign G[6] = in1[18] & in2[18];
    assign P[6] = in1[18] ^ in2[18];
    assign G[7] = in1[17] & in2[17];
    assign P[7] = in1[17] ^ in2[17];
    assign G[8] = in1[16] & in2[16];
    assign P[8] = in1[16] ^ in2[16];
    assign G[9] = in1[15] & in2[15];
    assign P[9] = in1[15] ^ in2[15];
    assign G[10] = in1[14] & in2[14];
    assign P[10] = in1[14] ^ in2[14];
    assign G[11] = in1[13] & in2[13];
    assign P[11] = in1[13] ^ in2[13];
    assign G[12] = in1[12] & in2[12];
    assign P[12] = in1[12] ^ in2[12];
    assign G[13] = in1[11] & in2[11];
    assign P[13] = in1[11] ^ in2[11];
    assign G[14] = in1[10] & in2[10];
    assign P[14] = in1[10] ^ in2[10];
    assign G[15] = in1[9] & in2[9];
    assign P[15] = in1[9] ^ in2[9];
    assign G[16] = in1[8] & in2[8];
    assign P[16] = in1[8] ^ in2[8];
    assign G[17] = in1[7] & in2[7];
    assign P[17] = in1[7] ^ in2[7];
    assign G[18] = in1[6] & in2[6];
    assign P[18] = in1[6] ^ in2[6];
    assign G[19] = in1[5] & in2[5];
    assign P[19] = in1[5] ^ in2[5];
    assign G[20] = in1[4] & in2[4];
    assign P[20] = in1[4] ^ in2[4];
    assign G[21] = in1[3] & in2[3];
    assign P[21] = in1[3] ^ in2[3];
    assign G[22] = in1[2] & in2[2];
    assign P[22] = in1[2] ^ in2[2];
    assign G[23] = in1[1] & in2[1];
    assign P[23] = in1[1] ^ in2[1];
    assign G[24] = in1[0] & in2[0];
    assign P[24] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign cout = G[24] | (P[24] & C[24]);
    assign sum = P ^ C;
endmodule

module CLA_24(output [23:0] sum, output cout, input [23:0] in1, input [23:0] in2);

    wire[23:0] G;
    wire[23:0] C;
    wire[23:0] P;

    assign G[0] = in1[23] & in2[23];
    assign P[0] = in1[23] ^ in2[23];
    assign G[1] = in1[22] & in2[22];
    assign P[1] = in1[22] ^ in2[22];
    assign G[2] = in1[21] & in2[21];
    assign P[2] = in1[21] ^ in2[21];
    assign G[3] = in1[20] & in2[20];
    assign P[3] = in1[20] ^ in2[20];
    assign G[4] = in1[19] & in2[19];
    assign P[4] = in1[19] ^ in2[19];
    assign G[5] = in1[18] & in2[18];
    assign P[5] = in1[18] ^ in2[18];
    assign G[6] = in1[17] & in2[17];
    assign P[6] = in1[17] ^ in2[17];
    assign G[7] = in1[16] & in2[16];
    assign P[7] = in1[16] ^ in2[16];
    assign G[8] = in1[15] & in2[15];
    assign P[8] = in1[15] ^ in2[15];
    assign G[9] = in1[14] & in2[14];
    assign P[9] = in1[14] ^ in2[14];
    assign G[10] = in1[13] & in2[13];
    assign P[10] = in1[13] ^ in2[13];
    assign G[11] = in1[12] & in2[12];
    assign P[11] = in1[12] ^ in2[12];
    assign G[12] = in1[11] & in2[11];
    assign P[12] = in1[11] ^ in2[11];
    assign G[13] = in1[10] & in2[10];
    assign P[13] = in1[10] ^ in2[10];
    assign G[14] = in1[9] & in2[9];
    assign P[14] = in1[9] ^ in2[9];
    assign G[15] = in1[8] & in2[8];
    assign P[15] = in1[8] ^ in2[8];
    assign G[16] = in1[7] & in2[7];
    assign P[16] = in1[7] ^ in2[7];
    assign G[17] = in1[6] & in2[6];
    assign P[17] = in1[6] ^ in2[6];
    assign G[18] = in1[5] & in2[5];
    assign P[18] = in1[5] ^ in2[5];
    assign G[19] = in1[4] & in2[4];
    assign P[19] = in1[4] ^ in2[4];
    assign G[20] = in1[3] & in2[3];
    assign P[20] = in1[3] ^ in2[3];
    assign G[21] = in1[2] & in2[2];
    assign P[21] = in1[2] ^ in2[2];
    assign G[22] = in1[1] & in2[1];
    assign P[22] = in1[1] ^ in2[1];
    assign G[23] = in1[0] & in2[0];
    assign P[23] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign cout = G[23] | (P[23] & C[23]);
    assign sum = P ^ C;
endmodule

module CLA_23(output [22:0] sum, output cout, input [22:0] in1, input [22:0] in2);

    wire[22:0] G;
    wire[22:0] C;
    wire[22:0] P;

    assign G[0] = in1[22] & in2[22];
    assign P[0] = in1[22] ^ in2[22];
    assign G[1] = in1[21] & in2[21];
    assign P[1] = in1[21] ^ in2[21];
    assign G[2] = in1[20] & in2[20];
    assign P[2] = in1[20] ^ in2[20];
    assign G[3] = in1[19] & in2[19];
    assign P[3] = in1[19] ^ in2[19];
    assign G[4] = in1[18] & in2[18];
    assign P[4] = in1[18] ^ in2[18];
    assign G[5] = in1[17] & in2[17];
    assign P[5] = in1[17] ^ in2[17];
    assign G[6] = in1[16] & in2[16];
    assign P[6] = in1[16] ^ in2[16];
    assign G[7] = in1[15] & in2[15];
    assign P[7] = in1[15] ^ in2[15];
    assign G[8] = in1[14] & in2[14];
    assign P[8] = in1[14] ^ in2[14];
    assign G[9] = in1[13] & in2[13];
    assign P[9] = in1[13] ^ in2[13];
    assign G[10] = in1[12] & in2[12];
    assign P[10] = in1[12] ^ in2[12];
    assign G[11] = in1[11] & in2[11];
    assign P[11] = in1[11] ^ in2[11];
    assign G[12] = in1[10] & in2[10];
    assign P[12] = in1[10] ^ in2[10];
    assign G[13] = in1[9] & in2[9];
    assign P[13] = in1[9] ^ in2[9];
    assign G[14] = in1[8] & in2[8];
    assign P[14] = in1[8] ^ in2[8];
    assign G[15] = in1[7] & in2[7];
    assign P[15] = in1[7] ^ in2[7];
    assign G[16] = in1[6] & in2[6];
    assign P[16] = in1[6] ^ in2[6];
    assign G[17] = in1[5] & in2[5];
    assign P[17] = in1[5] ^ in2[5];
    assign G[18] = in1[4] & in2[4];
    assign P[18] = in1[4] ^ in2[4];
    assign G[19] = in1[3] & in2[3];
    assign P[19] = in1[3] ^ in2[3];
    assign G[20] = in1[2] & in2[2];
    assign P[20] = in1[2] ^ in2[2];
    assign G[21] = in1[1] & in2[1];
    assign P[21] = in1[1] ^ in2[1];
    assign G[22] = in1[0] & in2[0];
    assign P[22] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign cout = G[22] | (P[22] & C[22]);
    assign sum = P ^ C;
endmodule

module CLA_22(output [21:0] sum, output cout, input [21:0] in1, input [21:0] in2);

    wire[21:0] G;
    wire[21:0] C;
    wire[21:0] P;

    assign G[0] = in1[21] & in2[21];
    assign P[0] = in1[21] ^ in2[21];
    assign G[1] = in1[20] & in2[20];
    assign P[1] = in1[20] ^ in2[20];
    assign G[2] = in1[19] & in2[19];
    assign P[2] = in1[19] ^ in2[19];
    assign G[3] = in1[18] & in2[18];
    assign P[3] = in1[18] ^ in2[18];
    assign G[4] = in1[17] & in2[17];
    assign P[4] = in1[17] ^ in2[17];
    assign G[5] = in1[16] & in2[16];
    assign P[5] = in1[16] ^ in2[16];
    assign G[6] = in1[15] & in2[15];
    assign P[6] = in1[15] ^ in2[15];
    assign G[7] = in1[14] & in2[14];
    assign P[7] = in1[14] ^ in2[14];
    assign G[8] = in1[13] & in2[13];
    assign P[8] = in1[13] ^ in2[13];
    assign G[9] = in1[12] & in2[12];
    assign P[9] = in1[12] ^ in2[12];
    assign G[10] = in1[11] & in2[11];
    assign P[10] = in1[11] ^ in2[11];
    assign G[11] = in1[10] & in2[10];
    assign P[11] = in1[10] ^ in2[10];
    assign G[12] = in1[9] & in2[9];
    assign P[12] = in1[9] ^ in2[9];
    assign G[13] = in1[8] & in2[8];
    assign P[13] = in1[8] ^ in2[8];
    assign G[14] = in1[7] & in2[7];
    assign P[14] = in1[7] ^ in2[7];
    assign G[15] = in1[6] & in2[6];
    assign P[15] = in1[6] ^ in2[6];
    assign G[16] = in1[5] & in2[5];
    assign P[16] = in1[5] ^ in2[5];
    assign G[17] = in1[4] & in2[4];
    assign P[17] = in1[4] ^ in2[4];
    assign G[18] = in1[3] & in2[3];
    assign P[18] = in1[3] ^ in2[3];
    assign G[19] = in1[2] & in2[2];
    assign P[19] = in1[2] ^ in2[2];
    assign G[20] = in1[1] & in2[1];
    assign P[20] = in1[1] ^ in2[1];
    assign G[21] = in1[0] & in2[0];
    assign P[21] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign cout = G[21] | (P[21] & C[21]);
    assign sum = P ^ C;
endmodule

module CLA_21(output [20:0] sum, output cout, input [20:0] in1, input [20:0] in2);

    wire[20:0] G;
    wire[20:0] C;
    wire[20:0] P;

    assign G[0] = in1[20] & in2[20];
    assign P[0] = in1[20] ^ in2[20];
    assign G[1] = in1[19] & in2[19];
    assign P[1] = in1[19] ^ in2[19];
    assign G[2] = in1[18] & in2[18];
    assign P[2] = in1[18] ^ in2[18];
    assign G[3] = in1[17] & in2[17];
    assign P[3] = in1[17] ^ in2[17];
    assign G[4] = in1[16] & in2[16];
    assign P[4] = in1[16] ^ in2[16];
    assign G[5] = in1[15] & in2[15];
    assign P[5] = in1[15] ^ in2[15];
    assign G[6] = in1[14] & in2[14];
    assign P[6] = in1[14] ^ in2[14];
    assign G[7] = in1[13] & in2[13];
    assign P[7] = in1[13] ^ in2[13];
    assign G[8] = in1[12] & in2[12];
    assign P[8] = in1[12] ^ in2[12];
    assign G[9] = in1[11] & in2[11];
    assign P[9] = in1[11] ^ in2[11];
    assign G[10] = in1[10] & in2[10];
    assign P[10] = in1[10] ^ in2[10];
    assign G[11] = in1[9] & in2[9];
    assign P[11] = in1[9] ^ in2[9];
    assign G[12] = in1[8] & in2[8];
    assign P[12] = in1[8] ^ in2[8];
    assign G[13] = in1[7] & in2[7];
    assign P[13] = in1[7] ^ in2[7];
    assign G[14] = in1[6] & in2[6];
    assign P[14] = in1[6] ^ in2[6];
    assign G[15] = in1[5] & in2[5];
    assign P[15] = in1[5] ^ in2[5];
    assign G[16] = in1[4] & in2[4];
    assign P[16] = in1[4] ^ in2[4];
    assign G[17] = in1[3] & in2[3];
    assign P[17] = in1[3] ^ in2[3];
    assign G[18] = in1[2] & in2[2];
    assign P[18] = in1[2] ^ in2[2];
    assign G[19] = in1[1] & in2[1];
    assign P[19] = in1[1] ^ in2[1];
    assign G[20] = in1[0] & in2[0];
    assign P[20] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign cout = G[20] | (P[20] & C[20]);
    assign sum = P ^ C;
endmodule

module CLA_20(output [19:0] sum, output cout, input [19:0] in1, input [19:0] in2);

    wire[19:0] G;
    wire[19:0] C;
    wire[19:0] P;

    assign G[0] = in1[19] & in2[19];
    assign P[0] = in1[19] ^ in2[19];
    assign G[1] = in1[18] & in2[18];
    assign P[1] = in1[18] ^ in2[18];
    assign G[2] = in1[17] & in2[17];
    assign P[2] = in1[17] ^ in2[17];
    assign G[3] = in1[16] & in2[16];
    assign P[3] = in1[16] ^ in2[16];
    assign G[4] = in1[15] & in2[15];
    assign P[4] = in1[15] ^ in2[15];
    assign G[5] = in1[14] & in2[14];
    assign P[5] = in1[14] ^ in2[14];
    assign G[6] = in1[13] & in2[13];
    assign P[6] = in1[13] ^ in2[13];
    assign G[7] = in1[12] & in2[12];
    assign P[7] = in1[12] ^ in2[12];
    assign G[8] = in1[11] & in2[11];
    assign P[8] = in1[11] ^ in2[11];
    assign G[9] = in1[10] & in2[10];
    assign P[9] = in1[10] ^ in2[10];
    assign G[10] = in1[9] & in2[9];
    assign P[10] = in1[9] ^ in2[9];
    assign G[11] = in1[8] & in2[8];
    assign P[11] = in1[8] ^ in2[8];
    assign G[12] = in1[7] & in2[7];
    assign P[12] = in1[7] ^ in2[7];
    assign G[13] = in1[6] & in2[6];
    assign P[13] = in1[6] ^ in2[6];
    assign G[14] = in1[5] & in2[5];
    assign P[14] = in1[5] ^ in2[5];
    assign G[15] = in1[4] & in2[4];
    assign P[15] = in1[4] ^ in2[4];
    assign G[16] = in1[3] & in2[3];
    assign P[16] = in1[3] ^ in2[3];
    assign G[17] = in1[2] & in2[2];
    assign P[17] = in1[2] ^ in2[2];
    assign G[18] = in1[1] & in2[1];
    assign P[18] = in1[1] ^ in2[1];
    assign G[19] = in1[0] & in2[0];
    assign P[19] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign cout = G[19] | (P[19] & C[19]);
    assign sum = P ^ C;
endmodule

module CLA_19(output [18:0] sum, output cout, input [18:0] in1, input [18:0] in2);

    wire[18:0] G;
    wire[18:0] C;
    wire[18:0] P;

    assign G[0] = in1[18] & in2[18];
    assign P[0] = in1[18] ^ in2[18];
    assign G[1] = in1[17] & in2[17];
    assign P[1] = in1[17] ^ in2[17];
    assign G[2] = in1[16] & in2[16];
    assign P[2] = in1[16] ^ in2[16];
    assign G[3] = in1[15] & in2[15];
    assign P[3] = in1[15] ^ in2[15];
    assign G[4] = in1[14] & in2[14];
    assign P[4] = in1[14] ^ in2[14];
    assign G[5] = in1[13] & in2[13];
    assign P[5] = in1[13] ^ in2[13];
    assign G[6] = in1[12] & in2[12];
    assign P[6] = in1[12] ^ in2[12];
    assign G[7] = in1[11] & in2[11];
    assign P[7] = in1[11] ^ in2[11];
    assign G[8] = in1[10] & in2[10];
    assign P[8] = in1[10] ^ in2[10];
    assign G[9] = in1[9] & in2[9];
    assign P[9] = in1[9] ^ in2[9];
    assign G[10] = in1[8] & in2[8];
    assign P[10] = in1[8] ^ in2[8];
    assign G[11] = in1[7] & in2[7];
    assign P[11] = in1[7] ^ in2[7];
    assign G[12] = in1[6] & in2[6];
    assign P[12] = in1[6] ^ in2[6];
    assign G[13] = in1[5] & in2[5];
    assign P[13] = in1[5] ^ in2[5];
    assign G[14] = in1[4] & in2[4];
    assign P[14] = in1[4] ^ in2[4];
    assign G[15] = in1[3] & in2[3];
    assign P[15] = in1[3] ^ in2[3];
    assign G[16] = in1[2] & in2[2];
    assign P[16] = in1[2] ^ in2[2];
    assign G[17] = in1[1] & in2[1];
    assign P[17] = in1[1] ^ in2[1];
    assign G[18] = in1[0] & in2[0];
    assign P[18] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign cout = G[18] | (P[18] & C[18]);
    assign sum = P ^ C;
endmodule

module CLA_18(output [17:0] sum, output cout, input [17:0] in1, input [17:0] in2);

    wire[17:0] G;
    wire[17:0] C;
    wire[17:0] P;

    assign G[0] = in1[17] & in2[17];
    assign P[0] = in1[17] ^ in2[17];
    assign G[1] = in1[16] & in2[16];
    assign P[1] = in1[16] ^ in2[16];
    assign G[2] = in1[15] & in2[15];
    assign P[2] = in1[15] ^ in2[15];
    assign G[3] = in1[14] & in2[14];
    assign P[3] = in1[14] ^ in2[14];
    assign G[4] = in1[13] & in2[13];
    assign P[4] = in1[13] ^ in2[13];
    assign G[5] = in1[12] & in2[12];
    assign P[5] = in1[12] ^ in2[12];
    assign G[6] = in1[11] & in2[11];
    assign P[6] = in1[11] ^ in2[11];
    assign G[7] = in1[10] & in2[10];
    assign P[7] = in1[10] ^ in2[10];
    assign G[8] = in1[9] & in2[9];
    assign P[8] = in1[9] ^ in2[9];
    assign G[9] = in1[8] & in2[8];
    assign P[9] = in1[8] ^ in2[8];
    assign G[10] = in1[7] & in2[7];
    assign P[10] = in1[7] ^ in2[7];
    assign G[11] = in1[6] & in2[6];
    assign P[11] = in1[6] ^ in2[6];
    assign G[12] = in1[5] & in2[5];
    assign P[12] = in1[5] ^ in2[5];
    assign G[13] = in1[4] & in2[4];
    assign P[13] = in1[4] ^ in2[4];
    assign G[14] = in1[3] & in2[3];
    assign P[14] = in1[3] ^ in2[3];
    assign G[15] = in1[2] & in2[2];
    assign P[15] = in1[2] ^ in2[2];
    assign G[16] = in1[1] & in2[1];
    assign P[16] = in1[1] ^ in2[1];
    assign G[17] = in1[0] & in2[0];
    assign P[17] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign cout = G[17] | (P[17] & C[17]);
    assign sum = P ^ C;
endmodule

module CLA_17(output [16:0] sum, output cout, input [16:0] in1, input [16:0] in2);

    wire[16:0] G;
    wire[16:0] C;
    wire[16:0] P;

    assign G[0] = in1[16] & in2[16];
    assign P[0] = in1[16] ^ in2[16];
    assign G[1] = in1[15] & in2[15];
    assign P[1] = in1[15] ^ in2[15];
    assign G[2] = in1[14] & in2[14];
    assign P[2] = in1[14] ^ in2[14];
    assign G[3] = in1[13] & in2[13];
    assign P[3] = in1[13] ^ in2[13];
    assign G[4] = in1[12] & in2[12];
    assign P[4] = in1[12] ^ in2[12];
    assign G[5] = in1[11] & in2[11];
    assign P[5] = in1[11] ^ in2[11];
    assign G[6] = in1[10] & in2[10];
    assign P[6] = in1[10] ^ in2[10];
    assign G[7] = in1[9] & in2[9];
    assign P[7] = in1[9] ^ in2[9];
    assign G[8] = in1[8] & in2[8];
    assign P[8] = in1[8] ^ in2[8];
    assign G[9] = in1[7] & in2[7];
    assign P[9] = in1[7] ^ in2[7];
    assign G[10] = in1[6] & in2[6];
    assign P[10] = in1[6] ^ in2[6];
    assign G[11] = in1[5] & in2[5];
    assign P[11] = in1[5] ^ in2[5];
    assign G[12] = in1[4] & in2[4];
    assign P[12] = in1[4] ^ in2[4];
    assign G[13] = in1[3] & in2[3];
    assign P[13] = in1[3] ^ in2[3];
    assign G[14] = in1[2] & in2[2];
    assign P[14] = in1[2] ^ in2[2];
    assign G[15] = in1[1] & in2[1];
    assign P[15] = in1[1] ^ in2[1];
    assign G[16] = in1[0] & in2[0];
    assign P[16] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign cout = G[16] | (P[16] & C[16]);
    assign sum = P ^ C;
endmodule

module CLA_16(output [15:0] sum, output cout, input [15:0] in1, input [15:0] in2);

    wire[15:0] G;
    wire[15:0] C;
    wire[15:0] P;

    assign G[0] = in1[15] & in2[15];
    assign P[0] = in1[15] ^ in2[15];
    assign G[1] = in1[14] & in2[14];
    assign P[1] = in1[14] ^ in2[14];
    assign G[2] = in1[13] & in2[13];
    assign P[2] = in1[13] ^ in2[13];
    assign G[3] = in1[12] & in2[12];
    assign P[3] = in1[12] ^ in2[12];
    assign G[4] = in1[11] & in2[11];
    assign P[4] = in1[11] ^ in2[11];
    assign G[5] = in1[10] & in2[10];
    assign P[5] = in1[10] ^ in2[10];
    assign G[6] = in1[9] & in2[9];
    assign P[6] = in1[9] ^ in2[9];
    assign G[7] = in1[8] & in2[8];
    assign P[7] = in1[8] ^ in2[8];
    assign G[8] = in1[7] & in2[7];
    assign P[8] = in1[7] ^ in2[7];
    assign G[9] = in1[6] & in2[6];
    assign P[9] = in1[6] ^ in2[6];
    assign G[10] = in1[5] & in2[5];
    assign P[10] = in1[5] ^ in2[5];
    assign G[11] = in1[4] & in2[4];
    assign P[11] = in1[4] ^ in2[4];
    assign G[12] = in1[3] & in2[3];
    assign P[12] = in1[3] ^ in2[3];
    assign G[13] = in1[2] & in2[2];
    assign P[13] = in1[2] ^ in2[2];
    assign G[14] = in1[1] & in2[1];
    assign P[14] = in1[1] ^ in2[1];
    assign G[15] = in1[0] & in2[0];
    assign P[15] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign cout = G[15] | (P[15] & C[15]);
    assign sum = P ^ C;
endmodule

module CLA_15(output [14:0] sum, output cout, input [14:0] in1, input [14:0] in2);

    wire[14:0] G;
    wire[14:0] C;
    wire[14:0] P;

    assign G[0] = in1[14] & in2[14];
    assign P[0] = in1[14] ^ in2[14];
    assign G[1] = in1[13] & in2[13];
    assign P[1] = in1[13] ^ in2[13];
    assign G[2] = in1[12] & in2[12];
    assign P[2] = in1[12] ^ in2[12];
    assign G[3] = in1[11] & in2[11];
    assign P[3] = in1[11] ^ in2[11];
    assign G[4] = in1[10] & in2[10];
    assign P[4] = in1[10] ^ in2[10];
    assign G[5] = in1[9] & in2[9];
    assign P[5] = in1[9] ^ in2[9];
    assign G[6] = in1[8] & in2[8];
    assign P[6] = in1[8] ^ in2[8];
    assign G[7] = in1[7] & in2[7];
    assign P[7] = in1[7] ^ in2[7];
    assign G[8] = in1[6] & in2[6];
    assign P[8] = in1[6] ^ in2[6];
    assign G[9] = in1[5] & in2[5];
    assign P[9] = in1[5] ^ in2[5];
    assign G[10] = in1[4] & in2[4];
    assign P[10] = in1[4] ^ in2[4];
    assign G[11] = in1[3] & in2[3];
    assign P[11] = in1[3] ^ in2[3];
    assign G[12] = in1[2] & in2[2];
    assign P[12] = in1[2] ^ in2[2];
    assign G[13] = in1[1] & in2[1];
    assign P[13] = in1[1] ^ in2[1];
    assign G[14] = in1[0] & in2[0];
    assign P[14] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign cout = G[14] | (P[14] & C[14]);
    assign sum = P ^ C;
endmodule

module CLA_14(output [13:0] sum, output cout, input [13:0] in1, input [13:0] in2);

    wire[13:0] G;
    wire[13:0] C;
    wire[13:0] P;

    assign G[0] = in1[13] & in2[13];
    assign P[0] = in1[13] ^ in2[13];
    assign G[1] = in1[12] & in2[12];
    assign P[1] = in1[12] ^ in2[12];
    assign G[2] = in1[11] & in2[11];
    assign P[2] = in1[11] ^ in2[11];
    assign G[3] = in1[10] & in2[10];
    assign P[3] = in1[10] ^ in2[10];
    assign G[4] = in1[9] & in2[9];
    assign P[4] = in1[9] ^ in2[9];
    assign G[5] = in1[8] & in2[8];
    assign P[5] = in1[8] ^ in2[8];
    assign G[6] = in1[7] & in2[7];
    assign P[6] = in1[7] ^ in2[7];
    assign G[7] = in1[6] & in2[6];
    assign P[7] = in1[6] ^ in2[6];
    assign G[8] = in1[5] & in2[5];
    assign P[8] = in1[5] ^ in2[5];
    assign G[9] = in1[4] & in2[4];
    assign P[9] = in1[4] ^ in2[4];
    assign G[10] = in1[3] & in2[3];
    assign P[10] = in1[3] ^ in2[3];
    assign G[11] = in1[2] & in2[2];
    assign P[11] = in1[2] ^ in2[2];
    assign G[12] = in1[1] & in2[1];
    assign P[12] = in1[1] ^ in2[1];
    assign G[13] = in1[0] & in2[0];
    assign P[13] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign cout = G[13] | (P[13] & C[13]);
    assign sum = P ^ C;
endmodule

module CLA_13(output [12:0] sum, output cout, input [12:0] in1, input [12:0] in2);

    wire[12:0] G;
    wire[12:0] C;
    wire[12:0] P;

    assign G[0] = in1[12] & in2[12];
    assign P[0] = in1[12] ^ in2[12];
    assign G[1] = in1[11] & in2[11];
    assign P[1] = in1[11] ^ in2[11];
    assign G[2] = in1[10] & in2[10];
    assign P[2] = in1[10] ^ in2[10];
    assign G[3] = in1[9] & in2[9];
    assign P[3] = in1[9] ^ in2[9];
    assign G[4] = in1[8] & in2[8];
    assign P[4] = in1[8] ^ in2[8];
    assign G[5] = in1[7] & in2[7];
    assign P[5] = in1[7] ^ in2[7];
    assign G[6] = in1[6] & in2[6];
    assign P[6] = in1[6] ^ in2[6];
    assign G[7] = in1[5] & in2[5];
    assign P[7] = in1[5] ^ in2[5];
    assign G[8] = in1[4] & in2[4];
    assign P[8] = in1[4] ^ in2[4];
    assign G[9] = in1[3] & in2[3];
    assign P[9] = in1[3] ^ in2[3];
    assign G[10] = in1[2] & in2[2];
    assign P[10] = in1[2] ^ in2[2];
    assign G[11] = in1[1] & in2[1];
    assign P[11] = in1[1] ^ in2[1];
    assign G[12] = in1[0] & in2[0];
    assign P[12] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign cout = G[12] | (P[12] & C[12]);
    assign sum = P ^ C;
endmodule

module CLA_12(output [11:0] sum, output cout, input [11:0] in1, input [11:0] in2);

    wire[11:0] G;
    wire[11:0] C;
    wire[11:0] P;

    assign G[0] = in1[11] & in2[11];
    assign P[0] = in1[11] ^ in2[11];
    assign G[1] = in1[10] & in2[10];
    assign P[1] = in1[10] ^ in2[10];
    assign G[2] = in1[9] & in2[9];
    assign P[2] = in1[9] ^ in2[9];
    assign G[3] = in1[8] & in2[8];
    assign P[3] = in1[8] ^ in2[8];
    assign G[4] = in1[7] & in2[7];
    assign P[4] = in1[7] ^ in2[7];
    assign G[5] = in1[6] & in2[6];
    assign P[5] = in1[6] ^ in2[6];
    assign G[6] = in1[5] & in2[5];
    assign P[6] = in1[5] ^ in2[5];
    assign G[7] = in1[4] & in2[4];
    assign P[7] = in1[4] ^ in2[4];
    assign G[8] = in1[3] & in2[3];
    assign P[8] = in1[3] ^ in2[3];
    assign G[9] = in1[2] & in2[2];
    assign P[9] = in1[2] ^ in2[2];
    assign G[10] = in1[1] & in2[1];
    assign P[10] = in1[1] ^ in2[1];
    assign G[11] = in1[0] & in2[0];
    assign P[11] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign cout = G[11] | (P[11] & C[11]);
    assign sum = P ^ C;
endmodule

module CLA_11(output [10:0] sum, output cout, input [10:0] in1, input [10:0] in2);

    wire[10:0] G;
    wire[10:0] C;
    wire[10:0] P;

    assign G[0] = in1[10] & in2[10];
    assign P[0] = in1[10] ^ in2[10];
    assign G[1] = in1[9] & in2[9];
    assign P[1] = in1[9] ^ in2[9];
    assign G[2] = in1[8] & in2[8];
    assign P[2] = in1[8] ^ in2[8];
    assign G[3] = in1[7] & in2[7];
    assign P[3] = in1[7] ^ in2[7];
    assign G[4] = in1[6] & in2[6];
    assign P[4] = in1[6] ^ in2[6];
    assign G[5] = in1[5] & in2[5];
    assign P[5] = in1[5] ^ in2[5];
    assign G[6] = in1[4] & in2[4];
    assign P[6] = in1[4] ^ in2[4];
    assign G[7] = in1[3] & in2[3];
    assign P[7] = in1[3] ^ in2[3];
    assign G[8] = in1[2] & in2[2];
    assign P[8] = in1[2] ^ in2[2];
    assign G[9] = in1[1] & in2[1];
    assign P[9] = in1[1] ^ in2[1];
    assign G[10] = in1[0] & in2[0];
    assign P[10] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign cout = G[10] | (P[10] & C[10]);
    assign sum = P ^ C;
endmodule

module CLA_10(output [9:0] sum, output cout, input [9:0] in1, input [9:0] in2);

    wire[9:0] G;
    wire[9:0] C;
    wire[9:0] P;

    assign G[0] = in1[9] & in2[9];
    assign P[0] = in1[9] ^ in2[9];
    assign G[1] = in1[8] & in2[8];
    assign P[1] = in1[8] ^ in2[8];
    assign G[2] = in1[7] & in2[7];
    assign P[2] = in1[7] ^ in2[7];
    assign G[3] = in1[6] & in2[6];
    assign P[3] = in1[6] ^ in2[6];
    assign G[4] = in1[5] & in2[5];
    assign P[4] = in1[5] ^ in2[5];
    assign G[5] = in1[4] & in2[4];
    assign P[5] = in1[4] ^ in2[4];
    assign G[6] = in1[3] & in2[3];
    assign P[6] = in1[3] ^ in2[3];
    assign G[7] = in1[2] & in2[2];
    assign P[7] = in1[2] ^ in2[2];
    assign G[8] = in1[1] & in2[1];
    assign P[8] = in1[1] ^ in2[1];
    assign G[9] = in1[0] & in2[0];
    assign P[9] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign cout = G[9] | (P[9] & C[9]);
    assign sum = P ^ C;
endmodule

module CLA_9(output [8:0] sum, output cout, input [8:0] in1, input [8:0] in2);

    wire[8:0] G;
    wire[8:0] C;
    wire[8:0] P;

    assign G[0] = in1[8] & in2[8];
    assign P[0] = in1[8] ^ in2[8];
    assign G[1] = in1[7] & in2[7];
    assign P[1] = in1[7] ^ in2[7];
    assign G[2] = in1[6] & in2[6];
    assign P[2] = in1[6] ^ in2[6];
    assign G[3] = in1[5] & in2[5];
    assign P[3] = in1[5] ^ in2[5];
    assign G[4] = in1[4] & in2[4];
    assign P[4] = in1[4] ^ in2[4];
    assign G[5] = in1[3] & in2[3];
    assign P[5] = in1[3] ^ in2[3];
    assign G[6] = in1[2] & in2[2];
    assign P[6] = in1[2] ^ in2[2];
    assign G[7] = in1[1] & in2[1];
    assign P[7] = in1[1] ^ in2[1];
    assign G[8] = in1[0] & in2[0];
    assign P[8] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign cout = G[8] | (P[8] & C[8]);
    assign sum = P ^ C;
endmodule

module CLA_8(output [7:0] sum, output cout, input [7:0] in1, input [7:0] in2);

    wire[7:0] G;
    wire[7:0] C;
    wire[7:0] P;

    assign G[0] = in1[7] & in2[7];
    assign P[0] = in1[7] ^ in2[7];
    assign G[1] = in1[6] & in2[6];
    assign P[1] = in1[6] ^ in2[6];
    assign G[2] = in1[5] & in2[5];
    assign P[2] = in1[5] ^ in2[5];
    assign G[3] = in1[4] & in2[4];
    assign P[3] = in1[4] ^ in2[4];
    assign G[4] = in1[3] & in2[3];
    assign P[4] = in1[3] ^ in2[3];
    assign G[5] = in1[2] & in2[2];
    assign P[5] = in1[2] ^ in2[2];
    assign G[6] = in1[1] & in2[1];
    assign P[6] = in1[1] ^ in2[1];
    assign G[7] = in1[0] & in2[0];
    assign P[7] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign cout = G[7] | (P[7] & C[7]);
    assign sum = P ^ C;
endmodule

module CLA_7(output [6:0] sum, output cout, input [6:0] in1, input [6:0] in2);

    wire[6:0] G;
    wire[6:0] C;
    wire[6:0] P;

    assign G[0] = in1[6] & in2[6];
    assign P[0] = in1[6] ^ in2[6];
    assign G[1] = in1[5] & in2[5];
    assign P[1] = in1[5] ^ in2[5];
    assign G[2] = in1[4] & in2[4];
    assign P[2] = in1[4] ^ in2[4];
    assign G[3] = in1[3] & in2[3];
    assign P[3] = in1[3] ^ in2[3];
    assign G[4] = in1[2] & in2[2];
    assign P[4] = in1[2] ^ in2[2];
    assign G[5] = in1[1] & in2[1];
    assign P[5] = in1[1] ^ in2[1];
    assign G[6] = in1[0] & in2[0];
    assign P[6] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign cout = G[6] | (P[6] & C[6]);
    assign sum = P ^ C;
endmodule

module CLA_6(output [5:0] sum, output cout, input [5:0] in1, input [5:0] in2);

    wire[5:0] G;
    wire[5:0] C;
    wire[5:0] P;

    assign G[0] = in1[5] & in2[5];
    assign P[0] = in1[5] ^ in2[5];
    assign G[1] = in1[4] & in2[4];
    assign P[1] = in1[4] ^ in2[4];
    assign G[2] = in1[3] & in2[3];
    assign P[2] = in1[3] ^ in2[3];
    assign G[3] = in1[2] & in2[2];
    assign P[3] = in1[2] ^ in2[2];
    assign G[4] = in1[1] & in2[1];
    assign P[4] = in1[1] ^ in2[1];
    assign G[5] = in1[0] & in2[0];
    assign P[5] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign cout = G[5] | (P[5] & C[5]);
    assign sum = P ^ C;
endmodule

module CLA_5(output [4:0] sum, output cout, input [4:0] in1, input [4:0] in2);

    wire[4:0] G;
    wire[4:0] C;
    wire[4:0] P;

    assign G[0] = in1[4] & in2[4];
    assign P[0] = in1[4] ^ in2[4];
    assign G[1] = in1[3] & in2[3];
    assign P[1] = in1[3] ^ in2[3];
    assign G[2] = in1[2] & in2[2];
    assign P[2] = in1[2] ^ in2[2];
    assign G[3] = in1[1] & in2[1];
    assign P[3] = in1[1] ^ in2[1];
    assign G[4] = in1[0] & in2[0];
    assign P[4] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign cout = G[4] | (P[4] & C[4]);
    assign sum = P ^ C;
endmodule

module CLA_4(output [3:0] sum, output cout, input [3:0] in1, input [3:0] in2);

    wire[3:0] G;
    wire[3:0] C;
    wire[3:0] P;

    assign G[0] = in1[3] & in2[3];
    assign P[0] = in1[3] ^ in2[3];
    assign G[1] = in1[2] & in2[2];
    assign P[1] = in1[2] ^ in2[2];
    assign G[2] = in1[1] & in2[1];
    assign P[2] = in1[1] ^ in2[1];
    assign G[3] = in1[0] & in2[0];
    assign P[3] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA_3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2);

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in1[2] & in2[2];
    assign P[0] = in1[2] ^ in2[2];
    assign G[1] = in1[1] & in2[1];
    assign P[1] = in1[1] ^ in2[1];
    assign G[2] = in1[0] & in2[0];
    assign P[2] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA_2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2);

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in1[1] & in2[1];
    assign P[0] = in1[1] ^ in2[1];
    assign G[1] = in1[0] & in2[0];
    assign P[1] = in1[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule

