module multiplier_64bits_version10(product, A, B);

    output [127:0] product;
    input [63:0] A, B;

    wire [63:0] pp0;
    wire [63:0] pp1;
    wire [63:0] pp2;
    wire [63:0] pp3;
    wire [63:0] pp4;
    wire [63:0] pp5;
    wire [63:0] pp6;
    wire [63:0] pp7;
    wire [63:0] pp8;
    wire [63:0] pp9;
    wire [63:0] pp10;
    wire [63:0] pp11;
    wire [63:0] pp12;
    wire [63:0] pp13;
    wire [63:0] pp14;
    wire [63:0] pp15;
    wire [63:0] pp16;
    wire [63:0] pp17;
    wire [63:0] pp18;
    wire [63:0] pp19;
    wire [63:0] pp20;
    wire [63:0] pp21;
    wire [63:0] pp22;
    wire [63:0] pp23;
    wire [63:0] pp24;
    wire [63:0] pp25;
    wire [63:0] pp26;
    wire [63:0] pp27;
    wire [63:0] pp28;
    wire [63:0] pp29;
    wire [63:0] pp30;
    wire [63:0] pp31;
    wire [63:0] pp32;
    wire [63:0] pp33;
    wire [63:0] pp34;
    wire [63:0] pp35;
    wire [63:0] pp36;
    wire [63:0] pp37;
    wire [63:0] pp38;
    wire [63:0] pp39;
    wire [63:0] pp40;
    wire [63:0] pp41;
    wire [63:0] pp42;
    wire [63:0] pp43;
    wire [63:0] pp44;
    wire [63:0] pp45;
    wire [63:0] pp46;
    wire [63:0] pp47;
    wire [63:0] pp48;
    wire [63:0] pp49;
    wire [63:0] pp50;
    wire [63:0] pp51;
    wire [63:0] pp52;
    wire [63:0] pp53;
    wire [63:0] pp54;
    wire [63:0] pp55;
    wire [63:0] pp56;
    wire [63:0] pp57;
    wire [63:0] pp58;
    wire [63:0] pp59;
    wire [63:0] pp60;
    wire [63:0] pp61;
    wire [63:0] pp62;
    wire [63:0] pp63;


    assign pp0 = A[0] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp1 = A[1] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp2 = A[2] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp3 = A[3] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp4 = A[4] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp5 = A[5] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp6 = A[6] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp7 = A[7] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp8 = A[8] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp9 = A[9] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp10 = A[10] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp11 = A[11] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp12 = A[12] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp13 = A[13] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp14 = A[14] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp15 = A[15] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp16 = A[16] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp17 = A[17] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp18 = A[18] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp19 = A[19] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp20 = A[20] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp21 = A[21] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp22 = A[22] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp23 = A[23] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp24 = A[24] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp25 = A[25] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp26 = A[26] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp27 = A[27] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp28 = A[28] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp29 = A[29] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp30 = A[30] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp31 = A[31] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp32 = A[32] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp33 = A[33] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp34 = A[34] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp35 = A[35] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp36 = A[36] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp37 = A[37] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp38 = A[38] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp39 = A[39] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp40 = A[40] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp41 = A[41] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp42 = A[42] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp43 = A[43] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp44 = A[44] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp45 = A[45] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp46 = A[46] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp47 = A[47] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp48 = A[48] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp49 = A[49] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp50 = A[50] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp51 = A[51] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp52 = A[52] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp53 = A[53] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp54 = A[54] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp55 = A[55] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp56 = A[56] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp57 = A[57] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp58 = A[58] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp59 = A[59] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp60 = A[60] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp61 = A[61] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp62 = A[62] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;
    assign pp63 = A[63] ? B: 64'b0000000000000000000000000000000000000000000000000000000000000000;


    /*Stage 1*/
    wire[63:0] s1, in1_1, in1_2;
    wire c1;
    assign in1_1 = {pp0[32],pp0[33],pp0[34],pp0[35],pp0[36],pp0[37],pp0[38],pp0[39],pp0[40],pp0[41],pp0[42],pp0[43],pp0[44],pp0[45],pp0[46],pp0[47],pp0[48],pp0[49],pp0[50],pp0[51],pp0[52],pp0[53],pp0[54],pp0[55],pp0[56],pp0[57],pp0[58],pp0[59],pp0[60],pp0[61],pp0[62],pp0[63],pp1[63],pp2[63],pp3[63],pp4[63],pp5[63],pp6[63],pp7[63],pp8[63],pp9[63],pp10[63],pp11[63],pp12[63],pp13[63],pp14[63],pp15[63],pp16[63],pp17[63],pp18[63],pp19[63],pp20[63],pp21[63],pp22[63],pp23[63],pp24[63],pp25[63],pp26[63],pp27[63],pp28[63],pp29[63],pp30[63],pp31[63],pp32[63]};
    assign in1_2 = {pp1[31],pp1[32],pp1[33],pp1[34],pp1[35],pp1[36],pp1[37],pp1[38],pp1[39],pp1[40],pp1[41],pp1[42],pp1[43],pp1[44],pp1[45],pp1[46],pp1[47],pp1[48],pp1[49],pp1[50],pp1[51],pp1[52],pp1[53],pp1[54],pp1[55],pp1[56],pp1[57],pp1[58],pp1[59],pp1[60],pp1[61],pp1[62],pp2[62],pp3[62],pp4[62],pp5[62],pp6[62],pp7[62],pp8[62],pp9[62],pp10[62],pp11[62],pp12[62],pp13[62],pp14[62],pp15[62],pp16[62],pp17[62],pp18[62],pp19[62],pp20[62],pp21[62],pp22[62],pp23[62],pp24[62],pp25[62],pp26[62],pp27[62],pp28[62],pp29[62],pp30[62],pp31[62],pp32[62],pp33[62]};
    CLA_64 KS_1(s1, c1, in1_1, in1_2);
    wire[61:0] s2, in2_1, in2_2;
    wire c2;
    assign in2_1 = {pp2[31],pp2[32],pp2[33],pp2[34],pp2[35],pp2[36],pp2[37],pp2[38],pp2[39],pp2[40],pp2[41],pp2[42],pp2[43],pp2[44],pp2[45],pp2[46],pp2[47],pp2[48],pp2[49],pp2[50],pp2[51],pp2[52],pp2[53],pp2[54],pp2[55],pp2[56],pp2[57],pp2[58],pp2[59],pp2[60],pp2[61],pp3[61],pp4[61],pp5[61],pp6[61],pp7[61],pp8[61],pp9[61],pp10[61],pp11[61],pp12[61],pp13[61],pp14[61],pp15[61],pp16[61],pp17[61],pp18[61],pp19[61],pp20[61],pp21[61],pp22[61],pp23[61],pp24[61],pp25[61],pp26[61],pp27[61],pp28[61],pp29[61],pp30[61],pp31[61],pp32[61],pp33[61]};
    assign in2_2 = {pp3[30],pp3[31],pp3[32],pp3[33],pp3[34],pp3[35],pp3[36],pp3[37],pp3[38],pp3[39],pp3[40],pp3[41],pp3[42],pp3[43],pp3[44],pp3[45],pp3[46],pp3[47],pp3[48],pp3[49],pp3[50],pp3[51],pp3[52],pp3[53],pp3[54],pp3[55],pp3[56],pp3[57],pp3[58],pp3[59],pp3[60],pp4[60],pp5[60],pp6[60],pp7[60],pp8[60],pp9[60],pp10[60],pp11[60],pp12[60],pp13[60],pp14[60],pp15[60],pp16[60],pp17[60],pp18[60],pp19[60],pp20[60],pp21[60],pp22[60],pp23[60],pp24[60],pp25[60],pp26[60],pp27[60],pp28[60],pp29[60],pp30[60],pp31[60],pp32[60],pp33[60],pp34[60]};
    CLA_62 KS_2(s2, c2, in2_1, in2_2);
    wire[59:0] s3, in3_1, in3_2;
    wire c3;
    assign in3_1 = {pp4[30],pp4[31],pp4[32],pp4[33],pp4[34],pp4[35],pp4[36],pp4[37],pp4[38],pp4[39],pp4[40],pp4[41],pp4[42],pp4[43],pp4[44],pp4[45],pp4[46],pp4[47],pp4[48],pp4[49],pp4[50],pp4[51],pp4[52],pp4[53],pp4[54],pp4[55],pp4[56],pp4[57],pp4[58],pp4[59],pp5[59],pp6[59],pp7[59],pp8[59],pp9[59],pp10[59],pp11[59],pp12[59],pp13[59],pp14[59],pp15[59],pp16[59],pp17[59],pp18[59],pp19[59],pp20[59],pp21[59],pp22[59],pp23[59],pp24[59],pp25[59],pp26[59],pp27[59],pp28[59],pp29[59],pp30[59],pp31[59],pp32[59],pp33[59],pp34[59]};
    assign in3_2 = {pp5[29],pp5[30],pp5[31],pp5[32],pp5[33],pp5[34],pp5[35],pp5[36],pp5[37],pp5[38],pp5[39],pp5[40],pp5[41],pp5[42],pp5[43],pp5[44],pp5[45],pp5[46],pp5[47],pp5[48],pp5[49],pp5[50],pp5[51],pp5[52],pp5[53],pp5[54],pp5[55],pp5[56],pp5[57],pp5[58],pp6[58],pp7[58],pp8[58],pp9[58],pp10[58],pp11[58],pp12[58],pp13[58],pp14[58],pp15[58],pp16[58],pp17[58],pp18[58],pp19[58],pp20[58],pp21[58],pp22[58],pp23[58],pp24[58],pp25[58],pp26[58],pp27[58],pp28[58],pp29[58],pp30[58],pp31[58],pp32[58],pp33[58],pp34[58],pp35[58]};
    CLA_60 KS_3(s3, c3, in3_1, in3_2);
    wire[57:0] s4, in4_1, in4_2;
    wire c4;
    assign in4_1 = {pp6[29],pp6[30],pp6[31],pp6[32],pp6[33],pp6[34],pp6[35],pp6[36],pp6[37],pp6[38],pp6[39],pp6[40],pp6[41],pp6[42],pp6[43],pp6[44],pp6[45],pp6[46],pp6[47],pp6[48],pp6[49],pp6[50],pp6[51],pp6[52],pp6[53],pp6[54],pp6[55],pp6[56],pp6[57],pp7[57],pp8[57],pp9[57],pp10[57],pp11[57],pp12[57],pp13[57],pp14[57],pp15[57],pp16[57],pp17[57],pp18[57],pp19[57],pp20[57],pp21[57],pp22[57],pp23[57],pp24[57],pp25[57],pp26[57],pp27[57],pp28[57],pp29[57],pp30[57],pp31[57],pp32[57],pp33[57],pp34[57],pp35[57]};
    assign in4_2 = {pp7[28],pp7[29],pp7[30],pp7[31],pp7[32],pp7[33],pp7[34],pp7[35],pp7[36],pp7[37],pp7[38],pp7[39],pp7[40],pp7[41],pp7[42],pp7[43],pp7[44],pp7[45],pp7[46],pp7[47],pp7[48],pp7[49],pp7[50],pp7[51],pp7[52],pp7[53],pp7[54],pp7[55],pp7[56],pp8[56],pp9[56],pp10[56],pp11[56],pp12[56],pp13[56],pp14[56],pp15[56],pp16[56],pp17[56],pp18[56],pp19[56],pp20[56],pp21[56],pp22[56],pp23[56],pp24[56],pp25[56],pp26[56],pp27[56],pp28[56],pp29[56],pp30[56],pp31[56],pp32[56],pp33[56],pp34[56],pp35[56],pp36[56]};
    CLA_58 KS_4(s4, c4, in4_1, in4_2);
    wire[55:0] s5, in5_1, in5_2;
    wire c5;
    assign in5_1 = {pp8[28],pp8[29],pp8[30],pp8[31],pp8[32],pp8[33],pp8[34],pp8[35],pp8[36],pp8[37],pp8[38],pp8[39],pp8[40],pp8[41],pp8[42],pp8[43],pp8[44],pp8[45],pp8[46],pp8[47],pp8[48],pp8[49],pp8[50],pp8[51],pp8[52],pp8[53],pp8[54],pp8[55],pp9[55],pp10[55],pp11[55],pp12[55],pp13[55],pp14[55],pp15[55],pp16[55],pp17[55],pp18[55],pp19[55],pp20[55],pp21[55],pp22[55],pp23[55],pp24[55],pp25[55],pp26[55],pp27[55],pp28[55],pp29[55],pp30[55],pp31[55],pp32[55],pp33[55],pp34[55],pp35[55],pp36[55]};
    assign in5_2 = {pp9[27],pp9[28],pp9[29],pp9[30],pp9[31],pp9[32],pp9[33],pp9[34],pp9[35],pp9[36],pp9[37],pp9[38],pp9[39],pp9[40],pp9[41],pp9[42],pp9[43],pp9[44],pp9[45],pp9[46],pp9[47],pp9[48],pp9[49],pp9[50],pp9[51],pp9[52],pp9[53],pp9[54],pp10[54],pp11[54],pp12[54],pp13[54],pp14[54],pp15[54],pp16[54],pp17[54],pp18[54],pp19[54],pp20[54],pp21[54],pp22[54],pp23[54],pp24[54],pp25[54],pp26[54],pp27[54],pp28[54],pp29[54],pp30[54],pp31[54],pp32[54],pp33[54],pp34[54],pp35[54],pp36[54],pp37[54]};
    CLA_56 KS_5(s5, c5, in5_1, in5_2);
    wire[53:0] s6, in6_1, in6_2;
    wire c6;
    assign in6_1 = {pp10[27],pp10[28],pp10[29],pp10[30],pp10[31],pp10[32],pp10[33],pp10[34],pp10[35],pp10[36],pp10[37],pp10[38],pp10[39],pp10[40],pp10[41],pp10[42],pp10[43],pp10[44],pp10[45],pp10[46],pp10[47],pp10[48],pp10[49],pp10[50],pp10[51],pp10[52],pp10[53],pp11[53],pp12[53],pp13[53],pp14[53],pp15[53],pp16[53],pp17[53],pp18[53],pp19[53],pp20[53],pp21[53],pp22[53],pp23[53],pp24[53],pp25[53],pp26[53],pp27[53],pp28[53],pp29[53],pp30[53],pp31[53],pp32[53],pp33[53],pp34[53],pp35[53],pp36[53],pp37[53]};
    assign in6_2 = {pp11[26],pp11[27],pp11[28],pp11[29],pp11[30],pp11[31],pp11[32],pp11[33],pp11[34],pp11[35],pp11[36],pp11[37],pp11[38],pp11[39],pp11[40],pp11[41],pp11[42],pp11[43],pp11[44],pp11[45],pp11[46],pp11[47],pp11[48],pp11[49],pp11[50],pp11[51],pp11[52],pp12[52],pp13[52],pp14[52],pp15[52],pp16[52],pp17[52],pp18[52],pp19[52],pp20[52],pp21[52],pp22[52],pp23[52],pp24[52],pp25[52],pp26[52],pp27[52],pp28[52],pp29[52],pp30[52],pp31[52],pp32[52],pp33[52],pp34[52],pp35[52],pp36[52],pp37[52],pp38[52]};
    CLA_54 KS_6(s6, c6, in6_1, in6_2);
    wire[51:0] s7, in7_1, in7_2;
    wire c7;
    assign in7_1 = {pp12[26],pp12[27],pp12[28],pp12[29],pp12[30],pp12[31],pp12[32],pp12[33],pp12[34],pp12[35],pp12[36],pp12[37],pp12[38],pp12[39],pp12[40],pp12[41],pp12[42],pp12[43],pp12[44],pp12[45],pp12[46],pp12[47],pp12[48],pp12[49],pp12[50],pp12[51],pp13[51],pp14[51],pp15[51],pp16[51],pp17[51],pp18[51],pp19[51],pp20[51],pp21[51],pp22[51],pp23[51],pp24[51],pp25[51],pp26[51],pp27[51],pp28[51],pp29[51],pp30[51],pp31[51],pp32[51],pp33[51],pp34[51],pp35[51],pp36[51],pp37[51],pp38[51]};
    assign in7_2 = {pp13[25],pp13[26],pp13[27],pp13[28],pp13[29],pp13[30],pp13[31],pp13[32],pp13[33],pp13[34],pp13[35],pp13[36],pp13[37],pp13[38],pp13[39],pp13[40],pp13[41],pp13[42],pp13[43],pp13[44],pp13[45],pp13[46],pp13[47],pp13[48],pp13[49],pp13[50],pp14[50],pp15[50],pp16[50],pp17[50],pp18[50],pp19[50],pp20[50],pp21[50],pp22[50],pp23[50],pp24[50],pp25[50],pp26[50],pp27[50],pp28[50],pp29[50],pp30[50],pp31[50],pp32[50],pp33[50],pp34[50],pp35[50],pp36[50],pp37[50],pp38[50],pp39[50]};
    CLA_52 KS_7(s7, c7, in7_1, in7_2);
    wire[49:0] s8, in8_1, in8_2;
    wire c8;
    assign in8_1 = {pp14[25],pp14[26],pp14[27],pp14[28],pp14[29],pp14[30],pp14[31],pp14[32],pp14[33],pp14[34],pp14[35],pp14[36],pp14[37],pp14[38],pp14[39],pp14[40],pp14[41],pp14[42],pp14[43],pp14[44],pp14[45],pp14[46],pp14[47],pp14[48],pp14[49],pp15[49],pp16[49],pp17[49],pp18[49],pp19[49],pp20[49],pp21[49],pp22[49],pp23[49],pp24[49],pp25[49],pp26[49],pp27[49],pp28[49],pp29[49],pp30[49],pp31[49],pp32[49],pp33[49],pp34[49],pp35[49],pp36[49],pp37[49],pp38[49],pp39[49]};
    assign in8_2 = {pp15[24],pp15[25],pp15[26],pp15[27],pp15[28],pp15[29],pp15[30],pp15[31],pp15[32],pp15[33],pp15[34],pp15[35],pp15[36],pp15[37],pp15[38],pp15[39],pp15[40],pp15[41],pp15[42],pp15[43],pp15[44],pp15[45],pp15[46],pp15[47],pp15[48],pp16[48],pp17[48],pp18[48],pp19[48],pp20[48],pp21[48],pp22[48],pp23[48],pp24[48],pp25[48],pp26[48],pp27[48],pp28[48],pp29[48],pp30[48],pp31[48],pp32[48],pp33[48],pp34[48],pp35[48],pp36[48],pp37[48],pp38[48],pp39[48],pp40[48]};
    CLA_50 KS_8(s8, c8, in8_1, in8_2);
    wire[47:0] s9, in9_1, in9_2;
    wire c9;
    assign in9_1 = {pp16[24],pp16[25],pp16[26],pp16[27],pp16[28],pp16[29],pp16[30],pp16[31],pp16[32],pp16[33],pp16[34],pp16[35],pp16[36],pp16[37],pp16[38],pp16[39],pp16[40],pp16[41],pp16[42],pp16[43],pp16[44],pp16[45],pp16[46],pp16[47],pp17[47],pp18[47],pp19[47],pp20[47],pp21[47],pp22[47],pp23[47],pp24[47],pp25[47],pp26[47],pp27[47],pp28[47],pp29[47],pp30[47],pp31[47],pp32[47],pp33[47],pp34[47],pp35[47],pp36[47],pp37[47],pp38[47],pp39[47],pp40[47]};
    assign in9_2 = {pp17[23],pp17[24],pp17[25],pp17[26],pp17[27],pp17[28],pp17[29],pp17[30],pp17[31],pp17[32],pp17[33],pp17[34],pp17[35],pp17[36],pp17[37],pp17[38],pp17[39],pp17[40],pp17[41],pp17[42],pp17[43],pp17[44],pp17[45],pp17[46],pp18[46],pp19[46],pp20[46],pp21[46],pp22[46],pp23[46],pp24[46],pp25[46],pp26[46],pp27[46],pp28[46],pp29[46],pp30[46],pp31[46],pp32[46],pp33[46],pp34[46],pp35[46],pp36[46],pp37[46],pp38[46],pp39[46],pp40[46],pp41[46]};
    CLA_48 KS_9(s9, c9, in9_1, in9_2);
    wire[45:0] s10, in10_1, in10_2;
    wire c10;
    assign in10_1 = {pp18[23],pp18[24],pp18[25],pp18[26],pp18[27],pp18[28],pp18[29],pp18[30],pp18[31],pp18[32],pp18[33],pp18[34],pp18[35],pp18[36],pp18[37],pp18[38],pp18[39],pp18[40],pp18[41],pp18[42],pp18[43],pp18[44],pp18[45],pp19[45],pp20[45],pp21[45],pp22[45],pp23[45],pp24[45],pp25[45],pp26[45],pp27[45],pp28[45],pp29[45],pp30[45],pp31[45],pp32[45],pp33[45],pp34[45],pp35[45],pp36[45],pp37[45],pp38[45],pp39[45],pp40[45],pp41[45]};
    assign in10_2 = {pp19[22],pp19[23],pp19[24],pp19[25],pp19[26],pp19[27],pp19[28],pp19[29],pp19[30],pp19[31],pp19[32],pp19[33],pp19[34],pp19[35],pp19[36],pp19[37],pp19[38],pp19[39],pp19[40],pp19[41],pp19[42],pp19[43],pp19[44],pp20[44],pp21[44],pp22[44],pp23[44],pp24[44],pp25[44],pp26[44],pp27[44],pp28[44],pp29[44],pp30[44],pp31[44],pp32[44],pp33[44],pp34[44],pp35[44],pp36[44],pp37[44],pp38[44],pp39[44],pp40[44],pp41[44],pp42[44]};
    CLA_46 KS_10(s10, c10, in10_1, in10_2);
    wire[43:0] s11, in11_1, in11_2;
    wire c11;
    assign in11_1 = {pp20[22],pp20[23],pp20[24],pp20[25],pp20[26],pp20[27],pp20[28],pp20[29],pp20[30],pp20[31],pp20[32],pp20[33],pp20[34],pp20[35],pp20[36],pp20[37],pp20[38],pp20[39],pp20[40],pp20[41],pp20[42],pp20[43],pp21[43],pp22[43],pp23[43],pp24[43],pp25[43],pp26[43],pp27[43],pp28[43],pp29[43],pp30[43],pp31[43],pp32[43],pp33[43],pp34[43],pp35[43],pp36[43],pp37[43],pp38[43],pp39[43],pp40[43],pp41[43],pp42[43]};
    assign in11_2 = {pp21[21],pp21[22],pp21[23],pp21[24],pp21[25],pp21[26],pp21[27],pp21[28],pp21[29],pp21[30],pp21[31],pp21[32],pp21[33],pp21[34],pp21[35],pp21[36],pp21[37],pp21[38],pp21[39],pp21[40],pp21[41],pp21[42],pp22[42],pp23[42],pp24[42],pp25[42],pp26[42],pp27[42],pp28[42],pp29[42],pp30[42],pp31[42],pp32[42],pp33[42],pp34[42],pp35[42],pp36[42],pp37[42],pp38[42],pp39[42],pp40[42],pp41[42],pp42[42],pp43[42]};
    CLA_44 KS_11(s11, c11, in11_1, in11_2);
    wire[41:0] s12, in12_1, in12_2;
    wire c12;
    assign in12_1 = {pp22[21],pp22[22],pp22[23],pp22[24],pp22[25],pp22[26],pp22[27],pp22[28],pp22[29],pp22[30],pp22[31],pp22[32],pp22[33],pp22[34],pp22[35],pp22[36],pp22[37],pp22[38],pp22[39],pp22[40],pp22[41],pp23[41],pp24[41],pp25[41],pp26[41],pp27[41],pp28[41],pp29[41],pp30[41],pp31[41],pp32[41],pp33[41],pp34[41],pp35[41],pp36[41],pp37[41],pp38[41],pp39[41],pp40[41],pp41[41],pp42[41],pp43[41]};
    assign in12_2 = {pp23[20],pp23[21],pp23[22],pp23[23],pp23[24],pp23[25],pp23[26],pp23[27],pp23[28],pp23[29],pp23[30],pp23[31],pp23[32],pp23[33],pp23[34],pp23[35],pp23[36],pp23[37],pp23[38],pp23[39],pp23[40],pp24[40],pp25[40],pp26[40],pp27[40],pp28[40],pp29[40],pp30[40],pp31[40],pp32[40],pp33[40],pp34[40],pp35[40],pp36[40],pp37[40],pp38[40],pp39[40],pp40[40],pp41[40],pp42[40],pp43[40],pp44[40]};
    CLA_42 KS_12(s12, c12, in12_1, in12_2);
    wire[39:0] s13, in13_1, in13_2;
    wire c13;
    assign in13_1 = {pp24[20],pp24[21],pp24[22],pp24[23],pp24[24],pp24[25],pp24[26],pp24[27],pp24[28],pp24[29],pp24[30],pp24[31],pp24[32],pp24[33],pp24[34],pp24[35],pp24[36],pp24[37],pp24[38],pp24[39],pp25[39],pp26[39],pp27[39],pp28[39],pp29[39],pp30[39],pp31[39],pp32[39],pp33[39],pp34[39],pp35[39],pp36[39],pp37[39],pp38[39],pp39[39],pp40[39],pp41[39],pp42[39],pp43[39],pp44[39]};
    assign in13_2 = {pp25[19],pp25[20],pp25[21],pp25[22],pp25[23],pp25[24],pp25[25],pp25[26],pp25[27],pp25[28],pp25[29],pp25[30],pp25[31],pp25[32],pp25[33],pp25[34],pp25[35],pp25[36],pp25[37],pp25[38],pp26[38],pp27[38],pp28[38],pp29[38],pp30[38],pp31[38],pp32[38],pp33[38],pp34[38],pp35[38],pp36[38],pp37[38],pp38[38],pp39[38],pp40[38],pp41[38],pp42[38],pp43[38],pp44[38],pp45[38]};
    CLA_40 KS_13(s13, c13, in13_1, in13_2);
    wire[37:0] s14, in14_1, in14_2;
    wire c14;
    assign in14_1 = {pp26[19],pp26[20],pp26[21],pp26[22],pp26[23],pp26[24],pp26[25],pp26[26],pp26[27],pp26[28],pp26[29],pp26[30],pp26[31],pp26[32],pp26[33],pp26[34],pp26[35],pp26[36],pp26[37],pp27[37],pp28[37],pp29[37],pp30[37],pp31[37],pp32[37],pp33[37],pp34[37],pp35[37],pp36[37],pp37[37],pp38[37],pp39[37],pp40[37],pp41[37],pp42[37],pp43[37],pp44[37],pp45[37]};
    assign in14_2 = {pp27[18],pp27[19],pp27[20],pp27[21],pp27[22],pp27[23],pp27[24],pp27[25],pp27[26],pp27[27],pp27[28],pp27[29],pp27[30],pp27[31],pp27[32],pp27[33],pp27[34],pp27[35],pp27[36],pp28[36],pp29[36],pp30[36],pp31[36],pp32[36],pp33[36],pp34[36],pp35[36],pp36[36],pp37[36],pp38[36],pp39[36],pp40[36],pp41[36],pp42[36],pp43[36],pp44[36],pp45[36],pp46[36]};
    CLA_38 KS_14(s14, c14, in14_1, in14_2);
    wire[35:0] s15, in15_1, in15_2;
    wire c15;
    assign in15_1 = {pp28[18],pp28[19],pp28[20],pp28[21],pp28[22],pp28[23],pp28[24],pp28[25],pp28[26],pp28[27],pp28[28],pp28[29],pp28[30],pp28[31],pp28[32],pp28[33],pp28[34],pp28[35],pp29[35],pp30[35],pp31[35],pp32[35],pp33[35],pp34[35],pp35[35],pp36[35],pp37[35],pp38[35],pp39[35],pp40[35],pp41[35],pp42[35],pp43[35],pp44[35],pp45[35],pp46[35]};
    assign in15_2 = {pp29[17],pp29[18],pp29[19],pp29[20],pp29[21],pp29[22],pp29[23],pp29[24],pp29[25],pp29[26],pp29[27],pp29[28],pp29[29],pp29[30],pp29[31],pp29[32],pp29[33],pp29[34],pp30[34],pp31[34],pp32[34],pp33[34],pp34[34],pp35[34],pp36[34],pp37[34],pp38[34],pp39[34],pp40[34],pp41[34],pp42[34],pp43[34],pp44[34],pp45[34],pp46[34],pp47[34]};
    CLA_36 KS_15(s15, c15, in15_1, in15_2);
    wire[33:0] s16, in16_1, in16_2;
    wire c16;
    assign in16_1 = {pp30[17],pp30[18],pp30[19],pp30[20],pp30[21],pp30[22],pp30[23],pp30[24],pp30[25],pp30[26],pp30[27],pp30[28],pp30[29],pp30[30],pp30[31],pp30[32],pp30[33],pp31[33],pp32[33],pp33[33],pp34[33],pp35[33],pp36[33],pp37[33],pp38[33],pp39[33],pp40[33],pp41[33],pp42[33],pp43[33],pp44[33],pp45[33],pp46[33],pp47[33]};
    assign in16_2 = {pp31[16],pp31[17],pp31[18],pp31[19],pp31[20],pp31[21],pp31[22],pp31[23],pp31[24],pp31[25],pp31[26],pp31[27],pp31[28],pp31[29],pp31[30],pp31[31],pp31[32],pp32[32],pp33[32],pp34[32],pp35[32],pp36[32],pp37[32],pp38[32],pp39[32],pp40[32],pp41[32],pp42[32],pp43[32],pp44[32],pp45[32],pp46[32],pp47[32],pp48[32]};
    CLA_34 KS_16(s16, c16, in16_1, in16_2);
    wire[31:0] s17, in17_1, in17_2;
    wire c17;
    assign in17_1 = {pp32[16],pp32[17],pp32[18],pp32[19],pp32[20],pp32[21],pp32[22],pp32[23],pp32[24],pp32[25],pp32[26],pp32[27],pp32[28],pp32[29],pp32[30],pp32[31],pp33[31],pp34[31],pp35[31],pp36[31],pp37[31],pp38[31],pp39[31],pp40[31],pp41[31],pp42[31],pp43[31],pp44[31],pp45[31],pp46[31],pp47[31],pp48[31]};
    assign in17_2 = {pp33[15],pp33[16],pp33[17],pp33[18],pp33[19],pp33[20],pp33[21],pp33[22],pp33[23],pp33[24],pp33[25],pp33[26],pp33[27],pp33[28],pp33[29],pp33[30],pp34[30],pp35[30],pp36[30],pp37[30],pp38[30],pp39[30],pp40[30],pp41[30],pp42[30],pp43[30],pp44[30],pp45[30],pp46[30],pp47[30],pp48[30],pp49[30]};
    CLA_32 KS_17(s17, c17, in17_1, in17_2);
    wire[29:0] s18, in18_1, in18_2;
    wire c18;
    assign in18_1 = {pp34[15],pp34[16],pp34[17],pp34[18],pp34[19],pp34[20],pp34[21],pp34[22],pp34[23],pp34[24],pp34[25],pp34[26],pp34[27],pp34[28],pp34[29],pp35[29],pp36[29],pp37[29],pp38[29],pp39[29],pp40[29],pp41[29],pp42[29],pp43[29],pp44[29],pp45[29],pp46[29],pp47[29],pp48[29],pp49[29]};
    assign in18_2 = {pp35[14],pp35[15],pp35[16],pp35[17],pp35[18],pp35[19],pp35[20],pp35[21],pp35[22],pp35[23],pp35[24],pp35[25],pp35[26],pp35[27],pp35[28],pp36[28],pp37[28],pp38[28],pp39[28],pp40[28],pp41[28],pp42[28],pp43[28],pp44[28],pp45[28],pp46[28],pp47[28],pp48[28],pp49[28],pp50[28]};
    CLA_30 KS_18(s18, c18, in18_1, in18_2);
    wire[27:0] s19, in19_1, in19_2;
    wire c19;
    assign in19_1 = {pp36[14],pp36[15],pp36[16],pp36[17],pp36[18],pp36[19],pp36[20],pp36[21],pp36[22],pp36[23],pp36[24],pp36[25],pp36[26],pp36[27],pp37[27],pp38[27],pp39[27],pp40[27],pp41[27],pp42[27],pp43[27],pp44[27],pp45[27],pp46[27],pp47[27],pp48[27],pp49[27],pp50[27]};
    assign in19_2 = {pp37[13],pp37[14],pp37[15],pp37[16],pp37[17],pp37[18],pp37[19],pp37[20],pp37[21],pp37[22],pp37[23],pp37[24],pp37[25],pp37[26],pp38[26],pp39[26],pp40[26],pp41[26],pp42[26],pp43[26],pp44[26],pp45[26],pp46[26],pp47[26],pp48[26],pp49[26],pp50[26],pp51[26]};
    CLA_28 KS_19(s19, c19, in19_1, in19_2);
    wire[25:0] s20, in20_1, in20_2;
    wire c20;
    assign in20_1 = {pp38[13],pp38[14],pp38[15],pp38[16],pp38[17],pp38[18],pp38[19],pp38[20],pp38[21],pp38[22],pp38[23],pp38[24],pp38[25],pp39[25],pp40[25],pp41[25],pp42[25],pp43[25],pp44[25],pp45[25],pp46[25],pp47[25],pp48[25],pp49[25],pp50[25],pp51[25]};
    assign in20_2 = {pp39[12],pp39[13],pp39[14],pp39[15],pp39[16],pp39[17],pp39[18],pp39[19],pp39[20],pp39[21],pp39[22],pp39[23],pp39[24],pp40[24],pp41[24],pp42[24],pp43[24],pp44[24],pp45[24],pp46[24],pp47[24],pp48[24],pp49[24],pp50[24],pp51[24],pp52[24]};
    CLA_26 KS_20(s20, c20, in20_1, in20_2);
    wire[23:0] s21, in21_1, in21_2;
    wire c21;
    assign in21_1 = {pp40[12],pp40[13],pp40[14],pp40[15],pp40[16],pp40[17],pp40[18],pp40[19],pp40[20],pp40[21],pp40[22],pp40[23],pp41[23],pp42[23],pp43[23],pp44[23],pp45[23],pp46[23],pp47[23],pp48[23],pp49[23],pp50[23],pp51[23],pp52[23]};
    assign in21_2 = {pp41[11],pp41[12],pp41[13],pp41[14],pp41[15],pp41[16],pp41[17],pp41[18],pp41[19],pp41[20],pp41[21],pp41[22],pp42[22],pp43[22],pp44[22],pp45[22],pp46[22],pp47[22],pp48[22],pp49[22],pp50[22],pp51[22],pp52[22],pp53[22]};
    CLA_24 KS_21(s21, c21, in21_1, in21_2);
    wire[21:0] s22, in22_1, in22_2;
    wire c22;
    assign in22_1 = {pp42[11],pp42[12],pp42[13],pp42[14],pp42[15],pp42[16],pp42[17],pp42[18],pp42[19],pp42[20],pp42[21],pp43[21],pp44[21],pp45[21],pp46[21],pp47[21],pp48[21],pp49[21],pp50[21],pp51[21],pp52[21],pp53[21]};
    assign in22_2 = {pp43[10],pp43[11],pp43[12],pp43[13],pp43[14],pp43[15],pp43[16],pp43[17],pp43[18],pp43[19],pp43[20],pp44[20],pp45[20],pp46[20],pp47[20],pp48[20],pp49[20],pp50[20],pp51[20],pp52[20],pp53[20],pp54[20]};
    CLA_22 KS_22(s22, c22, in22_1, in22_2);
    wire[19:0] s23, in23_1, in23_2;
    wire c23;
    assign in23_1 = {pp44[10],pp44[11],pp44[12],pp44[13],pp44[14],pp44[15],pp44[16],pp44[17],pp44[18],pp44[19],pp45[19],pp46[19],pp47[19],pp48[19],pp49[19],pp50[19],pp51[19],pp52[19],pp53[19],pp54[19]};
    assign in23_2 = {pp45[9],pp45[10],pp45[11],pp45[12],pp45[13],pp45[14],pp45[15],pp45[16],pp45[17],pp45[18],pp46[18],pp47[18],pp48[18],pp49[18],pp50[18],pp51[18],pp52[18],pp53[18],pp54[18],pp55[18]};
    CLA_20 KS_23(s23, c23, in23_1, in23_2);
    wire[17:0] s24, in24_1, in24_2;
    wire c24;
    assign in24_1 = {pp46[9],pp46[10],pp46[11],pp46[12],pp46[13],pp46[14],pp46[15],pp46[16],pp46[17],pp47[17],pp48[17],pp49[17],pp50[17],pp51[17],pp52[17],pp53[17],pp54[17],pp55[17]};
    assign in24_2 = {pp47[8],pp47[9],pp47[10],pp47[11],pp47[12],pp47[13],pp47[14],pp47[15],pp47[16],pp48[16],pp49[16],pp50[16],pp51[16],pp52[16],pp53[16],pp54[16],pp55[16],pp56[16]};
    CLA_18 KS_24(s24, c24, in24_1, in24_2);
    wire[15:0] s25, in25_1, in25_2;
    wire c25;
    assign in25_1 = {pp48[8],pp48[9],pp48[10],pp48[11],pp48[12],pp48[13],pp48[14],pp48[15],pp49[15],pp50[15],pp51[15],pp52[15],pp53[15],pp54[15],pp55[15],pp56[15]};
    assign in25_2 = {pp49[7],pp49[8],pp49[9],pp49[10],pp49[11],pp49[12],pp49[13],pp49[14],pp50[14],pp51[14],pp52[14],pp53[14],pp54[14],pp55[14],pp56[14],pp57[14]};
    CLA_16 KS_25(s25, c25, in25_1, in25_2);
    wire[13:0] s26, in26_1, in26_2;
    wire c26;
    assign in26_1 = {pp50[7],pp50[8],pp50[9],pp50[10],pp50[11],pp50[12],pp50[13],pp51[13],pp52[13],pp53[13],pp54[13],pp55[13],pp56[13],pp57[13]};
    assign in26_2 = {pp51[6],pp51[7],pp51[8],pp51[9],pp51[10],pp51[11],pp51[12],pp52[12],pp53[12],pp54[12],pp55[12],pp56[12],pp57[12],pp58[12]};
    CLA_14 KS_26(s26, c26, in26_1, in26_2);
    wire[11:0] s27, in27_1, in27_2;
    wire c27;
    assign in27_1 = {pp52[6],pp52[7],pp52[8],pp52[9],pp52[10],pp52[11],pp53[11],pp54[11],pp55[11],pp56[11],pp57[11],pp58[11]};
    assign in27_2 = {pp53[5],pp53[6],pp53[7],pp53[8],pp53[9],pp53[10],pp54[10],pp55[10],pp56[10],pp57[10],pp58[10],pp59[10]};
    CLA_12 KS_27(s27, c27, in27_1, in27_2);
    wire[9:0] s28, in28_1, in28_2;
    wire c28;
    assign in28_1 = {pp54[5],pp54[6],pp54[7],pp54[8],pp54[9],pp55[9],pp56[9],pp57[9],pp58[9],pp59[9]};
    assign in28_2 = {pp55[4],pp55[5],pp55[6],pp55[7],pp55[8],pp56[8],pp57[8],pp58[8],pp59[8],pp60[8]};
    CLA_10 KS_28(s28, c28, in28_1, in28_2);
    wire[7:0] s29, in29_1, in29_2;
    wire c29;
    assign in29_1 = {pp56[4],pp56[5],pp56[6],pp56[7],pp57[7],pp58[7],pp59[7],pp60[7]};
    assign in29_2 = {pp57[3],pp57[4],pp57[5],pp57[6],pp58[6],pp59[6],pp60[6],pp61[6]};
    CLA_8 KS_29(s29, c29, in29_1, in29_2);
    wire[5:0] s30, in30_1, in30_2;
    wire c30;
    assign in30_1 = {pp58[3],pp58[4],pp58[5],pp59[5],pp60[5],pp61[5]};
    assign in30_2 = {pp59[2],pp59[3],pp59[4],pp60[4],pp61[4],pp62[4]};
    CLA_6 KS_30(s30, c30, in30_1, in30_2);
    wire[3:0] s31, in31_1, in31_2;
    wire c31;
    assign in31_1 = {pp60[2],pp60[3],pp61[3],pp62[3]};
    assign in31_2 = {pp61[1],pp61[2],pp62[2],pp63[2]};
    CLA_4 KS_31(s31, c31, in31_1, in31_2);
    wire[1:0] s32, in32_1, in32_2;
    wire c32;
    assign in32_1 = {pp62[1],pp63[1]};
    assign in32_2 = {pp63[0],1'b0};
    CLA_2 KS_32(s32, c32, in32_1, in32_2);

    /*Stage 2*/
    wire[95:0] s33, in33_1, in33_2;
    wire c33;
    assign in33_1 = {pp0[16],pp0[17],pp0[18],pp0[19],pp0[20],pp0[21],pp0[22],pp0[23],pp0[24],pp0[25],pp0[26],pp0[27],pp0[28],pp0[29],pp0[30],pp0[31],pp2[30],pp4[29],pp6[28],pp8[27],pp10[26],pp12[25],pp14[24],pp16[23],pp18[22],pp20[21],pp22[20],pp24[19],pp26[18],pp28[17],pp30[16],pp32[15],pp34[14],pp36[13],pp38[12],pp40[11],pp42[10],pp44[9],pp46[8],pp48[7],pp50[6],pp52[5],pp54[4],pp56[3],pp58[2],pp60[1],pp62[0],s1[31],s1[32],s1[33],pp63[3],pp62[5],pp61[7],pp60[9],pp59[11],pp58[13],pp57[15],pp56[17],pp55[19],pp54[21],pp53[23],pp52[25],pp51[27],pp50[29],pp49[31],pp48[33],pp47[35],pp46[37],pp45[39],pp44[41],pp43[43],pp42[45],pp41[47],pp40[49],pp39[51],pp38[53],pp37[55],pp36[57],pp35[59],pp34[61],pp33[63],pp34[63],pp35[63],pp36[63],pp37[63],pp38[63],pp39[63],pp40[63],pp41[63],pp42[63],pp43[63],pp44[63],pp45[63],pp46[63],pp47[63],pp48[63]};
    assign in33_2 = {pp1[15],pp1[16],pp1[17],pp1[18],pp1[19],pp1[20],pp1[21],pp1[22],pp1[23],pp1[24],pp1[25],pp1[26],pp1[27],pp1[28],pp1[29],pp1[30],pp3[29],pp5[28],pp7[27],pp9[26],pp11[25],pp13[24],pp15[23],pp17[22],pp19[21],pp21[20],pp23[19],pp25[18],pp27[17],pp29[16],pp31[15],pp33[14],pp35[13],pp37[12],pp39[11],pp41[10],pp43[9],pp45[8],pp47[7],pp49[6],pp51[5],pp53[4],pp55[3],pp57[2],pp59[1],pp61[0],s1[30],s2[30],s2[31],s2[32],s1[34],pp63[4],pp62[6],pp61[8],pp60[10],pp59[12],pp58[14],pp57[16],pp56[18],pp55[20],pp54[22],pp53[24],pp52[26],pp51[28],pp50[30],pp49[32],pp48[34],pp47[36],pp46[38],pp45[40],pp44[42],pp43[44],pp42[46],pp41[48],pp40[50],pp39[52],pp38[54],pp37[56],pp36[58],pp35[60],pp34[62],pp35[62],pp36[62],pp37[62],pp38[62],pp39[62],pp40[62],pp41[62],pp42[62],pp43[62],pp44[62],pp45[62],pp46[62],pp47[62],pp48[62],pp49[62]};
    CLA_96 KS_33(s33, c33, in33_1, in33_2);
    wire[93:0] s34, in34_1, in34_2;
    wire c34;
    assign in34_1 = {pp2[15],pp2[16],pp2[17],pp2[18],pp2[19],pp2[20],pp2[21],pp2[22],pp2[23],pp2[24],pp2[25],pp2[26],pp2[27],pp2[28],pp2[29],pp4[28],pp6[27],pp8[26],pp10[25],pp12[24],pp14[23],pp16[22],pp18[21],pp20[20],pp22[19],pp24[18],pp26[17],pp28[16],pp30[15],pp32[14],pp34[13],pp36[12],pp38[11],pp40[10],pp42[9],pp44[8],pp46[7],pp48[6],pp50[5],pp52[4],pp54[3],pp56[2],pp58[1],pp60[0],s1[29],s2[29],s3[29],s3[30],s3[31],s2[33],s1[35],pp63[5],pp62[7],pp61[9],pp60[11],pp59[13],pp58[15],pp57[17],pp56[19],pp55[21],pp54[23],pp53[25],pp52[27],pp51[29],pp50[31],pp49[33],pp48[35],pp47[37],pp46[39],pp45[41],pp44[43],pp43[45],pp42[47],pp41[49],pp40[51],pp39[53],pp38[55],pp37[57],pp36[59],pp35[61],pp36[61],pp37[61],pp38[61],pp39[61],pp40[61],pp41[61],pp42[61],pp43[61],pp44[61],pp45[61],pp46[61],pp47[61],pp48[61],pp49[61]};
    assign in34_2 = {pp3[14],pp3[15],pp3[16],pp3[17],pp3[18],pp3[19],pp3[20],pp3[21],pp3[22],pp3[23],pp3[24],pp3[25],pp3[26],pp3[27],pp3[28],pp5[27],pp7[26],pp9[25],pp11[24],pp13[23],pp15[22],pp17[21],pp19[20],pp21[19],pp23[18],pp25[17],pp27[16],pp29[15],pp31[14],pp33[13],pp35[12],pp37[11],pp39[10],pp41[9],pp43[8],pp45[7],pp47[6],pp49[5],pp51[4],pp53[3],pp55[2],pp57[1],pp59[0],s1[28],s2[28],s3[28],s4[28],s4[29],s4[30],s3[32],s2[34],s1[36],pp63[6],pp62[8],pp61[10],pp60[12],pp59[14],pp58[16],pp57[18],pp56[20],pp55[22],pp54[24],pp53[26],pp52[28],pp51[30],pp50[32],pp49[34],pp48[36],pp47[38],pp46[40],pp45[42],pp44[44],pp43[46],pp42[48],pp41[50],pp40[52],pp39[54],pp38[56],pp37[58],pp36[60],pp37[60],pp38[60],pp39[60],pp40[60],pp41[60],pp42[60],pp43[60],pp44[60],pp45[60],pp46[60],pp47[60],pp48[60],pp49[60],pp50[60]};
    CLA_94 KS_34(s34, c34, in34_1, in34_2);
    wire[91:0] s35, in35_1, in35_2;
    wire c35;
    assign in35_1 = {pp4[14],pp4[15],pp4[16],pp4[17],pp4[18],pp4[19],pp4[20],pp4[21],pp4[22],pp4[23],pp4[24],pp4[25],pp4[26],pp4[27],pp6[26],pp8[25],pp10[24],pp12[23],pp14[22],pp16[21],pp18[20],pp20[19],pp22[18],pp24[17],pp26[16],pp28[15],pp30[14],pp32[13],pp34[12],pp36[11],pp38[10],pp40[9],pp42[8],pp44[7],pp46[6],pp48[5],pp50[4],pp52[3],pp54[2],pp56[1],pp58[0],s1[27],s2[27],s3[27],s4[27],s5[27],s5[28],s5[29],s4[31],s3[33],s2[35],s1[37],pp63[7],pp62[9],pp61[11],pp60[13],pp59[15],pp58[17],pp57[19],pp56[21],pp55[23],pp54[25],pp53[27],pp52[29],pp51[31],pp50[33],pp49[35],pp48[37],pp47[39],pp46[41],pp45[43],pp44[45],pp43[47],pp42[49],pp41[51],pp40[53],pp39[55],pp38[57],pp37[59],pp38[59],pp39[59],pp40[59],pp41[59],pp42[59],pp43[59],pp44[59],pp45[59],pp46[59],pp47[59],pp48[59],pp49[59],pp50[59]};
    assign in35_2 = {pp5[13],pp5[14],pp5[15],pp5[16],pp5[17],pp5[18],pp5[19],pp5[20],pp5[21],pp5[22],pp5[23],pp5[24],pp5[25],pp5[26],pp7[25],pp9[24],pp11[23],pp13[22],pp15[21],pp17[20],pp19[19],pp21[18],pp23[17],pp25[16],pp27[15],pp29[14],pp31[13],pp33[12],pp35[11],pp37[10],pp39[9],pp41[8],pp43[7],pp45[6],pp47[5],pp49[4],pp51[3],pp53[2],pp55[1],pp57[0],s1[26],s2[26],s3[26],s4[26],s5[26],s6[26],s6[27],s6[28],s5[30],s4[32],s3[34],s2[36],s1[38],pp63[8],pp62[10],pp61[12],pp60[14],pp59[16],pp58[18],pp57[20],pp56[22],pp55[24],pp54[26],pp53[28],pp52[30],pp51[32],pp50[34],pp49[36],pp48[38],pp47[40],pp46[42],pp45[44],pp44[46],pp43[48],pp42[50],pp41[52],pp40[54],pp39[56],pp38[58],pp39[58],pp40[58],pp41[58],pp42[58],pp43[58],pp44[58],pp45[58],pp46[58],pp47[58],pp48[58],pp49[58],pp50[58],pp51[58]};
    CLA_92 KS_35(s35, c35, in35_1, in35_2);
    wire[89:0] s36, in36_1, in36_2;
    wire c36;
    assign in36_1 = {pp6[13],pp6[14],pp6[15],pp6[16],pp6[17],pp6[18],pp6[19],pp6[20],pp6[21],pp6[22],pp6[23],pp6[24],pp6[25],pp8[24],pp10[23],pp12[22],pp14[21],pp16[20],pp18[19],pp20[18],pp22[17],pp24[16],pp26[15],pp28[14],pp30[13],pp32[12],pp34[11],pp36[10],pp38[9],pp40[8],pp42[7],pp44[6],pp46[5],pp48[4],pp50[3],pp52[2],pp54[1],pp56[0],s1[25],s2[25],s3[25],s4[25],s5[25],s6[25],s7[25],s7[26],s7[27],s6[29],s5[31],s4[33],s3[35],s2[37],s1[39],pp63[9],pp62[11],pp61[13],pp60[15],pp59[17],pp58[19],pp57[21],pp56[23],pp55[25],pp54[27],pp53[29],pp52[31],pp51[33],pp50[35],pp49[37],pp48[39],pp47[41],pp46[43],pp45[45],pp44[47],pp43[49],pp42[51],pp41[53],pp40[55],pp39[57],pp40[57],pp41[57],pp42[57],pp43[57],pp44[57],pp45[57],pp46[57],pp47[57],pp48[57],pp49[57],pp50[57],pp51[57]};
    assign in36_2 = {pp7[12],pp7[13],pp7[14],pp7[15],pp7[16],pp7[17],pp7[18],pp7[19],pp7[20],pp7[21],pp7[22],pp7[23],pp7[24],pp9[23],pp11[22],pp13[21],pp15[20],pp17[19],pp19[18],pp21[17],pp23[16],pp25[15],pp27[14],pp29[13],pp31[12],pp33[11],pp35[10],pp37[9],pp39[8],pp41[7],pp43[6],pp45[5],pp47[4],pp49[3],pp51[2],pp53[1],pp55[0],s1[24],s2[24],s3[24],s4[24],s5[24],s6[24],s7[24],s8[24],s8[25],s8[26],s7[28],s6[30],s5[32],s4[34],s3[36],s2[38],s1[40],pp63[10],pp62[12],pp61[14],pp60[16],pp59[18],pp58[20],pp57[22],pp56[24],pp55[26],pp54[28],pp53[30],pp52[32],pp51[34],pp50[36],pp49[38],pp48[40],pp47[42],pp46[44],pp45[46],pp44[48],pp43[50],pp42[52],pp41[54],pp40[56],pp41[56],pp42[56],pp43[56],pp44[56],pp45[56],pp46[56],pp47[56],pp48[56],pp49[56],pp50[56],pp51[56],pp52[56]};
    CLA_90 KS_36(s36, c36, in36_1, in36_2);
    wire[87:0] s37, in37_1, in37_2;
    wire c37;
    assign in37_1 = {pp8[12],pp8[13],pp8[14],pp8[15],pp8[16],pp8[17],pp8[18],pp8[19],pp8[20],pp8[21],pp8[22],pp8[23],pp10[22],pp12[21],pp14[20],pp16[19],pp18[18],pp20[17],pp22[16],pp24[15],pp26[14],pp28[13],pp30[12],pp32[11],pp34[10],pp36[9],pp38[8],pp40[7],pp42[6],pp44[5],pp46[4],pp48[3],pp50[2],pp52[1],pp54[0],s1[23],s2[23],s3[23],s4[23],s5[23],s6[23],s7[23],s8[23],s9[23],s9[24],s9[25],s8[27],s7[29],s6[31],s5[33],s4[35],s3[37],s2[39],s1[41],pp63[11],pp62[13],pp61[15],pp60[17],pp59[19],pp58[21],pp57[23],pp56[25],pp55[27],pp54[29],pp53[31],pp52[33],pp51[35],pp50[37],pp49[39],pp48[41],pp47[43],pp46[45],pp45[47],pp44[49],pp43[51],pp42[53],pp41[55],pp42[55],pp43[55],pp44[55],pp45[55],pp46[55],pp47[55],pp48[55],pp49[55],pp50[55],pp51[55],pp52[55]};
    assign in37_2 = {pp9[11],pp9[12],pp9[13],pp9[14],pp9[15],pp9[16],pp9[17],pp9[18],pp9[19],pp9[20],pp9[21],pp9[22],pp11[21],pp13[20],pp15[19],pp17[18],pp19[17],pp21[16],pp23[15],pp25[14],pp27[13],pp29[12],pp31[11],pp33[10],pp35[9],pp37[8],pp39[7],pp41[6],pp43[5],pp45[4],pp47[3],pp49[2],pp51[1],pp53[0],s1[22],s2[22],s3[22],s4[22],s5[22],s6[22],s7[22],s8[22],s9[22],s10[22],s10[23],s10[24],s9[26],s8[28],s7[30],s6[32],s5[34],s4[36],s3[38],s2[40],s1[42],pp63[12],pp62[14],pp61[16],pp60[18],pp59[20],pp58[22],pp57[24],pp56[26],pp55[28],pp54[30],pp53[32],pp52[34],pp51[36],pp50[38],pp49[40],pp48[42],pp47[44],pp46[46],pp45[48],pp44[50],pp43[52],pp42[54],pp43[54],pp44[54],pp45[54],pp46[54],pp47[54],pp48[54],pp49[54],pp50[54],pp51[54],pp52[54],pp53[54]};
    CLA_88 KS_37(s37, c37, in37_1, in37_2);
    wire[85:0] s38, in38_1, in38_2;
    wire c38;
    assign in38_1 = {pp10[11],pp10[12],pp10[13],pp10[14],pp10[15],pp10[16],pp10[17],pp10[18],pp10[19],pp10[20],pp10[21],pp12[20],pp14[19],pp16[18],pp18[17],pp20[16],pp22[15],pp24[14],pp26[13],pp28[12],pp30[11],pp32[10],pp34[9],pp36[8],pp38[7],pp40[6],pp42[5],pp44[4],pp46[3],pp48[2],pp50[1],pp52[0],s1[21],s2[21],s3[21],s4[21],s5[21],s6[21],s7[21],s8[21],s9[21],s10[21],s11[21],s11[22],s11[23],s10[25],s9[27],s8[29],s7[31],s6[33],s5[35],s4[37],s3[39],s2[41],s1[43],pp63[13],pp62[15],pp61[17],pp60[19],pp59[21],pp58[23],pp57[25],pp56[27],pp55[29],pp54[31],pp53[33],pp52[35],pp51[37],pp50[39],pp49[41],pp48[43],pp47[45],pp46[47],pp45[49],pp44[51],pp43[53],pp44[53],pp45[53],pp46[53],pp47[53],pp48[53],pp49[53],pp50[53],pp51[53],pp52[53],pp53[53]};
    assign in38_2 = {pp11[10],pp11[11],pp11[12],pp11[13],pp11[14],pp11[15],pp11[16],pp11[17],pp11[18],pp11[19],pp11[20],pp13[19],pp15[18],pp17[17],pp19[16],pp21[15],pp23[14],pp25[13],pp27[12],pp29[11],pp31[10],pp33[9],pp35[8],pp37[7],pp39[6],pp41[5],pp43[4],pp45[3],pp47[2],pp49[1],pp51[0],s1[20],s2[20],s3[20],s4[20],s5[20],s6[20],s7[20],s8[20],s9[20],s10[20],s11[20],s12[20],s12[21],s12[22],s11[24],s10[26],s9[28],s8[30],s7[32],s6[34],s5[36],s4[38],s3[40],s2[42],s1[44],pp63[14],pp62[16],pp61[18],pp60[20],pp59[22],pp58[24],pp57[26],pp56[28],pp55[30],pp54[32],pp53[34],pp52[36],pp51[38],pp50[40],pp49[42],pp48[44],pp47[46],pp46[48],pp45[50],pp44[52],pp45[52],pp46[52],pp47[52],pp48[52],pp49[52],pp50[52],pp51[52],pp52[52],pp53[52],pp54[52]};
    CLA_86 KS_38(s38, c38, in38_1, in38_2);
    wire[83:0] s39, in39_1, in39_2;
    wire c39;
    assign in39_1 = {pp12[10],pp12[11],pp12[12],pp12[13],pp12[14],pp12[15],pp12[16],pp12[17],pp12[18],pp12[19],pp14[18],pp16[17],pp18[16],pp20[15],pp22[14],pp24[13],pp26[12],pp28[11],pp30[10],pp32[9],pp34[8],pp36[7],pp38[6],pp40[5],pp42[4],pp44[3],pp46[2],pp48[1],pp50[0],s1[19],s2[19],s3[19],s4[19],s5[19],s6[19],s7[19],s8[19],s9[19],s10[19],s11[19],s12[19],s13[19],s13[20],s13[21],s12[23],s11[25],s10[27],s9[29],s8[31],s7[33],s6[35],s5[37],s4[39],s3[41],s2[43],s1[45],pp63[15],pp62[17],pp61[19],pp60[21],pp59[23],pp58[25],pp57[27],pp56[29],pp55[31],pp54[33],pp53[35],pp52[37],pp51[39],pp50[41],pp49[43],pp48[45],pp47[47],pp46[49],pp45[51],pp46[51],pp47[51],pp48[51],pp49[51],pp50[51],pp51[51],pp52[51],pp53[51],pp54[51]};
    assign in39_2 = {pp13[9],pp13[10],pp13[11],pp13[12],pp13[13],pp13[14],pp13[15],pp13[16],pp13[17],pp13[18],pp15[17],pp17[16],pp19[15],pp21[14],pp23[13],pp25[12],pp27[11],pp29[10],pp31[9],pp33[8],pp35[7],pp37[6],pp39[5],pp41[4],pp43[3],pp45[2],pp47[1],pp49[0],s1[18],s2[18],s3[18],s4[18],s5[18],s6[18],s7[18],s8[18],s9[18],s10[18],s11[18],s12[18],s13[18],s14[18],s14[19],s14[20],s13[22],s12[24],s11[26],s10[28],s9[30],s8[32],s7[34],s6[36],s5[38],s4[40],s3[42],s2[44],s1[46],pp63[16],pp62[18],pp61[20],pp60[22],pp59[24],pp58[26],pp57[28],pp56[30],pp55[32],pp54[34],pp53[36],pp52[38],pp51[40],pp50[42],pp49[44],pp48[46],pp47[48],pp46[50],pp47[50],pp48[50],pp49[50],pp50[50],pp51[50],pp52[50],pp53[50],pp54[50],pp55[50]};
    CLA_84 KS_39(s39, c39, in39_1, in39_2);
    wire[81:0] s40, in40_1, in40_2;
    wire c40;
    assign in40_1 = {pp14[9],pp14[10],pp14[11],pp14[12],pp14[13],pp14[14],pp14[15],pp14[16],pp14[17],pp16[16],pp18[15],pp20[14],pp22[13],pp24[12],pp26[11],pp28[10],pp30[9],pp32[8],pp34[7],pp36[6],pp38[5],pp40[4],pp42[3],pp44[2],pp46[1],pp48[0],s1[17],s2[17],s3[17],s4[17],s5[17],s6[17],s7[17],s8[17],s9[17],s10[17],s11[17],s12[17],s13[17],s14[17],s15[17],s15[18],s15[19],s14[21],s13[23],s12[25],s11[27],s10[29],s9[31],s8[33],s7[35],s6[37],s5[39],s4[41],s3[43],s2[45],s1[47],pp63[17],pp62[19],pp61[21],pp60[23],pp59[25],pp58[27],pp57[29],pp56[31],pp55[33],pp54[35],pp53[37],pp52[39],pp51[41],pp50[43],pp49[45],pp48[47],pp47[49],pp48[49],pp49[49],pp50[49],pp51[49],pp52[49],pp53[49],pp54[49],pp55[49]};
    assign in40_2 = {pp15[8],pp15[9],pp15[10],pp15[11],pp15[12],pp15[13],pp15[14],pp15[15],pp15[16],pp17[15],pp19[14],pp21[13],pp23[12],pp25[11],pp27[10],pp29[9],pp31[8],pp33[7],pp35[6],pp37[5],pp39[4],pp41[3],pp43[2],pp45[1],pp47[0],s1[16],s2[16],s3[16],s4[16],s5[16],s6[16],s7[16],s8[16],s9[16],s10[16],s11[16],s12[16],s13[16],s14[16],s15[16],s16[16],s16[17],s16[18],s15[20],s14[22],s13[24],s12[26],s11[28],s10[30],s9[32],s8[34],s7[36],s6[38],s5[40],s4[42],s3[44],s2[46],s1[48],pp63[18],pp62[20],pp61[22],pp60[24],pp59[26],pp58[28],pp57[30],pp56[32],pp55[34],pp54[36],pp53[38],pp52[40],pp51[42],pp50[44],pp49[46],pp48[48],pp49[48],pp50[48],pp51[48],pp52[48],pp53[48],pp54[48],pp55[48],pp56[48]};
    CLA_82 KS_40(s40, c40, in40_1, in40_2);
    wire[79:0] s41, in41_1, in41_2;
    wire c41;
    assign in41_1 = {pp16[8],pp16[9],pp16[10],pp16[11],pp16[12],pp16[13],pp16[14],pp16[15],pp18[14],pp20[13],pp22[12],pp24[11],pp26[10],pp28[9],pp30[8],pp32[7],pp34[6],pp36[5],pp38[4],pp40[3],pp42[2],pp44[1],pp46[0],s1[15],s2[15],s3[15],s4[15],s5[15],s6[15],s7[15],s8[15],s9[15],s10[15],s11[15],s12[15],s13[15],s14[15],s15[15],s16[15],s17[15],s17[16],s17[17],s16[19],s15[21],s14[23],s13[25],s12[27],s11[29],s10[31],s9[33],s8[35],s7[37],s6[39],s5[41],s4[43],s3[45],s2[47],s1[49],pp63[19],pp62[21],pp61[23],pp60[25],pp59[27],pp58[29],pp57[31],pp56[33],pp55[35],pp54[37],pp53[39],pp52[41],pp51[43],pp50[45],pp49[47],pp50[47],pp51[47],pp52[47],pp53[47],pp54[47],pp55[47],pp56[47]};
    assign in41_2 = {pp17[7],pp17[8],pp17[9],pp17[10],pp17[11],pp17[12],pp17[13],pp17[14],pp19[13],pp21[12],pp23[11],pp25[10],pp27[9],pp29[8],pp31[7],pp33[6],pp35[5],pp37[4],pp39[3],pp41[2],pp43[1],pp45[0],s1[14],s2[14],s3[14],s4[14],s5[14],s6[14],s7[14],s8[14],s9[14],s10[14],s11[14],s12[14],s13[14],s14[14],s15[14],s16[14],s17[14],s18[14],s18[15],s18[16],s17[18],s16[20],s15[22],s14[24],s13[26],s12[28],s11[30],s10[32],s9[34],s8[36],s7[38],s6[40],s5[42],s4[44],s3[46],s2[48],s1[50],pp63[20],pp62[22],pp61[24],pp60[26],pp59[28],pp58[30],pp57[32],pp56[34],pp55[36],pp54[38],pp53[40],pp52[42],pp51[44],pp50[46],pp51[46],pp52[46],pp53[46],pp54[46],pp55[46],pp56[46],pp57[46]};
    CLA_80 KS_41(s41, c41, in41_1, in41_2);
    wire[77:0] s42, in42_1, in42_2;
    wire c42;
    assign in42_1 = {pp18[7],pp18[8],pp18[9],pp18[10],pp18[11],pp18[12],pp18[13],pp20[12],pp22[11],pp24[10],pp26[9],pp28[8],pp30[7],pp32[6],pp34[5],pp36[4],pp38[3],pp40[2],pp42[1],pp44[0],s1[13],s2[13],s3[13],s4[13],s5[13],s6[13],s7[13],s8[13],s9[13],s10[13],s11[13],s12[13],s13[13],s14[13],s15[13],s16[13],s17[13],s18[13],s19[13],s19[14],s19[15],s18[17],s17[19],s16[21],s15[23],s14[25],s13[27],s12[29],s11[31],s10[33],s9[35],s8[37],s7[39],s6[41],s5[43],s4[45],s3[47],s2[49],s1[51],pp63[21],pp62[23],pp61[25],pp60[27],pp59[29],pp58[31],pp57[33],pp56[35],pp55[37],pp54[39],pp53[41],pp52[43],pp51[45],pp52[45],pp53[45],pp54[45],pp55[45],pp56[45],pp57[45]};
    assign in42_2 = {pp19[6],pp19[7],pp19[8],pp19[9],pp19[10],pp19[11],pp19[12],pp21[11],pp23[10],pp25[9],pp27[8],pp29[7],pp31[6],pp33[5],pp35[4],pp37[3],pp39[2],pp41[1],pp43[0],s1[12],s2[12],s3[12],s4[12],s5[12],s6[12],s7[12],s8[12],s9[12],s10[12],s11[12],s12[12],s13[12],s14[12],s15[12],s16[12],s17[12],s18[12],s19[12],s20[12],s20[13],s20[14],s19[16],s18[18],s17[20],s16[22],s15[24],s14[26],s13[28],s12[30],s11[32],s10[34],s9[36],s8[38],s7[40],s6[42],s5[44],s4[46],s3[48],s2[50],s1[52],pp63[22],pp62[24],pp61[26],pp60[28],pp59[30],pp58[32],pp57[34],pp56[36],pp55[38],pp54[40],pp53[42],pp52[44],pp53[44],pp54[44],pp55[44],pp56[44],pp57[44],pp58[44]};
    CLA_78 KS_42(s42, c42, in42_1, in42_2);
    wire[75:0] s43, in43_1, in43_2;
    wire c43;
    assign in43_1 = {pp20[6],pp20[7],pp20[8],pp20[9],pp20[10],pp20[11],pp22[10],pp24[9],pp26[8],pp28[7],pp30[6],pp32[5],pp34[4],pp36[3],pp38[2],pp40[1],pp42[0],s1[11],s2[11],s3[11],s4[11],s5[11],s6[11],s7[11],s8[11],s9[11],s10[11],s11[11],s12[11],s13[11],s14[11],s15[11],s16[11],s17[11],s18[11],s19[11],s20[11],s21[11],s21[12],s21[13],s20[15],s19[17],s18[19],s17[21],s16[23],s15[25],s14[27],s13[29],s12[31],s11[33],s10[35],s9[37],s8[39],s7[41],s6[43],s5[45],s4[47],s3[49],s2[51],s1[53],pp63[23],pp62[25],pp61[27],pp60[29],pp59[31],pp58[33],pp57[35],pp56[37],pp55[39],pp54[41],pp53[43],pp54[43],pp55[43],pp56[43],pp57[43],pp58[43]};
    assign in43_2 = {pp21[5],pp21[6],pp21[7],pp21[8],pp21[9],pp21[10],pp23[9],pp25[8],pp27[7],pp29[6],pp31[5],pp33[4],pp35[3],pp37[2],pp39[1],pp41[0],s1[10],s2[10],s3[10],s4[10],s5[10],s6[10],s7[10],s8[10],s9[10],s10[10],s11[10],s12[10],s13[10],s14[10],s15[10],s16[10],s17[10],s18[10],s19[10],s20[10],s21[10],s22[10],s22[11],s22[12],s21[14],s20[16],s19[18],s18[20],s17[22],s16[24],s15[26],s14[28],s13[30],s12[32],s11[34],s10[36],s9[38],s8[40],s7[42],s6[44],s5[46],s4[48],s3[50],s2[52],s1[54],pp63[24],pp62[26],pp61[28],pp60[30],pp59[32],pp58[34],pp57[36],pp56[38],pp55[40],pp54[42],pp55[42],pp56[42],pp57[42],pp58[42],pp59[42]};
    CLA_76 KS_43(s43, c43, in43_1, in43_2);
    wire[73:0] s44, in44_1, in44_2;
    wire c44;
    assign in44_1 = {pp22[5],pp22[6],pp22[7],pp22[8],pp22[9],pp24[8],pp26[7],pp28[6],pp30[5],pp32[4],pp34[3],pp36[2],pp38[1],pp40[0],s1[9],s2[9],s3[9],s4[9],s5[9],s6[9],s7[9],s8[9],s9[9],s10[9],s11[9],s12[9],s13[9],s14[9],s15[9],s16[9],s17[9],s18[9],s19[9],s20[9],s21[9],s22[9],s23[9],s23[10],s23[11],s22[13],s21[15],s20[17],s19[19],s18[21],s17[23],s16[25],s15[27],s14[29],s13[31],s12[33],s11[35],s10[37],s9[39],s8[41],s7[43],s6[45],s5[47],s4[49],s3[51],s2[53],s1[55],pp63[25],pp62[27],pp61[29],pp60[31],pp59[33],pp58[35],pp57[37],pp56[39],pp55[41],pp56[41],pp57[41],pp58[41],pp59[41]};
    assign in44_2 = {pp23[4],pp23[5],pp23[6],pp23[7],pp23[8],pp25[7],pp27[6],pp29[5],pp31[4],pp33[3],pp35[2],pp37[1],pp39[0],s1[8],s2[8],s3[8],s4[8],s5[8],s6[8],s7[8],s8[8],s9[8],s10[8],s11[8],s12[8],s13[8],s14[8],s15[8],s16[8],s17[8],s18[8],s19[8],s20[8],s21[8],s22[8],s23[8],s24[8],s24[9],s24[10],s23[12],s22[14],s21[16],s20[18],s19[20],s18[22],s17[24],s16[26],s15[28],s14[30],s13[32],s12[34],s11[36],s10[38],s9[40],s8[42],s7[44],s6[46],s5[48],s4[50],s3[52],s2[54],s1[56],pp63[26],pp62[28],pp61[30],pp60[32],pp59[34],pp58[36],pp57[38],pp56[40],pp57[40],pp58[40],pp59[40],pp60[40]};
    CLA_74 KS_44(s44, c44, in44_1, in44_2);
    wire[71:0] s45, in45_1, in45_2;
    wire c45;
    assign in45_1 = {pp24[4],pp24[5],pp24[6],pp24[7],pp26[6],pp28[5],pp30[4],pp32[3],pp34[2],pp36[1],pp38[0],s1[7],s2[7],s3[7],s4[7],s5[7],s6[7],s7[7],s8[7],s9[7],s10[7],s11[7],s12[7],s13[7],s14[7],s15[7],s16[7],s17[7],s18[7],s19[7],s20[7],s21[7],s22[7],s23[7],s24[7],s25[7],s25[8],s25[9],s24[11],s23[13],s22[15],s21[17],s20[19],s19[21],s18[23],s17[25],s16[27],s15[29],s14[31],s13[33],s12[35],s11[37],s10[39],s9[41],s8[43],s7[45],s6[47],s5[49],s4[51],s3[53],s2[55],s1[57],pp63[27],pp62[29],pp61[31],pp60[33],pp59[35],pp58[37],pp57[39],pp58[39],pp59[39],pp60[39]};
    assign in45_2 = {pp25[3],pp25[4],pp25[5],pp25[6],pp27[5],pp29[4],pp31[3],pp33[2],pp35[1],pp37[0],s1[6],s2[6],s3[6],s4[6],s5[6],s6[6],s7[6],s8[6],s9[6],s10[6],s11[6],s12[6],s13[6],s14[6],s15[6],s16[6],s17[6],s18[6],s19[6],s20[6],s21[6],s22[6],s23[6],s24[6],s25[6],s26[6],s26[7],s26[8],s25[10],s24[12],s23[14],s22[16],s21[18],s20[20],s19[22],s18[24],s17[26],s16[28],s15[30],s14[32],s13[34],s12[36],s11[38],s10[40],s9[42],s8[44],s7[46],s6[48],s5[50],s4[52],s3[54],s2[56],s1[58],pp63[28],pp62[30],pp61[32],pp60[34],pp59[36],pp58[38],pp59[38],pp60[38],pp61[38]};
    CLA_72 KS_45(s45, c45, in45_1, in45_2);
    wire[69:0] s46, in46_1, in46_2;
    wire c46;
    assign in46_1 = {pp26[3],pp26[4],pp26[5],pp28[4],pp30[3],pp32[2],pp34[1],pp36[0],s1[5],s2[5],s3[5],s4[5],s5[5],s6[5],s7[5],s8[5],s9[5],s10[5],s11[5],s12[5],s13[5],s14[5],s15[5],s16[5],s17[5],s18[5],s19[5],s20[5],s21[5],s22[5],s23[5],s24[5],s25[5],s26[5],s27[5],s27[6],s27[7],s26[9],s25[11],s24[13],s23[15],s22[17],s21[19],s20[21],s19[23],s18[25],s17[27],s16[29],s15[31],s14[33],s13[35],s12[37],s11[39],s10[41],s9[43],s8[45],s7[47],s6[49],s5[51],s4[53],s3[55],s2[57],s1[59],pp63[29],pp62[31],pp61[33],pp60[35],pp59[37],pp60[37],pp61[37]};
    assign in46_2 = {pp27[2],pp27[3],pp27[4],pp29[3],pp31[2],pp33[1],pp35[0],s1[4],s2[4],s3[4],s4[4],s5[4],s6[4],s7[4],s8[4],s9[4],s10[4],s11[4],s12[4],s13[4],s14[4],s15[4],s16[4],s17[4],s18[4],s19[4],s20[4],s21[4],s22[4],s23[4],s24[4],s25[4],s26[4],s27[4],s28[4],s28[5],s28[6],s27[8],s26[10],s25[12],s24[14],s23[16],s22[18],s21[20],s20[22],s19[24],s18[26],s17[28],s16[30],s15[32],s14[34],s13[36],s12[38],s11[40],s10[42],s9[44],s8[46],s7[48],s6[50],s5[52],s4[54],s3[56],s2[58],s1[60],pp63[30],pp62[32],pp61[34],pp60[36],pp61[36],pp62[36]};
    CLA_70 KS_46(s46, c46, in46_1, in46_2);
    wire[67:0] s47, in47_1, in47_2;
    wire c47;
    assign in47_1 = {pp28[2],pp28[3],pp30[2],pp32[1],pp34[0],s1[3],s2[3],s3[3],s4[3],s5[3],s6[3],s7[3],s8[3],s9[3],s10[3],s11[3],s12[3],s13[3],s14[3],s15[3],s16[3],s17[3],s18[3],s19[3],s20[3],s21[3],s22[3],s23[3],s24[3],s25[3],s26[3],s27[3],s28[3],s29[3],s29[4],s29[5],s28[7],s27[9],s26[11],s25[13],s24[15],s23[17],s22[19],s21[21],s20[23],s19[25],s18[27],s17[29],s16[31],s15[33],s14[35],s13[37],s12[39],s11[41],s10[43],s9[45],s8[47],s7[49],s6[51],s5[53],s4[55],s3[57],s2[59],s1[61],pp63[31],pp62[33],pp61[35],pp62[35]};
    assign in47_2 = {pp29[1],pp29[2],pp31[1],pp33[0],s1[2],s2[2],s3[2],s4[2],s5[2],s6[2],s7[2],s8[2],s9[2],s10[2],s11[2],s12[2],s13[2],s14[2],s15[2],s16[2],s17[2],s18[2],s19[2],s20[2],s21[2],s22[2],s23[2],s24[2],s25[2],s26[2],s27[2],s28[2],s29[2],s30[2],s30[3],s30[4],s29[6],s28[8],s27[10],s26[12],s25[14],s24[16],s23[18],s22[20],s21[22],s20[24],s19[26],s18[28],s17[30],s16[32],s15[34],s14[36],s13[38],s12[40],s11[42],s10[44],s9[46],s8[48],s7[50],s6[52],s5[54],s4[56],s3[58],s2[60],s1[62],pp63[32],pp62[34],pp63[34]};
    CLA_68 KS_47(s47, c47, in47_1, in47_2);
    wire[65:0] s48, in48_1, in48_2;
    wire c48;
    assign in48_1 = {pp30[1],pp32[0],s1[1],s2[1],s3[1],s4[1],s5[1],s6[1],s7[1],s8[1],s9[1],s10[1],s11[1],s12[1],s13[1],s14[1],s15[1],s16[1],s17[1],s18[1],s19[1],s20[1],s21[1],s22[1],s23[1],s24[1],s25[1],s26[1],s27[1],s28[1],s29[1],s30[1],s31[1],s31[2],s31[3],s30[5],s29[7],s28[9],s27[11],s26[13],s25[15],s24[17],s23[19],s22[21],s21[23],s20[25],s19[27],s18[29],s17[31],s16[33],s15[35],s14[37],s13[39],s12[41],s11[43],s10[45],s9[47],s8[49],s7[51],s6[53],s5[55],s4[57],s3[59],s2[61],s1[63],pp63[33]};
    assign in48_2 = {pp31[0],s1[0],s2[0],s3[0],s4[0],s5[0],s6[0],s7[0],s8[0],s9[0],s10[0],s11[0],s12[0],s13[0],s14[0],s15[0],s16[0],s17[0],s18[0],s19[0],s20[0],s21[0],s22[0],s23[0],s24[0],s25[0],s26[0],s27[0],s28[0],s29[0],s30[0],s31[0],s32[0],s32[1],c32,c31,c30,c29,c28,c27,c26,c25,c24,c23,c22,c21,c20,c19,c18,c17,c16,c15,c14,c13,c12,c11,c10,c9,c8,c7,c6,c5,c4,c3,c2,c1};
    CLA_66 KS_48(s48, c48, in48_1, in48_2);

    /*Stage 3*/
    wire[111:0] s49, in49_1, in49_2;
    wire c49;
    assign in49_1 = {pp0[8],pp0[9],pp0[10],pp0[11],pp0[12],pp0[13],pp0[14],pp0[15],pp2[14],pp4[13],pp6[12],pp8[11],pp10[10],pp12[9],pp14[8],pp16[7],pp18[6],pp20[5],pp22[4],pp24[3],pp26[2],pp28[1],pp30[0],s33[15],s33[16],s33[17],s33[18],s33[19],s33[20],s33[21],s33[22],s33[23],s33[24],s33[25],s33[26],s33[27],s33[28],s33[29],s33[30],s33[31],s33[32],s33[33],s33[34],s33[35],s33[36],s33[37],s33[38],s33[39],s33[40],s33[41],s33[42],s33[43],s33[44],s33[45],s33[46],s33[47],s33[48],s33[49],s33[50],s33[51],s33[52],s33[53],s33[54],s33[55],s33[56],s33[57],s33[58],s33[59],s33[60],s33[61],s33[62],s33[63],s33[64],s33[65],s33[66],s33[67],s33[68],s33[69],s33[70],s33[71],s33[72],s33[73],s33[74],s33[75],s33[76],s33[77],s33[78],s33[79],s33[80],s33[81],pp63[35],pp62[37],pp61[39],pp60[41],pp59[43],pp58[45],pp57[47],pp56[49],pp55[51],pp54[53],pp53[55],pp52[57],pp51[59],pp50[61],pp49[63],pp50[63],pp51[63],pp52[63],pp53[63],pp54[63],pp55[63],pp56[63]};
    assign in49_2 = {pp1[7],pp1[8],pp1[9],pp1[10],pp1[11],pp1[12],pp1[13],pp1[14],pp3[13],pp5[12],pp7[11],pp9[10],pp11[9],pp13[8],pp15[7],pp17[6],pp19[5],pp21[4],pp23[3],pp25[2],pp27[1],pp29[0],s33[14],s34[14],s34[15],s34[16],s34[17],s34[18],s34[19],s34[20],s34[21],s34[22],s34[23],s34[24],s34[25],s34[26],s34[27],s34[28],s34[29],s34[30],s34[31],s34[32],s34[33],s34[34],s34[35],s34[36],s34[37],s34[38],s34[39],s34[40],s34[41],s34[42],s34[43],s34[44],s34[45],s34[46],s34[47],s34[48],s34[49],s34[50],s34[51],s34[52],s34[53],s34[54],s34[55],s34[56],s34[57],s34[58],s34[59],s34[60],s34[61],s34[62],s34[63],s34[64],s34[65],s34[66],s34[67],s34[68],s34[69],s34[70],s34[71],s34[72],s34[73],s34[74],s34[75],s34[76],s34[77],s34[78],s34[79],s34[80],s33[82],pp63[36],pp62[38],pp61[40],pp60[42],pp59[44],pp58[46],pp57[48],pp56[50],pp55[52],pp54[54],pp53[56],pp52[58],pp51[60],pp50[62],pp51[62],pp52[62],pp53[62],pp54[62],pp55[62],pp56[62],pp57[62]};
    CLA_112 KS_49(s49, c49, in49_1, in49_2);
    wire[109:0] s50, in50_1, in50_2;
    wire c50;
    assign in50_1 = {pp2[7],pp2[8],pp2[9],pp2[10],pp2[11],pp2[12],pp2[13],pp4[12],pp6[11],pp8[10],pp10[9],pp12[8],pp14[7],pp16[6],pp18[5],pp20[4],pp22[3],pp24[2],pp26[1],pp28[0],s33[13],s34[13],s35[13],s35[14],s35[15],s35[16],s35[17],s35[18],s35[19],s35[20],s35[21],s35[22],s35[23],s35[24],s35[25],s35[26],s35[27],s35[28],s35[29],s35[30],s35[31],s35[32],s35[33],s35[34],s35[35],s35[36],s35[37],s35[38],s35[39],s35[40],s35[41],s35[42],s35[43],s35[44],s35[45],s35[46],s35[47],s35[48],s35[49],s35[50],s35[51],s35[52],s35[53],s35[54],s35[55],s35[56],s35[57],s35[58],s35[59],s35[60],s35[61],s35[62],s35[63],s35[64],s35[65],s35[66],s35[67],s35[68],s35[69],s35[70],s35[71],s35[72],s35[73],s35[74],s35[75],s35[76],s35[77],s35[78],s35[79],s34[81],s33[83],pp63[37],pp62[39],pp61[41],pp60[43],pp59[45],pp58[47],pp57[49],pp56[51],pp55[53],pp54[55],pp53[57],pp52[59],pp51[61],pp52[61],pp53[61],pp54[61],pp55[61],pp56[61],pp57[61]};
    assign in50_2 = {pp3[6],pp3[7],pp3[8],pp3[9],pp3[10],pp3[11],pp3[12],pp5[11],pp7[10],pp9[9],pp11[8],pp13[7],pp15[6],pp17[5],pp19[4],pp21[3],pp23[2],pp25[1],pp27[0],s33[12],s34[12],s35[12],s36[12],s36[13],s36[14],s36[15],s36[16],s36[17],s36[18],s36[19],s36[20],s36[21],s36[22],s36[23],s36[24],s36[25],s36[26],s36[27],s36[28],s36[29],s36[30],s36[31],s36[32],s36[33],s36[34],s36[35],s36[36],s36[37],s36[38],s36[39],s36[40],s36[41],s36[42],s36[43],s36[44],s36[45],s36[46],s36[47],s36[48],s36[49],s36[50],s36[51],s36[52],s36[53],s36[54],s36[55],s36[56],s36[57],s36[58],s36[59],s36[60],s36[61],s36[62],s36[63],s36[64],s36[65],s36[66],s36[67],s36[68],s36[69],s36[70],s36[71],s36[72],s36[73],s36[74],s36[75],s36[76],s36[77],s36[78],s35[80],s34[82],s33[84],pp63[38],pp62[40],pp61[42],pp60[44],pp59[46],pp58[48],pp57[50],pp56[52],pp55[54],pp54[56],pp53[58],pp52[60],pp53[60],pp54[60],pp55[60],pp56[60],pp57[60],pp58[60]};
    CLA_110 KS_50(s50, c50, in50_1, in50_2);
    wire[107:0] s51, in51_1, in51_2;
    wire c51;
    assign in51_1 = {pp4[6],pp4[7],pp4[8],pp4[9],pp4[10],pp4[11],pp6[10],pp8[9],pp10[8],pp12[7],pp14[6],pp16[5],pp18[4],pp20[3],pp22[2],pp24[1],pp26[0],s33[11],s34[11],s35[11],s36[11],s37[11],s37[12],s37[13],s37[14],s37[15],s37[16],s37[17],s37[18],s37[19],s37[20],s37[21],s37[22],s37[23],s37[24],s37[25],s37[26],s37[27],s37[28],s37[29],s37[30],s37[31],s37[32],s37[33],s37[34],s37[35],s37[36],s37[37],s37[38],s37[39],s37[40],s37[41],s37[42],s37[43],s37[44],s37[45],s37[46],s37[47],s37[48],s37[49],s37[50],s37[51],s37[52],s37[53],s37[54],s37[55],s37[56],s37[57],s37[58],s37[59],s37[60],s37[61],s37[62],s37[63],s37[64],s37[65],s37[66],s37[67],s37[68],s37[69],s37[70],s37[71],s37[72],s37[73],s37[74],s37[75],s37[76],s37[77],s36[79],s35[81],s34[83],s33[85],pp63[39],pp62[41],pp61[43],pp60[45],pp59[47],pp58[49],pp57[51],pp56[53],pp55[55],pp54[57],pp53[59],pp54[59],pp55[59],pp56[59],pp57[59],pp58[59]};
    assign in51_2 = {pp5[5],pp5[6],pp5[7],pp5[8],pp5[9],pp5[10],pp7[9],pp9[8],pp11[7],pp13[6],pp15[5],pp17[4],pp19[3],pp21[2],pp23[1],pp25[0],s33[10],s34[10],s35[10],s36[10],s37[10],s38[10],s38[11],s38[12],s38[13],s38[14],s38[15],s38[16],s38[17],s38[18],s38[19],s38[20],s38[21],s38[22],s38[23],s38[24],s38[25],s38[26],s38[27],s38[28],s38[29],s38[30],s38[31],s38[32],s38[33],s38[34],s38[35],s38[36],s38[37],s38[38],s38[39],s38[40],s38[41],s38[42],s38[43],s38[44],s38[45],s38[46],s38[47],s38[48],s38[49],s38[50],s38[51],s38[52],s38[53],s38[54],s38[55],s38[56],s38[57],s38[58],s38[59],s38[60],s38[61],s38[62],s38[63],s38[64],s38[65],s38[66],s38[67],s38[68],s38[69],s38[70],s38[71],s38[72],s38[73],s38[74],s38[75],s38[76],s37[78],s36[80],s35[82],s34[84],s33[86],pp63[40],pp62[42],pp61[44],pp60[46],pp59[48],pp58[50],pp57[52],pp56[54],pp55[56],pp54[58],pp55[58],pp56[58],pp57[58],pp58[58],pp59[58]};
    CLA_108 KS_51(s51, c51, in51_1, in51_2);
    wire[105:0] s52, in52_1, in52_2;
    wire c52;
    assign in52_1 = {pp6[5],pp6[6],pp6[7],pp6[8],pp6[9],pp8[8],pp10[7],pp12[6],pp14[5],pp16[4],pp18[3],pp20[2],pp22[1],pp24[0],s33[9],s34[9],s35[9],s36[9],s37[9],s38[9],s39[9],s39[10],s39[11],s39[12],s39[13],s39[14],s39[15],s39[16],s39[17],s39[18],s39[19],s39[20],s39[21],s39[22],s39[23],s39[24],s39[25],s39[26],s39[27],s39[28],s39[29],s39[30],s39[31],s39[32],s39[33],s39[34],s39[35],s39[36],s39[37],s39[38],s39[39],s39[40],s39[41],s39[42],s39[43],s39[44],s39[45],s39[46],s39[47],s39[48],s39[49],s39[50],s39[51],s39[52],s39[53],s39[54],s39[55],s39[56],s39[57],s39[58],s39[59],s39[60],s39[61],s39[62],s39[63],s39[64],s39[65],s39[66],s39[67],s39[68],s39[69],s39[70],s39[71],s39[72],s39[73],s39[74],s39[75],s38[77],s37[79],s36[81],s35[83],s34[85],s33[87],pp63[41],pp62[43],pp61[45],pp60[47],pp59[49],pp58[51],pp57[53],pp56[55],pp55[57],pp56[57],pp57[57],pp58[57],pp59[57]};
    assign in52_2 = {pp7[4],pp7[5],pp7[6],pp7[7],pp7[8],pp9[7],pp11[6],pp13[5],pp15[4],pp17[3],pp19[2],pp21[1],pp23[0],s33[8],s34[8],s35[8],s36[8],s37[8],s38[8],s39[8],s40[8],s40[9],s40[10],s40[11],s40[12],s40[13],s40[14],s40[15],s40[16],s40[17],s40[18],s40[19],s40[20],s40[21],s40[22],s40[23],s40[24],s40[25],s40[26],s40[27],s40[28],s40[29],s40[30],s40[31],s40[32],s40[33],s40[34],s40[35],s40[36],s40[37],s40[38],s40[39],s40[40],s40[41],s40[42],s40[43],s40[44],s40[45],s40[46],s40[47],s40[48],s40[49],s40[50],s40[51],s40[52],s40[53],s40[54],s40[55],s40[56],s40[57],s40[58],s40[59],s40[60],s40[61],s40[62],s40[63],s40[64],s40[65],s40[66],s40[67],s40[68],s40[69],s40[70],s40[71],s40[72],s40[73],s40[74],s39[76],s38[78],s37[80],s36[82],s35[84],s34[86],s33[88],pp63[42],pp62[44],pp61[46],pp60[48],pp59[50],pp58[52],pp57[54],pp56[56],pp57[56],pp58[56],pp59[56],pp60[56]};
    CLA_106 KS_52(s52, c52, in52_1, in52_2);
    wire[103:0] s53, in53_1, in53_2;
    wire c53;
    assign in53_1 = {pp8[4],pp8[5],pp8[6],pp8[7],pp10[6],pp12[5],pp14[4],pp16[3],pp18[2],pp20[1],pp22[0],s33[7],s34[7],s35[7],s36[7],s37[7],s38[7],s39[7],s40[7],s41[7],s41[8],s41[9],s41[10],s41[11],s41[12],s41[13],s41[14],s41[15],s41[16],s41[17],s41[18],s41[19],s41[20],s41[21],s41[22],s41[23],s41[24],s41[25],s41[26],s41[27],s41[28],s41[29],s41[30],s41[31],s41[32],s41[33],s41[34],s41[35],s41[36],s41[37],s41[38],s41[39],s41[40],s41[41],s41[42],s41[43],s41[44],s41[45],s41[46],s41[47],s41[48],s41[49],s41[50],s41[51],s41[52],s41[53],s41[54],s41[55],s41[56],s41[57],s41[58],s41[59],s41[60],s41[61],s41[62],s41[63],s41[64],s41[65],s41[66],s41[67],s41[68],s41[69],s41[70],s41[71],s41[72],s41[73],s40[75],s39[77],s38[79],s37[81],s36[83],s35[85],s34[87],s33[89],pp63[43],pp62[45],pp61[47],pp60[49],pp59[51],pp58[53],pp57[55],pp58[55],pp59[55],pp60[55]};
    assign in53_2 = {pp9[3],pp9[4],pp9[5],pp9[6],pp11[5],pp13[4],pp15[3],pp17[2],pp19[1],pp21[0],s33[6],s34[6],s35[6],s36[6],s37[6],s38[6],s39[6],s40[6],s41[6],s42[6],s42[7],s42[8],s42[9],s42[10],s42[11],s42[12],s42[13],s42[14],s42[15],s42[16],s42[17],s42[18],s42[19],s42[20],s42[21],s42[22],s42[23],s42[24],s42[25],s42[26],s42[27],s42[28],s42[29],s42[30],s42[31],s42[32],s42[33],s42[34],s42[35],s42[36],s42[37],s42[38],s42[39],s42[40],s42[41],s42[42],s42[43],s42[44],s42[45],s42[46],s42[47],s42[48],s42[49],s42[50],s42[51],s42[52],s42[53],s42[54],s42[55],s42[56],s42[57],s42[58],s42[59],s42[60],s42[61],s42[62],s42[63],s42[64],s42[65],s42[66],s42[67],s42[68],s42[69],s42[70],s42[71],s42[72],s41[74],s40[76],s39[78],s38[80],s37[82],s36[84],s35[86],s34[88],s33[90],pp63[44],pp62[46],pp61[48],pp60[50],pp59[52],pp58[54],pp59[54],pp60[54],pp61[54]};
    CLA_104 KS_53(s53, c53, in53_1, in53_2);
    wire[101:0] s54, in54_1, in54_2;
    wire c54;
    assign in54_1 = {pp10[3],pp10[4],pp10[5],pp12[4],pp14[3],pp16[2],pp18[1],pp20[0],s33[5],s34[5],s35[5],s36[5],s37[5],s38[5],s39[5],s40[5],s41[5],s42[5],s43[5],s43[6],s43[7],s43[8],s43[9],s43[10],s43[11],s43[12],s43[13],s43[14],s43[15],s43[16],s43[17],s43[18],s43[19],s43[20],s43[21],s43[22],s43[23],s43[24],s43[25],s43[26],s43[27],s43[28],s43[29],s43[30],s43[31],s43[32],s43[33],s43[34],s43[35],s43[36],s43[37],s43[38],s43[39],s43[40],s43[41],s43[42],s43[43],s43[44],s43[45],s43[46],s43[47],s43[48],s43[49],s43[50],s43[51],s43[52],s43[53],s43[54],s43[55],s43[56],s43[57],s43[58],s43[59],s43[60],s43[61],s43[62],s43[63],s43[64],s43[65],s43[66],s43[67],s43[68],s43[69],s43[70],s43[71],s42[73],s41[75],s40[77],s39[79],s38[81],s37[83],s36[85],s35[87],s34[89],s33[91],pp63[45],pp62[47],pp61[49],pp60[51],pp59[53],pp60[53],pp61[53]};
    assign in54_2 = {pp11[2],pp11[3],pp11[4],pp13[3],pp15[2],pp17[1],pp19[0],s33[4],s34[4],s35[4],s36[4],s37[4],s38[4],s39[4],s40[4],s41[4],s42[4],s43[4],s44[4],s44[5],s44[6],s44[7],s44[8],s44[9],s44[10],s44[11],s44[12],s44[13],s44[14],s44[15],s44[16],s44[17],s44[18],s44[19],s44[20],s44[21],s44[22],s44[23],s44[24],s44[25],s44[26],s44[27],s44[28],s44[29],s44[30],s44[31],s44[32],s44[33],s44[34],s44[35],s44[36],s44[37],s44[38],s44[39],s44[40],s44[41],s44[42],s44[43],s44[44],s44[45],s44[46],s44[47],s44[48],s44[49],s44[50],s44[51],s44[52],s44[53],s44[54],s44[55],s44[56],s44[57],s44[58],s44[59],s44[60],s44[61],s44[62],s44[63],s44[64],s44[65],s44[66],s44[67],s44[68],s44[69],s44[70],s43[72],s42[74],s41[76],s40[78],s39[80],s38[82],s37[84],s36[86],s35[88],s34[90],s33[92],pp63[46],pp62[48],pp61[50],pp60[52],pp61[52],pp62[52]};
    CLA_102 KS_54(s54, c54, in54_1, in54_2);
    wire[99:0] s55, in55_1, in55_2;
    wire c55;
    assign in55_1 = {pp12[2],pp12[3],pp14[2],pp16[1],pp18[0],s33[3],s34[3],s35[3],s36[3],s37[3],s38[3],s39[3],s40[3],s41[3],s42[3],s43[3],s44[3],s45[3],s45[4],s45[5],s45[6],s45[7],s45[8],s45[9],s45[10],s45[11],s45[12],s45[13],s45[14],s45[15],s45[16],s45[17],s45[18],s45[19],s45[20],s45[21],s45[22],s45[23],s45[24],s45[25],s45[26],s45[27],s45[28],s45[29],s45[30],s45[31],s45[32],s45[33],s45[34],s45[35],s45[36],s45[37],s45[38],s45[39],s45[40],s45[41],s45[42],s45[43],s45[44],s45[45],s45[46],s45[47],s45[48],s45[49],s45[50],s45[51],s45[52],s45[53],s45[54],s45[55],s45[56],s45[57],s45[58],s45[59],s45[60],s45[61],s45[62],s45[63],s45[64],s45[65],s45[66],s45[67],s45[68],s45[69],s44[71],s43[73],s42[75],s41[77],s40[79],s39[81],s38[83],s37[85],s36[87],s35[89],s34[91],s33[93],pp63[47],pp62[49],pp61[51],pp62[51]};
    assign in55_2 = {pp13[1],pp13[2],pp15[1],pp17[0],s33[2],s34[2],s35[2],s36[2],s37[2],s38[2],s39[2],s40[2],s41[2],s42[2],s43[2],s44[2],s45[2],s46[2],s46[3],s46[4],s46[5],s46[6],s46[7],s46[8],s46[9],s46[10],s46[11],s46[12],s46[13],s46[14],s46[15],s46[16],s46[17],s46[18],s46[19],s46[20],s46[21],s46[22],s46[23],s46[24],s46[25],s46[26],s46[27],s46[28],s46[29],s46[30],s46[31],s46[32],s46[33],s46[34],s46[35],s46[36],s46[37],s46[38],s46[39],s46[40],s46[41],s46[42],s46[43],s46[44],s46[45],s46[46],s46[47],s46[48],s46[49],s46[50],s46[51],s46[52],s46[53],s46[54],s46[55],s46[56],s46[57],s46[58],s46[59],s46[60],s46[61],s46[62],s46[63],s46[64],s46[65],s46[66],s46[67],s46[68],s45[70],s44[72],s43[74],s42[76],s41[78],s40[80],s39[82],s38[84],s37[86],s36[88],s35[90],s34[92],s33[94],pp63[48],pp62[50],pp63[50]};
    CLA_100 KS_55(s55, c55, in55_1, in55_2);
    wire[97:0] s56, in56_1, in56_2;
    wire c56;
    assign in56_1 = {pp14[1],pp16[0],s33[1],s34[1],s35[1],s36[1],s37[1],s38[1],s39[1],s40[1],s41[1],s42[1],s43[1],s44[1],s45[1],s46[1],s47[1],s47[2],s47[3],s47[4],s47[5],s47[6],s47[7],s47[8],s47[9],s47[10],s47[11],s47[12],s47[13],s47[14],s47[15],s47[16],s47[17],s47[18],s47[19],s47[20],s47[21],s47[22],s47[23],s47[24],s47[25],s47[26],s47[27],s47[28],s47[29],s47[30],s47[31],s47[32],s47[33],s47[34],s47[35],s47[36],s47[37],s47[38],s47[39],s47[40],s47[41],s47[42],s47[43],s47[44],s47[45],s47[46],s47[47],s47[48],s47[49],s47[50],s47[51],s47[52],s47[53],s47[54],s47[55],s47[56],s47[57],s47[58],s47[59],s47[60],s47[61],s47[62],s47[63],s47[64],s47[65],s47[66],s47[67],s46[69],s45[71],s44[73],s43[75],s42[77],s41[79],s40[81],s39[83],s38[85],s37[87],s36[89],s35[91],s34[93],s33[95],pp63[49]};
    assign in56_2 = {pp15[0],s33[0],s34[0],s35[0],s36[0],s37[0],s38[0],s39[0],s40[0],s41[0],s42[0],s43[0],s44[0],s45[0],s46[0],s47[0],s48[0],s48[1],s48[2],s48[3],s48[4],s48[5],s48[6],s48[7],s48[8],s48[9],s48[10],s48[11],s48[12],s48[13],s48[14],s48[15],s48[16],s48[17],s48[18],s48[19],s48[20],s48[21],s48[22],s48[23],s48[24],s48[25],s48[26],s48[27],s48[28],s48[29],s48[30],s48[31],s48[32],s48[33],s48[34],s48[35],s48[36],s48[37],s48[38],s48[39],s48[40],s48[41],s48[42],s48[43],s48[44],s48[45],s48[46],s48[47],s48[48],s48[49],s48[50],s48[51],s48[52],s48[53],s48[54],s48[55],s48[56],s48[57],s48[58],s48[59],s48[60],s48[61],s48[62],s48[63],s48[64],s48[65],c48,c47,c46,c45,c44,c43,c42,c41,c40,c39,c38,c37,c36,c35,c34,c33};
    CLA_98 KS_56(s56, c56, in56_1, in56_2);

    /*Stage 4*/
    wire[119:0] s57, in57_1, in57_2;
    wire c57;
    assign in57_1 = {pp0[4],pp0[5],pp0[6],pp0[7],pp2[6],pp4[5],pp6[4],pp8[3],pp10[2],pp12[1],pp14[0],s49[7],s49[8],s49[9],s49[10],s49[11],s49[12],s49[13],s49[14],s49[15],s49[16],s49[17],s49[18],s49[19],s49[20],s49[21],s49[22],s49[23],s49[24],s49[25],s49[26],s49[27],s49[28],s49[29],s49[30],s49[31],s49[32],s49[33],s49[34],s49[35],s49[36],s49[37],s49[38],s49[39],s49[40],s49[41],s49[42],s49[43],s49[44],s49[45],s49[46],s49[47],s49[48],s49[49],s49[50],s49[51],s49[52],s49[53],s49[54],s49[55],s49[56],s49[57],s49[58],s49[59],s49[60],s49[61],s49[62],s49[63],s49[64],s49[65],s49[66],s49[67],s49[68],s49[69],s49[70],s49[71],s49[72],s49[73],s49[74],s49[75],s49[76],s49[77],s49[78],s49[79],s49[80],s49[81],s49[82],s49[83],s49[84],s49[85],s49[86],s49[87],s49[88],s49[89],s49[90],s49[91],s49[92],s49[93],s49[94],s49[95],s49[96],s49[97],s49[98],s49[99],s49[100],s49[101],s49[102],s49[103],s49[104],s49[105],pp63[51],pp62[53],pp61[55],pp60[57],pp59[59],pp58[61],pp57[63],pp58[63],pp59[63],pp60[63]};
    assign in57_2 = {pp1[3],pp1[4],pp1[5],pp1[6],pp3[5],pp5[4],pp7[3],pp9[2],pp11[1],pp13[0],s49[6],s50[6],s50[7],s50[8],s50[9],s50[10],s50[11],s50[12],s50[13],s50[14],s50[15],s50[16],s50[17],s50[18],s50[19],s50[20],s50[21],s50[22],s50[23],s50[24],s50[25],s50[26],s50[27],s50[28],s50[29],s50[30],s50[31],s50[32],s50[33],s50[34],s50[35],s50[36],s50[37],s50[38],s50[39],s50[40],s50[41],s50[42],s50[43],s50[44],s50[45],s50[46],s50[47],s50[48],s50[49],s50[50],s50[51],s50[52],s50[53],s50[54],s50[55],s50[56],s50[57],s50[58],s50[59],s50[60],s50[61],s50[62],s50[63],s50[64],s50[65],s50[66],s50[67],s50[68],s50[69],s50[70],s50[71],s50[72],s50[73],s50[74],s50[75],s50[76],s50[77],s50[78],s50[79],s50[80],s50[81],s50[82],s50[83],s50[84],s50[85],s50[86],s50[87],s50[88],s50[89],s50[90],s50[91],s50[92],s50[93],s50[94],s50[95],s50[96],s50[97],s50[98],s50[99],s50[100],s50[101],s50[102],s50[103],s50[104],s49[106],pp63[52],pp62[54],pp61[56],pp60[58],pp59[60],pp58[62],pp59[62],pp60[62],pp61[62]};
    CLA_120 KS_57(s57, c57, in57_1, in57_2);
    wire[117:0] s58, in58_1, in58_2;
    wire c58;
    assign in58_1 = {pp2[3],pp2[4],pp2[5],pp4[4],pp6[3],pp8[2],pp10[1],pp12[0],s49[5],s50[5],s51[5],s51[6],s51[7],s51[8],s51[9],s51[10],s51[11],s51[12],s51[13],s51[14],s51[15],s51[16],s51[17],s51[18],s51[19],s51[20],s51[21],s51[22],s51[23],s51[24],s51[25],s51[26],s51[27],s51[28],s51[29],s51[30],s51[31],s51[32],s51[33],s51[34],s51[35],s51[36],s51[37],s51[38],s51[39],s51[40],s51[41],s51[42],s51[43],s51[44],s51[45],s51[46],s51[47],s51[48],s51[49],s51[50],s51[51],s51[52],s51[53],s51[54],s51[55],s51[56],s51[57],s51[58],s51[59],s51[60],s51[61],s51[62],s51[63],s51[64],s51[65],s51[66],s51[67],s51[68],s51[69],s51[70],s51[71],s51[72],s51[73],s51[74],s51[75],s51[76],s51[77],s51[78],s51[79],s51[80],s51[81],s51[82],s51[83],s51[84],s51[85],s51[86],s51[87],s51[88],s51[89],s51[90],s51[91],s51[92],s51[93],s51[94],s51[95],s51[96],s51[97],s51[98],s51[99],s51[100],s51[101],s51[102],s51[103],s50[105],s49[107],pp63[53],pp62[55],pp61[57],pp60[59],pp59[61],pp60[61],pp61[61]};
    assign in58_2 = {pp3[2],pp3[3],pp3[4],pp5[3],pp7[2],pp9[1],pp11[0],s49[4],s50[4],s51[4],s52[4],s52[5],s52[6],s52[7],s52[8],s52[9],s52[10],s52[11],s52[12],s52[13],s52[14],s52[15],s52[16],s52[17],s52[18],s52[19],s52[20],s52[21],s52[22],s52[23],s52[24],s52[25],s52[26],s52[27],s52[28],s52[29],s52[30],s52[31],s52[32],s52[33],s52[34],s52[35],s52[36],s52[37],s52[38],s52[39],s52[40],s52[41],s52[42],s52[43],s52[44],s52[45],s52[46],s52[47],s52[48],s52[49],s52[50],s52[51],s52[52],s52[53],s52[54],s52[55],s52[56],s52[57],s52[58],s52[59],s52[60],s52[61],s52[62],s52[63],s52[64],s52[65],s52[66],s52[67],s52[68],s52[69],s52[70],s52[71],s52[72],s52[73],s52[74],s52[75],s52[76],s52[77],s52[78],s52[79],s52[80],s52[81],s52[82],s52[83],s52[84],s52[85],s52[86],s52[87],s52[88],s52[89],s52[90],s52[91],s52[92],s52[93],s52[94],s52[95],s52[96],s52[97],s52[98],s52[99],s52[100],s52[101],s52[102],s51[104],s50[106],s49[108],pp63[54],pp62[56],pp61[58],pp60[60],pp61[60],pp62[60]};
    CLA_118 KS_58(s58, c58, in58_1, in58_2);
    wire[115:0] s59, in59_1, in59_2;
    wire c59;
    assign in59_1 = {pp4[2],pp4[3],pp6[2],pp8[1],pp10[0],s49[3],s50[3],s51[3],s52[3],s53[3],s53[4],s53[5],s53[6],s53[7],s53[8],s53[9],s53[10],s53[11],s53[12],s53[13],s53[14],s53[15],s53[16],s53[17],s53[18],s53[19],s53[20],s53[21],s53[22],s53[23],s53[24],s53[25],s53[26],s53[27],s53[28],s53[29],s53[30],s53[31],s53[32],s53[33],s53[34],s53[35],s53[36],s53[37],s53[38],s53[39],s53[40],s53[41],s53[42],s53[43],s53[44],s53[45],s53[46],s53[47],s53[48],s53[49],s53[50],s53[51],s53[52],s53[53],s53[54],s53[55],s53[56],s53[57],s53[58],s53[59],s53[60],s53[61],s53[62],s53[63],s53[64],s53[65],s53[66],s53[67],s53[68],s53[69],s53[70],s53[71],s53[72],s53[73],s53[74],s53[75],s53[76],s53[77],s53[78],s53[79],s53[80],s53[81],s53[82],s53[83],s53[84],s53[85],s53[86],s53[87],s53[88],s53[89],s53[90],s53[91],s53[92],s53[93],s53[94],s53[95],s53[96],s53[97],s53[98],s53[99],s53[100],s53[101],s52[103],s51[105],s50[107],s49[109],pp63[55],pp62[57],pp61[59],pp62[59]};
    assign in59_2 = {pp5[1],pp5[2],pp7[1],pp9[0],s49[2],s50[2],s51[2],s52[2],s53[2],s54[2],s54[3],s54[4],s54[5],s54[6],s54[7],s54[8],s54[9],s54[10],s54[11],s54[12],s54[13],s54[14],s54[15],s54[16],s54[17],s54[18],s54[19],s54[20],s54[21],s54[22],s54[23],s54[24],s54[25],s54[26],s54[27],s54[28],s54[29],s54[30],s54[31],s54[32],s54[33],s54[34],s54[35],s54[36],s54[37],s54[38],s54[39],s54[40],s54[41],s54[42],s54[43],s54[44],s54[45],s54[46],s54[47],s54[48],s54[49],s54[50],s54[51],s54[52],s54[53],s54[54],s54[55],s54[56],s54[57],s54[58],s54[59],s54[60],s54[61],s54[62],s54[63],s54[64],s54[65],s54[66],s54[67],s54[68],s54[69],s54[70],s54[71],s54[72],s54[73],s54[74],s54[75],s54[76],s54[77],s54[78],s54[79],s54[80],s54[81],s54[82],s54[83],s54[84],s54[85],s54[86],s54[87],s54[88],s54[89],s54[90],s54[91],s54[92],s54[93],s54[94],s54[95],s54[96],s54[97],s54[98],s54[99],s54[100],s53[102],s52[104],s51[106],s50[108],s49[110],pp63[56],pp62[58],pp63[58]};
    CLA_116 KS_59(s59, c59, in59_1, in59_2);
    wire[113:0] s60, in60_1, in60_2;
    wire c60;
    assign in60_1 = {pp6[1],pp8[0],s49[1],s50[1],s51[1],s52[1],s53[1],s54[1],s55[1],s55[2],s55[3],s55[4],s55[5],s55[6],s55[7],s55[8],s55[9],s55[10],s55[11],s55[12],s55[13],s55[14],s55[15],s55[16],s55[17],s55[18],s55[19],s55[20],s55[21],s55[22],s55[23],s55[24],s55[25],s55[26],s55[27],s55[28],s55[29],s55[30],s55[31],s55[32],s55[33],s55[34],s55[35],s55[36],s55[37],s55[38],s55[39],s55[40],s55[41],s55[42],s55[43],s55[44],s55[45],s55[46],s55[47],s55[48],s55[49],s55[50],s55[51],s55[52],s55[53],s55[54],s55[55],s55[56],s55[57],s55[58],s55[59],s55[60],s55[61],s55[62],s55[63],s55[64],s55[65],s55[66],s55[67],s55[68],s55[69],s55[70],s55[71],s55[72],s55[73],s55[74],s55[75],s55[76],s55[77],s55[78],s55[79],s55[80],s55[81],s55[82],s55[83],s55[84],s55[85],s55[86],s55[87],s55[88],s55[89],s55[90],s55[91],s55[92],s55[93],s55[94],s55[95],s55[96],s55[97],s55[98],s55[99],s54[101],s53[103],s52[105],s51[107],s50[109],s49[111],pp63[57]};
    assign in60_2 = {pp7[0],s49[0],s50[0],s51[0],s52[0],s53[0],s54[0],s55[0],s56[0],s56[1],s56[2],s56[3],s56[4],s56[5],s56[6],s56[7],s56[8],s56[9],s56[10],s56[11],s56[12],s56[13],s56[14],s56[15],s56[16],s56[17],s56[18],s56[19],s56[20],s56[21],s56[22],s56[23],s56[24],s56[25],s56[26],s56[27],s56[28],s56[29],s56[30],s56[31],s56[32],s56[33],s56[34],s56[35],s56[36],s56[37],s56[38],s56[39],s56[40],s56[41],s56[42],s56[43],s56[44],s56[45],s56[46],s56[47],s56[48],s56[49],s56[50],s56[51],s56[52],s56[53],s56[54],s56[55],s56[56],s56[57],s56[58],s56[59],s56[60],s56[61],s56[62],s56[63],s56[64],s56[65],s56[66],s56[67],s56[68],s56[69],s56[70],s56[71],s56[72],s56[73],s56[74],s56[75],s56[76],s56[77],s56[78],s56[79],s56[80],s56[81],s56[82],s56[83],s56[84],s56[85],s56[86],s56[87],s56[88],s56[89],s56[90],s56[91],s56[92],s56[93],s56[94],s56[95],s56[96],s56[97],c56,c55,c54,c53,c52,c51,c50,c49};
    CLA_114 KS_60(s60, c60, in60_1, in60_2);

    /*Stage 5*/
    wire[123:0] s61, in61_1, in61_2;
    wire c61;
    assign in61_1 = {pp0[2],pp0[3],pp2[2],pp4[1],pp6[0],s57[3],s57[4],s57[5],s57[6],s57[7],s57[8],s57[9],s57[10],s57[11],s57[12],s57[13],s57[14],s57[15],s57[16],s57[17],s57[18],s57[19],s57[20],s57[21],s57[22],s57[23],s57[24],s57[25],s57[26],s57[27],s57[28],s57[29],s57[30],s57[31],s57[32],s57[33],s57[34],s57[35],s57[36],s57[37],s57[38],s57[39],s57[40],s57[41],s57[42],s57[43],s57[44],s57[45],s57[46],s57[47],s57[48],s57[49],s57[50],s57[51],s57[52],s57[53],s57[54],s57[55],s57[56],s57[57],s57[58],s57[59],s57[60],s57[61],s57[62],s57[63],s57[64],s57[65],s57[66],s57[67],s57[68],s57[69],s57[70],s57[71],s57[72],s57[73],s57[74],s57[75],s57[76],s57[77],s57[78],s57[79],s57[80],s57[81],s57[82],s57[83],s57[84],s57[85],s57[86],s57[87],s57[88],s57[89],s57[90],s57[91],s57[92],s57[93],s57[94],s57[95],s57[96],s57[97],s57[98],s57[99],s57[100],s57[101],s57[102],s57[103],s57[104],s57[105],s57[106],s57[107],s57[108],s57[109],s57[110],s57[111],s57[112],s57[113],s57[114],s57[115],s57[116],s57[117],pp63[59],pp62[61],pp61[63],pp62[63]};
    assign in61_2 = {pp1[1],pp1[2],pp3[1],pp5[0],s57[2],s58[2],s58[3],s58[4],s58[5],s58[6],s58[7],s58[8],s58[9],s58[10],s58[11],s58[12],s58[13],s58[14],s58[15],s58[16],s58[17],s58[18],s58[19],s58[20],s58[21],s58[22],s58[23],s58[24],s58[25],s58[26],s58[27],s58[28],s58[29],s58[30],s58[31],s58[32],s58[33],s58[34],s58[35],s58[36],s58[37],s58[38],s58[39],s58[40],s58[41],s58[42],s58[43],s58[44],s58[45],s58[46],s58[47],s58[48],s58[49],s58[50],s58[51],s58[52],s58[53],s58[54],s58[55],s58[56],s58[57],s58[58],s58[59],s58[60],s58[61],s58[62],s58[63],s58[64],s58[65],s58[66],s58[67],s58[68],s58[69],s58[70],s58[71],s58[72],s58[73],s58[74],s58[75],s58[76],s58[77],s58[78],s58[79],s58[80],s58[81],s58[82],s58[83],s58[84],s58[85],s58[86],s58[87],s58[88],s58[89],s58[90],s58[91],s58[92],s58[93],s58[94],s58[95],s58[96],s58[97],s58[98],s58[99],s58[100],s58[101],s58[102],s58[103],s58[104],s58[105],s58[106],s58[107],s58[108],s58[109],s58[110],s58[111],s58[112],s58[113],s58[114],s58[115],s58[116],s57[118],pp63[60],pp62[62],pp63[62]};
    CLA_124 KS_61(s61, c61, in61_1, in61_2);
    wire[121:0] s62, in62_1, in62_2;
    wire c62;
    assign in62_1 = {pp2[1],pp4[0],s57[1],s58[1],s59[1],s59[2],s59[3],s59[4],s59[5],s59[6],s59[7],s59[8],s59[9],s59[10],s59[11],s59[12],s59[13],s59[14],s59[15],s59[16],s59[17],s59[18],s59[19],s59[20],s59[21],s59[22],s59[23],s59[24],s59[25],s59[26],s59[27],s59[28],s59[29],s59[30],s59[31],s59[32],s59[33],s59[34],s59[35],s59[36],s59[37],s59[38],s59[39],s59[40],s59[41],s59[42],s59[43],s59[44],s59[45],s59[46],s59[47],s59[48],s59[49],s59[50],s59[51],s59[52],s59[53],s59[54],s59[55],s59[56],s59[57],s59[58],s59[59],s59[60],s59[61],s59[62],s59[63],s59[64],s59[65],s59[66],s59[67],s59[68],s59[69],s59[70],s59[71],s59[72],s59[73],s59[74],s59[75],s59[76],s59[77],s59[78],s59[79],s59[80],s59[81],s59[82],s59[83],s59[84],s59[85],s59[86],s59[87],s59[88],s59[89],s59[90],s59[91],s59[92],s59[93],s59[94],s59[95],s59[96],s59[97],s59[98],s59[99],s59[100],s59[101],s59[102],s59[103],s59[104],s59[105],s59[106],s59[107],s59[108],s59[109],s59[110],s59[111],s59[112],s59[113],s59[114],s59[115],s58[117],s57[119],pp63[61]};
    assign in62_2 = {pp3[0],s57[0],s58[0],s59[0],s60[0],s60[1],s60[2],s60[3],s60[4],s60[5],s60[6],s60[7],s60[8],s60[9],s60[10],s60[11],s60[12],s60[13],s60[14],s60[15],s60[16],s60[17],s60[18],s60[19],s60[20],s60[21],s60[22],s60[23],s60[24],s60[25],s60[26],s60[27],s60[28],s60[29],s60[30],s60[31],s60[32],s60[33],s60[34],s60[35],s60[36],s60[37],s60[38],s60[39],s60[40],s60[41],s60[42],s60[43],s60[44],s60[45],s60[46],s60[47],s60[48],s60[49],s60[50],s60[51],s60[52],s60[53],s60[54],s60[55],s60[56],s60[57],s60[58],s60[59],s60[60],s60[61],s60[62],s60[63],s60[64],s60[65],s60[66],s60[67],s60[68],s60[69],s60[70],s60[71],s60[72],s60[73],s60[74],s60[75],s60[76],s60[77],s60[78],s60[79],s60[80],s60[81],s60[82],s60[83],s60[84],s60[85],s60[86],s60[87],s60[88],s60[89],s60[90],s60[91],s60[92],s60[93],s60[94],s60[95],s60[96],s60[97],s60[98],s60[99],s60[100],s60[101],s60[102],s60[103],s60[104],s60[105],s60[106],s60[107],s60[108],s60[109],s60[110],s60[111],s60[112],s60[113],c60,c59,c58,c57};
    CLA_122 KS_62(s62, c62, in62_1, in62_2);


    /*Final Stage 5*/
    wire[125:0] s, in_1, in_2;
    wire c;
    assign in_1 = {pp0[1],pp2[0],s61[1],s61[2],s61[3],s61[4],s61[5],s61[6],s61[7],s61[8],s61[9],s61[10],s61[11],s61[12],s61[13],s61[14],s61[15],s61[16],s61[17],s61[18],s61[19],s61[20],s61[21],s61[22],s61[23],s61[24],s61[25],s61[26],s61[27],s61[28],s61[29],s61[30],s61[31],s61[32],s61[33],s61[34],s61[35],s61[36],s61[37],s61[38],s61[39],s61[40],s61[41],s61[42],s61[43],s61[44],s61[45],s61[46],s61[47],s61[48],s61[49],s61[50],s61[51],s61[52],s61[53],s61[54],s61[55],s61[56],s61[57],s61[58],s61[59],s61[60],s61[61],s61[62],s61[63],s61[64],s61[65],s61[66],s61[67],s61[68],s61[69],s61[70],s61[71],s61[72],s61[73],s61[74],s61[75],s61[76],s61[77],s61[78],s61[79],s61[80],s61[81],s61[82],s61[83],s61[84],s61[85],s61[86],s61[87],s61[88],s61[89],s61[90],s61[91],s61[92],s61[93],s61[94],s61[95],s61[96],s61[97],s61[98],s61[99],s61[100],s61[101],s61[102],s61[103],s61[104],s61[105],s61[106],s61[107],s61[108],s61[109],s61[110],s61[111],s61[112],s61[113],s61[114],s61[115],s61[116],s61[117],s61[118],s61[119],s61[120],s61[121],s61[122],s61[123],pp63[63]};
    assign in_2 = {pp1[0],s61[0],s62[0],s62[1],s62[2],s62[3],s62[4],s62[5],s62[6],s62[7],s62[8],s62[9],s62[10],s62[11],s62[12],s62[13],s62[14],s62[15],s62[16],s62[17],s62[18],s62[19],s62[20],s62[21],s62[22],s62[23],s62[24],s62[25],s62[26],s62[27],s62[28],s62[29],s62[30],s62[31],s62[32],s62[33],s62[34],s62[35],s62[36],s62[37],s62[38],s62[39],s62[40],s62[41],s62[42],s62[43],s62[44],s62[45],s62[46],s62[47],s62[48],s62[49],s62[50],s62[51],s62[52],s62[53],s62[54],s62[55],s62[56],s62[57],s62[58],s62[59],s62[60],s62[61],s62[62],s62[63],s62[64],s62[65],s62[66],s62[67],s62[68],s62[69],s62[70],s62[71],s62[72],s62[73],s62[74],s62[75],s62[76],s62[77],s62[78],s62[79],s62[80],s62[81],s62[82],s62[83],s62[84],s62[85],s62[86],s62[87],s62[88],s62[89],s62[90],s62[91],s62[92],s62[93],s62[94],s62[95],s62[96],s62[97],s62[98],s62[99],s62[100],s62[101],s62[102],s62[103],s62[104],s62[105],s62[106],s62[107],s62[108],s62[109],s62[110],s62[111],s62[112],s62[113],s62[114],s62[115],s62[116],s62[117],s62[118],s62[119],s62[120],s62[121],c62,c61};
    CLA_126(s, c, in_1, in_2);

    assign product[0] = pp0[0];
    assign product[1] = s[0];
    assign product[2] = s[1];
    assign product[3] = s[2];
    assign product[4] = s[3];
    assign product[5] = s[4];
    assign product[6] = s[5];
    assign product[7] = s[6];
    assign product[8] = s[7];
    assign product[9] = s[8];
    assign product[10] = s[9];
    assign product[11] = s[10];
    assign product[12] = s[11];
    assign product[13] = s[12];
    assign product[14] = s[13];
    assign product[15] = s[14];
    assign product[16] = s[15];
    assign product[17] = s[16];
    assign product[18] = s[17];
    assign product[19] = s[18];
    assign product[20] = s[19];
    assign product[21] = s[20];
    assign product[22] = s[21];
    assign product[23] = s[22];
    assign product[24] = s[23];
    assign product[25] = s[24];
    assign product[26] = s[25];
    assign product[27] = s[26];
    assign product[28] = s[27];
    assign product[29] = s[28];
    assign product[30] = s[29];
    assign product[31] = s[30];
    assign product[32] = s[31];
    assign product[33] = s[32];
    assign product[34] = s[33];
    assign product[35] = s[34];
    assign product[36] = s[35];
    assign product[37] = s[36];
    assign product[38] = s[37];
    assign product[39] = s[38];
    assign product[40] = s[39];
    assign product[41] = s[40];
    assign product[42] = s[41];
    assign product[43] = s[42];
    assign product[44] = s[43];
    assign product[45] = s[44];
    assign product[46] = s[45];
    assign product[47] = s[46];
    assign product[48] = s[47];
    assign product[49] = s[48];
    assign product[50] = s[49];
    assign product[51] = s[50];
    assign product[52] = s[51];
    assign product[53] = s[52];
    assign product[54] = s[53];
    assign product[55] = s[54];
    assign product[56] = s[55];
    assign product[57] = s[56];
    assign product[58] = s[57];
    assign product[59] = s[58];
    assign product[60] = s[59];
    assign product[61] = s[60];
    assign product[62] = s[61];
    assign product[63] = s[62];
    assign product[64] = s[63];
    assign product[65] = s[64];
    assign product[66] = s[65];
    assign product[67] = s[66];
    assign product[68] = s[67];
    assign product[69] = s[68];
    assign product[70] = s[69];
    assign product[71] = s[70];
    assign product[72] = s[71];
    assign product[73] = s[72];
    assign product[74] = s[73];
    assign product[75] = s[74];
    assign product[76] = s[75];
    assign product[77] = s[76];
    assign product[78] = s[77];
    assign product[79] = s[78];
    assign product[80] = s[79];
    assign product[81] = s[80];
    assign product[82] = s[81];
    assign product[83] = s[82];
    assign product[84] = s[83];
    assign product[85] = s[84];
    assign product[86] = s[85];
    assign product[87] = s[86];
    assign product[88] = s[87];
    assign product[89] = s[88];
    assign product[90] = s[89];
    assign product[91] = s[90];
    assign product[92] = s[91];
    assign product[93] = s[92];
    assign product[94] = s[93];
    assign product[95] = s[94];
    assign product[96] = s[95];
    assign product[97] = s[96];
    assign product[98] = s[97];
    assign product[99] = s[98];
    assign product[100] = s[99];
    assign product[101] = s[100];
    assign product[102] = s[101];
    assign product[103] = s[102];
    assign product[104] = s[103];
    assign product[105] = s[104];
    assign product[106] = s[105];
    assign product[107] = s[106];
    assign product[108] = s[107];
    assign product[109] = s[108];
    assign product[110] = s[109];
    assign product[111] = s[110];
    assign product[112] = s[111];
    assign product[113] = s[112];
    assign product[114] = s[113];
    assign product[115] = s[114];
    assign product[116] = s[115];
    assign product[117] = s[116];
    assign product[118] = s[117];
    assign product[119] = s[118];
    assign product[120] = s[119];
    assign product[121] = s[120];
    assign product[122] = s[121];
    assign product[123] = s[122];
    assign product[124] = s[123];
    assign product[125] = s[124];
    assign product[126] = s[125];
    assign product[127] = c;
endmodule

module CLA256(output [255:0] sum, output cout, input [255:0] in1, input [255:0] in2;

    wire[255:0] G;
    wire[255:0] C;
    wire[255:0] P;

    assign G[0] = in[255] & in2[255];
    assign P[0] = in[255] ^ in2[255];
    assign G[1] = in[254] & in2[254];
    assign P[1] = in[254] ^ in2[254];
    assign G[2] = in[253] & in2[253];
    assign P[2] = in[253] ^ in2[253];
    assign G[3] = in[252] & in2[252];
    assign P[3] = in[252] ^ in2[252];
    assign G[4] = in[251] & in2[251];
    assign P[4] = in[251] ^ in2[251];
    assign G[5] = in[250] & in2[250];
    assign P[5] = in[250] ^ in2[250];
    assign G[6] = in[249] & in2[249];
    assign P[6] = in[249] ^ in2[249];
    assign G[7] = in[248] & in2[248];
    assign P[7] = in[248] ^ in2[248];
    assign G[8] = in[247] & in2[247];
    assign P[8] = in[247] ^ in2[247];
    assign G[9] = in[246] & in2[246];
    assign P[9] = in[246] ^ in2[246];
    assign G[10] = in[245] & in2[245];
    assign P[10] = in[245] ^ in2[245];
    assign G[11] = in[244] & in2[244];
    assign P[11] = in[244] ^ in2[244];
    assign G[12] = in[243] & in2[243];
    assign P[12] = in[243] ^ in2[243];
    assign G[13] = in[242] & in2[242];
    assign P[13] = in[242] ^ in2[242];
    assign G[14] = in[241] & in2[241];
    assign P[14] = in[241] ^ in2[241];
    assign G[15] = in[240] & in2[240];
    assign P[15] = in[240] ^ in2[240];
    assign G[16] = in[239] & in2[239];
    assign P[16] = in[239] ^ in2[239];
    assign G[17] = in[238] & in2[238];
    assign P[17] = in[238] ^ in2[238];
    assign G[18] = in[237] & in2[237];
    assign P[18] = in[237] ^ in2[237];
    assign G[19] = in[236] & in2[236];
    assign P[19] = in[236] ^ in2[236];
    assign G[20] = in[235] & in2[235];
    assign P[20] = in[235] ^ in2[235];
    assign G[21] = in[234] & in2[234];
    assign P[21] = in[234] ^ in2[234];
    assign G[22] = in[233] & in2[233];
    assign P[22] = in[233] ^ in2[233];
    assign G[23] = in[232] & in2[232];
    assign P[23] = in[232] ^ in2[232];
    assign G[24] = in[231] & in2[231];
    assign P[24] = in[231] ^ in2[231];
    assign G[25] = in[230] & in2[230];
    assign P[25] = in[230] ^ in2[230];
    assign G[26] = in[229] & in2[229];
    assign P[26] = in[229] ^ in2[229];
    assign G[27] = in[228] & in2[228];
    assign P[27] = in[228] ^ in2[228];
    assign G[28] = in[227] & in2[227];
    assign P[28] = in[227] ^ in2[227];
    assign G[29] = in[226] & in2[226];
    assign P[29] = in[226] ^ in2[226];
    assign G[30] = in[225] & in2[225];
    assign P[30] = in[225] ^ in2[225];
    assign G[31] = in[224] & in2[224];
    assign P[31] = in[224] ^ in2[224];
    assign G[32] = in[223] & in2[223];
    assign P[32] = in[223] ^ in2[223];
    assign G[33] = in[222] & in2[222];
    assign P[33] = in[222] ^ in2[222];
    assign G[34] = in[221] & in2[221];
    assign P[34] = in[221] ^ in2[221];
    assign G[35] = in[220] & in2[220];
    assign P[35] = in[220] ^ in2[220];
    assign G[36] = in[219] & in2[219];
    assign P[36] = in[219] ^ in2[219];
    assign G[37] = in[218] & in2[218];
    assign P[37] = in[218] ^ in2[218];
    assign G[38] = in[217] & in2[217];
    assign P[38] = in[217] ^ in2[217];
    assign G[39] = in[216] & in2[216];
    assign P[39] = in[216] ^ in2[216];
    assign G[40] = in[215] & in2[215];
    assign P[40] = in[215] ^ in2[215];
    assign G[41] = in[214] & in2[214];
    assign P[41] = in[214] ^ in2[214];
    assign G[42] = in[213] & in2[213];
    assign P[42] = in[213] ^ in2[213];
    assign G[43] = in[212] & in2[212];
    assign P[43] = in[212] ^ in2[212];
    assign G[44] = in[211] & in2[211];
    assign P[44] = in[211] ^ in2[211];
    assign G[45] = in[210] & in2[210];
    assign P[45] = in[210] ^ in2[210];
    assign G[46] = in[209] & in2[209];
    assign P[46] = in[209] ^ in2[209];
    assign G[47] = in[208] & in2[208];
    assign P[47] = in[208] ^ in2[208];
    assign G[48] = in[207] & in2[207];
    assign P[48] = in[207] ^ in2[207];
    assign G[49] = in[206] & in2[206];
    assign P[49] = in[206] ^ in2[206];
    assign G[50] = in[205] & in2[205];
    assign P[50] = in[205] ^ in2[205];
    assign G[51] = in[204] & in2[204];
    assign P[51] = in[204] ^ in2[204];
    assign G[52] = in[203] & in2[203];
    assign P[52] = in[203] ^ in2[203];
    assign G[53] = in[202] & in2[202];
    assign P[53] = in[202] ^ in2[202];
    assign G[54] = in[201] & in2[201];
    assign P[54] = in[201] ^ in2[201];
    assign G[55] = in[200] & in2[200];
    assign P[55] = in[200] ^ in2[200];
    assign G[56] = in[199] & in2[199];
    assign P[56] = in[199] ^ in2[199];
    assign G[57] = in[198] & in2[198];
    assign P[57] = in[198] ^ in2[198];
    assign G[58] = in[197] & in2[197];
    assign P[58] = in[197] ^ in2[197];
    assign G[59] = in[196] & in2[196];
    assign P[59] = in[196] ^ in2[196];
    assign G[60] = in[195] & in2[195];
    assign P[60] = in[195] ^ in2[195];
    assign G[61] = in[194] & in2[194];
    assign P[61] = in[194] ^ in2[194];
    assign G[62] = in[193] & in2[193];
    assign P[62] = in[193] ^ in2[193];
    assign G[63] = in[192] & in2[192];
    assign P[63] = in[192] ^ in2[192];
    assign G[64] = in[191] & in2[191];
    assign P[64] = in[191] ^ in2[191];
    assign G[65] = in[190] & in2[190];
    assign P[65] = in[190] ^ in2[190];
    assign G[66] = in[189] & in2[189];
    assign P[66] = in[189] ^ in2[189];
    assign G[67] = in[188] & in2[188];
    assign P[67] = in[188] ^ in2[188];
    assign G[68] = in[187] & in2[187];
    assign P[68] = in[187] ^ in2[187];
    assign G[69] = in[186] & in2[186];
    assign P[69] = in[186] ^ in2[186];
    assign G[70] = in[185] & in2[185];
    assign P[70] = in[185] ^ in2[185];
    assign G[71] = in[184] & in2[184];
    assign P[71] = in[184] ^ in2[184];
    assign G[72] = in[183] & in2[183];
    assign P[72] = in[183] ^ in2[183];
    assign G[73] = in[182] & in2[182];
    assign P[73] = in[182] ^ in2[182];
    assign G[74] = in[181] & in2[181];
    assign P[74] = in[181] ^ in2[181];
    assign G[75] = in[180] & in2[180];
    assign P[75] = in[180] ^ in2[180];
    assign G[76] = in[179] & in2[179];
    assign P[76] = in[179] ^ in2[179];
    assign G[77] = in[178] & in2[178];
    assign P[77] = in[178] ^ in2[178];
    assign G[78] = in[177] & in2[177];
    assign P[78] = in[177] ^ in2[177];
    assign G[79] = in[176] & in2[176];
    assign P[79] = in[176] ^ in2[176];
    assign G[80] = in[175] & in2[175];
    assign P[80] = in[175] ^ in2[175];
    assign G[81] = in[174] & in2[174];
    assign P[81] = in[174] ^ in2[174];
    assign G[82] = in[173] & in2[173];
    assign P[82] = in[173] ^ in2[173];
    assign G[83] = in[172] & in2[172];
    assign P[83] = in[172] ^ in2[172];
    assign G[84] = in[171] & in2[171];
    assign P[84] = in[171] ^ in2[171];
    assign G[85] = in[170] & in2[170];
    assign P[85] = in[170] ^ in2[170];
    assign G[86] = in[169] & in2[169];
    assign P[86] = in[169] ^ in2[169];
    assign G[87] = in[168] & in2[168];
    assign P[87] = in[168] ^ in2[168];
    assign G[88] = in[167] & in2[167];
    assign P[88] = in[167] ^ in2[167];
    assign G[89] = in[166] & in2[166];
    assign P[89] = in[166] ^ in2[166];
    assign G[90] = in[165] & in2[165];
    assign P[90] = in[165] ^ in2[165];
    assign G[91] = in[164] & in2[164];
    assign P[91] = in[164] ^ in2[164];
    assign G[92] = in[163] & in2[163];
    assign P[92] = in[163] ^ in2[163];
    assign G[93] = in[162] & in2[162];
    assign P[93] = in[162] ^ in2[162];
    assign G[94] = in[161] & in2[161];
    assign P[94] = in[161] ^ in2[161];
    assign G[95] = in[160] & in2[160];
    assign P[95] = in[160] ^ in2[160];
    assign G[96] = in[159] & in2[159];
    assign P[96] = in[159] ^ in2[159];
    assign G[97] = in[158] & in2[158];
    assign P[97] = in[158] ^ in2[158];
    assign G[98] = in[157] & in2[157];
    assign P[98] = in[157] ^ in2[157];
    assign G[99] = in[156] & in2[156];
    assign P[99] = in[156] ^ in2[156];
    assign G[100] = in[155] & in2[155];
    assign P[100] = in[155] ^ in2[155];
    assign G[101] = in[154] & in2[154];
    assign P[101] = in[154] ^ in2[154];
    assign G[102] = in[153] & in2[153];
    assign P[102] = in[153] ^ in2[153];
    assign G[103] = in[152] & in2[152];
    assign P[103] = in[152] ^ in2[152];
    assign G[104] = in[151] & in2[151];
    assign P[104] = in[151] ^ in2[151];
    assign G[105] = in[150] & in2[150];
    assign P[105] = in[150] ^ in2[150];
    assign G[106] = in[149] & in2[149];
    assign P[106] = in[149] ^ in2[149];
    assign G[107] = in[148] & in2[148];
    assign P[107] = in[148] ^ in2[148];
    assign G[108] = in[147] & in2[147];
    assign P[108] = in[147] ^ in2[147];
    assign G[109] = in[146] & in2[146];
    assign P[109] = in[146] ^ in2[146];
    assign G[110] = in[145] & in2[145];
    assign P[110] = in[145] ^ in2[145];
    assign G[111] = in[144] & in2[144];
    assign P[111] = in[144] ^ in2[144];
    assign G[112] = in[143] & in2[143];
    assign P[112] = in[143] ^ in2[143];
    assign G[113] = in[142] & in2[142];
    assign P[113] = in[142] ^ in2[142];
    assign G[114] = in[141] & in2[141];
    assign P[114] = in[141] ^ in2[141];
    assign G[115] = in[140] & in2[140];
    assign P[115] = in[140] ^ in2[140];
    assign G[116] = in[139] & in2[139];
    assign P[116] = in[139] ^ in2[139];
    assign G[117] = in[138] & in2[138];
    assign P[117] = in[138] ^ in2[138];
    assign G[118] = in[137] & in2[137];
    assign P[118] = in[137] ^ in2[137];
    assign G[119] = in[136] & in2[136];
    assign P[119] = in[136] ^ in2[136];
    assign G[120] = in[135] & in2[135];
    assign P[120] = in[135] ^ in2[135];
    assign G[121] = in[134] & in2[134];
    assign P[121] = in[134] ^ in2[134];
    assign G[122] = in[133] & in2[133];
    assign P[122] = in[133] ^ in2[133];
    assign G[123] = in[132] & in2[132];
    assign P[123] = in[132] ^ in2[132];
    assign G[124] = in[131] & in2[131];
    assign P[124] = in[131] ^ in2[131];
    assign G[125] = in[130] & in2[130];
    assign P[125] = in[130] ^ in2[130];
    assign G[126] = in[129] & in2[129];
    assign P[126] = in[129] ^ in2[129];
    assign G[127] = in[128] & in2[128];
    assign P[127] = in[128] ^ in2[128];
    assign G[128] = in[127] & in2[127];
    assign P[128] = in[127] ^ in2[127];
    assign G[129] = in[126] & in2[126];
    assign P[129] = in[126] ^ in2[126];
    assign G[130] = in[125] & in2[125];
    assign P[130] = in[125] ^ in2[125];
    assign G[131] = in[124] & in2[124];
    assign P[131] = in[124] ^ in2[124];
    assign G[132] = in[123] & in2[123];
    assign P[132] = in[123] ^ in2[123];
    assign G[133] = in[122] & in2[122];
    assign P[133] = in[122] ^ in2[122];
    assign G[134] = in[121] & in2[121];
    assign P[134] = in[121] ^ in2[121];
    assign G[135] = in[120] & in2[120];
    assign P[135] = in[120] ^ in2[120];
    assign G[136] = in[119] & in2[119];
    assign P[136] = in[119] ^ in2[119];
    assign G[137] = in[118] & in2[118];
    assign P[137] = in[118] ^ in2[118];
    assign G[138] = in[117] & in2[117];
    assign P[138] = in[117] ^ in2[117];
    assign G[139] = in[116] & in2[116];
    assign P[139] = in[116] ^ in2[116];
    assign G[140] = in[115] & in2[115];
    assign P[140] = in[115] ^ in2[115];
    assign G[141] = in[114] & in2[114];
    assign P[141] = in[114] ^ in2[114];
    assign G[142] = in[113] & in2[113];
    assign P[142] = in[113] ^ in2[113];
    assign G[143] = in[112] & in2[112];
    assign P[143] = in[112] ^ in2[112];
    assign G[144] = in[111] & in2[111];
    assign P[144] = in[111] ^ in2[111];
    assign G[145] = in[110] & in2[110];
    assign P[145] = in[110] ^ in2[110];
    assign G[146] = in[109] & in2[109];
    assign P[146] = in[109] ^ in2[109];
    assign G[147] = in[108] & in2[108];
    assign P[147] = in[108] ^ in2[108];
    assign G[148] = in[107] & in2[107];
    assign P[148] = in[107] ^ in2[107];
    assign G[149] = in[106] & in2[106];
    assign P[149] = in[106] ^ in2[106];
    assign G[150] = in[105] & in2[105];
    assign P[150] = in[105] ^ in2[105];
    assign G[151] = in[104] & in2[104];
    assign P[151] = in[104] ^ in2[104];
    assign G[152] = in[103] & in2[103];
    assign P[152] = in[103] ^ in2[103];
    assign G[153] = in[102] & in2[102];
    assign P[153] = in[102] ^ in2[102];
    assign G[154] = in[101] & in2[101];
    assign P[154] = in[101] ^ in2[101];
    assign G[155] = in[100] & in2[100];
    assign P[155] = in[100] ^ in2[100];
    assign G[156] = in[99] & in2[99];
    assign P[156] = in[99] ^ in2[99];
    assign G[157] = in[98] & in2[98];
    assign P[157] = in[98] ^ in2[98];
    assign G[158] = in[97] & in2[97];
    assign P[158] = in[97] ^ in2[97];
    assign G[159] = in[96] & in2[96];
    assign P[159] = in[96] ^ in2[96];
    assign G[160] = in[95] & in2[95];
    assign P[160] = in[95] ^ in2[95];
    assign G[161] = in[94] & in2[94];
    assign P[161] = in[94] ^ in2[94];
    assign G[162] = in[93] & in2[93];
    assign P[162] = in[93] ^ in2[93];
    assign G[163] = in[92] & in2[92];
    assign P[163] = in[92] ^ in2[92];
    assign G[164] = in[91] & in2[91];
    assign P[164] = in[91] ^ in2[91];
    assign G[165] = in[90] & in2[90];
    assign P[165] = in[90] ^ in2[90];
    assign G[166] = in[89] & in2[89];
    assign P[166] = in[89] ^ in2[89];
    assign G[167] = in[88] & in2[88];
    assign P[167] = in[88] ^ in2[88];
    assign G[168] = in[87] & in2[87];
    assign P[168] = in[87] ^ in2[87];
    assign G[169] = in[86] & in2[86];
    assign P[169] = in[86] ^ in2[86];
    assign G[170] = in[85] & in2[85];
    assign P[170] = in[85] ^ in2[85];
    assign G[171] = in[84] & in2[84];
    assign P[171] = in[84] ^ in2[84];
    assign G[172] = in[83] & in2[83];
    assign P[172] = in[83] ^ in2[83];
    assign G[173] = in[82] & in2[82];
    assign P[173] = in[82] ^ in2[82];
    assign G[174] = in[81] & in2[81];
    assign P[174] = in[81] ^ in2[81];
    assign G[175] = in[80] & in2[80];
    assign P[175] = in[80] ^ in2[80];
    assign G[176] = in[79] & in2[79];
    assign P[176] = in[79] ^ in2[79];
    assign G[177] = in[78] & in2[78];
    assign P[177] = in[78] ^ in2[78];
    assign G[178] = in[77] & in2[77];
    assign P[178] = in[77] ^ in2[77];
    assign G[179] = in[76] & in2[76];
    assign P[179] = in[76] ^ in2[76];
    assign G[180] = in[75] & in2[75];
    assign P[180] = in[75] ^ in2[75];
    assign G[181] = in[74] & in2[74];
    assign P[181] = in[74] ^ in2[74];
    assign G[182] = in[73] & in2[73];
    assign P[182] = in[73] ^ in2[73];
    assign G[183] = in[72] & in2[72];
    assign P[183] = in[72] ^ in2[72];
    assign G[184] = in[71] & in2[71];
    assign P[184] = in[71] ^ in2[71];
    assign G[185] = in[70] & in2[70];
    assign P[185] = in[70] ^ in2[70];
    assign G[186] = in[69] & in2[69];
    assign P[186] = in[69] ^ in2[69];
    assign G[187] = in[68] & in2[68];
    assign P[187] = in[68] ^ in2[68];
    assign G[188] = in[67] & in2[67];
    assign P[188] = in[67] ^ in2[67];
    assign G[189] = in[66] & in2[66];
    assign P[189] = in[66] ^ in2[66];
    assign G[190] = in[65] & in2[65];
    assign P[190] = in[65] ^ in2[65];
    assign G[191] = in[64] & in2[64];
    assign P[191] = in[64] ^ in2[64];
    assign G[192] = in[63] & in2[63];
    assign P[192] = in[63] ^ in2[63];
    assign G[193] = in[62] & in2[62];
    assign P[193] = in[62] ^ in2[62];
    assign G[194] = in[61] & in2[61];
    assign P[194] = in[61] ^ in2[61];
    assign G[195] = in[60] & in2[60];
    assign P[195] = in[60] ^ in2[60];
    assign G[196] = in[59] & in2[59];
    assign P[196] = in[59] ^ in2[59];
    assign G[197] = in[58] & in2[58];
    assign P[197] = in[58] ^ in2[58];
    assign G[198] = in[57] & in2[57];
    assign P[198] = in[57] ^ in2[57];
    assign G[199] = in[56] & in2[56];
    assign P[199] = in[56] ^ in2[56];
    assign G[200] = in[55] & in2[55];
    assign P[200] = in[55] ^ in2[55];
    assign G[201] = in[54] & in2[54];
    assign P[201] = in[54] ^ in2[54];
    assign G[202] = in[53] & in2[53];
    assign P[202] = in[53] ^ in2[53];
    assign G[203] = in[52] & in2[52];
    assign P[203] = in[52] ^ in2[52];
    assign G[204] = in[51] & in2[51];
    assign P[204] = in[51] ^ in2[51];
    assign G[205] = in[50] & in2[50];
    assign P[205] = in[50] ^ in2[50];
    assign G[206] = in[49] & in2[49];
    assign P[206] = in[49] ^ in2[49];
    assign G[207] = in[48] & in2[48];
    assign P[207] = in[48] ^ in2[48];
    assign G[208] = in[47] & in2[47];
    assign P[208] = in[47] ^ in2[47];
    assign G[209] = in[46] & in2[46];
    assign P[209] = in[46] ^ in2[46];
    assign G[210] = in[45] & in2[45];
    assign P[210] = in[45] ^ in2[45];
    assign G[211] = in[44] & in2[44];
    assign P[211] = in[44] ^ in2[44];
    assign G[212] = in[43] & in2[43];
    assign P[212] = in[43] ^ in2[43];
    assign G[213] = in[42] & in2[42];
    assign P[213] = in[42] ^ in2[42];
    assign G[214] = in[41] & in2[41];
    assign P[214] = in[41] ^ in2[41];
    assign G[215] = in[40] & in2[40];
    assign P[215] = in[40] ^ in2[40];
    assign G[216] = in[39] & in2[39];
    assign P[216] = in[39] ^ in2[39];
    assign G[217] = in[38] & in2[38];
    assign P[217] = in[38] ^ in2[38];
    assign G[218] = in[37] & in2[37];
    assign P[218] = in[37] ^ in2[37];
    assign G[219] = in[36] & in2[36];
    assign P[219] = in[36] ^ in2[36];
    assign G[220] = in[35] & in2[35];
    assign P[220] = in[35] ^ in2[35];
    assign G[221] = in[34] & in2[34];
    assign P[221] = in[34] ^ in2[34];
    assign G[222] = in[33] & in2[33];
    assign P[222] = in[33] ^ in2[33];
    assign G[223] = in[32] & in2[32];
    assign P[223] = in[32] ^ in2[32];
    assign G[224] = in[31] & in2[31];
    assign P[224] = in[31] ^ in2[31];
    assign G[225] = in[30] & in2[30];
    assign P[225] = in[30] ^ in2[30];
    assign G[226] = in[29] & in2[29];
    assign P[226] = in[29] ^ in2[29];
    assign G[227] = in[28] & in2[28];
    assign P[227] = in[28] ^ in2[28];
    assign G[228] = in[27] & in2[27];
    assign P[228] = in[27] ^ in2[27];
    assign G[229] = in[26] & in2[26];
    assign P[229] = in[26] ^ in2[26];
    assign G[230] = in[25] & in2[25];
    assign P[230] = in[25] ^ in2[25];
    assign G[231] = in[24] & in2[24];
    assign P[231] = in[24] ^ in2[24];
    assign G[232] = in[23] & in2[23];
    assign P[232] = in[23] ^ in2[23];
    assign G[233] = in[22] & in2[22];
    assign P[233] = in[22] ^ in2[22];
    assign G[234] = in[21] & in2[21];
    assign P[234] = in[21] ^ in2[21];
    assign G[235] = in[20] & in2[20];
    assign P[235] = in[20] ^ in2[20];
    assign G[236] = in[19] & in2[19];
    assign P[236] = in[19] ^ in2[19];
    assign G[237] = in[18] & in2[18];
    assign P[237] = in[18] ^ in2[18];
    assign G[238] = in[17] & in2[17];
    assign P[238] = in[17] ^ in2[17];
    assign G[239] = in[16] & in2[16];
    assign P[239] = in[16] ^ in2[16];
    assign G[240] = in[15] & in2[15];
    assign P[240] = in[15] ^ in2[15];
    assign G[241] = in[14] & in2[14];
    assign P[241] = in[14] ^ in2[14];
    assign G[242] = in[13] & in2[13];
    assign P[242] = in[13] ^ in2[13];
    assign G[243] = in[12] & in2[12];
    assign P[243] = in[12] ^ in2[12];
    assign G[244] = in[11] & in2[11];
    assign P[244] = in[11] ^ in2[11];
    assign G[245] = in[10] & in2[10];
    assign P[245] = in[10] ^ in2[10];
    assign G[246] = in[9] & in2[9];
    assign P[246] = in[9] ^ in2[9];
    assign G[247] = in[8] & in2[8];
    assign P[247] = in[8] ^ in2[8];
    assign G[248] = in[7] & in2[7];
    assign P[248] = in[7] ^ in2[7];
    assign G[249] = in[6] & in2[6];
    assign P[249] = in[6] ^ in2[6];
    assign G[250] = in[5] & in2[5];
    assign P[250] = in[5] ^ in2[5];
    assign G[251] = in[4] & in2[4];
    assign P[251] = in[4] ^ in2[4];
    assign G[252] = in[3] & in2[3];
    assign P[252] = in[3] ^ in2[3];
    assign G[253] = in[2] & in2[2];
    assign P[253] = in[2] ^ in2[2];
    assign G[254] = in[1] & in2[1];
    assign P[254] = in[1] ^ in2[1];
    assign G[255] = in[0] & in2[0];
    assign P[255] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign C[252] = G[251] | (P[251] & C[251]);
    assign C[253] = G[252] | (P[252] & C[252]);
    assign C[254] = G[253] | (P[253] & C[253]);
    assign C[255] = G[254] | (P[254] & C[254]);
    assign cout = G[255] | (P[255] & C[255]);
    assign sum = P ^ C;
endmodule

module CLA255(output [254:0] sum, output cout, input [254:0] in1, input [254:0] in2;

    wire[254:0] G;
    wire[254:0] C;
    wire[254:0] P;

    assign G[0] = in[254] & in2[254];
    assign P[0] = in[254] ^ in2[254];
    assign G[1] = in[253] & in2[253];
    assign P[1] = in[253] ^ in2[253];
    assign G[2] = in[252] & in2[252];
    assign P[2] = in[252] ^ in2[252];
    assign G[3] = in[251] & in2[251];
    assign P[3] = in[251] ^ in2[251];
    assign G[4] = in[250] & in2[250];
    assign P[4] = in[250] ^ in2[250];
    assign G[5] = in[249] & in2[249];
    assign P[5] = in[249] ^ in2[249];
    assign G[6] = in[248] & in2[248];
    assign P[6] = in[248] ^ in2[248];
    assign G[7] = in[247] & in2[247];
    assign P[7] = in[247] ^ in2[247];
    assign G[8] = in[246] & in2[246];
    assign P[8] = in[246] ^ in2[246];
    assign G[9] = in[245] & in2[245];
    assign P[9] = in[245] ^ in2[245];
    assign G[10] = in[244] & in2[244];
    assign P[10] = in[244] ^ in2[244];
    assign G[11] = in[243] & in2[243];
    assign P[11] = in[243] ^ in2[243];
    assign G[12] = in[242] & in2[242];
    assign P[12] = in[242] ^ in2[242];
    assign G[13] = in[241] & in2[241];
    assign P[13] = in[241] ^ in2[241];
    assign G[14] = in[240] & in2[240];
    assign P[14] = in[240] ^ in2[240];
    assign G[15] = in[239] & in2[239];
    assign P[15] = in[239] ^ in2[239];
    assign G[16] = in[238] & in2[238];
    assign P[16] = in[238] ^ in2[238];
    assign G[17] = in[237] & in2[237];
    assign P[17] = in[237] ^ in2[237];
    assign G[18] = in[236] & in2[236];
    assign P[18] = in[236] ^ in2[236];
    assign G[19] = in[235] & in2[235];
    assign P[19] = in[235] ^ in2[235];
    assign G[20] = in[234] & in2[234];
    assign P[20] = in[234] ^ in2[234];
    assign G[21] = in[233] & in2[233];
    assign P[21] = in[233] ^ in2[233];
    assign G[22] = in[232] & in2[232];
    assign P[22] = in[232] ^ in2[232];
    assign G[23] = in[231] & in2[231];
    assign P[23] = in[231] ^ in2[231];
    assign G[24] = in[230] & in2[230];
    assign P[24] = in[230] ^ in2[230];
    assign G[25] = in[229] & in2[229];
    assign P[25] = in[229] ^ in2[229];
    assign G[26] = in[228] & in2[228];
    assign P[26] = in[228] ^ in2[228];
    assign G[27] = in[227] & in2[227];
    assign P[27] = in[227] ^ in2[227];
    assign G[28] = in[226] & in2[226];
    assign P[28] = in[226] ^ in2[226];
    assign G[29] = in[225] & in2[225];
    assign P[29] = in[225] ^ in2[225];
    assign G[30] = in[224] & in2[224];
    assign P[30] = in[224] ^ in2[224];
    assign G[31] = in[223] & in2[223];
    assign P[31] = in[223] ^ in2[223];
    assign G[32] = in[222] & in2[222];
    assign P[32] = in[222] ^ in2[222];
    assign G[33] = in[221] & in2[221];
    assign P[33] = in[221] ^ in2[221];
    assign G[34] = in[220] & in2[220];
    assign P[34] = in[220] ^ in2[220];
    assign G[35] = in[219] & in2[219];
    assign P[35] = in[219] ^ in2[219];
    assign G[36] = in[218] & in2[218];
    assign P[36] = in[218] ^ in2[218];
    assign G[37] = in[217] & in2[217];
    assign P[37] = in[217] ^ in2[217];
    assign G[38] = in[216] & in2[216];
    assign P[38] = in[216] ^ in2[216];
    assign G[39] = in[215] & in2[215];
    assign P[39] = in[215] ^ in2[215];
    assign G[40] = in[214] & in2[214];
    assign P[40] = in[214] ^ in2[214];
    assign G[41] = in[213] & in2[213];
    assign P[41] = in[213] ^ in2[213];
    assign G[42] = in[212] & in2[212];
    assign P[42] = in[212] ^ in2[212];
    assign G[43] = in[211] & in2[211];
    assign P[43] = in[211] ^ in2[211];
    assign G[44] = in[210] & in2[210];
    assign P[44] = in[210] ^ in2[210];
    assign G[45] = in[209] & in2[209];
    assign P[45] = in[209] ^ in2[209];
    assign G[46] = in[208] & in2[208];
    assign P[46] = in[208] ^ in2[208];
    assign G[47] = in[207] & in2[207];
    assign P[47] = in[207] ^ in2[207];
    assign G[48] = in[206] & in2[206];
    assign P[48] = in[206] ^ in2[206];
    assign G[49] = in[205] & in2[205];
    assign P[49] = in[205] ^ in2[205];
    assign G[50] = in[204] & in2[204];
    assign P[50] = in[204] ^ in2[204];
    assign G[51] = in[203] & in2[203];
    assign P[51] = in[203] ^ in2[203];
    assign G[52] = in[202] & in2[202];
    assign P[52] = in[202] ^ in2[202];
    assign G[53] = in[201] & in2[201];
    assign P[53] = in[201] ^ in2[201];
    assign G[54] = in[200] & in2[200];
    assign P[54] = in[200] ^ in2[200];
    assign G[55] = in[199] & in2[199];
    assign P[55] = in[199] ^ in2[199];
    assign G[56] = in[198] & in2[198];
    assign P[56] = in[198] ^ in2[198];
    assign G[57] = in[197] & in2[197];
    assign P[57] = in[197] ^ in2[197];
    assign G[58] = in[196] & in2[196];
    assign P[58] = in[196] ^ in2[196];
    assign G[59] = in[195] & in2[195];
    assign P[59] = in[195] ^ in2[195];
    assign G[60] = in[194] & in2[194];
    assign P[60] = in[194] ^ in2[194];
    assign G[61] = in[193] & in2[193];
    assign P[61] = in[193] ^ in2[193];
    assign G[62] = in[192] & in2[192];
    assign P[62] = in[192] ^ in2[192];
    assign G[63] = in[191] & in2[191];
    assign P[63] = in[191] ^ in2[191];
    assign G[64] = in[190] & in2[190];
    assign P[64] = in[190] ^ in2[190];
    assign G[65] = in[189] & in2[189];
    assign P[65] = in[189] ^ in2[189];
    assign G[66] = in[188] & in2[188];
    assign P[66] = in[188] ^ in2[188];
    assign G[67] = in[187] & in2[187];
    assign P[67] = in[187] ^ in2[187];
    assign G[68] = in[186] & in2[186];
    assign P[68] = in[186] ^ in2[186];
    assign G[69] = in[185] & in2[185];
    assign P[69] = in[185] ^ in2[185];
    assign G[70] = in[184] & in2[184];
    assign P[70] = in[184] ^ in2[184];
    assign G[71] = in[183] & in2[183];
    assign P[71] = in[183] ^ in2[183];
    assign G[72] = in[182] & in2[182];
    assign P[72] = in[182] ^ in2[182];
    assign G[73] = in[181] & in2[181];
    assign P[73] = in[181] ^ in2[181];
    assign G[74] = in[180] & in2[180];
    assign P[74] = in[180] ^ in2[180];
    assign G[75] = in[179] & in2[179];
    assign P[75] = in[179] ^ in2[179];
    assign G[76] = in[178] & in2[178];
    assign P[76] = in[178] ^ in2[178];
    assign G[77] = in[177] & in2[177];
    assign P[77] = in[177] ^ in2[177];
    assign G[78] = in[176] & in2[176];
    assign P[78] = in[176] ^ in2[176];
    assign G[79] = in[175] & in2[175];
    assign P[79] = in[175] ^ in2[175];
    assign G[80] = in[174] & in2[174];
    assign P[80] = in[174] ^ in2[174];
    assign G[81] = in[173] & in2[173];
    assign P[81] = in[173] ^ in2[173];
    assign G[82] = in[172] & in2[172];
    assign P[82] = in[172] ^ in2[172];
    assign G[83] = in[171] & in2[171];
    assign P[83] = in[171] ^ in2[171];
    assign G[84] = in[170] & in2[170];
    assign P[84] = in[170] ^ in2[170];
    assign G[85] = in[169] & in2[169];
    assign P[85] = in[169] ^ in2[169];
    assign G[86] = in[168] & in2[168];
    assign P[86] = in[168] ^ in2[168];
    assign G[87] = in[167] & in2[167];
    assign P[87] = in[167] ^ in2[167];
    assign G[88] = in[166] & in2[166];
    assign P[88] = in[166] ^ in2[166];
    assign G[89] = in[165] & in2[165];
    assign P[89] = in[165] ^ in2[165];
    assign G[90] = in[164] & in2[164];
    assign P[90] = in[164] ^ in2[164];
    assign G[91] = in[163] & in2[163];
    assign P[91] = in[163] ^ in2[163];
    assign G[92] = in[162] & in2[162];
    assign P[92] = in[162] ^ in2[162];
    assign G[93] = in[161] & in2[161];
    assign P[93] = in[161] ^ in2[161];
    assign G[94] = in[160] & in2[160];
    assign P[94] = in[160] ^ in2[160];
    assign G[95] = in[159] & in2[159];
    assign P[95] = in[159] ^ in2[159];
    assign G[96] = in[158] & in2[158];
    assign P[96] = in[158] ^ in2[158];
    assign G[97] = in[157] & in2[157];
    assign P[97] = in[157] ^ in2[157];
    assign G[98] = in[156] & in2[156];
    assign P[98] = in[156] ^ in2[156];
    assign G[99] = in[155] & in2[155];
    assign P[99] = in[155] ^ in2[155];
    assign G[100] = in[154] & in2[154];
    assign P[100] = in[154] ^ in2[154];
    assign G[101] = in[153] & in2[153];
    assign P[101] = in[153] ^ in2[153];
    assign G[102] = in[152] & in2[152];
    assign P[102] = in[152] ^ in2[152];
    assign G[103] = in[151] & in2[151];
    assign P[103] = in[151] ^ in2[151];
    assign G[104] = in[150] & in2[150];
    assign P[104] = in[150] ^ in2[150];
    assign G[105] = in[149] & in2[149];
    assign P[105] = in[149] ^ in2[149];
    assign G[106] = in[148] & in2[148];
    assign P[106] = in[148] ^ in2[148];
    assign G[107] = in[147] & in2[147];
    assign P[107] = in[147] ^ in2[147];
    assign G[108] = in[146] & in2[146];
    assign P[108] = in[146] ^ in2[146];
    assign G[109] = in[145] & in2[145];
    assign P[109] = in[145] ^ in2[145];
    assign G[110] = in[144] & in2[144];
    assign P[110] = in[144] ^ in2[144];
    assign G[111] = in[143] & in2[143];
    assign P[111] = in[143] ^ in2[143];
    assign G[112] = in[142] & in2[142];
    assign P[112] = in[142] ^ in2[142];
    assign G[113] = in[141] & in2[141];
    assign P[113] = in[141] ^ in2[141];
    assign G[114] = in[140] & in2[140];
    assign P[114] = in[140] ^ in2[140];
    assign G[115] = in[139] & in2[139];
    assign P[115] = in[139] ^ in2[139];
    assign G[116] = in[138] & in2[138];
    assign P[116] = in[138] ^ in2[138];
    assign G[117] = in[137] & in2[137];
    assign P[117] = in[137] ^ in2[137];
    assign G[118] = in[136] & in2[136];
    assign P[118] = in[136] ^ in2[136];
    assign G[119] = in[135] & in2[135];
    assign P[119] = in[135] ^ in2[135];
    assign G[120] = in[134] & in2[134];
    assign P[120] = in[134] ^ in2[134];
    assign G[121] = in[133] & in2[133];
    assign P[121] = in[133] ^ in2[133];
    assign G[122] = in[132] & in2[132];
    assign P[122] = in[132] ^ in2[132];
    assign G[123] = in[131] & in2[131];
    assign P[123] = in[131] ^ in2[131];
    assign G[124] = in[130] & in2[130];
    assign P[124] = in[130] ^ in2[130];
    assign G[125] = in[129] & in2[129];
    assign P[125] = in[129] ^ in2[129];
    assign G[126] = in[128] & in2[128];
    assign P[126] = in[128] ^ in2[128];
    assign G[127] = in[127] & in2[127];
    assign P[127] = in[127] ^ in2[127];
    assign G[128] = in[126] & in2[126];
    assign P[128] = in[126] ^ in2[126];
    assign G[129] = in[125] & in2[125];
    assign P[129] = in[125] ^ in2[125];
    assign G[130] = in[124] & in2[124];
    assign P[130] = in[124] ^ in2[124];
    assign G[131] = in[123] & in2[123];
    assign P[131] = in[123] ^ in2[123];
    assign G[132] = in[122] & in2[122];
    assign P[132] = in[122] ^ in2[122];
    assign G[133] = in[121] & in2[121];
    assign P[133] = in[121] ^ in2[121];
    assign G[134] = in[120] & in2[120];
    assign P[134] = in[120] ^ in2[120];
    assign G[135] = in[119] & in2[119];
    assign P[135] = in[119] ^ in2[119];
    assign G[136] = in[118] & in2[118];
    assign P[136] = in[118] ^ in2[118];
    assign G[137] = in[117] & in2[117];
    assign P[137] = in[117] ^ in2[117];
    assign G[138] = in[116] & in2[116];
    assign P[138] = in[116] ^ in2[116];
    assign G[139] = in[115] & in2[115];
    assign P[139] = in[115] ^ in2[115];
    assign G[140] = in[114] & in2[114];
    assign P[140] = in[114] ^ in2[114];
    assign G[141] = in[113] & in2[113];
    assign P[141] = in[113] ^ in2[113];
    assign G[142] = in[112] & in2[112];
    assign P[142] = in[112] ^ in2[112];
    assign G[143] = in[111] & in2[111];
    assign P[143] = in[111] ^ in2[111];
    assign G[144] = in[110] & in2[110];
    assign P[144] = in[110] ^ in2[110];
    assign G[145] = in[109] & in2[109];
    assign P[145] = in[109] ^ in2[109];
    assign G[146] = in[108] & in2[108];
    assign P[146] = in[108] ^ in2[108];
    assign G[147] = in[107] & in2[107];
    assign P[147] = in[107] ^ in2[107];
    assign G[148] = in[106] & in2[106];
    assign P[148] = in[106] ^ in2[106];
    assign G[149] = in[105] & in2[105];
    assign P[149] = in[105] ^ in2[105];
    assign G[150] = in[104] & in2[104];
    assign P[150] = in[104] ^ in2[104];
    assign G[151] = in[103] & in2[103];
    assign P[151] = in[103] ^ in2[103];
    assign G[152] = in[102] & in2[102];
    assign P[152] = in[102] ^ in2[102];
    assign G[153] = in[101] & in2[101];
    assign P[153] = in[101] ^ in2[101];
    assign G[154] = in[100] & in2[100];
    assign P[154] = in[100] ^ in2[100];
    assign G[155] = in[99] & in2[99];
    assign P[155] = in[99] ^ in2[99];
    assign G[156] = in[98] & in2[98];
    assign P[156] = in[98] ^ in2[98];
    assign G[157] = in[97] & in2[97];
    assign P[157] = in[97] ^ in2[97];
    assign G[158] = in[96] & in2[96];
    assign P[158] = in[96] ^ in2[96];
    assign G[159] = in[95] & in2[95];
    assign P[159] = in[95] ^ in2[95];
    assign G[160] = in[94] & in2[94];
    assign P[160] = in[94] ^ in2[94];
    assign G[161] = in[93] & in2[93];
    assign P[161] = in[93] ^ in2[93];
    assign G[162] = in[92] & in2[92];
    assign P[162] = in[92] ^ in2[92];
    assign G[163] = in[91] & in2[91];
    assign P[163] = in[91] ^ in2[91];
    assign G[164] = in[90] & in2[90];
    assign P[164] = in[90] ^ in2[90];
    assign G[165] = in[89] & in2[89];
    assign P[165] = in[89] ^ in2[89];
    assign G[166] = in[88] & in2[88];
    assign P[166] = in[88] ^ in2[88];
    assign G[167] = in[87] & in2[87];
    assign P[167] = in[87] ^ in2[87];
    assign G[168] = in[86] & in2[86];
    assign P[168] = in[86] ^ in2[86];
    assign G[169] = in[85] & in2[85];
    assign P[169] = in[85] ^ in2[85];
    assign G[170] = in[84] & in2[84];
    assign P[170] = in[84] ^ in2[84];
    assign G[171] = in[83] & in2[83];
    assign P[171] = in[83] ^ in2[83];
    assign G[172] = in[82] & in2[82];
    assign P[172] = in[82] ^ in2[82];
    assign G[173] = in[81] & in2[81];
    assign P[173] = in[81] ^ in2[81];
    assign G[174] = in[80] & in2[80];
    assign P[174] = in[80] ^ in2[80];
    assign G[175] = in[79] & in2[79];
    assign P[175] = in[79] ^ in2[79];
    assign G[176] = in[78] & in2[78];
    assign P[176] = in[78] ^ in2[78];
    assign G[177] = in[77] & in2[77];
    assign P[177] = in[77] ^ in2[77];
    assign G[178] = in[76] & in2[76];
    assign P[178] = in[76] ^ in2[76];
    assign G[179] = in[75] & in2[75];
    assign P[179] = in[75] ^ in2[75];
    assign G[180] = in[74] & in2[74];
    assign P[180] = in[74] ^ in2[74];
    assign G[181] = in[73] & in2[73];
    assign P[181] = in[73] ^ in2[73];
    assign G[182] = in[72] & in2[72];
    assign P[182] = in[72] ^ in2[72];
    assign G[183] = in[71] & in2[71];
    assign P[183] = in[71] ^ in2[71];
    assign G[184] = in[70] & in2[70];
    assign P[184] = in[70] ^ in2[70];
    assign G[185] = in[69] & in2[69];
    assign P[185] = in[69] ^ in2[69];
    assign G[186] = in[68] & in2[68];
    assign P[186] = in[68] ^ in2[68];
    assign G[187] = in[67] & in2[67];
    assign P[187] = in[67] ^ in2[67];
    assign G[188] = in[66] & in2[66];
    assign P[188] = in[66] ^ in2[66];
    assign G[189] = in[65] & in2[65];
    assign P[189] = in[65] ^ in2[65];
    assign G[190] = in[64] & in2[64];
    assign P[190] = in[64] ^ in2[64];
    assign G[191] = in[63] & in2[63];
    assign P[191] = in[63] ^ in2[63];
    assign G[192] = in[62] & in2[62];
    assign P[192] = in[62] ^ in2[62];
    assign G[193] = in[61] & in2[61];
    assign P[193] = in[61] ^ in2[61];
    assign G[194] = in[60] & in2[60];
    assign P[194] = in[60] ^ in2[60];
    assign G[195] = in[59] & in2[59];
    assign P[195] = in[59] ^ in2[59];
    assign G[196] = in[58] & in2[58];
    assign P[196] = in[58] ^ in2[58];
    assign G[197] = in[57] & in2[57];
    assign P[197] = in[57] ^ in2[57];
    assign G[198] = in[56] & in2[56];
    assign P[198] = in[56] ^ in2[56];
    assign G[199] = in[55] & in2[55];
    assign P[199] = in[55] ^ in2[55];
    assign G[200] = in[54] & in2[54];
    assign P[200] = in[54] ^ in2[54];
    assign G[201] = in[53] & in2[53];
    assign P[201] = in[53] ^ in2[53];
    assign G[202] = in[52] & in2[52];
    assign P[202] = in[52] ^ in2[52];
    assign G[203] = in[51] & in2[51];
    assign P[203] = in[51] ^ in2[51];
    assign G[204] = in[50] & in2[50];
    assign P[204] = in[50] ^ in2[50];
    assign G[205] = in[49] & in2[49];
    assign P[205] = in[49] ^ in2[49];
    assign G[206] = in[48] & in2[48];
    assign P[206] = in[48] ^ in2[48];
    assign G[207] = in[47] & in2[47];
    assign P[207] = in[47] ^ in2[47];
    assign G[208] = in[46] & in2[46];
    assign P[208] = in[46] ^ in2[46];
    assign G[209] = in[45] & in2[45];
    assign P[209] = in[45] ^ in2[45];
    assign G[210] = in[44] & in2[44];
    assign P[210] = in[44] ^ in2[44];
    assign G[211] = in[43] & in2[43];
    assign P[211] = in[43] ^ in2[43];
    assign G[212] = in[42] & in2[42];
    assign P[212] = in[42] ^ in2[42];
    assign G[213] = in[41] & in2[41];
    assign P[213] = in[41] ^ in2[41];
    assign G[214] = in[40] & in2[40];
    assign P[214] = in[40] ^ in2[40];
    assign G[215] = in[39] & in2[39];
    assign P[215] = in[39] ^ in2[39];
    assign G[216] = in[38] & in2[38];
    assign P[216] = in[38] ^ in2[38];
    assign G[217] = in[37] & in2[37];
    assign P[217] = in[37] ^ in2[37];
    assign G[218] = in[36] & in2[36];
    assign P[218] = in[36] ^ in2[36];
    assign G[219] = in[35] & in2[35];
    assign P[219] = in[35] ^ in2[35];
    assign G[220] = in[34] & in2[34];
    assign P[220] = in[34] ^ in2[34];
    assign G[221] = in[33] & in2[33];
    assign P[221] = in[33] ^ in2[33];
    assign G[222] = in[32] & in2[32];
    assign P[222] = in[32] ^ in2[32];
    assign G[223] = in[31] & in2[31];
    assign P[223] = in[31] ^ in2[31];
    assign G[224] = in[30] & in2[30];
    assign P[224] = in[30] ^ in2[30];
    assign G[225] = in[29] & in2[29];
    assign P[225] = in[29] ^ in2[29];
    assign G[226] = in[28] & in2[28];
    assign P[226] = in[28] ^ in2[28];
    assign G[227] = in[27] & in2[27];
    assign P[227] = in[27] ^ in2[27];
    assign G[228] = in[26] & in2[26];
    assign P[228] = in[26] ^ in2[26];
    assign G[229] = in[25] & in2[25];
    assign P[229] = in[25] ^ in2[25];
    assign G[230] = in[24] & in2[24];
    assign P[230] = in[24] ^ in2[24];
    assign G[231] = in[23] & in2[23];
    assign P[231] = in[23] ^ in2[23];
    assign G[232] = in[22] & in2[22];
    assign P[232] = in[22] ^ in2[22];
    assign G[233] = in[21] & in2[21];
    assign P[233] = in[21] ^ in2[21];
    assign G[234] = in[20] & in2[20];
    assign P[234] = in[20] ^ in2[20];
    assign G[235] = in[19] & in2[19];
    assign P[235] = in[19] ^ in2[19];
    assign G[236] = in[18] & in2[18];
    assign P[236] = in[18] ^ in2[18];
    assign G[237] = in[17] & in2[17];
    assign P[237] = in[17] ^ in2[17];
    assign G[238] = in[16] & in2[16];
    assign P[238] = in[16] ^ in2[16];
    assign G[239] = in[15] & in2[15];
    assign P[239] = in[15] ^ in2[15];
    assign G[240] = in[14] & in2[14];
    assign P[240] = in[14] ^ in2[14];
    assign G[241] = in[13] & in2[13];
    assign P[241] = in[13] ^ in2[13];
    assign G[242] = in[12] & in2[12];
    assign P[242] = in[12] ^ in2[12];
    assign G[243] = in[11] & in2[11];
    assign P[243] = in[11] ^ in2[11];
    assign G[244] = in[10] & in2[10];
    assign P[244] = in[10] ^ in2[10];
    assign G[245] = in[9] & in2[9];
    assign P[245] = in[9] ^ in2[9];
    assign G[246] = in[8] & in2[8];
    assign P[246] = in[8] ^ in2[8];
    assign G[247] = in[7] & in2[7];
    assign P[247] = in[7] ^ in2[7];
    assign G[248] = in[6] & in2[6];
    assign P[248] = in[6] ^ in2[6];
    assign G[249] = in[5] & in2[5];
    assign P[249] = in[5] ^ in2[5];
    assign G[250] = in[4] & in2[4];
    assign P[250] = in[4] ^ in2[4];
    assign G[251] = in[3] & in2[3];
    assign P[251] = in[3] ^ in2[3];
    assign G[252] = in[2] & in2[2];
    assign P[252] = in[2] ^ in2[2];
    assign G[253] = in[1] & in2[1];
    assign P[253] = in[1] ^ in2[1];
    assign G[254] = in[0] & in2[0];
    assign P[254] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign C[252] = G[251] | (P[251] & C[251]);
    assign C[253] = G[252] | (P[252] & C[252]);
    assign C[254] = G[253] | (P[253] & C[253]);
    assign cout = G[254] | (P[254] & C[254]);
    assign sum = P ^ C;
endmodule

module CLA254(output [253:0] sum, output cout, input [253:0] in1, input [253:0] in2;

    wire[253:0] G;
    wire[253:0] C;
    wire[253:0] P;

    assign G[0] = in[253] & in2[253];
    assign P[0] = in[253] ^ in2[253];
    assign G[1] = in[252] & in2[252];
    assign P[1] = in[252] ^ in2[252];
    assign G[2] = in[251] & in2[251];
    assign P[2] = in[251] ^ in2[251];
    assign G[3] = in[250] & in2[250];
    assign P[3] = in[250] ^ in2[250];
    assign G[4] = in[249] & in2[249];
    assign P[4] = in[249] ^ in2[249];
    assign G[5] = in[248] & in2[248];
    assign P[5] = in[248] ^ in2[248];
    assign G[6] = in[247] & in2[247];
    assign P[6] = in[247] ^ in2[247];
    assign G[7] = in[246] & in2[246];
    assign P[7] = in[246] ^ in2[246];
    assign G[8] = in[245] & in2[245];
    assign P[8] = in[245] ^ in2[245];
    assign G[9] = in[244] & in2[244];
    assign P[9] = in[244] ^ in2[244];
    assign G[10] = in[243] & in2[243];
    assign P[10] = in[243] ^ in2[243];
    assign G[11] = in[242] & in2[242];
    assign P[11] = in[242] ^ in2[242];
    assign G[12] = in[241] & in2[241];
    assign P[12] = in[241] ^ in2[241];
    assign G[13] = in[240] & in2[240];
    assign P[13] = in[240] ^ in2[240];
    assign G[14] = in[239] & in2[239];
    assign P[14] = in[239] ^ in2[239];
    assign G[15] = in[238] & in2[238];
    assign P[15] = in[238] ^ in2[238];
    assign G[16] = in[237] & in2[237];
    assign P[16] = in[237] ^ in2[237];
    assign G[17] = in[236] & in2[236];
    assign P[17] = in[236] ^ in2[236];
    assign G[18] = in[235] & in2[235];
    assign P[18] = in[235] ^ in2[235];
    assign G[19] = in[234] & in2[234];
    assign P[19] = in[234] ^ in2[234];
    assign G[20] = in[233] & in2[233];
    assign P[20] = in[233] ^ in2[233];
    assign G[21] = in[232] & in2[232];
    assign P[21] = in[232] ^ in2[232];
    assign G[22] = in[231] & in2[231];
    assign P[22] = in[231] ^ in2[231];
    assign G[23] = in[230] & in2[230];
    assign P[23] = in[230] ^ in2[230];
    assign G[24] = in[229] & in2[229];
    assign P[24] = in[229] ^ in2[229];
    assign G[25] = in[228] & in2[228];
    assign P[25] = in[228] ^ in2[228];
    assign G[26] = in[227] & in2[227];
    assign P[26] = in[227] ^ in2[227];
    assign G[27] = in[226] & in2[226];
    assign P[27] = in[226] ^ in2[226];
    assign G[28] = in[225] & in2[225];
    assign P[28] = in[225] ^ in2[225];
    assign G[29] = in[224] & in2[224];
    assign P[29] = in[224] ^ in2[224];
    assign G[30] = in[223] & in2[223];
    assign P[30] = in[223] ^ in2[223];
    assign G[31] = in[222] & in2[222];
    assign P[31] = in[222] ^ in2[222];
    assign G[32] = in[221] & in2[221];
    assign P[32] = in[221] ^ in2[221];
    assign G[33] = in[220] & in2[220];
    assign P[33] = in[220] ^ in2[220];
    assign G[34] = in[219] & in2[219];
    assign P[34] = in[219] ^ in2[219];
    assign G[35] = in[218] & in2[218];
    assign P[35] = in[218] ^ in2[218];
    assign G[36] = in[217] & in2[217];
    assign P[36] = in[217] ^ in2[217];
    assign G[37] = in[216] & in2[216];
    assign P[37] = in[216] ^ in2[216];
    assign G[38] = in[215] & in2[215];
    assign P[38] = in[215] ^ in2[215];
    assign G[39] = in[214] & in2[214];
    assign P[39] = in[214] ^ in2[214];
    assign G[40] = in[213] & in2[213];
    assign P[40] = in[213] ^ in2[213];
    assign G[41] = in[212] & in2[212];
    assign P[41] = in[212] ^ in2[212];
    assign G[42] = in[211] & in2[211];
    assign P[42] = in[211] ^ in2[211];
    assign G[43] = in[210] & in2[210];
    assign P[43] = in[210] ^ in2[210];
    assign G[44] = in[209] & in2[209];
    assign P[44] = in[209] ^ in2[209];
    assign G[45] = in[208] & in2[208];
    assign P[45] = in[208] ^ in2[208];
    assign G[46] = in[207] & in2[207];
    assign P[46] = in[207] ^ in2[207];
    assign G[47] = in[206] & in2[206];
    assign P[47] = in[206] ^ in2[206];
    assign G[48] = in[205] & in2[205];
    assign P[48] = in[205] ^ in2[205];
    assign G[49] = in[204] & in2[204];
    assign P[49] = in[204] ^ in2[204];
    assign G[50] = in[203] & in2[203];
    assign P[50] = in[203] ^ in2[203];
    assign G[51] = in[202] & in2[202];
    assign P[51] = in[202] ^ in2[202];
    assign G[52] = in[201] & in2[201];
    assign P[52] = in[201] ^ in2[201];
    assign G[53] = in[200] & in2[200];
    assign P[53] = in[200] ^ in2[200];
    assign G[54] = in[199] & in2[199];
    assign P[54] = in[199] ^ in2[199];
    assign G[55] = in[198] & in2[198];
    assign P[55] = in[198] ^ in2[198];
    assign G[56] = in[197] & in2[197];
    assign P[56] = in[197] ^ in2[197];
    assign G[57] = in[196] & in2[196];
    assign P[57] = in[196] ^ in2[196];
    assign G[58] = in[195] & in2[195];
    assign P[58] = in[195] ^ in2[195];
    assign G[59] = in[194] & in2[194];
    assign P[59] = in[194] ^ in2[194];
    assign G[60] = in[193] & in2[193];
    assign P[60] = in[193] ^ in2[193];
    assign G[61] = in[192] & in2[192];
    assign P[61] = in[192] ^ in2[192];
    assign G[62] = in[191] & in2[191];
    assign P[62] = in[191] ^ in2[191];
    assign G[63] = in[190] & in2[190];
    assign P[63] = in[190] ^ in2[190];
    assign G[64] = in[189] & in2[189];
    assign P[64] = in[189] ^ in2[189];
    assign G[65] = in[188] & in2[188];
    assign P[65] = in[188] ^ in2[188];
    assign G[66] = in[187] & in2[187];
    assign P[66] = in[187] ^ in2[187];
    assign G[67] = in[186] & in2[186];
    assign P[67] = in[186] ^ in2[186];
    assign G[68] = in[185] & in2[185];
    assign P[68] = in[185] ^ in2[185];
    assign G[69] = in[184] & in2[184];
    assign P[69] = in[184] ^ in2[184];
    assign G[70] = in[183] & in2[183];
    assign P[70] = in[183] ^ in2[183];
    assign G[71] = in[182] & in2[182];
    assign P[71] = in[182] ^ in2[182];
    assign G[72] = in[181] & in2[181];
    assign P[72] = in[181] ^ in2[181];
    assign G[73] = in[180] & in2[180];
    assign P[73] = in[180] ^ in2[180];
    assign G[74] = in[179] & in2[179];
    assign P[74] = in[179] ^ in2[179];
    assign G[75] = in[178] & in2[178];
    assign P[75] = in[178] ^ in2[178];
    assign G[76] = in[177] & in2[177];
    assign P[76] = in[177] ^ in2[177];
    assign G[77] = in[176] & in2[176];
    assign P[77] = in[176] ^ in2[176];
    assign G[78] = in[175] & in2[175];
    assign P[78] = in[175] ^ in2[175];
    assign G[79] = in[174] & in2[174];
    assign P[79] = in[174] ^ in2[174];
    assign G[80] = in[173] & in2[173];
    assign P[80] = in[173] ^ in2[173];
    assign G[81] = in[172] & in2[172];
    assign P[81] = in[172] ^ in2[172];
    assign G[82] = in[171] & in2[171];
    assign P[82] = in[171] ^ in2[171];
    assign G[83] = in[170] & in2[170];
    assign P[83] = in[170] ^ in2[170];
    assign G[84] = in[169] & in2[169];
    assign P[84] = in[169] ^ in2[169];
    assign G[85] = in[168] & in2[168];
    assign P[85] = in[168] ^ in2[168];
    assign G[86] = in[167] & in2[167];
    assign P[86] = in[167] ^ in2[167];
    assign G[87] = in[166] & in2[166];
    assign P[87] = in[166] ^ in2[166];
    assign G[88] = in[165] & in2[165];
    assign P[88] = in[165] ^ in2[165];
    assign G[89] = in[164] & in2[164];
    assign P[89] = in[164] ^ in2[164];
    assign G[90] = in[163] & in2[163];
    assign P[90] = in[163] ^ in2[163];
    assign G[91] = in[162] & in2[162];
    assign P[91] = in[162] ^ in2[162];
    assign G[92] = in[161] & in2[161];
    assign P[92] = in[161] ^ in2[161];
    assign G[93] = in[160] & in2[160];
    assign P[93] = in[160] ^ in2[160];
    assign G[94] = in[159] & in2[159];
    assign P[94] = in[159] ^ in2[159];
    assign G[95] = in[158] & in2[158];
    assign P[95] = in[158] ^ in2[158];
    assign G[96] = in[157] & in2[157];
    assign P[96] = in[157] ^ in2[157];
    assign G[97] = in[156] & in2[156];
    assign P[97] = in[156] ^ in2[156];
    assign G[98] = in[155] & in2[155];
    assign P[98] = in[155] ^ in2[155];
    assign G[99] = in[154] & in2[154];
    assign P[99] = in[154] ^ in2[154];
    assign G[100] = in[153] & in2[153];
    assign P[100] = in[153] ^ in2[153];
    assign G[101] = in[152] & in2[152];
    assign P[101] = in[152] ^ in2[152];
    assign G[102] = in[151] & in2[151];
    assign P[102] = in[151] ^ in2[151];
    assign G[103] = in[150] & in2[150];
    assign P[103] = in[150] ^ in2[150];
    assign G[104] = in[149] & in2[149];
    assign P[104] = in[149] ^ in2[149];
    assign G[105] = in[148] & in2[148];
    assign P[105] = in[148] ^ in2[148];
    assign G[106] = in[147] & in2[147];
    assign P[106] = in[147] ^ in2[147];
    assign G[107] = in[146] & in2[146];
    assign P[107] = in[146] ^ in2[146];
    assign G[108] = in[145] & in2[145];
    assign P[108] = in[145] ^ in2[145];
    assign G[109] = in[144] & in2[144];
    assign P[109] = in[144] ^ in2[144];
    assign G[110] = in[143] & in2[143];
    assign P[110] = in[143] ^ in2[143];
    assign G[111] = in[142] & in2[142];
    assign P[111] = in[142] ^ in2[142];
    assign G[112] = in[141] & in2[141];
    assign P[112] = in[141] ^ in2[141];
    assign G[113] = in[140] & in2[140];
    assign P[113] = in[140] ^ in2[140];
    assign G[114] = in[139] & in2[139];
    assign P[114] = in[139] ^ in2[139];
    assign G[115] = in[138] & in2[138];
    assign P[115] = in[138] ^ in2[138];
    assign G[116] = in[137] & in2[137];
    assign P[116] = in[137] ^ in2[137];
    assign G[117] = in[136] & in2[136];
    assign P[117] = in[136] ^ in2[136];
    assign G[118] = in[135] & in2[135];
    assign P[118] = in[135] ^ in2[135];
    assign G[119] = in[134] & in2[134];
    assign P[119] = in[134] ^ in2[134];
    assign G[120] = in[133] & in2[133];
    assign P[120] = in[133] ^ in2[133];
    assign G[121] = in[132] & in2[132];
    assign P[121] = in[132] ^ in2[132];
    assign G[122] = in[131] & in2[131];
    assign P[122] = in[131] ^ in2[131];
    assign G[123] = in[130] & in2[130];
    assign P[123] = in[130] ^ in2[130];
    assign G[124] = in[129] & in2[129];
    assign P[124] = in[129] ^ in2[129];
    assign G[125] = in[128] & in2[128];
    assign P[125] = in[128] ^ in2[128];
    assign G[126] = in[127] & in2[127];
    assign P[126] = in[127] ^ in2[127];
    assign G[127] = in[126] & in2[126];
    assign P[127] = in[126] ^ in2[126];
    assign G[128] = in[125] & in2[125];
    assign P[128] = in[125] ^ in2[125];
    assign G[129] = in[124] & in2[124];
    assign P[129] = in[124] ^ in2[124];
    assign G[130] = in[123] & in2[123];
    assign P[130] = in[123] ^ in2[123];
    assign G[131] = in[122] & in2[122];
    assign P[131] = in[122] ^ in2[122];
    assign G[132] = in[121] & in2[121];
    assign P[132] = in[121] ^ in2[121];
    assign G[133] = in[120] & in2[120];
    assign P[133] = in[120] ^ in2[120];
    assign G[134] = in[119] & in2[119];
    assign P[134] = in[119] ^ in2[119];
    assign G[135] = in[118] & in2[118];
    assign P[135] = in[118] ^ in2[118];
    assign G[136] = in[117] & in2[117];
    assign P[136] = in[117] ^ in2[117];
    assign G[137] = in[116] & in2[116];
    assign P[137] = in[116] ^ in2[116];
    assign G[138] = in[115] & in2[115];
    assign P[138] = in[115] ^ in2[115];
    assign G[139] = in[114] & in2[114];
    assign P[139] = in[114] ^ in2[114];
    assign G[140] = in[113] & in2[113];
    assign P[140] = in[113] ^ in2[113];
    assign G[141] = in[112] & in2[112];
    assign P[141] = in[112] ^ in2[112];
    assign G[142] = in[111] & in2[111];
    assign P[142] = in[111] ^ in2[111];
    assign G[143] = in[110] & in2[110];
    assign P[143] = in[110] ^ in2[110];
    assign G[144] = in[109] & in2[109];
    assign P[144] = in[109] ^ in2[109];
    assign G[145] = in[108] & in2[108];
    assign P[145] = in[108] ^ in2[108];
    assign G[146] = in[107] & in2[107];
    assign P[146] = in[107] ^ in2[107];
    assign G[147] = in[106] & in2[106];
    assign P[147] = in[106] ^ in2[106];
    assign G[148] = in[105] & in2[105];
    assign P[148] = in[105] ^ in2[105];
    assign G[149] = in[104] & in2[104];
    assign P[149] = in[104] ^ in2[104];
    assign G[150] = in[103] & in2[103];
    assign P[150] = in[103] ^ in2[103];
    assign G[151] = in[102] & in2[102];
    assign P[151] = in[102] ^ in2[102];
    assign G[152] = in[101] & in2[101];
    assign P[152] = in[101] ^ in2[101];
    assign G[153] = in[100] & in2[100];
    assign P[153] = in[100] ^ in2[100];
    assign G[154] = in[99] & in2[99];
    assign P[154] = in[99] ^ in2[99];
    assign G[155] = in[98] & in2[98];
    assign P[155] = in[98] ^ in2[98];
    assign G[156] = in[97] & in2[97];
    assign P[156] = in[97] ^ in2[97];
    assign G[157] = in[96] & in2[96];
    assign P[157] = in[96] ^ in2[96];
    assign G[158] = in[95] & in2[95];
    assign P[158] = in[95] ^ in2[95];
    assign G[159] = in[94] & in2[94];
    assign P[159] = in[94] ^ in2[94];
    assign G[160] = in[93] & in2[93];
    assign P[160] = in[93] ^ in2[93];
    assign G[161] = in[92] & in2[92];
    assign P[161] = in[92] ^ in2[92];
    assign G[162] = in[91] & in2[91];
    assign P[162] = in[91] ^ in2[91];
    assign G[163] = in[90] & in2[90];
    assign P[163] = in[90] ^ in2[90];
    assign G[164] = in[89] & in2[89];
    assign P[164] = in[89] ^ in2[89];
    assign G[165] = in[88] & in2[88];
    assign P[165] = in[88] ^ in2[88];
    assign G[166] = in[87] & in2[87];
    assign P[166] = in[87] ^ in2[87];
    assign G[167] = in[86] & in2[86];
    assign P[167] = in[86] ^ in2[86];
    assign G[168] = in[85] & in2[85];
    assign P[168] = in[85] ^ in2[85];
    assign G[169] = in[84] & in2[84];
    assign P[169] = in[84] ^ in2[84];
    assign G[170] = in[83] & in2[83];
    assign P[170] = in[83] ^ in2[83];
    assign G[171] = in[82] & in2[82];
    assign P[171] = in[82] ^ in2[82];
    assign G[172] = in[81] & in2[81];
    assign P[172] = in[81] ^ in2[81];
    assign G[173] = in[80] & in2[80];
    assign P[173] = in[80] ^ in2[80];
    assign G[174] = in[79] & in2[79];
    assign P[174] = in[79] ^ in2[79];
    assign G[175] = in[78] & in2[78];
    assign P[175] = in[78] ^ in2[78];
    assign G[176] = in[77] & in2[77];
    assign P[176] = in[77] ^ in2[77];
    assign G[177] = in[76] & in2[76];
    assign P[177] = in[76] ^ in2[76];
    assign G[178] = in[75] & in2[75];
    assign P[178] = in[75] ^ in2[75];
    assign G[179] = in[74] & in2[74];
    assign P[179] = in[74] ^ in2[74];
    assign G[180] = in[73] & in2[73];
    assign P[180] = in[73] ^ in2[73];
    assign G[181] = in[72] & in2[72];
    assign P[181] = in[72] ^ in2[72];
    assign G[182] = in[71] & in2[71];
    assign P[182] = in[71] ^ in2[71];
    assign G[183] = in[70] & in2[70];
    assign P[183] = in[70] ^ in2[70];
    assign G[184] = in[69] & in2[69];
    assign P[184] = in[69] ^ in2[69];
    assign G[185] = in[68] & in2[68];
    assign P[185] = in[68] ^ in2[68];
    assign G[186] = in[67] & in2[67];
    assign P[186] = in[67] ^ in2[67];
    assign G[187] = in[66] & in2[66];
    assign P[187] = in[66] ^ in2[66];
    assign G[188] = in[65] & in2[65];
    assign P[188] = in[65] ^ in2[65];
    assign G[189] = in[64] & in2[64];
    assign P[189] = in[64] ^ in2[64];
    assign G[190] = in[63] & in2[63];
    assign P[190] = in[63] ^ in2[63];
    assign G[191] = in[62] & in2[62];
    assign P[191] = in[62] ^ in2[62];
    assign G[192] = in[61] & in2[61];
    assign P[192] = in[61] ^ in2[61];
    assign G[193] = in[60] & in2[60];
    assign P[193] = in[60] ^ in2[60];
    assign G[194] = in[59] & in2[59];
    assign P[194] = in[59] ^ in2[59];
    assign G[195] = in[58] & in2[58];
    assign P[195] = in[58] ^ in2[58];
    assign G[196] = in[57] & in2[57];
    assign P[196] = in[57] ^ in2[57];
    assign G[197] = in[56] & in2[56];
    assign P[197] = in[56] ^ in2[56];
    assign G[198] = in[55] & in2[55];
    assign P[198] = in[55] ^ in2[55];
    assign G[199] = in[54] & in2[54];
    assign P[199] = in[54] ^ in2[54];
    assign G[200] = in[53] & in2[53];
    assign P[200] = in[53] ^ in2[53];
    assign G[201] = in[52] & in2[52];
    assign P[201] = in[52] ^ in2[52];
    assign G[202] = in[51] & in2[51];
    assign P[202] = in[51] ^ in2[51];
    assign G[203] = in[50] & in2[50];
    assign P[203] = in[50] ^ in2[50];
    assign G[204] = in[49] & in2[49];
    assign P[204] = in[49] ^ in2[49];
    assign G[205] = in[48] & in2[48];
    assign P[205] = in[48] ^ in2[48];
    assign G[206] = in[47] & in2[47];
    assign P[206] = in[47] ^ in2[47];
    assign G[207] = in[46] & in2[46];
    assign P[207] = in[46] ^ in2[46];
    assign G[208] = in[45] & in2[45];
    assign P[208] = in[45] ^ in2[45];
    assign G[209] = in[44] & in2[44];
    assign P[209] = in[44] ^ in2[44];
    assign G[210] = in[43] & in2[43];
    assign P[210] = in[43] ^ in2[43];
    assign G[211] = in[42] & in2[42];
    assign P[211] = in[42] ^ in2[42];
    assign G[212] = in[41] & in2[41];
    assign P[212] = in[41] ^ in2[41];
    assign G[213] = in[40] & in2[40];
    assign P[213] = in[40] ^ in2[40];
    assign G[214] = in[39] & in2[39];
    assign P[214] = in[39] ^ in2[39];
    assign G[215] = in[38] & in2[38];
    assign P[215] = in[38] ^ in2[38];
    assign G[216] = in[37] & in2[37];
    assign P[216] = in[37] ^ in2[37];
    assign G[217] = in[36] & in2[36];
    assign P[217] = in[36] ^ in2[36];
    assign G[218] = in[35] & in2[35];
    assign P[218] = in[35] ^ in2[35];
    assign G[219] = in[34] & in2[34];
    assign P[219] = in[34] ^ in2[34];
    assign G[220] = in[33] & in2[33];
    assign P[220] = in[33] ^ in2[33];
    assign G[221] = in[32] & in2[32];
    assign P[221] = in[32] ^ in2[32];
    assign G[222] = in[31] & in2[31];
    assign P[222] = in[31] ^ in2[31];
    assign G[223] = in[30] & in2[30];
    assign P[223] = in[30] ^ in2[30];
    assign G[224] = in[29] & in2[29];
    assign P[224] = in[29] ^ in2[29];
    assign G[225] = in[28] & in2[28];
    assign P[225] = in[28] ^ in2[28];
    assign G[226] = in[27] & in2[27];
    assign P[226] = in[27] ^ in2[27];
    assign G[227] = in[26] & in2[26];
    assign P[227] = in[26] ^ in2[26];
    assign G[228] = in[25] & in2[25];
    assign P[228] = in[25] ^ in2[25];
    assign G[229] = in[24] & in2[24];
    assign P[229] = in[24] ^ in2[24];
    assign G[230] = in[23] & in2[23];
    assign P[230] = in[23] ^ in2[23];
    assign G[231] = in[22] & in2[22];
    assign P[231] = in[22] ^ in2[22];
    assign G[232] = in[21] & in2[21];
    assign P[232] = in[21] ^ in2[21];
    assign G[233] = in[20] & in2[20];
    assign P[233] = in[20] ^ in2[20];
    assign G[234] = in[19] & in2[19];
    assign P[234] = in[19] ^ in2[19];
    assign G[235] = in[18] & in2[18];
    assign P[235] = in[18] ^ in2[18];
    assign G[236] = in[17] & in2[17];
    assign P[236] = in[17] ^ in2[17];
    assign G[237] = in[16] & in2[16];
    assign P[237] = in[16] ^ in2[16];
    assign G[238] = in[15] & in2[15];
    assign P[238] = in[15] ^ in2[15];
    assign G[239] = in[14] & in2[14];
    assign P[239] = in[14] ^ in2[14];
    assign G[240] = in[13] & in2[13];
    assign P[240] = in[13] ^ in2[13];
    assign G[241] = in[12] & in2[12];
    assign P[241] = in[12] ^ in2[12];
    assign G[242] = in[11] & in2[11];
    assign P[242] = in[11] ^ in2[11];
    assign G[243] = in[10] & in2[10];
    assign P[243] = in[10] ^ in2[10];
    assign G[244] = in[9] & in2[9];
    assign P[244] = in[9] ^ in2[9];
    assign G[245] = in[8] & in2[8];
    assign P[245] = in[8] ^ in2[8];
    assign G[246] = in[7] & in2[7];
    assign P[246] = in[7] ^ in2[7];
    assign G[247] = in[6] & in2[6];
    assign P[247] = in[6] ^ in2[6];
    assign G[248] = in[5] & in2[5];
    assign P[248] = in[5] ^ in2[5];
    assign G[249] = in[4] & in2[4];
    assign P[249] = in[4] ^ in2[4];
    assign G[250] = in[3] & in2[3];
    assign P[250] = in[3] ^ in2[3];
    assign G[251] = in[2] & in2[2];
    assign P[251] = in[2] ^ in2[2];
    assign G[252] = in[1] & in2[1];
    assign P[252] = in[1] ^ in2[1];
    assign G[253] = in[0] & in2[0];
    assign P[253] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign C[252] = G[251] | (P[251] & C[251]);
    assign C[253] = G[252] | (P[252] & C[252]);
    assign cout = G[253] | (P[253] & C[253]);
    assign sum = P ^ C;
endmodule

module CLA253(output [252:0] sum, output cout, input [252:0] in1, input [252:0] in2;

    wire[252:0] G;
    wire[252:0] C;
    wire[252:0] P;

    assign G[0] = in[252] & in2[252];
    assign P[0] = in[252] ^ in2[252];
    assign G[1] = in[251] & in2[251];
    assign P[1] = in[251] ^ in2[251];
    assign G[2] = in[250] & in2[250];
    assign P[2] = in[250] ^ in2[250];
    assign G[3] = in[249] & in2[249];
    assign P[3] = in[249] ^ in2[249];
    assign G[4] = in[248] & in2[248];
    assign P[4] = in[248] ^ in2[248];
    assign G[5] = in[247] & in2[247];
    assign P[5] = in[247] ^ in2[247];
    assign G[6] = in[246] & in2[246];
    assign P[6] = in[246] ^ in2[246];
    assign G[7] = in[245] & in2[245];
    assign P[7] = in[245] ^ in2[245];
    assign G[8] = in[244] & in2[244];
    assign P[8] = in[244] ^ in2[244];
    assign G[9] = in[243] & in2[243];
    assign P[9] = in[243] ^ in2[243];
    assign G[10] = in[242] & in2[242];
    assign P[10] = in[242] ^ in2[242];
    assign G[11] = in[241] & in2[241];
    assign P[11] = in[241] ^ in2[241];
    assign G[12] = in[240] & in2[240];
    assign P[12] = in[240] ^ in2[240];
    assign G[13] = in[239] & in2[239];
    assign P[13] = in[239] ^ in2[239];
    assign G[14] = in[238] & in2[238];
    assign P[14] = in[238] ^ in2[238];
    assign G[15] = in[237] & in2[237];
    assign P[15] = in[237] ^ in2[237];
    assign G[16] = in[236] & in2[236];
    assign P[16] = in[236] ^ in2[236];
    assign G[17] = in[235] & in2[235];
    assign P[17] = in[235] ^ in2[235];
    assign G[18] = in[234] & in2[234];
    assign P[18] = in[234] ^ in2[234];
    assign G[19] = in[233] & in2[233];
    assign P[19] = in[233] ^ in2[233];
    assign G[20] = in[232] & in2[232];
    assign P[20] = in[232] ^ in2[232];
    assign G[21] = in[231] & in2[231];
    assign P[21] = in[231] ^ in2[231];
    assign G[22] = in[230] & in2[230];
    assign P[22] = in[230] ^ in2[230];
    assign G[23] = in[229] & in2[229];
    assign P[23] = in[229] ^ in2[229];
    assign G[24] = in[228] & in2[228];
    assign P[24] = in[228] ^ in2[228];
    assign G[25] = in[227] & in2[227];
    assign P[25] = in[227] ^ in2[227];
    assign G[26] = in[226] & in2[226];
    assign P[26] = in[226] ^ in2[226];
    assign G[27] = in[225] & in2[225];
    assign P[27] = in[225] ^ in2[225];
    assign G[28] = in[224] & in2[224];
    assign P[28] = in[224] ^ in2[224];
    assign G[29] = in[223] & in2[223];
    assign P[29] = in[223] ^ in2[223];
    assign G[30] = in[222] & in2[222];
    assign P[30] = in[222] ^ in2[222];
    assign G[31] = in[221] & in2[221];
    assign P[31] = in[221] ^ in2[221];
    assign G[32] = in[220] & in2[220];
    assign P[32] = in[220] ^ in2[220];
    assign G[33] = in[219] & in2[219];
    assign P[33] = in[219] ^ in2[219];
    assign G[34] = in[218] & in2[218];
    assign P[34] = in[218] ^ in2[218];
    assign G[35] = in[217] & in2[217];
    assign P[35] = in[217] ^ in2[217];
    assign G[36] = in[216] & in2[216];
    assign P[36] = in[216] ^ in2[216];
    assign G[37] = in[215] & in2[215];
    assign P[37] = in[215] ^ in2[215];
    assign G[38] = in[214] & in2[214];
    assign P[38] = in[214] ^ in2[214];
    assign G[39] = in[213] & in2[213];
    assign P[39] = in[213] ^ in2[213];
    assign G[40] = in[212] & in2[212];
    assign P[40] = in[212] ^ in2[212];
    assign G[41] = in[211] & in2[211];
    assign P[41] = in[211] ^ in2[211];
    assign G[42] = in[210] & in2[210];
    assign P[42] = in[210] ^ in2[210];
    assign G[43] = in[209] & in2[209];
    assign P[43] = in[209] ^ in2[209];
    assign G[44] = in[208] & in2[208];
    assign P[44] = in[208] ^ in2[208];
    assign G[45] = in[207] & in2[207];
    assign P[45] = in[207] ^ in2[207];
    assign G[46] = in[206] & in2[206];
    assign P[46] = in[206] ^ in2[206];
    assign G[47] = in[205] & in2[205];
    assign P[47] = in[205] ^ in2[205];
    assign G[48] = in[204] & in2[204];
    assign P[48] = in[204] ^ in2[204];
    assign G[49] = in[203] & in2[203];
    assign P[49] = in[203] ^ in2[203];
    assign G[50] = in[202] & in2[202];
    assign P[50] = in[202] ^ in2[202];
    assign G[51] = in[201] & in2[201];
    assign P[51] = in[201] ^ in2[201];
    assign G[52] = in[200] & in2[200];
    assign P[52] = in[200] ^ in2[200];
    assign G[53] = in[199] & in2[199];
    assign P[53] = in[199] ^ in2[199];
    assign G[54] = in[198] & in2[198];
    assign P[54] = in[198] ^ in2[198];
    assign G[55] = in[197] & in2[197];
    assign P[55] = in[197] ^ in2[197];
    assign G[56] = in[196] & in2[196];
    assign P[56] = in[196] ^ in2[196];
    assign G[57] = in[195] & in2[195];
    assign P[57] = in[195] ^ in2[195];
    assign G[58] = in[194] & in2[194];
    assign P[58] = in[194] ^ in2[194];
    assign G[59] = in[193] & in2[193];
    assign P[59] = in[193] ^ in2[193];
    assign G[60] = in[192] & in2[192];
    assign P[60] = in[192] ^ in2[192];
    assign G[61] = in[191] & in2[191];
    assign P[61] = in[191] ^ in2[191];
    assign G[62] = in[190] & in2[190];
    assign P[62] = in[190] ^ in2[190];
    assign G[63] = in[189] & in2[189];
    assign P[63] = in[189] ^ in2[189];
    assign G[64] = in[188] & in2[188];
    assign P[64] = in[188] ^ in2[188];
    assign G[65] = in[187] & in2[187];
    assign P[65] = in[187] ^ in2[187];
    assign G[66] = in[186] & in2[186];
    assign P[66] = in[186] ^ in2[186];
    assign G[67] = in[185] & in2[185];
    assign P[67] = in[185] ^ in2[185];
    assign G[68] = in[184] & in2[184];
    assign P[68] = in[184] ^ in2[184];
    assign G[69] = in[183] & in2[183];
    assign P[69] = in[183] ^ in2[183];
    assign G[70] = in[182] & in2[182];
    assign P[70] = in[182] ^ in2[182];
    assign G[71] = in[181] & in2[181];
    assign P[71] = in[181] ^ in2[181];
    assign G[72] = in[180] & in2[180];
    assign P[72] = in[180] ^ in2[180];
    assign G[73] = in[179] & in2[179];
    assign P[73] = in[179] ^ in2[179];
    assign G[74] = in[178] & in2[178];
    assign P[74] = in[178] ^ in2[178];
    assign G[75] = in[177] & in2[177];
    assign P[75] = in[177] ^ in2[177];
    assign G[76] = in[176] & in2[176];
    assign P[76] = in[176] ^ in2[176];
    assign G[77] = in[175] & in2[175];
    assign P[77] = in[175] ^ in2[175];
    assign G[78] = in[174] & in2[174];
    assign P[78] = in[174] ^ in2[174];
    assign G[79] = in[173] & in2[173];
    assign P[79] = in[173] ^ in2[173];
    assign G[80] = in[172] & in2[172];
    assign P[80] = in[172] ^ in2[172];
    assign G[81] = in[171] & in2[171];
    assign P[81] = in[171] ^ in2[171];
    assign G[82] = in[170] & in2[170];
    assign P[82] = in[170] ^ in2[170];
    assign G[83] = in[169] & in2[169];
    assign P[83] = in[169] ^ in2[169];
    assign G[84] = in[168] & in2[168];
    assign P[84] = in[168] ^ in2[168];
    assign G[85] = in[167] & in2[167];
    assign P[85] = in[167] ^ in2[167];
    assign G[86] = in[166] & in2[166];
    assign P[86] = in[166] ^ in2[166];
    assign G[87] = in[165] & in2[165];
    assign P[87] = in[165] ^ in2[165];
    assign G[88] = in[164] & in2[164];
    assign P[88] = in[164] ^ in2[164];
    assign G[89] = in[163] & in2[163];
    assign P[89] = in[163] ^ in2[163];
    assign G[90] = in[162] & in2[162];
    assign P[90] = in[162] ^ in2[162];
    assign G[91] = in[161] & in2[161];
    assign P[91] = in[161] ^ in2[161];
    assign G[92] = in[160] & in2[160];
    assign P[92] = in[160] ^ in2[160];
    assign G[93] = in[159] & in2[159];
    assign P[93] = in[159] ^ in2[159];
    assign G[94] = in[158] & in2[158];
    assign P[94] = in[158] ^ in2[158];
    assign G[95] = in[157] & in2[157];
    assign P[95] = in[157] ^ in2[157];
    assign G[96] = in[156] & in2[156];
    assign P[96] = in[156] ^ in2[156];
    assign G[97] = in[155] & in2[155];
    assign P[97] = in[155] ^ in2[155];
    assign G[98] = in[154] & in2[154];
    assign P[98] = in[154] ^ in2[154];
    assign G[99] = in[153] & in2[153];
    assign P[99] = in[153] ^ in2[153];
    assign G[100] = in[152] & in2[152];
    assign P[100] = in[152] ^ in2[152];
    assign G[101] = in[151] & in2[151];
    assign P[101] = in[151] ^ in2[151];
    assign G[102] = in[150] & in2[150];
    assign P[102] = in[150] ^ in2[150];
    assign G[103] = in[149] & in2[149];
    assign P[103] = in[149] ^ in2[149];
    assign G[104] = in[148] & in2[148];
    assign P[104] = in[148] ^ in2[148];
    assign G[105] = in[147] & in2[147];
    assign P[105] = in[147] ^ in2[147];
    assign G[106] = in[146] & in2[146];
    assign P[106] = in[146] ^ in2[146];
    assign G[107] = in[145] & in2[145];
    assign P[107] = in[145] ^ in2[145];
    assign G[108] = in[144] & in2[144];
    assign P[108] = in[144] ^ in2[144];
    assign G[109] = in[143] & in2[143];
    assign P[109] = in[143] ^ in2[143];
    assign G[110] = in[142] & in2[142];
    assign P[110] = in[142] ^ in2[142];
    assign G[111] = in[141] & in2[141];
    assign P[111] = in[141] ^ in2[141];
    assign G[112] = in[140] & in2[140];
    assign P[112] = in[140] ^ in2[140];
    assign G[113] = in[139] & in2[139];
    assign P[113] = in[139] ^ in2[139];
    assign G[114] = in[138] & in2[138];
    assign P[114] = in[138] ^ in2[138];
    assign G[115] = in[137] & in2[137];
    assign P[115] = in[137] ^ in2[137];
    assign G[116] = in[136] & in2[136];
    assign P[116] = in[136] ^ in2[136];
    assign G[117] = in[135] & in2[135];
    assign P[117] = in[135] ^ in2[135];
    assign G[118] = in[134] & in2[134];
    assign P[118] = in[134] ^ in2[134];
    assign G[119] = in[133] & in2[133];
    assign P[119] = in[133] ^ in2[133];
    assign G[120] = in[132] & in2[132];
    assign P[120] = in[132] ^ in2[132];
    assign G[121] = in[131] & in2[131];
    assign P[121] = in[131] ^ in2[131];
    assign G[122] = in[130] & in2[130];
    assign P[122] = in[130] ^ in2[130];
    assign G[123] = in[129] & in2[129];
    assign P[123] = in[129] ^ in2[129];
    assign G[124] = in[128] & in2[128];
    assign P[124] = in[128] ^ in2[128];
    assign G[125] = in[127] & in2[127];
    assign P[125] = in[127] ^ in2[127];
    assign G[126] = in[126] & in2[126];
    assign P[126] = in[126] ^ in2[126];
    assign G[127] = in[125] & in2[125];
    assign P[127] = in[125] ^ in2[125];
    assign G[128] = in[124] & in2[124];
    assign P[128] = in[124] ^ in2[124];
    assign G[129] = in[123] & in2[123];
    assign P[129] = in[123] ^ in2[123];
    assign G[130] = in[122] & in2[122];
    assign P[130] = in[122] ^ in2[122];
    assign G[131] = in[121] & in2[121];
    assign P[131] = in[121] ^ in2[121];
    assign G[132] = in[120] & in2[120];
    assign P[132] = in[120] ^ in2[120];
    assign G[133] = in[119] & in2[119];
    assign P[133] = in[119] ^ in2[119];
    assign G[134] = in[118] & in2[118];
    assign P[134] = in[118] ^ in2[118];
    assign G[135] = in[117] & in2[117];
    assign P[135] = in[117] ^ in2[117];
    assign G[136] = in[116] & in2[116];
    assign P[136] = in[116] ^ in2[116];
    assign G[137] = in[115] & in2[115];
    assign P[137] = in[115] ^ in2[115];
    assign G[138] = in[114] & in2[114];
    assign P[138] = in[114] ^ in2[114];
    assign G[139] = in[113] & in2[113];
    assign P[139] = in[113] ^ in2[113];
    assign G[140] = in[112] & in2[112];
    assign P[140] = in[112] ^ in2[112];
    assign G[141] = in[111] & in2[111];
    assign P[141] = in[111] ^ in2[111];
    assign G[142] = in[110] & in2[110];
    assign P[142] = in[110] ^ in2[110];
    assign G[143] = in[109] & in2[109];
    assign P[143] = in[109] ^ in2[109];
    assign G[144] = in[108] & in2[108];
    assign P[144] = in[108] ^ in2[108];
    assign G[145] = in[107] & in2[107];
    assign P[145] = in[107] ^ in2[107];
    assign G[146] = in[106] & in2[106];
    assign P[146] = in[106] ^ in2[106];
    assign G[147] = in[105] & in2[105];
    assign P[147] = in[105] ^ in2[105];
    assign G[148] = in[104] & in2[104];
    assign P[148] = in[104] ^ in2[104];
    assign G[149] = in[103] & in2[103];
    assign P[149] = in[103] ^ in2[103];
    assign G[150] = in[102] & in2[102];
    assign P[150] = in[102] ^ in2[102];
    assign G[151] = in[101] & in2[101];
    assign P[151] = in[101] ^ in2[101];
    assign G[152] = in[100] & in2[100];
    assign P[152] = in[100] ^ in2[100];
    assign G[153] = in[99] & in2[99];
    assign P[153] = in[99] ^ in2[99];
    assign G[154] = in[98] & in2[98];
    assign P[154] = in[98] ^ in2[98];
    assign G[155] = in[97] & in2[97];
    assign P[155] = in[97] ^ in2[97];
    assign G[156] = in[96] & in2[96];
    assign P[156] = in[96] ^ in2[96];
    assign G[157] = in[95] & in2[95];
    assign P[157] = in[95] ^ in2[95];
    assign G[158] = in[94] & in2[94];
    assign P[158] = in[94] ^ in2[94];
    assign G[159] = in[93] & in2[93];
    assign P[159] = in[93] ^ in2[93];
    assign G[160] = in[92] & in2[92];
    assign P[160] = in[92] ^ in2[92];
    assign G[161] = in[91] & in2[91];
    assign P[161] = in[91] ^ in2[91];
    assign G[162] = in[90] & in2[90];
    assign P[162] = in[90] ^ in2[90];
    assign G[163] = in[89] & in2[89];
    assign P[163] = in[89] ^ in2[89];
    assign G[164] = in[88] & in2[88];
    assign P[164] = in[88] ^ in2[88];
    assign G[165] = in[87] & in2[87];
    assign P[165] = in[87] ^ in2[87];
    assign G[166] = in[86] & in2[86];
    assign P[166] = in[86] ^ in2[86];
    assign G[167] = in[85] & in2[85];
    assign P[167] = in[85] ^ in2[85];
    assign G[168] = in[84] & in2[84];
    assign P[168] = in[84] ^ in2[84];
    assign G[169] = in[83] & in2[83];
    assign P[169] = in[83] ^ in2[83];
    assign G[170] = in[82] & in2[82];
    assign P[170] = in[82] ^ in2[82];
    assign G[171] = in[81] & in2[81];
    assign P[171] = in[81] ^ in2[81];
    assign G[172] = in[80] & in2[80];
    assign P[172] = in[80] ^ in2[80];
    assign G[173] = in[79] & in2[79];
    assign P[173] = in[79] ^ in2[79];
    assign G[174] = in[78] & in2[78];
    assign P[174] = in[78] ^ in2[78];
    assign G[175] = in[77] & in2[77];
    assign P[175] = in[77] ^ in2[77];
    assign G[176] = in[76] & in2[76];
    assign P[176] = in[76] ^ in2[76];
    assign G[177] = in[75] & in2[75];
    assign P[177] = in[75] ^ in2[75];
    assign G[178] = in[74] & in2[74];
    assign P[178] = in[74] ^ in2[74];
    assign G[179] = in[73] & in2[73];
    assign P[179] = in[73] ^ in2[73];
    assign G[180] = in[72] & in2[72];
    assign P[180] = in[72] ^ in2[72];
    assign G[181] = in[71] & in2[71];
    assign P[181] = in[71] ^ in2[71];
    assign G[182] = in[70] & in2[70];
    assign P[182] = in[70] ^ in2[70];
    assign G[183] = in[69] & in2[69];
    assign P[183] = in[69] ^ in2[69];
    assign G[184] = in[68] & in2[68];
    assign P[184] = in[68] ^ in2[68];
    assign G[185] = in[67] & in2[67];
    assign P[185] = in[67] ^ in2[67];
    assign G[186] = in[66] & in2[66];
    assign P[186] = in[66] ^ in2[66];
    assign G[187] = in[65] & in2[65];
    assign P[187] = in[65] ^ in2[65];
    assign G[188] = in[64] & in2[64];
    assign P[188] = in[64] ^ in2[64];
    assign G[189] = in[63] & in2[63];
    assign P[189] = in[63] ^ in2[63];
    assign G[190] = in[62] & in2[62];
    assign P[190] = in[62] ^ in2[62];
    assign G[191] = in[61] & in2[61];
    assign P[191] = in[61] ^ in2[61];
    assign G[192] = in[60] & in2[60];
    assign P[192] = in[60] ^ in2[60];
    assign G[193] = in[59] & in2[59];
    assign P[193] = in[59] ^ in2[59];
    assign G[194] = in[58] & in2[58];
    assign P[194] = in[58] ^ in2[58];
    assign G[195] = in[57] & in2[57];
    assign P[195] = in[57] ^ in2[57];
    assign G[196] = in[56] & in2[56];
    assign P[196] = in[56] ^ in2[56];
    assign G[197] = in[55] & in2[55];
    assign P[197] = in[55] ^ in2[55];
    assign G[198] = in[54] & in2[54];
    assign P[198] = in[54] ^ in2[54];
    assign G[199] = in[53] & in2[53];
    assign P[199] = in[53] ^ in2[53];
    assign G[200] = in[52] & in2[52];
    assign P[200] = in[52] ^ in2[52];
    assign G[201] = in[51] & in2[51];
    assign P[201] = in[51] ^ in2[51];
    assign G[202] = in[50] & in2[50];
    assign P[202] = in[50] ^ in2[50];
    assign G[203] = in[49] & in2[49];
    assign P[203] = in[49] ^ in2[49];
    assign G[204] = in[48] & in2[48];
    assign P[204] = in[48] ^ in2[48];
    assign G[205] = in[47] & in2[47];
    assign P[205] = in[47] ^ in2[47];
    assign G[206] = in[46] & in2[46];
    assign P[206] = in[46] ^ in2[46];
    assign G[207] = in[45] & in2[45];
    assign P[207] = in[45] ^ in2[45];
    assign G[208] = in[44] & in2[44];
    assign P[208] = in[44] ^ in2[44];
    assign G[209] = in[43] & in2[43];
    assign P[209] = in[43] ^ in2[43];
    assign G[210] = in[42] & in2[42];
    assign P[210] = in[42] ^ in2[42];
    assign G[211] = in[41] & in2[41];
    assign P[211] = in[41] ^ in2[41];
    assign G[212] = in[40] & in2[40];
    assign P[212] = in[40] ^ in2[40];
    assign G[213] = in[39] & in2[39];
    assign P[213] = in[39] ^ in2[39];
    assign G[214] = in[38] & in2[38];
    assign P[214] = in[38] ^ in2[38];
    assign G[215] = in[37] & in2[37];
    assign P[215] = in[37] ^ in2[37];
    assign G[216] = in[36] & in2[36];
    assign P[216] = in[36] ^ in2[36];
    assign G[217] = in[35] & in2[35];
    assign P[217] = in[35] ^ in2[35];
    assign G[218] = in[34] & in2[34];
    assign P[218] = in[34] ^ in2[34];
    assign G[219] = in[33] & in2[33];
    assign P[219] = in[33] ^ in2[33];
    assign G[220] = in[32] & in2[32];
    assign P[220] = in[32] ^ in2[32];
    assign G[221] = in[31] & in2[31];
    assign P[221] = in[31] ^ in2[31];
    assign G[222] = in[30] & in2[30];
    assign P[222] = in[30] ^ in2[30];
    assign G[223] = in[29] & in2[29];
    assign P[223] = in[29] ^ in2[29];
    assign G[224] = in[28] & in2[28];
    assign P[224] = in[28] ^ in2[28];
    assign G[225] = in[27] & in2[27];
    assign P[225] = in[27] ^ in2[27];
    assign G[226] = in[26] & in2[26];
    assign P[226] = in[26] ^ in2[26];
    assign G[227] = in[25] & in2[25];
    assign P[227] = in[25] ^ in2[25];
    assign G[228] = in[24] & in2[24];
    assign P[228] = in[24] ^ in2[24];
    assign G[229] = in[23] & in2[23];
    assign P[229] = in[23] ^ in2[23];
    assign G[230] = in[22] & in2[22];
    assign P[230] = in[22] ^ in2[22];
    assign G[231] = in[21] & in2[21];
    assign P[231] = in[21] ^ in2[21];
    assign G[232] = in[20] & in2[20];
    assign P[232] = in[20] ^ in2[20];
    assign G[233] = in[19] & in2[19];
    assign P[233] = in[19] ^ in2[19];
    assign G[234] = in[18] & in2[18];
    assign P[234] = in[18] ^ in2[18];
    assign G[235] = in[17] & in2[17];
    assign P[235] = in[17] ^ in2[17];
    assign G[236] = in[16] & in2[16];
    assign P[236] = in[16] ^ in2[16];
    assign G[237] = in[15] & in2[15];
    assign P[237] = in[15] ^ in2[15];
    assign G[238] = in[14] & in2[14];
    assign P[238] = in[14] ^ in2[14];
    assign G[239] = in[13] & in2[13];
    assign P[239] = in[13] ^ in2[13];
    assign G[240] = in[12] & in2[12];
    assign P[240] = in[12] ^ in2[12];
    assign G[241] = in[11] & in2[11];
    assign P[241] = in[11] ^ in2[11];
    assign G[242] = in[10] & in2[10];
    assign P[242] = in[10] ^ in2[10];
    assign G[243] = in[9] & in2[9];
    assign P[243] = in[9] ^ in2[9];
    assign G[244] = in[8] & in2[8];
    assign P[244] = in[8] ^ in2[8];
    assign G[245] = in[7] & in2[7];
    assign P[245] = in[7] ^ in2[7];
    assign G[246] = in[6] & in2[6];
    assign P[246] = in[6] ^ in2[6];
    assign G[247] = in[5] & in2[5];
    assign P[247] = in[5] ^ in2[5];
    assign G[248] = in[4] & in2[4];
    assign P[248] = in[4] ^ in2[4];
    assign G[249] = in[3] & in2[3];
    assign P[249] = in[3] ^ in2[3];
    assign G[250] = in[2] & in2[2];
    assign P[250] = in[2] ^ in2[2];
    assign G[251] = in[1] & in2[1];
    assign P[251] = in[1] ^ in2[1];
    assign G[252] = in[0] & in2[0];
    assign P[252] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign C[252] = G[251] | (P[251] & C[251]);
    assign cout = G[252] | (P[252] & C[252]);
    assign sum = P ^ C;
endmodule

module CLA252(output [251:0] sum, output cout, input [251:0] in1, input [251:0] in2;

    wire[251:0] G;
    wire[251:0] C;
    wire[251:0] P;

    assign G[0] = in[251] & in2[251];
    assign P[0] = in[251] ^ in2[251];
    assign G[1] = in[250] & in2[250];
    assign P[1] = in[250] ^ in2[250];
    assign G[2] = in[249] & in2[249];
    assign P[2] = in[249] ^ in2[249];
    assign G[3] = in[248] & in2[248];
    assign P[3] = in[248] ^ in2[248];
    assign G[4] = in[247] & in2[247];
    assign P[4] = in[247] ^ in2[247];
    assign G[5] = in[246] & in2[246];
    assign P[5] = in[246] ^ in2[246];
    assign G[6] = in[245] & in2[245];
    assign P[6] = in[245] ^ in2[245];
    assign G[7] = in[244] & in2[244];
    assign P[7] = in[244] ^ in2[244];
    assign G[8] = in[243] & in2[243];
    assign P[8] = in[243] ^ in2[243];
    assign G[9] = in[242] & in2[242];
    assign P[9] = in[242] ^ in2[242];
    assign G[10] = in[241] & in2[241];
    assign P[10] = in[241] ^ in2[241];
    assign G[11] = in[240] & in2[240];
    assign P[11] = in[240] ^ in2[240];
    assign G[12] = in[239] & in2[239];
    assign P[12] = in[239] ^ in2[239];
    assign G[13] = in[238] & in2[238];
    assign P[13] = in[238] ^ in2[238];
    assign G[14] = in[237] & in2[237];
    assign P[14] = in[237] ^ in2[237];
    assign G[15] = in[236] & in2[236];
    assign P[15] = in[236] ^ in2[236];
    assign G[16] = in[235] & in2[235];
    assign P[16] = in[235] ^ in2[235];
    assign G[17] = in[234] & in2[234];
    assign P[17] = in[234] ^ in2[234];
    assign G[18] = in[233] & in2[233];
    assign P[18] = in[233] ^ in2[233];
    assign G[19] = in[232] & in2[232];
    assign P[19] = in[232] ^ in2[232];
    assign G[20] = in[231] & in2[231];
    assign P[20] = in[231] ^ in2[231];
    assign G[21] = in[230] & in2[230];
    assign P[21] = in[230] ^ in2[230];
    assign G[22] = in[229] & in2[229];
    assign P[22] = in[229] ^ in2[229];
    assign G[23] = in[228] & in2[228];
    assign P[23] = in[228] ^ in2[228];
    assign G[24] = in[227] & in2[227];
    assign P[24] = in[227] ^ in2[227];
    assign G[25] = in[226] & in2[226];
    assign P[25] = in[226] ^ in2[226];
    assign G[26] = in[225] & in2[225];
    assign P[26] = in[225] ^ in2[225];
    assign G[27] = in[224] & in2[224];
    assign P[27] = in[224] ^ in2[224];
    assign G[28] = in[223] & in2[223];
    assign P[28] = in[223] ^ in2[223];
    assign G[29] = in[222] & in2[222];
    assign P[29] = in[222] ^ in2[222];
    assign G[30] = in[221] & in2[221];
    assign P[30] = in[221] ^ in2[221];
    assign G[31] = in[220] & in2[220];
    assign P[31] = in[220] ^ in2[220];
    assign G[32] = in[219] & in2[219];
    assign P[32] = in[219] ^ in2[219];
    assign G[33] = in[218] & in2[218];
    assign P[33] = in[218] ^ in2[218];
    assign G[34] = in[217] & in2[217];
    assign P[34] = in[217] ^ in2[217];
    assign G[35] = in[216] & in2[216];
    assign P[35] = in[216] ^ in2[216];
    assign G[36] = in[215] & in2[215];
    assign P[36] = in[215] ^ in2[215];
    assign G[37] = in[214] & in2[214];
    assign P[37] = in[214] ^ in2[214];
    assign G[38] = in[213] & in2[213];
    assign P[38] = in[213] ^ in2[213];
    assign G[39] = in[212] & in2[212];
    assign P[39] = in[212] ^ in2[212];
    assign G[40] = in[211] & in2[211];
    assign P[40] = in[211] ^ in2[211];
    assign G[41] = in[210] & in2[210];
    assign P[41] = in[210] ^ in2[210];
    assign G[42] = in[209] & in2[209];
    assign P[42] = in[209] ^ in2[209];
    assign G[43] = in[208] & in2[208];
    assign P[43] = in[208] ^ in2[208];
    assign G[44] = in[207] & in2[207];
    assign P[44] = in[207] ^ in2[207];
    assign G[45] = in[206] & in2[206];
    assign P[45] = in[206] ^ in2[206];
    assign G[46] = in[205] & in2[205];
    assign P[46] = in[205] ^ in2[205];
    assign G[47] = in[204] & in2[204];
    assign P[47] = in[204] ^ in2[204];
    assign G[48] = in[203] & in2[203];
    assign P[48] = in[203] ^ in2[203];
    assign G[49] = in[202] & in2[202];
    assign P[49] = in[202] ^ in2[202];
    assign G[50] = in[201] & in2[201];
    assign P[50] = in[201] ^ in2[201];
    assign G[51] = in[200] & in2[200];
    assign P[51] = in[200] ^ in2[200];
    assign G[52] = in[199] & in2[199];
    assign P[52] = in[199] ^ in2[199];
    assign G[53] = in[198] & in2[198];
    assign P[53] = in[198] ^ in2[198];
    assign G[54] = in[197] & in2[197];
    assign P[54] = in[197] ^ in2[197];
    assign G[55] = in[196] & in2[196];
    assign P[55] = in[196] ^ in2[196];
    assign G[56] = in[195] & in2[195];
    assign P[56] = in[195] ^ in2[195];
    assign G[57] = in[194] & in2[194];
    assign P[57] = in[194] ^ in2[194];
    assign G[58] = in[193] & in2[193];
    assign P[58] = in[193] ^ in2[193];
    assign G[59] = in[192] & in2[192];
    assign P[59] = in[192] ^ in2[192];
    assign G[60] = in[191] & in2[191];
    assign P[60] = in[191] ^ in2[191];
    assign G[61] = in[190] & in2[190];
    assign P[61] = in[190] ^ in2[190];
    assign G[62] = in[189] & in2[189];
    assign P[62] = in[189] ^ in2[189];
    assign G[63] = in[188] & in2[188];
    assign P[63] = in[188] ^ in2[188];
    assign G[64] = in[187] & in2[187];
    assign P[64] = in[187] ^ in2[187];
    assign G[65] = in[186] & in2[186];
    assign P[65] = in[186] ^ in2[186];
    assign G[66] = in[185] & in2[185];
    assign P[66] = in[185] ^ in2[185];
    assign G[67] = in[184] & in2[184];
    assign P[67] = in[184] ^ in2[184];
    assign G[68] = in[183] & in2[183];
    assign P[68] = in[183] ^ in2[183];
    assign G[69] = in[182] & in2[182];
    assign P[69] = in[182] ^ in2[182];
    assign G[70] = in[181] & in2[181];
    assign P[70] = in[181] ^ in2[181];
    assign G[71] = in[180] & in2[180];
    assign P[71] = in[180] ^ in2[180];
    assign G[72] = in[179] & in2[179];
    assign P[72] = in[179] ^ in2[179];
    assign G[73] = in[178] & in2[178];
    assign P[73] = in[178] ^ in2[178];
    assign G[74] = in[177] & in2[177];
    assign P[74] = in[177] ^ in2[177];
    assign G[75] = in[176] & in2[176];
    assign P[75] = in[176] ^ in2[176];
    assign G[76] = in[175] & in2[175];
    assign P[76] = in[175] ^ in2[175];
    assign G[77] = in[174] & in2[174];
    assign P[77] = in[174] ^ in2[174];
    assign G[78] = in[173] & in2[173];
    assign P[78] = in[173] ^ in2[173];
    assign G[79] = in[172] & in2[172];
    assign P[79] = in[172] ^ in2[172];
    assign G[80] = in[171] & in2[171];
    assign P[80] = in[171] ^ in2[171];
    assign G[81] = in[170] & in2[170];
    assign P[81] = in[170] ^ in2[170];
    assign G[82] = in[169] & in2[169];
    assign P[82] = in[169] ^ in2[169];
    assign G[83] = in[168] & in2[168];
    assign P[83] = in[168] ^ in2[168];
    assign G[84] = in[167] & in2[167];
    assign P[84] = in[167] ^ in2[167];
    assign G[85] = in[166] & in2[166];
    assign P[85] = in[166] ^ in2[166];
    assign G[86] = in[165] & in2[165];
    assign P[86] = in[165] ^ in2[165];
    assign G[87] = in[164] & in2[164];
    assign P[87] = in[164] ^ in2[164];
    assign G[88] = in[163] & in2[163];
    assign P[88] = in[163] ^ in2[163];
    assign G[89] = in[162] & in2[162];
    assign P[89] = in[162] ^ in2[162];
    assign G[90] = in[161] & in2[161];
    assign P[90] = in[161] ^ in2[161];
    assign G[91] = in[160] & in2[160];
    assign P[91] = in[160] ^ in2[160];
    assign G[92] = in[159] & in2[159];
    assign P[92] = in[159] ^ in2[159];
    assign G[93] = in[158] & in2[158];
    assign P[93] = in[158] ^ in2[158];
    assign G[94] = in[157] & in2[157];
    assign P[94] = in[157] ^ in2[157];
    assign G[95] = in[156] & in2[156];
    assign P[95] = in[156] ^ in2[156];
    assign G[96] = in[155] & in2[155];
    assign P[96] = in[155] ^ in2[155];
    assign G[97] = in[154] & in2[154];
    assign P[97] = in[154] ^ in2[154];
    assign G[98] = in[153] & in2[153];
    assign P[98] = in[153] ^ in2[153];
    assign G[99] = in[152] & in2[152];
    assign P[99] = in[152] ^ in2[152];
    assign G[100] = in[151] & in2[151];
    assign P[100] = in[151] ^ in2[151];
    assign G[101] = in[150] & in2[150];
    assign P[101] = in[150] ^ in2[150];
    assign G[102] = in[149] & in2[149];
    assign P[102] = in[149] ^ in2[149];
    assign G[103] = in[148] & in2[148];
    assign P[103] = in[148] ^ in2[148];
    assign G[104] = in[147] & in2[147];
    assign P[104] = in[147] ^ in2[147];
    assign G[105] = in[146] & in2[146];
    assign P[105] = in[146] ^ in2[146];
    assign G[106] = in[145] & in2[145];
    assign P[106] = in[145] ^ in2[145];
    assign G[107] = in[144] & in2[144];
    assign P[107] = in[144] ^ in2[144];
    assign G[108] = in[143] & in2[143];
    assign P[108] = in[143] ^ in2[143];
    assign G[109] = in[142] & in2[142];
    assign P[109] = in[142] ^ in2[142];
    assign G[110] = in[141] & in2[141];
    assign P[110] = in[141] ^ in2[141];
    assign G[111] = in[140] & in2[140];
    assign P[111] = in[140] ^ in2[140];
    assign G[112] = in[139] & in2[139];
    assign P[112] = in[139] ^ in2[139];
    assign G[113] = in[138] & in2[138];
    assign P[113] = in[138] ^ in2[138];
    assign G[114] = in[137] & in2[137];
    assign P[114] = in[137] ^ in2[137];
    assign G[115] = in[136] & in2[136];
    assign P[115] = in[136] ^ in2[136];
    assign G[116] = in[135] & in2[135];
    assign P[116] = in[135] ^ in2[135];
    assign G[117] = in[134] & in2[134];
    assign P[117] = in[134] ^ in2[134];
    assign G[118] = in[133] & in2[133];
    assign P[118] = in[133] ^ in2[133];
    assign G[119] = in[132] & in2[132];
    assign P[119] = in[132] ^ in2[132];
    assign G[120] = in[131] & in2[131];
    assign P[120] = in[131] ^ in2[131];
    assign G[121] = in[130] & in2[130];
    assign P[121] = in[130] ^ in2[130];
    assign G[122] = in[129] & in2[129];
    assign P[122] = in[129] ^ in2[129];
    assign G[123] = in[128] & in2[128];
    assign P[123] = in[128] ^ in2[128];
    assign G[124] = in[127] & in2[127];
    assign P[124] = in[127] ^ in2[127];
    assign G[125] = in[126] & in2[126];
    assign P[125] = in[126] ^ in2[126];
    assign G[126] = in[125] & in2[125];
    assign P[126] = in[125] ^ in2[125];
    assign G[127] = in[124] & in2[124];
    assign P[127] = in[124] ^ in2[124];
    assign G[128] = in[123] & in2[123];
    assign P[128] = in[123] ^ in2[123];
    assign G[129] = in[122] & in2[122];
    assign P[129] = in[122] ^ in2[122];
    assign G[130] = in[121] & in2[121];
    assign P[130] = in[121] ^ in2[121];
    assign G[131] = in[120] & in2[120];
    assign P[131] = in[120] ^ in2[120];
    assign G[132] = in[119] & in2[119];
    assign P[132] = in[119] ^ in2[119];
    assign G[133] = in[118] & in2[118];
    assign P[133] = in[118] ^ in2[118];
    assign G[134] = in[117] & in2[117];
    assign P[134] = in[117] ^ in2[117];
    assign G[135] = in[116] & in2[116];
    assign P[135] = in[116] ^ in2[116];
    assign G[136] = in[115] & in2[115];
    assign P[136] = in[115] ^ in2[115];
    assign G[137] = in[114] & in2[114];
    assign P[137] = in[114] ^ in2[114];
    assign G[138] = in[113] & in2[113];
    assign P[138] = in[113] ^ in2[113];
    assign G[139] = in[112] & in2[112];
    assign P[139] = in[112] ^ in2[112];
    assign G[140] = in[111] & in2[111];
    assign P[140] = in[111] ^ in2[111];
    assign G[141] = in[110] & in2[110];
    assign P[141] = in[110] ^ in2[110];
    assign G[142] = in[109] & in2[109];
    assign P[142] = in[109] ^ in2[109];
    assign G[143] = in[108] & in2[108];
    assign P[143] = in[108] ^ in2[108];
    assign G[144] = in[107] & in2[107];
    assign P[144] = in[107] ^ in2[107];
    assign G[145] = in[106] & in2[106];
    assign P[145] = in[106] ^ in2[106];
    assign G[146] = in[105] & in2[105];
    assign P[146] = in[105] ^ in2[105];
    assign G[147] = in[104] & in2[104];
    assign P[147] = in[104] ^ in2[104];
    assign G[148] = in[103] & in2[103];
    assign P[148] = in[103] ^ in2[103];
    assign G[149] = in[102] & in2[102];
    assign P[149] = in[102] ^ in2[102];
    assign G[150] = in[101] & in2[101];
    assign P[150] = in[101] ^ in2[101];
    assign G[151] = in[100] & in2[100];
    assign P[151] = in[100] ^ in2[100];
    assign G[152] = in[99] & in2[99];
    assign P[152] = in[99] ^ in2[99];
    assign G[153] = in[98] & in2[98];
    assign P[153] = in[98] ^ in2[98];
    assign G[154] = in[97] & in2[97];
    assign P[154] = in[97] ^ in2[97];
    assign G[155] = in[96] & in2[96];
    assign P[155] = in[96] ^ in2[96];
    assign G[156] = in[95] & in2[95];
    assign P[156] = in[95] ^ in2[95];
    assign G[157] = in[94] & in2[94];
    assign P[157] = in[94] ^ in2[94];
    assign G[158] = in[93] & in2[93];
    assign P[158] = in[93] ^ in2[93];
    assign G[159] = in[92] & in2[92];
    assign P[159] = in[92] ^ in2[92];
    assign G[160] = in[91] & in2[91];
    assign P[160] = in[91] ^ in2[91];
    assign G[161] = in[90] & in2[90];
    assign P[161] = in[90] ^ in2[90];
    assign G[162] = in[89] & in2[89];
    assign P[162] = in[89] ^ in2[89];
    assign G[163] = in[88] & in2[88];
    assign P[163] = in[88] ^ in2[88];
    assign G[164] = in[87] & in2[87];
    assign P[164] = in[87] ^ in2[87];
    assign G[165] = in[86] & in2[86];
    assign P[165] = in[86] ^ in2[86];
    assign G[166] = in[85] & in2[85];
    assign P[166] = in[85] ^ in2[85];
    assign G[167] = in[84] & in2[84];
    assign P[167] = in[84] ^ in2[84];
    assign G[168] = in[83] & in2[83];
    assign P[168] = in[83] ^ in2[83];
    assign G[169] = in[82] & in2[82];
    assign P[169] = in[82] ^ in2[82];
    assign G[170] = in[81] & in2[81];
    assign P[170] = in[81] ^ in2[81];
    assign G[171] = in[80] & in2[80];
    assign P[171] = in[80] ^ in2[80];
    assign G[172] = in[79] & in2[79];
    assign P[172] = in[79] ^ in2[79];
    assign G[173] = in[78] & in2[78];
    assign P[173] = in[78] ^ in2[78];
    assign G[174] = in[77] & in2[77];
    assign P[174] = in[77] ^ in2[77];
    assign G[175] = in[76] & in2[76];
    assign P[175] = in[76] ^ in2[76];
    assign G[176] = in[75] & in2[75];
    assign P[176] = in[75] ^ in2[75];
    assign G[177] = in[74] & in2[74];
    assign P[177] = in[74] ^ in2[74];
    assign G[178] = in[73] & in2[73];
    assign P[178] = in[73] ^ in2[73];
    assign G[179] = in[72] & in2[72];
    assign P[179] = in[72] ^ in2[72];
    assign G[180] = in[71] & in2[71];
    assign P[180] = in[71] ^ in2[71];
    assign G[181] = in[70] & in2[70];
    assign P[181] = in[70] ^ in2[70];
    assign G[182] = in[69] & in2[69];
    assign P[182] = in[69] ^ in2[69];
    assign G[183] = in[68] & in2[68];
    assign P[183] = in[68] ^ in2[68];
    assign G[184] = in[67] & in2[67];
    assign P[184] = in[67] ^ in2[67];
    assign G[185] = in[66] & in2[66];
    assign P[185] = in[66] ^ in2[66];
    assign G[186] = in[65] & in2[65];
    assign P[186] = in[65] ^ in2[65];
    assign G[187] = in[64] & in2[64];
    assign P[187] = in[64] ^ in2[64];
    assign G[188] = in[63] & in2[63];
    assign P[188] = in[63] ^ in2[63];
    assign G[189] = in[62] & in2[62];
    assign P[189] = in[62] ^ in2[62];
    assign G[190] = in[61] & in2[61];
    assign P[190] = in[61] ^ in2[61];
    assign G[191] = in[60] & in2[60];
    assign P[191] = in[60] ^ in2[60];
    assign G[192] = in[59] & in2[59];
    assign P[192] = in[59] ^ in2[59];
    assign G[193] = in[58] & in2[58];
    assign P[193] = in[58] ^ in2[58];
    assign G[194] = in[57] & in2[57];
    assign P[194] = in[57] ^ in2[57];
    assign G[195] = in[56] & in2[56];
    assign P[195] = in[56] ^ in2[56];
    assign G[196] = in[55] & in2[55];
    assign P[196] = in[55] ^ in2[55];
    assign G[197] = in[54] & in2[54];
    assign P[197] = in[54] ^ in2[54];
    assign G[198] = in[53] & in2[53];
    assign P[198] = in[53] ^ in2[53];
    assign G[199] = in[52] & in2[52];
    assign P[199] = in[52] ^ in2[52];
    assign G[200] = in[51] & in2[51];
    assign P[200] = in[51] ^ in2[51];
    assign G[201] = in[50] & in2[50];
    assign P[201] = in[50] ^ in2[50];
    assign G[202] = in[49] & in2[49];
    assign P[202] = in[49] ^ in2[49];
    assign G[203] = in[48] & in2[48];
    assign P[203] = in[48] ^ in2[48];
    assign G[204] = in[47] & in2[47];
    assign P[204] = in[47] ^ in2[47];
    assign G[205] = in[46] & in2[46];
    assign P[205] = in[46] ^ in2[46];
    assign G[206] = in[45] & in2[45];
    assign P[206] = in[45] ^ in2[45];
    assign G[207] = in[44] & in2[44];
    assign P[207] = in[44] ^ in2[44];
    assign G[208] = in[43] & in2[43];
    assign P[208] = in[43] ^ in2[43];
    assign G[209] = in[42] & in2[42];
    assign P[209] = in[42] ^ in2[42];
    assign G[210] = in[41] & in2[41];
    assign P[210] = in[41] ^ in2[41];
    assign G[211] = in[40] & in2[40];
    assign P[211] = in[40] ^ in2[40];
    assign G[212] = in[39] & in2[39];
    assign P[212] = in[39] ^ in2[39];
    assign G[213] = in[38] & in2[38];
    assign P[213] = in[38] ^ in2[38];
    assign G[214] = in[37] & in2[37];
    assign P[214] = in[37] ^ in2[37];
    assign G[215] = in[36] & in2[36];
    assign P[215] = in[36] ^ in2[36];
    assign G[216] = in[35] & in2[35];
    assign P[216] = in[35] ^ in2[35];
    assign G[217] = in[34] & in2[34];
    assign P[217] = in[34] ^ in2[34];
    assign G[218] = in[33] & in2[33];
    assign P[218] = in[33] ^ in2[33];
    assign G[219] = in[32] & in2[32];
    assign P[219] = in[32] ^ in2[32];
    assign G[220] = in[31] & in2[31];
    assign P[220] = in[31] ^ in2[31];
    assign G[221] = in[30] & in2[30];
    assign P[221] = in[30] ^ in2[30];
    assign G[222] = in[29] & in2[29];
    assign P[222] = in[29] ^ in2[29];
    assign G[223] = in[28] & in2[28];
    assign P[223] = in[28] ^ in2[28];
    assign G[224] = in[27] & in2[27];
    assign P[224] = in[27] ^ in2[27];
    assign G[225] = in[26] & in2[26];
    assign P[225] = in[26] ^ in2[26];
    assign G[226] = in[25] & in2[25];
    assign P[226] = in[25] ^ in2[25];
    assign G[227] = in[24] & in2[24];
    assign P[227] = in[24] ^ in2[24];
    assign G[228] = in[23] & in2[23];
    assign P[228] = in[23] ^ in2[23];
    assign G[229] = in[22] & in2[22];
    assign P[229] = in[22] ^ in2[22];
    assign G[230] = in[21] & in2[21];
    assign P[230] = in[21] ^ in2[21];
    assign G[231] = in[20] & in2[20];
    assign P[231] = in[20] ^ in2[20];
    assign G[232] = in[19] & in2[19];
    assign P[232] = in[19] ^ in2[19];
    assign G[233] = in[18] & in2[18];
    assign P[233] = in[18] ^ in2[18];
    assign G[234] = in[17] & in2[17];
    assign P[234] = in[17] ^ in2[17];
    assign G[235] = in[16] & in2[16];
    assign P[235] = in[16] ^ in2[16];
    assign G[236] = in[15] & in2[15];
    assign P[236] = in[15] ^ in2[15];
    assign G[237] = in[14] & in2[14];
    assign P[237] = in[14] ^ in2[14];
    assign G[238] = in[13] & in2[13];
    assign P[238] = in[13] ^ in2[13];
    assign G[239] = in[12] & in2[12];
    assign P[239] = in[12] ^ in2[12];
    assign G[240] = in[11] & in2[11];
    assign P[240] = in[11] ^ in2[11];
    assign G[241] = in[10] & in2[10];
    assign P[241] = in[10] ^ in2[10];
    assign G[242] = in[9] & in2[9];
    assign P[242] = in[9] ^ in2[9];
    assign G[243] = in[8] & in2[8];
    assign P[243] = in[8] ^ in2[8];
    assign G[244] = in[7] & in2[7];
    assign P[244] = in[7] ^ in2[7];
    assign G[245] = in[6] & in2[6];
    assign P[245] = in[6] ^ in2[6];
    assign G[246] = in[5] & in2[5];
    assign P[246] = in[5] ^ in2[5];
    assign G[247] = in[4] & in2[4];
    assign P[247] = in[4] ^ in2[4];
    assign G[248] = in[3] & in2[3];
    assign P[248] = in[3] ^ in2[3];
    assign G[249] = in[2] & in2[2];
    assign P[249] = in[2] ^ in2[2];
    assign G[250] = in[1] & in2[1];
    assign P[250] = in[1] ^ in2[1];
    assign G[251] = in[0] & in2[0];
    assign P[251] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign C[251] = G[250] | (P[250] & C[250]);
    assign cout = G[251] | (P[251] & C[251]);
    assign sum = P ^ C;
endmodule

module CLA251(output [250:0] sum, output cout, input [250:0] in1, input [250:0] in2;

    wire[250:0] G;
    wire[250:0] C;
    wire[250:0] P;

    assign G[0] = in[250] & in2[250];
    assign P[0] = in[250] ^ in2[250];
    assign G[1] = in[249] & in2[249];
    assign P[1] = in[249] ^ in2[249];
    assign G[2] = in[248] & in2[248];
    assign P[2] = in[248] ^ in2[248];
    assign G[3] = in[247] & in2[247];
    assign P[3] = in[247] ^ in2[247];
    assign G[4] = in[246] & in2[246];
    assign P[4] = in[246] ^ in2[246];
    assign G[5] = in[245] & in2[245];
    assign P[5] = in[245] ^ in2[245];
    assign G[6] = in[244] & in2[244];
    assign P[6] = in[244] ^ in2[244];
    assign G[7] = in[243] & in2[243];
    assign P[7] = in[243] ^ in2[243];
    assign G[8] = in[242] & in2[242];
    assign P[8] = in[242] ^ in2[242];
    assign G[9] = in[241] & in2[241];
    assign P[9] = in[241] ^ in2[241];
    assign G[10] = in[240] & in2[240];
    assign P[10] = in[240] ^ in2[240];
    assign G[11] = in[239] & in2[239];
    assign P[11] = in[239] ^ in2[239];
    assign G[12] = in[238] & in2[238];
    assign P[12] = in[238] ^ in2[238];
    assign G[13] = in[237] & in2[237];
    assign P[13] = in[237] ^ in2[237];
    assign G[14] = in[236] & in2[236];
    assign P[14] = in[236] ^ in2[236];
    assign G[15] = in[235] & in2[235];
    assign P[15] = in[235] ^ in2[235];
    assign G[16] = in[234] & in2[234];
    assign P[16] = in[234] ^ in2[234];
    assign G[17] = in[233] & in2[233];
    assign P[17] = in[233] ^ in2[233];
    assign G[18] = in[232] & in2[232];
    assign P[18] = in[232] ^ in2[232];
    assign G[19] = in[231] & in2[231];
    assign P[19] = in[231] ^ in2[231];
    assign G[20] = in[230] & in2[230];
    assign P[20] = in[230] ^ in2[230];
    assign G[21] = in[229] & in2[229];
    assign P[21] = in[229] ^ in2[229];
    assign G[22] = in[228] & in2[228];
    assign P[22] = in[228] ^ in2[228];
    assign G[23] = in[227] & in2[227];
    assign P[23] = in[227] ^ in2[227];
    assign G[24] = in[226] & in2[226];
    assign P[24] = in[226] ^ in2[226];
    assign G[25] = in[225] & in2[225];
    assign P[25] = in[225] ^ in2[225];
    assign G[26] = in[224] & in2[224];
    assign P[26] = in[224] ^ in2[224];
    assign G[27] = in[223] & in2[223];
    assign P[27] = in[223] ^ in2[223];
    assign G[28] = in[222] & in2[222];
    assign P[28] = in[222] ^ in2[222];
    assign G[29] = in[221] & in2[221];
    assign P[29] = in[221] ^ in2[221];
    assign G[30] = in[220] & in2[220];
    assign P[30] = in[220] ^ in2[220];
    assign G[31] = in[219] & in2[219];
    assign P[31] = in[219] ^ in2[219];
    assign G[32] = in[218] & in2[218];
    assign P[32] = in[218] ^ in2[218];
    assign G[33] = in[217] & in2[217];
    assign P[33] = in[217] ^ in2[217];
    assign G[34] = in[216] & in2[216];
    assign P[34] = in[216] ^ in2[216];
    assign G[35] = in[215] & in2[215];
    assign P[35] = in[215] ^ in2[215];
    assign G[36] = in[214] & in2[214];
    assign P[36] = in[214] ^ in2[214];
    assign G[37] = in[213] & in2[213];
    assign P[37] = in[213] ^ in2[213];
    assign G[38] = in[212] & in2[212];
    assign P[38] = in[212] ^ in2[212];
    assign G[39] = in[211] & in2[211];
    assign P[39] = in[211] ^ in2[211];
    assign G[40] = in[210] & in2[210];
    assign P[40] = in[210] ^ in2[210];
    assign G[41] = in[209] & in2[209];
    assign P[41] = in[209] ^ in2[209];
    assign G[42] = in[208] & in2[208];
    assign P[42] = in[208] ^ in2[208];
    assign G[43] = in[207] & in2[207];
    assign P[43] = in[207] ^ in2[207];
    assign G[44] = in[206] & in2[206];
    assign P[44] = in[206] ^ in2[206];
    assign G[45] = in[205] & in2[205];
    assign P[45] = in[205] ^ in2[205];
    assign G[46] = in[204] & in2[204];
    assign P[46] = in[204] ^ in2[204];
    assign G[47] = in[203] & in2[203];
    assign P[47] = in[203] ^ in2[203];
    assign G[48] = in[202] & in2[202];
    assign P[48] = in[202] ^ in2[202];
    assign G[49] = in[201] & in2[201];
    assign P[49] = in[201] ^ in2[201];
    assign G[50] = in[200] & in2[200];
    assign P[50] = in[200] ^ in2[200];
    assign G[51] = in[199] & in2[199];
    assign P[51] = in[199] ^ in2[199];
    assign G[52] = in[198] & in2[198];
    assign P[52] = in[198] ^ in2[198];
    assign G[53] = in[197] & in2[197];
    assign P[53] = in[197] ^ in2[197];
    assign G[54] = in[196] & in2[196];
    assign P[54] = in[196] ^ in2[196];
    assign G[55] = in[195] & in2[195];
    assign P[55] = in[195] ^ in2[195];
    assign G[56] = in[194] & in2[194];
    assign P[56] = in[194] ^ in2[194];
    assign G[57] = in[193] & in2[193];
    assign P[57] = in[193] ^ in2[193];
    assign G[58] = in[192] & in2[192];
    assign P[58] = in[192] ^ in2[192];
    assign G[59] = in[191] & in2[191];
    assign P[59] = in[191] ^ in2[191];
    assign G[60] = in[190] & in2[190];
    assign P[60] = in[190] ^ in2[190];
    assign G[61] = in[189] & in2[189];
    assign P[61] = in[189] ^ in2[189];
    assign G[62] = in[188] & in2[188];
    assign P[62] = in[188] ^ in2[188];
    assign G[63] = in[187] & in2[187];
    assign P[63] = in[187] ^ in2[187];
    assign G[64] = in[186] & in2[186];
    assign P[64] = in[186] ^ in2[186];
    assign G[65] = in[185] & in2[185];
    assign P[65] = in[185] ^ in2[185];
    assign G[66] = in[184] & in2[184];
    assign P[66] = in[184] ^ in2[184];
    assign G[67] = in[183] & in2[183];
    assign P[67] = in[183] ^ in2[183];
    assign G[68] = in[182] & in2[182];
    assign P[68] = in[182] ^ in2[182];
    assign G[69] = in[181] & in2[181];
    assign P[69] = in[181] ^ in2[181];
    assign G[70] = in[180] & in2[180];
    assign P[70] = in[180] ^ in2[180];
    assign G[71] = in[179] & in2[179];
    assign P[71] = in[179] ^ in2[179];
    assign G[72] = in[178] & in2[178];
    assign P[72] = in[178] ^ in2[178];
    assign G[73] = in[177] & in2[177];
    assign P[73] = in[177] ^ in2[177];
    assign G[74] = in[176] & in2[176];
    assign P[74] = in[176] ^ in2[176];
    assign G[75] = in[175] & in2[175];
    assign P[75] = in[175] ^ in2[175];
    assign G[76] = in[174] & in2[174];
    assign P[76] = in[174] ^ in2[174];
    assign G[77] = in[173] & in2[173];
    assign P[77] = in[173] ^ in2[173];
    assign G[78] = in[172] & in2[172];
    assign P[78] = in[172] ^ in2[172];
    assign G[79] = in[171] & in2[171];
    assign P[79] = in[171] ^ in2[171];
    assign G[80] = in[170] & in2[170];
    assign P[80] = in[170] ^ in2[170];
    assign G[81] = in[169] & in2[169];
    assign P[81] = in[169] ^ in2[169];
    assign G[82] = in[168] & in2[168];
    assign P[82] = in[168] ^ in2[168];
    assign G[83] = in[167] & in2[167];
    assign P[83] = in[167] ^ in2[167];
    assign G[84] = in[166] & in2[166];
    assign P[84] = in[166] ^ in2[166];
    assign G[85] = in[165] & in2[165];
    assign P[85] = in[165] ^ in2[165];
    assign G[86] = in[164] & in2[164];
    assign P[86] = in[164] ^ in2[164];
    assign G[87] = in[163] & in2[163];
    assign P[87] = in[163] ^ in2[163];
    assign G[88] = in[162] & in2[162];
    assign P[88] = in[162] ^ in2[162];
    assign G[89] = in[161] & in2[161];
    assign P[89] = in[161] ^ in2[161];
    assign G[90] = in[160] & in2[160];
    assign P[90] = in[160] ^ in2[160];
    assign G[91] = in[159] & in2[159];
    assign P[91] = in[159] ^ in2[159];
    assign G[92] = in[158] & in2[158];
    assign P[92] = in[158] ^ in2[158];
    assign G[93] = in[157] & in2[157];
    assign P[93] = in[157] ^ in2[157];
    assign G[94] = in[156] & in2[156];
    assign P[94] = in[156] ^ in2[156];
    assign G[95] = in[155] & in2[155];
    assign P[95] = in[155] ^ in2[155];
    assign G[96] = in[154] & in2[154];
    assign P[96] = in[154] ^ in2[154];
    assign G[97] = in[153] & in2[153];
    assign P[97] = in[153] ^ in2[153];
    assign G[98] = in[152] & in2[152];
    assign P[98] = in[152] ^ in2[152];
    assign G[99] = in[151] & in2[151];
    assign P[99] = in[151] ^ in2[151];
    assign G[100] = in[150] & in2[150];
    assign P[100] = in[150] ^ in2[150];
    assign G[101] = in[149] & in2[149];
    assign P[101] = in[149] ^ in2[149];
    assign G[102] = in[148] & in2[148];
    assign P[102] = in[148] ^ in2[148];
    assign G[103] = in[147] & in2[147];
    assign P[103] = in[147] ^ in2[147];
    assign G[104] = in[146] & in2[146];
    assign P[104] = in[146] ^ in2[146];
    assign G[105] = in[145] & in2[145];
    assign P[105] = in[145] ^ in2[145];
    assign G[106] = in[144] & in2[144];
    assign P[106] = in[144] ^ in2[144];
    assign G[107] = in[143] & in2[143];
    assign P[107] = in[143] ^ in2[143];
    assign G[108] = in[142] & in2[142];
    assign P[108] = in[142] ^ in2[142];
    assign G[109] = in[141] & in2[141];
    assign P[109] = in[141] ^ in2[141];
    assign G[110] = in[140] & in2[140];
    assign P[110] = in[140] ^ in2[140];
    assign G[111] = in[139] & in2[139];
    assign P[111] = in[139] ^ in2[139];
    assign G[112] = in[138] & in2[138];
    assign P[112] = in[138] ^ in2[138];
    assign G[113] = in[137] & in2[137];
    assign P[113] = in[137] ^ in2[137];
    assign G[114] = in[136] & in2[136];
    assign P[114] = in[136] ^ in2[136];
    assign G[115] = in[135] & in2[135];
    assign P[115] = in[135] ^ in2[135];
    assign G[116] = in[134] & in2[134];
    assign P[116] = in[134] ^ in2[134];
    assign G[117] = in[133] & in2[133];
    assign P[117] = in[133] ^ in2[133];
    assign G[118] = in[132] & in2[132];
    assign P[118] = in[132] ^ in2[132];
    assign G[119] = in[131] & in2[131];
    assign P[119] = in[131] ^ in2[131];
    assign G[120] = in[130] & in2[130];
    assign P[120] = in[130] ^ in2[130];
    assign G[121] = in[129] & in2[129];
    assign P[121] = in[129] ^ in2[129];
    assign G[122] = in[128] & in2[128];
    assign P[122] = in[128] ^ in2[128];
    assign G[123] = in[127] & in2[127];
    assign P[123] = in[127] ^ in2[127];
    assign G[124] = in[126] & in2[126];
    assign P[124] = in[126] ^ in2[126];
    assign G[125] = in[125] & in2[125];
    assign P[125] = in[125] ^ in2[125];
    assign G[126] = in[124] & in2[124];
    assign P[126] = in[124] ^ in2[124];
    assign G[127] = in[123] & in2[123];
    assign P[127] = in[123] ^ in2[123];
    assign G[128] = in[122] & in2[122];
    assign P[128] = in[122] ^ in2[122];
    assign G[129] = in[121] & in2[121];
    assign P[129] = in[121] ^ in2[121];
    assign G[130] = in[120] & in2[120];
    assign P[130] = in[120] ^ in2[120];
    assign G[131] = in[119] & in2[119];
    assign P[131] = in[119] ^ in2[119];
    assign G[132] = in[118] & in2[118];
    assign P[132] = in[118] ^ in2[118];
    assign G[133] = in[117] & in2[117];
    assign P[133] = in[117] ^ in2[117];
    assign G[134] = in[116] & in2[116];
    assign P[134] = in[116] ^ in2[116];
    assign G[135] = in[115] & in2[115];
    assign P[135] = in[115] ^ in2[115];
    assign G[136] = in[114] & in2[114];
    assign P[136] = in[114] ^ in2[114];
    assign G[137] = in[113] & in2[113];
    assign P[137] = in[113] ^ in2[113];
    assign G[138] = in[112] & in2[112];
    assign P[138] = in[112] ^ in2[112];
    assign G[139] = in[111] & in2[111];
    assign P[139] = in[111] ^ in2[111];
    assign G[140] = in[110] & in2[110];
    assign P[140] = in[110] ^ in2[110];
    assign G[141] = in[109] & in2[109];
    assign P[141] = in[109] ^ in2[109];
    assign G[142] = in[108] & in2[108];
    assign P[142] = in[108] ^ in2[108];
    assign G[143] = in[107] & in2[107];
    assign P[143] = in[107] ^ in2[107];
    assign G[144] = in[106] & in2[106];
    assign P[144] = in[106] ^ in2[106];
    assign G[145] = in[105] & in2[105];
    assign P[145] = in[105] ^ in2[105];
    assign G[146] = in[104] & in2[104];
    assign P[146] = in[104] ^ in2[104];
    assign G[147] = in[103] & in2[103];
    assign P[147] = in[103] ^ in2[103];
    assign G[148] = in[102] & in2[102];
    assign P[148] = in[102] ^ in2[102];
    assign G[149] = in[101] & in2[101];
    assign P[149] = in[101] ^ in2[101];
    assign G[150] = in[100] & in2[100];
    assign P[150] = in[100] ^ in2[100];
    assign G[151] = in[99] & in2[99];
    assign P[151] = in[99] ^ in2[99];
    assign G[152] = in[98] & in2[98];
    assign P[152] = in[98] ^ in2[98];
    assign G[153] = in[97] & in2[97];
    assign P[153] = in[97] ^ in2[97];
    assign G[154] = in[96] & in2[96];
    assign P[154] = in[96] ^ in2[96];
    assign G[155] = in[95] & in2[95];
    assign P[155] = in[95] ^ in2[95];
    assign G[156] = in[94] & in2[94];
    assign P[156] = in[94] ^ in2[94];
    assign G[157] = in[93] & in2[93];
    assign P[157] = in[93] ^ in2[93];
    assign G[158] = in[92] & in2[92];
    assign P[158] = in[92] ^ in2[92];
    assign G[159] = in[91] & in2[91];
    assign P[159] = in[91] ^ in2[91];
    assign G[160] = in[90] & in2[90];
    assign P[160] = in[90] ^ in2[90];
    assign G[161] = in[89] & in2[89];
    assign P[161] = in[89] ^ in2[89];
    assign G[162] = in[88] & in2[88];
    assign P[162] = in[88] ^ in2[88];
    assign G[163] = in[87] & in2[87];
    assign P[163] = in[87] ^ in2[87];
    assign G[164] = in[86] & in2[86];
    assign P[164] = in[86] ^ in2[86];
    assign G[165] = in[85] & in2[85];
    assign P[165] = in[85] ^ in2[85];
    assign G[166] = in[84] & in2[84];
    assign P[166] = in[84] ^ in2[84];
    assign G[167] = in[83] & in2[83];
    assign P[167] = in[83] ^ in2[83];
    assign G[168] = in[82] & in2[82];
    assign P[168] = in[82] ^ in2[82];
    assign G[169] = in[81] & in2[81];
    assign P[169] = in[81] ^ in2[81];
    assign G[170] = in[80] & in2[80];
    assign P[170] = in[80] ^ in2[80];
    assign G[171] = in[79] & in2[79];
    assign P[171] = in[79] ^ in2[79];
    assign G[172] = in[78] & in2[78];
    assign P[172] = in[78] ^ in2[78];
    assign G[173] = in[77] & in2[77];
    assign P[173] = in[77] ^ in2[77];
    assign G[174] = in[76] & in2[76];
    assign P[174] = in[76] ^ in2[76];
    assign G[175] = in[75] & in2[75];
    assign P[175] = in[75] ^ in2[75];
    assign G[176] = in[74] & in2[74];
    assign P[176] = in[74] ^ in2[74];
    assign G[177] = in[73] & in2[73];
    assign P[177] = in[73] ^ in2[73];
    assign G[178] = in[72] & in2[72];
    assign P[178] = in[72] ^ in2[72];
    assign G[179] = in[71] & in2[71];
    assign P[179] = in[71] ^ in2[71];
    assign G[180] = in[70] & in2[70];
    assign P[180] = in[70] ^ in2[70];
    assign G[181] = in[69] & in2[69];
    assign P[181] = in[69] ^ in2[69];
    assign G[182] = in[68] & in2[68];
    assign P[182] = in[68] ^ in2[68];
    assign G[183] = in[67] & in2[67];
    assign P[183] = in[67] ^ in2[67];
    assign G[184] = in[66] & in2[66];
    assign P[184] = in[66] ^ in2[66];
    assign G[185] = in[65] & in2[65];
    assign P[185] = in[65] ^ in2[65];
    assign G[186] = in[64] & in2[64];
    assign P[186] = in[64] ^ in2[64];
    assign G[187] = in[63] & in2[63];
    assign P[187] = in[63] ^ in2[63];
    assign G[188] = in[62] & in2[62];
    assign P[188] = in[62] ^ in2[62];
    assign G[189] = in[61] & in2[61];
    assign P[189] = in[61] ^ in2[61];
    assign G[190] = in[60] & in2[60];
    assign P[190] = in[60] ^ in2[60];
    assign G[191] = in[59] & in2[59];
    assign P[191] = in[59] ^ in2[59];
    assign G[192] = in[58] & in2[58];
    assign P[192] = in[58] ^ in2[58];
    assign G[193] = in[57] & in2[57];
    assign P[193] = in[57] ^ in2[57];
    assign G[194] = in[56] & in2[56];
    assign P[194] = in[56] ^ in2[56];
    assign G[195] = in[55] & in2[55];
    assign P[195] = in[55] ^ in2[55];
    assign G[196] = in[54] & in2[54];
    assign P[196] = in[54] ^ in2[54];
    assign G[197] = in[53] & in2[53];
    assign P[197] = in[53] ^ in2[53];
    assign G[198] = in[52] & in2[52];
    assign P[198] = in[52] ^ in2[52];
    assign G[199] = in[51] & in2[51];
    assign P[199] = in[51] ^ in2[51];
    assign G[200] = in[50] & in2[50];
    assign P[200] = in[50] ^ in2[50];
    assign G[201] = in[49] & in2[49];
    assign P[201] = in[49] ^ in2[49];
    assign G[202] = in[48] & in2[48];
    assign P[202] = in[48] ^ in2[48];
    assign G[203] = in[47] & in2[47];
    assign P[203] = in[47] ^ in2[47];
    assign G[204] = in[46] & in2[46];
    assign P[204] = in[46] ^ in2[46];
    assign G[205] = in[45] & in2[45];
    assign P[205] = in[45] ^ in2[45];
    assign G[206] = in[44] & in2[44];
    assign P[206] = in[44] ^ in2[44];
    assign G[207] = in[43] & in2[43];
    assign P[207] = in[43] ^ in2[43];
    assign G[208] = in[42] & in2[42];
    assign P[208] = in[42] ^ in2[42];
    assign G[209] = in[41] & in2[41];
    assign P[209] = in[41] ^ in2[41];
    assign G[210] = in[40] & in2[40];
    assign P[210] = in[40] ^ in2[40];
    assign G[211] = in[39] & in2[39];
    assign P[211] = in[39] ^ in2[39];
    assign G[212] = in[38] & in2[38];
    assign P[212] = in[38] ^ in2[38];
    assign G[213] = in[37] & in2[37];
    assign P[213] = in[37] ^ in2[37];
    assign G[214] = in[36] & in2[36];
    assign P[214] = in[36] ^ in2[36];
    assign G[215] = in[35] & in2[35];
    assign P[215] = in[35] ^ in2[35];
    assign G[216] = in[34] & in2[34];
    assign P[216] = in[34] ^ in2[34];
    assign G[217] = in[33] & in2[33];
    assign P[217] = in[33] ^ in2[33];
    assign G[218] = in[32] & in2[32];
    assign P[218] = in[32] ^ in2[32];
    assign G[219] = in[31] & in2[31];
    assign P[219] = in[31] ^ in2[31];
    assign G[220] = in[30] & in2[30];
    assign P[220] = in[30] ^ in2[30];
    assign G[221] = in[29] & in2[29];
    assign P[221] = in[29] ^ in2[29];
    assign G[222] = in[28] & in2[28];
    assign P[222] = in[28] ^ in2[28];
    assign G[223] = in[27] & in2[27];
    assign P[223] = in[27] ^ in2[27];
    assign G[224] = in[26] & in2[26];
    assign P[224] = in[26] ^ in2[26];
    assign G[225] = in[25] & in2[25];
    assign P[225] = in[25] ^ in2[25];
    assign G[226] = in[24] & in2[24];
    assign P[226] = in[24] ^ in2[24];
    assign G[227] = in[23] & in2[23];
    assign P[227] = in[23] ^ in2[23];
    assign G[228] = in[22] & in2[22];
    assign P[228] = in[22] ^ in2[22];
    assign G[229] = in[21] & in2[21];
    assign P[229] = in[21] ^ in2[21];
    assign G[230] = in[20] & in2[20];
    assign P[230] = in[20] ^ in2[20];
    assign G[231] = in[19] & in2[19];
    assign P[231] = in[19] ^ in2[19];
    assign G[232] = in[18] & in2[18];
    assign P[232] = in[18] ^ in2[18];
    assign G[233] = in[17] & in2[17];
    assign P[233] = in[17] ^ in2[17];
    assign G[234] = in[16] & in2[16];
    assign P[234] = in[16] ^ in2[16];
    assign G[235] = in[15] & in2[15];
    assign P[235] = in[15] ^ in2[15];
    assign G[236] = in[14] & in2[14];
    assign P[236] = in[14] ^ in2[14];
    assign G[237] = in[13] & in2[13];
    assign P[237] = in[13] ^ in2[13];
    assign G[238] = in[12] & in2[12];
    assign P[238] = in[12] ^ in2[12];
    assign G[239] = in[11] & in2[11];
    assign P[239] = in[11] ^ in2[11];
    assign G[240] = in[10] & in2[10];
    assign P[240] = in[10] ^ in2[10];
    assign G[241] = in[9] & in2[9];
    assign P[241] = in[9] ^ in2[9];
    assign G[242] = in[8] & in2[8];
    assign P[242] = in[8] ^ in2[8];
    assign G[243] = in[7] & in2[7];
    assign P[243] = in[7] ^ in2[7];
    assign G[244] = in[6] & in2[6];
    assign P[244] = in[6] ^ in2[6];
    assign G[245] = in[5] & in2[5];
    assign P[245] = in[5] ^ in2[5];
    assign G[246] = in[4] & in2[4];
    assign P[246] = in[4] ^ in2[4];
    assign G[247] = in[3] & in2[3];
    assign P[247] = in[3] ^ in2[3];
    assign G[248] = in[2] & in2[2];
    assign P[248] = in[2] ^ in2[2];
    assign G[249] = in[1] & in2[1];
    assign P[249] = in[1] ^ in2[1];
    assign G[250] = in[0] & in2[0];
    assign P[250] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign C[250] = G[249] | (P[249] & C[249]);
    assign cout = G[250] | (P[250] & C[250]);
    assign sum = P ^ C;
endmodule

module CLA250(output [249:0] sum, output cout, input [249:0] in1, input [249:0] in2;

    wire[249:0] G;
    wire[249:0] C;
    wire[249:0] P;

    assign G[0] = in[249] & in2[249];
    assign P[0] = in[249] ^ in2[249];
    assign G[1] = in[248] & in2[248];
    assign P[1] = in[248] ^ in2[248];
    assign G[2] = in[247] & in2[247];
    assign P[2] = in[247] ^ in2[247];
    assign G[3] = in[246] & in2[246];
    assign P[3] = in[246] ^ in2[246];
    assign G[4] = in[245] & in2[245];
    assign P[4] = in[245] ^ in2[245];
    assign G[5] = in[244] & in2[244];
    assign P[5] = in[244] ^ in2[244];
    assign G[6] = in[243] & in2[243];
    assign P[6] = in[243] ^ in2[243];
    assign G[7] = in[242] & in2[242];
    assign P[7] = in[242] ^ in2[242];
    assign G[8] = in[241] & in2[241];
    assign P[8] = in[241] ^ in2[241];
    assign G[9] = in[240] & in2[240];
    assign P[9] = in[240] ^ in2[240];
    assign G[10] = in[239] & in2[239];
    assign P[10] = in[239] ^ in2[239];
    assign G[11] = in[238] & in2[238];
    assign P[11] = in[238] ^ in2[238];
    assign G[12] = in[237] & in2[237];
    assign P[12] = in[237] ^ in2[237];
    assign G[13] = in[236] & in2[236];
    assign P[13] = in[236] ^ in2[236];
    assign G[14] = in[235] & in2[235];
    assign P[14] = in[235] ^ in2[235];
    assign G[15] = in[234] & in2[234];
    assign P[15] = in[234] ^ in2[234];
    assign G[16] = in[233] & in2[233];
    assign P[16] = in[233] ^ in2[233];
    assign G[17] = in[232] & in2[232];
    assign P[17] = in[232] ^ in2[232];
    assign G[18] = in[231] & in2[231];
    assign P[18] = in[231] ^ in2[231];
    assign G[19] = in[230] & in2[230];
    assign P[19] = in[230] ^ in2[230];
    assign G[20] = in[229] & in2[229];
    assign P[20] = in[229] ^ in2[229];
    assign G[21] = in[228] & in2[228];
    assign P[21] = in[228] ^ in2[228];
    assign G[22] = in[227] & in2[227];
    assign P[22] = in[227] ^ in2[227];
    assign G[23] = in[226] & in2[226];
    assign P[23] = in[226] ^ in2[226];
    assign G[24] = in[225] & in2[225];
    assign P[24] = in[225] ^ in2[225];
    assign G[25] = in[224] & in2[224];
    assign P[25] = in[224] ^ in2[224];
    assign G[26] = in[223] & in2[223];
    assign P[26] = in[223] ^ in2[223];
    assign G[27] = in[222] & in2[222];
    assign P[27] = in[222] ^ in2[222];
    assign G[28] = in[221] & in2[221];
    assign P[28] = in[221] ^ in2[221];
    assign G[29] = in[220] & in2[220];
    assign P[29] = in[220] ^ in2[220];
    assign G[30] = in[219] & in2[219];
    assign P[30] = in[219] ^ in2[219];
    assign G[31] = in[218] & in2[218];
    assign P[31] = in[218] ^ in2[218];
    assign G[32] = in[217] & in2[217];
    assign P[32] = in[217] ^ in2[217];
    assign G[33] = in[216] & in2[216];
    assign P[33] = in[216] ^ in2[216];
    assign G[34] = in[215] & in2[215];
    assign P[34] = in[215] ^ in2[215];
    assign G[35] = in[214] & in2[214];
    assign P[35] = in[214] ^ in2[214];
    assign G[36] = in[213] & in2[213];
    assign P[36] = in[213] ^ in2[213];
    assign G[37] = in[212] & in2[212];
    assign P[37] = in[212] ^ in2[212];
    assign G[38] = in[211] & in2[211];
    assign P[38] = in[211] ^ in2[211];
    assign G[39] = in[210] & in2[210];
    assign P[39] = in[210] ^ in2[210];
    assign G[40] = in[209] & in2[209];
    assign P[40] = in[209] ^ in2[209];
    assign G[41] = in[208] & in2[208];
    assign P[41] = in[208] ^ in2[208];
    assign G[42] = in[207] & in2[207];
    assign P[42] = in[207] ^ in2[207];
    assign G[43] = in[206] & in2[206];
    assign P[43] = in[206] ^ in2[206];
    assign G[44] = in[205] & in2[205];
    assign P[44] = in[205] ^ in2[205];
    assign G[45] = in[204] & in2[204];
    assign P[45] = in[204] ^ in2[204];
    assign G[46] = in[203] & in2[203];
    assign P[46] = in[203] ^ in2[203];
    assign G[47] = in[202] & in2[202];
    assign P[47] = in[202] ^ in2[202];
    assign G[48] = in[201] & in2[201];
    assign P[48] = in[201] ^ in2[201];
    assign G[49] = in[200] & in2[200];
    assign P[49] = in[200] ^ in2[200];
    assign G[50] = in[199] & in2[199];
    assign P[50] = in[199] ^ in2[199];
    assign G[51] = in[198] & in2[198];
    assign P[51] = in[198] ^ in2[198];
    assign G[52] = in[197] & in2[197];
    assign P[52] = in[197] ^ in2[197];
    assign G[53] = in[196] & in2[196];
    assign P[53] = in[196] ^ in2[196];
    assign G[54] = in[195] & in2[195];
    assign P[54] = in[195] ^ in2[195];
    assign G[55] = in[194] & in2[194];
    assign P[55] = in[194] ^ in2[194];
    assign G[56] = in[193] & in2[193];
    assign P[56] = in[193] ^ in2[193];
    assign G[57] = in[192] & in2[192];
    assign P[57] = in[192] ^ in2[192];
    assign G[58] = in[191] & in2[191];
    assign P[58] = in[191] ^ in2[191];
    assign G[59] = in[190] & in2[190];
    assign P[59] = in[190] ^ in2[190];
    assign G[60] = in[189] & in2[189];
    assign P[60] = in[189] ^ in2[189];
    assign G[61] = in[188] & in2[188];
    assign P[61] = in[188] ^ in2[188];
    assign G[62] = in[187] & in2[187];
    assign P[62] = in[187] ^ in2[187];
    assign G[63] = in[186] & in2[186];
    assign P[63] = in[186] ^ in2[186];
    assign G[64] = in[185] & in2[185];
    assign P[64] = in[185] ^ in2[185];
    assign G[65] = in[184] & in2[184];
    assign P[65] = in[184] ^ in2[184];
    assign G[66] = in[183] & in2[183];
    assign P[66] = in[183] ^ in2[183];
    assign G[67] = in[182] & in2[182];
    assign P[67] = in[182] ^ in2[182];
    assign G[68] = in[181] & in2[181];
    assign P[68] = in[181] ^ in2[181];
    assign G[69] = in[180] & in2[180];
    assign P[69] = in[180] ^ in2[180];
    assign G[70] = in[179] & in2[179];
    assign P[70] = in[179] ^ in2[179];
    assign G[71] = in[178] & in2[178];
    assign P[71] = in[178] ^ in2[178];
    assign G[72] = in[177] & in2[177];
    assign P[72] = in[177] ^ in2[177];
    assign G[73] = in[176] & in2[176];
    assign P[73] = in[176] ^ in2[176];
    assign G[74] = in[175] & in2[175];
    assign P[74] = in[175] ^ in2[175];
    assign G[75] = in[174] & in2[174];
    assign P[75] = in[174] ^ in2[174];
    assign G[76] = in[173] & in2[173];
    assign P[76] = in[173] ^ in2[173];
    assign G[77] = in[172] & in2[172];
    assign P[77] = in[172] ^ in2[172];
    assign G[78] = in[171] & in2[171];
    assign P[78] = in[171] ^ in2[171];
    assign G[79] = in[170] & in2[170];
    assign P[79] = in[170] ^ in2[170];
    assign G[80] = in[169] & in2[169];
    assign P[80] = in[169] ^ in2[169];
    assign G[81] = in[168] & in2[168];
    assign P[81] = in[168] ^ in2[168];
    assign G[82] = in[167] & in2[167];
    assign P[82] = in[167] ^ in2[167];
    assign G[83] = in[166] & in2[166];
    assign P[83] = in[166] ^ in2[166];
    assign G[84] = in[165] & in2[165];
    assign P[84] = in[165] ^ in2[165];
    assign G[85] = in[164] & in2[164];
    assign P[85] = in[164] ^ in2[164];
    assign G[86] = in[163] & in2[163];
    assign P[86] = in[163] ^ in2[163];
    assign G[87] = in[162] & in2[162];
    assign P[87] = in[162] ^ in2[162];
    assign G[88] = in[161] & in2[161];
    assign P[88] = in[161] ^ in2[161];
    assign G[89] = in[160] & in2[160];
    assign P[89] = in[160] ^ in2[160];
    assign G[90] = in[159] & in2[159];
    assign P[90] = in[159] ^ in2[159];
    assign G[91] = in[158] & in2[158];
    assign P[91] = in[158] ^ in2[158];
    assign G[92] = in[157] & in2[157];
    assign P[92] = in[157] ^ in2[157];
    assign G[93] = in[156] & in2[156];
    assign P[93] = in[156] ^ in2[156];
    assign G[94] = in[155] & in2[155];
    assign P[94] = in[155] ^ in2[155];
    assign G[95] = in[154] & in2[154];
    assign P[95] = in[154] ^ in2[154];
    assign G[96] = in[153] & in2[153];
    assign P[96] = in[153] ^ in2[153];
    assign G[97] = in[152] & in2[152];
    assign P[97] = in[152] ^ in2[152];
    assign G[98] = in[151] & in2[151];
    assign P[98] = in[151] ^ in2[151];
    assign G[99] = in[150] & in2[150];
    assign P[99] = in[150] ^ in2[150];
    assign G[100] = in[149] & in2[149];
    assign P[100] = in[149] ^ in2[149];
    assign G[101] = in[148] & in2[148];
    assign P[101] = in[148] ^ in2[148];
    assign G[102] = in[147] & in2[147];
    assign P[102] = in[147] ^ in2[147];
    assign G[103] = in[146] & in2[146];
    assign P[103] = in[146] ^ in2[146];
    assign G[104] = in[145] & in2[145];
    assign P[104] = in[145] ^ in2[145];
    assign G[105] = in[144] & in2[144];
    assign P[105] = in[144] ^ in2[144];
    assign G[106] = in[143] & in2[143];
    assign P[106] = in[143] ^ in2[143];
    assign G[107] = in[142] & in2[142];
    assign P[107] = in[142] ^ in2[142];
    assign G[108] = in[141] & in2[141];
    assign P[108] = in[141] ^ in2[141];
    assign G[109] = in[140] & in2[140];
    assign P[109] = in[140] ^ in2[140];
    assign G[110] = in[139] & in2[139];
    assign P[110] = in[139] ^ in2[139];
    assign G[111] = in[138] & in2[138];
    assign P[111] = in[138] ^ in2[138];
    assign G[112] = in[137] & in2[137];
    assign P[112] = in[137] ^ in2[137];
    assign G[113] = in[136] & in2[136];
    assign P[113] = in[136] ^ in2[136];
    assign G[114] = in[135] & in2[135];
    assign P[114] = in[135] ^ in2[135];
    assign G[115] = in[134] & in2[134];
    assign P[115] = in[134] ^ in2[134];
    assign G[116] = in[133] & in2[133];
    assign P[116] = in[133] ^ in2[133];
    assign G[117] = in[132] & in2[132];
    assign P[117] = in[132] ^ in2[132];
    assign G[118] = in[131] & in2[131];
    assign P[118] = in[131] ^ in2[131];
    assign G[119] = in[130] & in2[130];
    assign P[119] = in[130] ^ in2[130];
    assign G[120] = in[129] & in2[129];
    assign P[120] = in[129] ^ in2[129];
    assign G[121] = in[128] & in2[128];
    assign P[121] = in[128] ^ in2[128];
    assign G[122] = in[127] & in2[127];
    assign P[122] = in[127] ^ in2[127];
    assign G[123] = in[126] & in2[126];
    assign P[123] = in[126] ^ in2[126];
    assign G[124] = in[125] & in2[125];
    assign P[124] = in[125] ^ in2[125];
    assign G[125] = in[124] & in2[124];
    assign P[125] = in[124] ^ in2[124];
    assign G[126] = in[123] & in2[123];
    assign P[126] = in[123] ^ in2[123];
    assign G[127] = in[122] & in2[122];
    assign P[127] = in[122] ^ in2[122];
    assign G[128] = in[121] & in2[121];
    assign P[128] = in[121] ^ in2[121];
    assign G[129] = in[120] & in2[120];
    assign P[129] = in[120] ^ in2[120];
    assign G[130] = in[119] & in2[119];
    assign P[130] = in[119] ^ in2[119];
    assign G[131] = in[118] & in2[118];
    assign P[131] = in[118] ^ in2[118];
    assign G[132] = in[117] & in2[117];
    assign P[132] = in[117] ^ in2[117];
    assign G[133] = in[116] & in2[116];
    assign P[133] = in[116] ^ in2[116];
    assign G[134] = in[115] & in2[115];
    assign P[134] = in[115] ^ in2[115];
    assign G[135] = in[114] & in2[114];
    assign P[135] = in[114] ^ in2[114];
    assign G[136] = in[113] & in2[113];
    assign P[136] = in[113] ^ in2[113];
    assign G[137] = in[112] & in2[112];
    assign P[137] = in[112] ^ in2[112];
    assign G[138] = in[111] & in2[111];
    assign P[138] = in[111] ^ in2[111];
    assign G[139] = in[110] & in2[110];
    assign P[139] = in[110] ^ in2[110];
    assign G[140] = in[109] & in2[109];
    assign P[140] = in[109] ^ in2[109];
    assign G[141] = in[108] & in2[108];
    assign P[141] = in[108] ^ in2[108];
    assign G[142] = in[107] & in2[107];
    assign P[142] = in[107] ^ in2[107];
    assign G[143] = in[106] & in2[106];
    assign P[143] = in[106] ^ in2[106];
    assign G[144] = in[105] & in2[105];
    assign P[144] = in[105] ^ in2[105];
    assign G[145] = in[104] & in2[104];
    assign P[145] = in[104] ^ in2[104];
    assign G[146] = in[103] & in2[103];
    assign P[146] = in[103] ^ in2[103];
    assign G[147] = in[102] & in2[102];
    assign P[147] = in[102] ^ in2[102];
    assign G[148] = in[101] & in2[101];
    assign P[148] = in[101] ^ in2[101];
    assign G[149] = in[100] & in2[100];
    assign P[149] = in[100] ^ in2[100];
    assign G[150] = in[99] & in2[99];
    assign P[150] = in[99] ^ in2[99];
    assign G[151] = in[98] & in2[98];
    assign P[151] = in[98] ^ in2[98];
    assign G[152] = in[97] & in2[97];
    assign P[152] = in[97] ^ in2[97];
    assign G[153] = in[96] & in2[96];
    assign P[153] = in[96] ^ in2[96];
    assign G[154] = in[95] & in2[95];
    assign P[154] = in[95] ^ in2[95];
    assign G[155] = in[94] & in2[94];
    assign P[155] = in[94] ^ in2[94];
    assign G[156] = in[93] & in2[93];
    assign P[156] = in[93] ^ in2[93];
    assign G[157] = in[92] & in2[92];
    assign P[157] = in[92] ^ in2[92];
    assign G[158] = in[91] & in2[91];
    assign P[158] = in[91] ^ in2[91];
    assign G[159] = in[90] & in2[90];
    assign P[159] = in[90] ^ in2[90];
    assign G[160] = in[89] & in2[89];
    assign P[160] = in[89] ^ in2[89];
    assign G[161] = in[88] & in2[88];
    assign P[161] = in[88] ^ in2[88];
    assign G[162] = in[87] & in2[87];
    assign P[162] = in[87] ^ in2[87];
    assign G[163] = in[86] & in2[86];
    assign P[163] = in[86] ^ in2[86];
    assign G[164] = in[85] & in2[85];
    assign P[164] = in[85] ^ in2[85];
    assign G[165] = in[84] & in2[84];
    assign P[165] = in[84] ^ in2[84];
    assign G[166] = in[83] & in2[83];
    assign P[166] = in[83] ^ in2[83];
    assign G[167] = in[82] & in2[82];
    assign P[167] = in[82] ^ in2[82];
    assign G[168] = in[81] & in2[81];
    assign P[168] = in[81] ^ in2[81];
    assign G[169] = in[80] & in2[80];
    assign P[169] = in[80] ^ in2[80];
    assign G[170] = in[79] & in2[79];
    assign P[170] = in[79] ^ in2[79];
    assign G[171] = in[78] & in2[78];
    assign P[171] = in[78] ^ in2[78];
    assign G[172] = in[77] & in2[77];
    assign P[172] = in[77] ^ in2[77];
    assign G[173] = in[76] & in2[76];
    assign P[173] = in[76] ^ in2[76];
    assign G[174] = in[75] & in2[75];
    assign P[174] = in[75] ^ in2[75];
    assign G[175] = in[74] & in2[74];
    assign P[175] = in[74] ^ in2[74];
    assign G[176] = in[73] & in2[73];
    assign P[176] = in[73] ^ in2[73];
    assign G[177] = in[72] & in2[72];
    assign P[177] = in[72] ^ in2[72];
    assign G[178] = in[71] & in2[71];
    assign P[178] = in[71] ^ in2[71];
    assign G[179] = in[70] & in2[70];
    assign P[179] = in[70] ^ in2[70];
    assign G[180] = in[69] & in2[69];
    assign P[180] = in[69] ^ in2[69];
    assign G[181] = in[68] & in2[68];
    assign P[181] = in[68] ^ in2[68];
    assign G[182] = in[67] & in2[67];
    assign P[182] = in[67] ^ in2[67];
    assign G[183] = in[66] & in2[66];
    assign P[183] = in[66] ^ in2[66];
    assign G[184] = in[65] & in2[65];
    assign P[184] = in[65] ^ in2[65];
    assign G[185] = in[64] & in2[64];
    assign P[185] = in[64] ^ in2[64];
    assign G[186] = in[63] & in2[63];
    assign P[186] = in[63] ^ in2[63];
    assign G[187] = in[62] & in2[62];
    assign P[187] = in[62] ^ in2[62];
    assign G[188] = in[61] & in2[61];
    assign P[188] = in[61] ^ in2[61];
    assign G[189] = in[60] & in2[60];
    assign P[189] = in[60] ^ in2[60];
    assign G[190] = in[59] & in2[59];
    assign P[190] = in[59] ^ in2[59];
    assign G[191] = in[58] & in2[58];
    assign P[191] = in[58] ^ in2[58];
    assign G[192] = in[57] & in2[57];
    assign P[192] = in[57] ^ in2[57];
    assign G[193] = in[56] & in2[56];
    assign P[193] = in[56] ^ in2[56];
    assign G[194] = in[55] & in2[55];
    assign P[194] = in[55] ^ in2[55];
    assign G[195] = in[54] & in2[54];
    assign P[195] = in[54] ^ in2[54];
    assign G[196] = in[53] & in2[53];
    assign P[196] = in[53] ^ in2[53];
    assign G[197] = in[52] & in2[52];
    assign P[197] = in[52] ^ in2[52];
    assign G[198] = in[51] & in2[51];
    assign P[198] = in[51] ^ in2[51];
    assign G[199] = in[50] & in2[50];
    assign P[199] = in[50] ^ in2[50];
    assign G[200] = in[49] & in2[49];
    assign P[200] = in[49] ^ in2[49];
    assign G[201] = in[48] & in2[48];
    assign P[201] = in[48] ^ in2[48];
    assign G[202] = in[47] & in2[47];
    assign P[202] = in[47] ^ in2[47];
    assign G[203] = in[46] & in2[46];
    assign P[203] = in[46] ^ in2[46];
    assign G[204] = in[45] & in2[45];
    assign P[204] = in[45] ^ in2[45];
    assign G[205] = in[44] & in2[44];
    assign P[205] = in[44] ^ in2[44];
    assign G[206] = in[43] & in2[43];
    assign P[206] = in[43] ^ in2[43];
    assign G[207] = in[42] & in2[42];
    assign P[207] = in[42] ^ in2[42];
    assign G[208] = in[41] & in2[41];
    assign P[208] = in[41] ^ in2[41];
    assign G[209] = in[40] & in2[40];
    assign P[209] = in[40] ^ in2[40];
    assign G[210] = in[39] & in2[39];
    assign P[210] = in[39] ^ in2[39];
    assign G[211] = in[38] & in2[38];
    assign P[211] = in[38] ^ in2[38];
    assign G[212] = in[37] & in2[37];
    assign P[212] = in[37] ^ in2[37];
    assign G[213] = in[36] & in2[36];
    assign P[213] = in[36] ^ in2[36];
    assign G[214] = in[35] & in2[35];
    assign P[214] = in[35] ^ in2[35];
    assign G[215] = in[34] & in2[34];
    assign P[215] = in[34] ^ in2[34];
    assign G[216] = in[33] & in2[33];
    assign P[216] = in[33] ^ in2[33];
    assign G[217] = in[32] & in2[32];
    assign P[217] = in[32] ^ in2[32];
    assign G[218] = in[31] & in2[31];
    assign P[218] = in[31] ^ in2[31];
    assign G[219] = in[30] & in2[30];
    assign P[219] = in[30] ^ in2[30];
    assign G[220] = in[29] & in2[29];
    assign P[220] = in[29] ^ in2[29];
    assign G[221] = in[28] & in2[28];
    assign P[221] = in[28] ^ in2[28];
    assign G[222] = in[27] & in2[27];
    assign P[222] = in[27] ^ in2[27];
    assign G[223] = in[26] & in2[26];
    assign P[223] = in[26] ^ in2[26];
    assign G[224] = in[25] & in2[25];
    assign P[224] = in[25] ^ in2[25];
    assign G[225] = in[24] & in2[24];
    assign P[225] = in[24] ^ in2[24];
    assign G[226] = in[23] & in2[23];
    assign P[226] = in[23] ^ in2[23];
    assign G[227] = in[22] & in2[22];
    assign P[227] = in[22] ^ in2[22];
    assign G[228] = in[21] & in2[21];
    assign P[228] = in[21] ^ in2[21];
    assign G[229] = in[20] & in2[20];
    assign P[229] = in[20] ^ in2[20];
    assign G[230] = in[19] & in2[19];
    assign P[230] = in[19] ^ in2[19];
    assign G[231] = in[18] & in2[18];
    assign P[231] = in[18] ^ in2[18];
    assign G[232] = in[17] & in2[17];
    assign P[232] = in[17] ^ in2[17];
    assign G[233] = in[16] & in2[16];
    assign P[233] = in[16] ^ in2[16];
    assign G[234] = in[15] & in2[15];
    assign P[234] = in[15] ^ in2[15];
    assign G[235] = in[14] & in2[14];
    assign P[235] = in[14] ^ in2[14];
    assign G[236] = in[13] & in2[13];
    assign P[236] = in[13] ^ in2[13];
    assign G[237] = in[12] & in2[12];
    assign P[237] = in[12] ^ in2[12];
    assign G[238] = in[11] & in2[11];
    assign P[238] = in[11] ^ in2[11];
    assign G[239] = in[10] & in2[10];
    assign P[239] = in[10] ^ in2[10];
    assign G[240] = in[9] & in2[9];
    assign P[240] = in[9] ^ in2[9];
    assign G[241] = in[8] & in2[8];
    assign P[241] = in[8] ^ in2[8];
    assign G[242] = in[7] & in2[7];
    assign P[242] = in[7] ^ in2[7];
    assign G[243] = in[6] & in2[6];
    assign P[243] = in[6] ^ in2[6];
    assign G[244] = in[5] & in2[5];
    assign P[244] = in[5] ^ in2[5];
    assign G[245] = in[4] & in2[4];
    assign P[245] = in[4] ^ in2[4];
    assign G[246] = in[3] & in2[3];
    assign P[246] = in[3] ^ in2[3];
    assign G[247] = in[2] & in2[2];
    assign P[247] = in[2] ^ in2[2];
    assign G[248] = in[1] & in2[1];
    assign P[248] = in[1] ^ in2[1];
    assign G[249] = in[0] & in2[0];
    assign P[249] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign C[249] = G[248] | (P[248] & C[248]);
    assign cout = G[249] | (P[249] & C[249]);
    assign sum = P ^ C;
endmodule

module CLA249(output [248:0] sum, output cout, input [248:0] in1, input [248:0] in2;

    wire[248:0] G;
    wire[248:0] C;
    wire[248:0] P;

    assign G[0] = in[248] & in2[248];
    assign P[0] = in[248] ^ in2[248];
    assign G[1] = in[247] & in2[247];
    assign P[1] = in[247] ^ in2[247];
    assign G[2] = in[246] & in2[246];
    assign P[2] = in[246] ^ in2[246];
    assign G[3] = in[245] & in2[245];
    assign P[3] = in[245] ^ in2[245];
    assign G[4] = in[244] & in2[244];
    assign P[4] = in[244] ^ in2[244];
    assign G[5] = in[243] & in2[243];
    assign P[5] = in[243] ^ in2[243];
    assign G[6] = in[242] & in2[242];
    assign P[6] = in[242] ^ in2[242];
    assign G[7] = in[241] & in2[241];
    assign P[7] = in[241] ^ in2[241];
    assign G[8] = in[240] & in2[240];
    assign P[8] = in[240] ^ in2[240];
    assign G[9] = in[239] & in2[239];
    assign P[9] = in[239] ^ in2[239];
    assign G[10] = in[238] & in2[238];
    assign P[10] = in[238] ^ in2[238];
    assign G[11] = in[237] & in2[237];
    assign P[11] = in[237] ^ in2[237];
    assign G[12] = in[236] & in2[236];
    assign P[12] = in[236] ^ in2[236];
    assign G[13] = in[235] & in2[235];
    assign P[13] = in[235] ^ in2[235];
    assign G[14] = in[234] & in2[234];
    assign P[14] = in[234] ^ in2[234];
    assign G[15] = in[233] & in2[233];
    assign P[15] = in[233] ^ in2[233];
    assign G[16] = in[232] & in2[232];
    assign P[16] = in[232] ^ in2[232];
    assign G[17] = in[231] & in2[231];
    assign P[17] = in[231] ^ in2[231];
    assign G[18] = in[230] & in2[230];
    assign P[18] = in[230] ^ in2[230];
    assign G[19] = in[229] & in2[229];
    assign P[19] = in[229] ^ in2[229];
    assign G[20] = in[228] & in2[228];
    assign P[20] = in[228] ^ in2[228];
    assign G[21] = in[227] & in2[227];
    assign P[21] = in[227] ^ in2[227];
    assign G[22] = in[226] & in2[226];
    assign P[22] = in[226] ^ in2[226];
    assign G[23] = in[225] & in2[225];
    assign P[23] = in[225] ^ in2[225];
    assign G[24] = in[224] & in2[224];
    assign P[24] = in[224] ^ in2[224];
    assign G[25] = in[223] & in2[223];
    assign P[25] = in[223] ^ in2[223];
    assign G[26] = in[222] & in2[222];
    assign P[26] = in[222] ^ in2[222];
    assign G[27] = in[221] & in2[221];
    assign P[27] = in[221] ^ in2[221];
    assign G[28] = in[220] & in2[220];
    assign P[28] = in[220] ^ in2[220];
    assign G[29] = in[219] & in2[219];
    assign P[29] = in[219] ^ in2[219];
    assign G[30] = in[218] & in2[218];
    assign P[30] = in[218] ^ in2[218];
    assign G[31] = in[217] & in2[217];
    assign P[31] = in[217] ^ in2[217];
    assign G[32] = in[216] & in2[216];
    assign P[32] = in[216] ^ in2[216];
    assign G[33] = in[215] & in2[215];
    assign P[33] = in[215] ^ in2[215];
    assign G[34] = in[214] & in2[214];
    assign P[34] = in[214] ^ in2[214];
    assign G[35] = in[213] & in2[213];
    assign P[35] = in[213] ^ in2[213];
    assign G[36] = in[212] & in2[212];
    assign P[36] = in[212] ^ in2[212];
    assign G[37] = in[211] & in2[211];
    assign P[37] = in[211] ^ in2[211];
    assign G[38] = in[210] & in2[210];
    assign P[38] = in[210] ^ in2[210];
    assign G[39] = in[209] & in2[209];
    assign P[39] = in[209] ^ in2[209];
    assign G[40] = in[208] & in2[208];
    assign P[40] = in[208] ^ in2[208];
    assign G[41] = in[207] & in2[207];
    assign P[41] = in[207] ^ in2[207];
    assign G[42] = in[206] & in2[206];
    assign P[42] = in[206] ^ in2[206];
    assign G[43] = in[205] & in2[205];
    assign P[43] = in[205] ^ in2[205];
    assign G[44] = in[204] & in2[204];
    assign P[44] = in[204] ^ in2[204];
    assign G[45] = in[203] & in2[203];
    assign P[45] = in[203] ^ in2[203];
    assign G[46] = in[202] & in2[202];
    assign P[46] = in[202] ^ in2[202];
    assign G[47] = in[201] & in2[201];
    assign P[47] = in[201] ^ in2[201];
    assign G[48] = in[200] & in2[200];
    assign P[48] = in[200] ^ in2[200];
    assign G[49] = in[199] & in2[199];
    assign P[49] = in[199] ^ in2[199];
    assign G[50] = in[198] & in2[198];
    assign P[50] = in[198] ^ in2[198];
    assign G[51] = in[197] & in2[197];
    assign P[51] = in[197] ^ in2[197];
    assign G[52] = in[196] & in2[196];
    assign P[52] = in[196] ^ in2[196];
    assign G[53] = in[195] & in2[195];
    assign P[53] = in[195] ^ in2[195];
    assign G[54] = in[194] & in2[194];
    assign P[54] = in[194] ^ in2[194];
    assign G[55] = in[193] & in2[193];
    assign P[55] = in[193] ^ in2[193];
    assign G[56] = in[192] & in2[192];
    assign P[56] = in[192] ^ in2[192];
    assign G[57] = in[191] & in2[191];
    assign P[57] = in[191] ^ in2[191];
    assign G[58] = in[190] & in2[190];
    assign P[58] = in[190] ^ in2[190];
    assign G[59] = in[189] & in2[189];
    assign P[59] = in[189] ^ in2[189];
    assign G[60] = in[188] & in2[188];
    assign P[60] = in[188] ^ in2[188];
    assign G[61] = in[187] & in2[187];
    assign P[61] = in[187] ^ in2[187];
    assign G[62] = in[186] & in2[186];
    assign P[62] = in[186] ^ in2[186];
    assign G[63] = in[185] & in2[185];
    assign P[63] = in[185] ^ in2[185];
    assign G[64] = in[184] & in2[184];
    assign P[64] = in[184] ^ in2[184];
    assign G[65] = in[183] & in2[183];
    assign P[65] = in[183] ^ in2[183];
    assign G[66] = in[182] & in2[182];
    assign P[66] = in[182] ^ in2[182];
    assign G[67] = in[181] & in2[181];
    assign P[67] = in[181] ^ in2[181];
    assign G[68] = in[180] & in2[180];
    assign P[68] = in[180] ^ in2[180];
    assign G[69] = in[179] & in2[179];
    assign P[69] = in[179] ^ in2[179];
    assign G[70] = in[178] & in2[178];
    assign P[70] = in[178] ^ in2[178];
    assign G[71] = in[177] & in2[177];
    assign P[71] = in[177] ^ in2[177];
    assign G[72] = in[176] & in2[176];
    assign P[72] = in[176] ^ in2[176];
    assign G[73] = in[175] & in2[175];
    assign P[73] = in[175] ^ in2[175];
    assign G[74] = in[174] & in2[174];
    assign P[74] = in[174] ^ in2[174];
    assign G[75] = in[173] & in2[173];
    assign P[75] = in[173] ^ in2[173];
    assign G[76] = in[172] & in2[172];
    assign P[76] = in[172] ^ in2[172];
    assign G[77] = in[171] & in2[171];
    assign P[77] = in[171] ^ in2[171];
    assign G[78] = in[170] & in2[170];
    assign P[78] = in[170] ^ in2[170];
    assign G[79] = in[169] & in2[169];
    assign P[79] = in[169] ^ in2[169];
    assign G[80] = in[168] & in2[168];
    assign P[80] = in[168] ^ in2[168];
    assign G[81] = in[167] & in2[167];
    assign P[81] = in[167] ^ in2[167];
    assign G[82] = in[166] & in2[166];
    assign P[82] = in[166] ^ in2[166];
    assign G[83] = in[165] & in2[165];
    assign P[83] = in[165] ^ in2[165];
    assign G[84] = in[164] & in2[164];
    assign P[84] = in[164] ^ in2[164];
    assign G[85] = in[163] & in2[163];
    assign P[85] = in[163] ^ in2[163];
    assign G[86] = in[162] & in2[162];
    assign P[86] = in[162] ^ in2[162];
    assign G[87] = in[161] & in2[161];
    assign P[87] = in[161] ^ in2[161];
    assign G[88] = in[160] & in2[160];
    assign P[88] = in[160] ^ in2[160];
    assign G[89] = in[159] & in2[159];
    assign P[89] = in[159] ^ in2[159];
    assign G[90] = in[158] & in2[158];
    assign P[90] = in[158] ^ in2[158];
    assign G[91] = in[157] & in2[157];
    assign P[91] = in[157] ^ in2[157];
    assign G[92] = in[156] & in2[156];
    assign P[92] = in[156] ^ in2[156];
    assign G[93] = in[155] & in2[155];
    assign P[93] = in[155] ^ in2[155];
    assign G[94] = in[154] & in2[154];
    assign P[94] = in[154] ^ in2[154];
    assign G[95] = in[153] & in2[153];
    assign P[95] = in[153] ^ in2[153];
    assign G[96] = in[152] & in2[152];
    assign P[96] = in[152] ^ in2[152];
    assign G[97] = in[151] & in2[151];
    assign P[97] = in[151] ^ in2[151];
    assign G[98] = in[150] & in2[150];
    assign P[98] = in[150] ^ in2[150];
    assign G[99] = in[149] & in2[149];
    assign P[99] = in[149] ^ in2[149];
    assign G[100] = in[148] & in2[148];
    assign P[100] = in[148] ^ in2[148];
    assign G[101] = in[147] & in2[147];
    assign P[101] = in[147] ^ in2[147];
    assign G[102] = in[146] & in2[146];
    assign P[102] = in[146] ^ in2[146];
    assign G[103] = in[145] & in2[145];
    assign P[103] = in[145] ^ in2[145];
    assign G[104] = in[144] & in2[144];
    assign P[104] = in[144] ^ in2[144];
    assign G[105] = in[143] & in2[143];
    assign P[105] = in[143] ^ in2[143];
    assign G[106] = in[142] & in2[142];
    assign P[106] = in[142] ^ in2[142];
    assign G[107] = in[141] & in2[141];
    assign P[107] = in[141] ^ in2[141];
    assign G[108] = in[140] & in2[140];
    assign P[108] = in[140] ^ in2[140];
    assign G[109] = in[139] & in2[139];
    assign P[109] = in[139] ^ in2[139];
    assign G[110] = in[138] & in2[138];
    assign P[110] = in[138] ^ in2[138];
    assign G[111] = in[137] & in2[137];
    assign P[111] = in[137] ^ in2[137];
    assign G[112] = in[136] & in2[136];
    assign P[112] = in[136] ^ in2[136];
    assign G[113] = in[135] & in2[135];
    assign P[113] = in[135] ^ in2[135];
    assign G[114] = in[134] & in2[134];
    assign P[114] = in[134] ^ in2[134];
    assign G[115] = in[133] & in2[133];
    assign P[115] = in[133] ^ in2[133];
    assign G[116] = in[132] & in2[132];
    assign P[116] = in[132] ^ in2[132];
    assign G[117] = in[131] & in2[131];
    assign P[117] = in[131] ^ in2[131];
    assign G[118] = in[130] & in2[130];
    assign P[118] = in[130] ^ in2[130];
    assign G[119] = in[129] & in2[129];
    assign P[119] = in[129] ^ in2[129];
    assign G[120] = in[128] & in2[128];
    assign P[120] = in[128] ^ in2[128];
    assign G[121] = in[127] & in2[127];
    assign P[121] = in[127] ^ in2[127];
    assign G[122] = in[126] & in2[126];
    assign P[122] = in[126] ^ in2[126];
    assign G[123] = in[125] & in2[125];
    assign P[123] = in[125] ^ in2[125];
    assign G[124] = in[124] & in2[124];
    assign P[124] = in[124] ^ in2[124];
    assign G[125] = in[123] & in2[123];
    assign P[125] = in[123] ^ in2[123];
    assign G[126] = in[122] & in2[122];
    assign P[126] = in[122] ^ in2[122];
    assign G[127] = in[121] & in2[121];
    assign P[127] = in[121] ^ in2[121];
    assign G[128] = in[120] & in2[120];
    assign P[128] = in[120] ^ in2[120];
    assign G[129] = in[119] & in2[119];
    assign P[129] = in[119] ^ in2[119];
    assign G[130] = in[118] & in2[118];
    assign P[130] = in[118] ^ in2[118];
    assign G[131] = in[117] & in2[117];
    assign P[131] = in[117] ^ in2[117];
    assign G[132] = in[116] & in2[116];
    assign P[132] = in[116] ^ in2[116];
    assign G[133] = in[115] & in2[115];
    assign P[133] = in[115] ^ in2[115];
    assign G[134] = in[114] & in2[114];
    assign P[134] = in[114] ^ in2[114];
    assign G[135] = in[113] & in2[113];
    assign P[135] = in[113] ^ in2[113];
    assign G[136] = in[112] & in2[112];
    assign P[136] = in[112] ^ in2[112];
    assign G[137] = in[111] & in2[111];
    assign P[137] = in[111] ^ in2[111];
    assign G[138] = in[110] & in2[110];
    assign P[138] = in[110] ^ in2[110];
    assign G[139] = in[109] & in2[109];
    assign P[139] = in[109] ^ in2[109];
    assign G[140] = in[108] & in2[108];
    assign P[140] = in[108] ^ in2[108];
    assign G[141] = in[107] & in2[107];
    assign P[141] = in[107] ^ in2[107];
    assign G[142] = in[106] & in2[106];
    assign P[142] = in[106] ^ in2[106];
    assign G[143] = in[105] & in2[105];
    assign P[143] = in[105] ^ in2[105];
    assign G[144] = in[104] & in2[104];
    assign P[144] = in[104] ^ in2[104];
    assign G[145] = in[103] & in2[103];
    assign P[145] = in[103] ^ in2[103];
    assign G[146] = in[102] & in2[102];
    assign P[146] = in[102] ^ in2[102];
    assign G[147] = in[101] & in2[101];
    assign P[147] = in[101] ^ in2[101];
    assign G[148] = in[100] & in2[100];
    assign P[148] = in[100] ^ in2[100];
    assign G[149] = in[99] & in2[99];
    assign P[149] = in[99] ^ in2[99];
    assign G[150] = in[98] & in2[98];
    assign P[150] = in[98] ^ in2[98];
    assign G[151] = in[97] & in2[97];
    assign P[151] = in[97] ^ in2[97];
    assign G[152] = in[96] & in2[96];
    assign P[152] = in[96] ^ in2[96];
    assign G[153] = in[95] & in2[95];
    assign P[153] = in[95] ^ in2[95];
    assign G[154] = in[94] & in2[94];
    assign P[154] = in[94] ^ in2[94];
    assign G[155] = in[93] & in2[93];
    assign P[155] = in[93] ^ in2[93];
    assign G[156] = in[92] & in2[92];
    assign P[156] = in[92] ^ in2[92];
    assign G[157] = in[91] & in2[91];
    assign P[157] = in[91] ^ in2[91];
    assign G[158] = in[90] & in2[90];
    assign P[158] = in[90] ^ in2[90];
    assign G[159] = in[89] & in2[89];
    assign P[159] = in[89] ^ in2[89];
    assign G[160] = in[88] & in2[88];
    assign P[160] = in[88] ^ in2[88];
    assign G[161] = in[87] & in2[87];
    assign P[161] = in[87] ^ in2[87];
    assign G[162] = in[86] & in2[86];
    assign P[162] = in[86] ^ in2[86];
    assign G[163] = in[85] & in2[85];
    assign P[163] = in[85] ^ in2[85];
    assign G[164] = in[84] & in2[84];
    assign P[164] = in[84] ^ in2[84];
    assign G[165] = in[83] & in2[83];
    assign P[165] = in[83] ^ in2[83];
    assign G[166] = in[82] & in2[82];
    assign P[166] = in[82] ^ in2[82];
    assign G[167] = in[81] & in2[81];
    assign P[167] = in[81] ^ in2[81];
    assign G[168] = in[80] & in2[80];
    assign P[168] = in[80] ^ in2[80];
    assign G[169] = in[79] & in2[79];
    assign P[169] = in[79] ^ in2[79];
    assign G[170] = in[78] & in2[78];
    assign P[170] = in[78] ^ in2[78];
    assign G[171] = in[77] & in2[77];
    assign P[171] = in[77] ^ in2[77];
    assign G[172] = in[76] & in2[76];
    assign P[172] = in[76] ^ in2[76];
    assign G[173] = in[75] & in2[75];
    assign P[173] = in[75] ^ in2[75];
    assign G[174] = in[74] & in2[74];
    assign P[174] = in[74] ^ in2[74];
    assign G[175] = in[73] & in2[73];
    assign P[175] = in[73] ^ in2[73];
    assign G[176] = in[72] & in2[72];
    assign P[176] = in[72] ^ in2[72];
    assign G[177] = in[71] & in2[71];
    assign P[177] = in[71] ^ in2[71];
    assign G[178] = in[70] & in2[70];
    assign P[178] = in[70] ^ in2[70];
    assign G[179] = in[69] & in2[69];
    assign P[179] = in[69] ^ in2[69];
    assign G[180] = in[68] & in2[68];
    assign P[180] = in[68] ^ in2[68];
    assign G[181] = in[67] & in2[67];
    assign P[181] = in[67] ^ in2[67];
    assign G[182] = in[66] & in2[66];
    assign P[182] = in[66] ^ in2[66];
    assign G[183] = in[65] & in2[65];
    assign P[183] = in[65] ^ in2[65];
    assign G[184] = in[64] & in2[64];
    assign P[184] = in[64] ^ in2[64];
    assign G[185] = in[63] & in2[63];
    assign P[185] = in[63] ^ in2[63];
    assign G[186] = in[62] & in2[62];
    assign P[186] = in[62] ^ in2[62];
    assign G[187] = in[61] & in2[61];
    assign P[187] = in[61] ^ in2[61];
    assign G[188] = in[60] & in2[60];
    assign P[188] = in[60] ^ in2[60];
    assign G[189] = in[59] & in2[59];
    assign P[189] = in[59] ^ in2[59];
    assign G[190] = in[58] & in2[58];
    assign P[190] = in[58] ^ in2[58];
    assign G[191] = in[57] & in2[57];
    assign P[191] = in[57] ^ in2[57];
    assign G[192] = in[56] & in2[56];
    assign P[192] = in[56] ^ in2[56];
    assign G[193] = in[55] & in2[55];
    assign P[193] = in[55] ^ in2[55];
    assign G[194] = in[54] & in2[54];
    assign P[194] = in[54] ^ in2[54];
    assign G[195] = in[53] & in2[53];
    assign P[195] = in[53] ^ in2[53];
    assign G[196] = in[52] & in2[52];
    assign P[196] = in[52] ^ in2[52];
    assign G[197] = in[51] & in2[51];
    assign P[197] = in[51] ^ in2[51];
    assign G[198] = in[50] & in2[50];
    assign P[198] = in[50] ^ in2[50];
    assign G[199] = in[49] & in2[49];
    assign P[199] = in[49] ^ in2[49];
    assign G[200] = in[48] & in2[48];
    assign P[200] = in[48] ^ in2[48];
    assign G[201] = in[47] & in2[47];
    assign P[201] = in[47] ^ in2[47];
    assign G[202] = in[46] & in2[46];
    assign P[202] = in[46] ^ in2[46];
    assign G[203] = in[45] & in2[45];
    assign P[203] = in[45] ^ in2[45];
    assign G[204] = in[44] & in2[44];
    assign P[204] = in[44] ^ in2[44];
    assign G[205] = in[43] & in2[43];
    assign P[205] = in[43] ^ in2[43];
    assign G[206] = in[42] & in2[42];
    assign P[206] = in[42] ^ in2[42];
    assign G[207] = in[41] & in2[41];
    assign P[207] = in[41] ^ in2[41];
    assign G[208] = in[40] & in2[40];
    assign P[208] = in[40] ^ in2[40];
    assign G[209] = in[39] & in2[39];
    assign P[209] = in[39] ^ in2[39];
    assign G[210] = in[38] & in2[38];
    assign P[210] = in[38] ^ in2[38];
    assign G[211] = in[37] & in2[37];
    assign P[211] = in[37] ^ in2[37];
    assign G[212] = in[36] & in2[36];
    assign P[212] = in[36] ^ in2[36];
    assign G[213] = in[35] & in2[35];
    assign P[213] = in[35] ^ in2[35];
    assign G[214] = in[34] & in2[34];
    assign P[214] = in[34] ^ in2[34];
    assign G[215] = in[33] & in2[33];
    assign P[215] = in[33] ^ in2[33];
    assign G[216] = in[32] & in2[32];
    assign P[216] = in[32] ^ in2[32];
    assign G[217] = in[31] & in2[31];
    assign P[217] = in[31] ^ in2[31];
    assign G[218] = in[30] & in2[30];
    assign P[218] = in[30] ^ in2[30];
    assign G[219] = in[29] & in2[29];
    assign P[219] = in[29] ^ in2[29];
    assign G[220] = in[28] & in2[28];
    assign P[220] = in[28] ^ in2[28];
    assign G[221] = in[27] & in2[27];
    assign P[221] = in[27] ^ in2[27];
    assign G[222] = in[26] & in2[26];
    assign P[222] = in[26] ^ in2[26];
    assign G[223] = in[25] & in2[25];
    assign P[223] = in[25] ^ in2[25];
    assign G[224] = in[24] & in2[24];
    assign P[224] = in[24] ^ in2[24];
    assign G[225] = in[23] & in2[23];
    assign P[225] = in[23] ^ in2[23];
    assign G[226] = in[22] & in2[22];
    assign P[226] = in[22] ^ in2[22];
    assign G[227] = in[21] & in2[21];
    assign P[227] = in[21] ^ in2[21];
    assign G[228] = in[20] & in2[20];
    assign P[228] = in[20] ^ in2[20];
    assign G[229] = in[19] & in2[19];
    assign P[229] = in[19] ^ in2[19];
    assign G[230] = in[18] & in2[18];
    assign P[230] = in[18] ^ in2[18];
    assign G[231] = in[17] & in2[17];
    assign P[231] = in[17] ^ in2[17];
    assign G[232] = in[16] & in2[16];
    assign P[232] = in[16] ^ in2[16];
    assign G[233] = in[15] & in2[15];
    assign P[233] = in[15] ^ in2[15];
    assign G[234] = in[14] & in2[14];
    assign P[234] = in[14] ^ in2[14];
    assign G[235] = in[13] & in2[13];
    assign P[235] = in[13] ^ in2[13];
    assign G[236] = in[12] & in2[12];
    assign P[236] = in[12] ^ in2[12];
    assign G[237] = in[11] & in2[11];
    assign P[237] = in[11] ^ in2[11];
    assign G[238] = in[10] & in2[10];
    assign P[238] = in[10] ^ in2[10];
    assign G[239] = in[9] & in2[9];
    assign P[239] = in[9] ^ in2[9];
    assign G[240] = in[8] & in2[8];
    assign P[240] = in[8] ^ in2[8];
    assign G[241] = in[7] & in2[7];
    assign P[241] = in[7] ^ in2[7];
    assign G[242] = in[6] & in2[6];
    assign P[242] = in[6] ^ in2[6];
    assign G[243] = in[5] & in2[5];
    assign P[243] = in[5] ^ in2[5];
    assign G[244] = in[4] & in2[4];
    assign P[244] = in[4] ^ in2[4];
    assign G[245] = in[3] & in2[3];
    assign P[245] = in[3] ^ in2[3];
    assign G[246] = in[2] & in2[2];
    assign P[246] = in[2] ^ in2[2];
    assign G[247] = in[1] & in2[1];
    assign P[247] = in[1] ^ in2[1];
    assign G[248] = in[0] & in2[0];
    assign P[248] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign C[248] = G[247] | (P[247] & C[247]);
    assign cout = G[248] | (P[248] & C[248]);
    assign sum = P ^ C;
endmodule

module CLA248(output [247:0] sum, output cout, input [247:0] in1, input [247:0] in2;

    wire[247:0] G;
    wire[247:0] C;
    wire[247:0] P;

    assign G[0] = in[247] & in2[247];
    assign P[0] = in[247] ^ in2[247];
    assign G[1] = in[246] & in2[246];
    assign P[1] = in[246] ^ in2[246];
    assign G[2] = in[245] & in2[245];
    assign P[2] = in[245] ^ in2[245];
    assign G[3] = in[244] & in2[244];
    assign P[3] = in[244] ^ in2[244];
    assign G[4] = in[243] & in2[243];
    assign P[4] = in[243] ^ in2[243];
    assign G[5] = in[242] & in2[242];
    assign P[5] = in[242] ^ in2[242];
    assign G[6] = in[241] & in2[241];
    assign P[6] = in[241] ^ in2[241];
    assign G[7] = in[240] & in2[240];
    assign P[7] = in[240] ^ in2[240];
    assign G[8] = in[239] & in2[239];
    assign P[8] = in[239] ^ in2[239];
    assign G[9] = in[238] & in2[238];
    assign P[9] = in[238] ^ in2[238];
    assign G[10] = in[237] & in2[237];
    assign P[10] = in[237] ^ in2[237];
    assign G[11] = in[236] & in2[236];
    assign P[11] = in[236] ^ in2[236];
    assign G[12] = in[235] & in2[235];
    assign P[12] = in[235] ^ in2[235];
    assign G[13] = in[234] & in2[234];
    assign P[13] = in[234] ^ in2[234];
    assign G[14] = in[233] & in2[233];
    assign P[14] = in[233] ^ in2[233];
    assign G[15] = in[232] & in2[232];
    assign P[15] = in[232] ^ in2[232];
    assign G[16] = in[231] & in2[231];
    assign P[16] = in[231] ^ in2[231];
    assign G[17] = in[230] & in2[230];
    assign P[17] = in[230] ^ in2[230];
    assign G[18] = in[229] & in2[229];
    assign P[18] = in[229] ^ in2[229];
    assign G[19] = in[228] & in2[228];
    assign P[19] = in[228] ^ in2[228];
    assign G[20] = in[227] & in2[227];
    assign P[20] = in[227] ^ in2[227];
    assign G[21] = in[226] & in2[226];
    assign P[21] = in[226] ^ in2[226];
    assign G[22] = in[225] & in2[225];
    assign P[22] = in[225] ^ in2[225];
    assign G[23] = in[224] & in2[224];
    assign P[23] = in[224] ^ in2[224];
    assign G[24] = in[223] & in2[223];
    assign P[24] = in[223] ^ in2[223];
    assign G[25] = in[222] & in2[222];
    assign P[25] = in[222] ^ in2[222];
    assign G[26] = in[221] & in2[221];
    assign P[26] = in[221] ^ in2[221];
    assign G[27] = in[220] & in2[220];
    assign P[27] = in[220] ^ in2[220];
    assign G[28] = in[219] & in2[219];
    assign P[28] = in[219] ^ in2[219];
    assign G[29] = in[218] & in2[218];
    assign P[29] = in[218] ^ in2[218];
    assign G[30] = in[217] & in2[217];
    assign P[30] = in[217] ^ in2[217];
    assign G[31] = in[216] & in2[216];
    assign P[31] = in[216] ^ in2[216];
    assign G[32] = in[215] & in2[215];
    assign P[32] = in[215] ^ in2[215];
    assign G[33] = in[214] & in2[214];
    assign P[33] = in[214] ^ in2[214];
    assign G[34] = in[213] & in2[213];
    assign P[34] = in[213] ^ in2[213];
    assign G[35] = in[212] & in2[212];
    assign P[35] = in[212] ^ in2[212];
    assign G[36] = in[211] & in2[211];
    assign P[36] = in[211] ^ in2[211];
    assign G[37] = in[210] & in2[210];
    assign P[37] = in[210] ^ in2[210];
    assign G[38] = in[209] & in2[209];
    assign P[38] = in[209] ^ in2[209];
    assign G[39] = in[208] & in2[208];
    assign P[39] = in[208] ^ in2[208];
    assign G[40] = in[207] & in2[207];
    assign P[40] = in[207] ^ in2[207];
    assign G[41] = in[206] & in2[206];
    assign P[41] = in[206] ^ in2[206];
    assign G[42] = in[205] & in2[205];
    assign P[42] = in[205] ^ in2[205];
    assign G[43] = in[204] & in2[204];
    assign P[43] = in[204] ^ in2[204];
    assign G[44] = in[203] & in2[203];
    assign P[44] = in[203] ^ in2[203];
    assign G[45] = in[202] & in2[202];
    assign P[45] = in[202] ^ in2[202];
    assign G[46] = in[201] & in2[201];
    assign P[46] = in[201] ^ in2[201];
    assign G[47] = in[200] & in2[200];
    assign P[47] = in[200] ^ in2[200];
    assign G[48] = in[199] & in2[199];
    assign P[48] = in[199] ^ in2[199];
    assign G[49] = in[198] & in2[198];
    assign P[49] = in[198] ^ in2[198];
    assign G[50] = in[197] & in2[197];
    assign P[50] = in[197] ^ in2[197];
    assign G[51] = in[196] & in2[196];
    assign P[51] = in[196] ^ in2[196];
    assign G[52] = in[195] & in2[195];
    assign P[52] = in[195] ^ in2[195];
    assign G[53] = in[194] & in2[194];
    assign P[53] = in[194] ^ in2[194];
    assign G[54] = in[193] & in2[193];
    assign P[54] = in[193] ^ in2[193];
    assign G[55] = in[192] & in2[192];
    assign P[55] = in[192] ^ in2[192];
    assign G[56] = in[191] & in2[191];
    assign P[56] = in[191] ^ in2[191];
    assign G[57] = in[190] & in2[190];
    assign P[57] = in[190] ^ in2[190];
    assign G[58] = in[189] & in2[189];
    assign P[58] = in[189] ^ in2[189];
    assign G[59] = in[188] & in2[188];
    assign P[59] = in[188] ^ in2[188];
    assign G[60] = in[187] & in2[187];
    assign P[60] = in[187] ^ in2[187];
    assign G[61] = in[186] & in2[186];
    assign P[61] = in[186] ^ in2[186];
    assign G[62] = in[185] & in2[185];
    assign P[62] = in[185] ^ in2[185];
    assign G[63] = in[184] & in2[184];
    assign P[63] = in[184] ^ in2[184];
    assign G[64] = in[183] & in2[183];
    assign P[64] = in[183] ^ in2[183];
    assign G[65] = in[182] & in2[182];
    assign P[65] = in[182] ^ in2[182];
    assign G[66] = in[181] & in2[181];
    assign P[66] = in[181] ^ in2[181];
    assign G[67] = in[180] & in2[180];
    assign P[67] = in[180] ^ in2[180];
    assign G[68] = in[179] & in2[179];
    assign P[68] = in[179] ^ in2[179];
    assign G[69] = in[178] & in2[178];
    assign P[69] = in[178] ^ in2[178];
    assign G[70] = in[177] & in2[177];
    assign P[70] = in[177] ^ in2[177];
    assign G[71] = in[176] & in2[176];
    assign P[71] = in[176] ^ in2[176];
    assign G[72] = in[175] & in2[175];
    assign P[72] = in[175] ^ in2[175];
    assign G[73] = in[174] & in2[174];
    assign P[73] = in[174] ^ in2[174];
    assign G[74] = in[173] & in2[173];
    assign P[74] = in[173] ^ in2[173];
    assign G[75] = in[172] & in2[172];
    assign P[75] = in[172] ^ in2[172];
    assign G[76] = in[171] & in2[171];
    assign P[76] = in[171] ^ in2[171];
    assign G[77] = in[170] & in2[170];
    assign P[77] = in[170] ^ in2[170];
    assign G[78] = in[169] & in2[169];
    assign P[78] = in[169] ^ in2[169];
    assign G[79] = in[168] & in2[168];
    assign P[79] = in[168] ^ in2[168];
    assign G[80] = in[167] & in2[167];
    assign P[80] = in[167] ^ in2[167];
    assign G[81] = in[166] & in2[166];
    assign P[81] = in[166] ^ in2[166];
    assign G[82] = in[165] & in2[165];
    assign P[82] = in[165] ^ in2[165];
    assign G[83] = in[164] & in2[164];
    assign P[83] = in[164] ^ in2[164];
    assign G[84] = in[163] & in2[163];
    assign P[84] = in[163] ^ in2[163];
    assign G[85] = in[162] & in2[162];
    assign P[85] = in[162] ^ in2[162];
    assign G[86] = in[161] & in2[161];
    assign P[86] = in[161] ^ in2[161];
    assign G[87] = in[160] & in2[160];
    assign P[87] = in[160] ^ in2[160];
    assign G[88] = in[159] & in2[159];
    assign P[88] = in[159] ^ in2[159];
    assign G[89] = in[158] & in2[158];
    assign P[89] = in[158] ^ in2[158];
    assign G[90] = in[157] & in2[157];
    assign P[90] = in[157] ^ in2[157];
    assign G[91] = in[156] & in2[156];
    assign P[91] = in[156] ^ in2[156];
    assign G[92] = in[155] & in2[155];
    assign P[92] = in[155] ^ in2[155];
    assign G[93] = in[154] & in2[154];
    assign P[93] = in[154] ^ in2[154];
    assign G[94] = in[153] & in2[153];
    assign P[94] = in[153] ^ in2[153];
    assign G[95] = in[152] & in2[152];
    assign P[95] = in[152] ^ in2[152];
    assign G[96] = in[151] & in2[151];
    assign P[96] = in[151] ^ in2[151];
    assign G[97] = in[150] & in2[150];
    assign P[97] = in[150] ^ in2[150];
    assign G[98] = in[149] & in2[149];
    assign P[98] = in[149] ^ in2[149];
    assign G[99] = in[148] & in2[148];
    assign P[99] = in[148] ^ in2[148];
    assign G[100] = in[147] & in2[147];
    assign P[100] = in[147] ^ in2[147];
    assign G[101] = in[146] & in2[146];
    assign P[101] = in[146] ^ in2[146];
    assign G[102] = in[145] & in2[145];
    assign P[102] = in[145] ^ in2[145];
    assign G[103] = in[144] & in2[144];
    assign P[103] = in[144] ^ in2[144];
    assign G[104] = in[143] & in2[143];
    assign P[104] = in[143] ^ in2[143];
    assign G[105] = in[142] & in2[142];
    assign P[105] = in[142] ^ in2[142];
    assign G[106] = in[141] & in2[141];
    assign P[106] = in[141] ^ in2[141];
    assign G[107] = in[140] & in2[140];
    assign P[107] = in[140] ^ in2[140];
    assign G[108] = in[139] & in2[139];
    assign P[108] = in[139] ^ in2[139];
    assign G[109] = in[138] & in2[138];
    assign P[109] = in[138] ^ in2[138];
    assign G[110] = in[137] & in2[137];
    assign P[110] = in[137] ^ in2[137];
    assign G[111] = in[136] & in2[136];
    assign P[111] = in[136] ^ in2[136];
    assign G[112] = in[135] & in2[135];
    assign P[112] = in[135] ^ in2[135];
    assign G[113] = in[134] & in2[134];
    assign P[113] = in[134] ^ in2[134];
    assign G[114] = in[133] & in2[133];
    assign P[114] = in[133] ^ in2[133];
    assign G[115] = in[132] & in2[132];
    assign P[115] = in[132] ^ in2[132];
    assign G[116] = in[131] & in2[131];
    assign P[116] = in[131] ^ in2[131];
    assign G[117] = in[130] & in2[130];
    assign P[117] = in[130] ^ in2[130];
    assign G[118] = in[129] & in2[129];
    assign P[118] = in[129] ^ in2[129];
    assign G[119] = in[128] & in2[128];
    assign P[119] = in[128] ^ in2[128];
    assign G[120] = in[127] & in2[127];
    assign P[120] = in[127] ^ in2[127];
    assign G[121] = in[126] & in2[126];
    assign P[121] = in[126] ^ in2[126];
    assign G[122] = in[125] & in2[125];
    assign P[122] = in[125] ^ in2[125];
    assign G[123] = in[124] & in2[124];
    assign P[123] = in[124] ^ in2[124];
    assign G[124] = in[123] & in2[123];
    assign P[124] = in[123] ^ in2[123];
    assign G[125] = in[122] & in2[122];
    assign P[125] = in[122] ^ in2[122];
    assign G[126] = in[121] & in2[121];
    assign P[126] = in[121] ^ in2[121];
    assign G[127] = in[120] & in2[120];
    assign P[127] = in[120] ^ in2[120];
    assign G[128] = in[119] & in2[119];
    assign P[128] = in[119] ^ in2[119];
    assign G[129] = in[118] & in2[118];
    assign P[129] = in[118] ^ in2[118];
    assign G[130] = in[117] & in2[117];
    assign P[130] = in[117] ^ in2[117];
    assign G[131] = in[116] & in2[116];
    assign P[131] = in[116] ^ in2[116];
    assign G[132] = in[115] & in2[115];
    assign P[132] = in[115] ^ in2[115];
    assign G[133] = in[114] & in2[114];
    assign P[133] = in[114] ^ in2[114];
    assign G[134] = in[113] & in2[113];
    assign P[134] = in[113] ^ in2[113];
    assign G[135] = in[112] & in2[112];
    assign P[135] = in[112] ^ in2[112];
    assign G[136] = in[111] & in2[111];
    assign P[136] = in[111] ^ in2[111];
    assign G[137] = in[110] & in2[110];
    assign P[137] = in[110] ^ in2[110];
    assign G[138] = in[109] & in2[109];
    assign P[138] = in[109] ^ in2[109];
    assign G[139] = in[108] & in2[108];
    assign P[139] = in[108] ^ in2[108];
    assign G[140] = in[107] & in2[107];
    assign P[140] = in[107] ^ in2[107];
    assign G[141] = in[106] & in2[106];
    assign P[141] = in[106] ^ in2[106];
    assign G[142] = in[105] & in2[105];
    assign P[142] = in[105] ^ in2[105];
    assign G[143] = in[104] & in2[104];
    assign P[143] = in[104] ^ in2[104];
    assign G[144] = in[103] & in2[103];
    assign P[144] = in[103] ^ in2[103];
    assign G[145] = in[102] & in2[102];
    assign P[145] = in[102] ^ in2[102];
    assign G[146] = in[101] & in2[101];
    assign P[146] = in[101] ^ in2[101];
    assign G[147] = in[100] & in2[100];
    assign P[147] = in[100] ^ in2[100];
    assign G[148] = in[99] & in2[99];
    assign P[148] = in[99] ^ in2[99];
    assign G[149] = in[98] & in2[98];
    assign P[149] = in[98] ^ in2[98];
    assign G[150] = in[97] & in2[97];
    assign P[150] = in[97] ^ in2[97];
    assign G[151] = in[96] & in2[96];
    assign P[151] = in[96] ^ in2[96];
    assign G[152] = in[95] & in2[95];
    assign P[152] = in[95] ^ in2[95];
    assign G[153] = in[94] & in2[94];
    assign P[153] = in[94] ^ in2[94];
    assign G[154] = in[93] & in2[93];
    assign P[154] = in[93] ^ in2[93];
    assign G[155] = in[92] & in2[92];
    assign P[155] = in[92] ^ in2[92];
    assign G[156] = in[91] & in2[91];
    assign P[156] = in[91] ^ in2[91];
    assign G[157] = in[90] & in2[90];
    assign P[157] = in[90] ^ in2[90];
    assign G[158] = in[89] & in2[89];
    assign P[158] = in[89] ^ in2[89];
    assign G[159] = in[88] & in2[88];
    assign P[159] = in[88] ^ in2[88];
    assign G[160] = in[87] & in2[87];
    assign P[160] = in[87] ^ in2[87];
    assign G[161] = in[86] & in2[86];
    assign P[161] = in[86] ^ in2[86];
    assign G[162] = in[85] & in2[85];
    assign P[162] = in[85] ^ in2[85];
    assign G[163] = in[84] & in2[84];
    assign P[163] = in[84] ^ in2[84];
    assign G[164] = in[83] & in2[83];
    assign P[164] = in[83] ^ in2[83];
    assign G[165] = in[82] & in2[82];
    assign P[165] = in[82] ^ in2[82];
    assign G[166] = in[81] & in2[81];
    assign P[166] = in[81] ^ in2[81];
    assign G[167] = in[80] & in2[80];
    assign P[167] = in[80] ^ in2[80];
    assign G[168] = in[79] & in2[79];
    assign P[168] = in[79] ^ in2[79];
    assign G[169] = in[78] & in2[78];
    assign P[169] = in[78] ^ in2[78];
    assign G[170] = in[77] & in2[77];
    assign P[170] = in[77] ^ in2[77];
    assign G[171] = in[76] & in2[76];
    assign P[171] = in[76] ^ in2[76];
    assign G[172] = in[75] & in2[75];
    assign P[172] = in[75] ^ in2[75];
    assign G[173] = in[74] & in2[74];
    assign P[173] = in[74] ^ in2[74];
    assign G[174] = in[73] & in2[73];
    assign P[174] = in[73] ^ in2[73];
    assign G[175] = in[72] & in2[72];
    assign P[175] = in[72] ^ in2[72];
    assign G[176] = in[71] & in2[71];
    assign P[176] = in[71] ^ in2[71];
    assign G[177] = in[70] & in2[70];
    assign P[177] = in[70] ^ in2[70];
    assign G[178] = in[69] & in2[69];
    assign P[178] = in[69] ^ in2[69];
    assign G[179] = in[68] & in2[68];
    assign P[179] = in[68] ^ in2[68];
    assign G[180] = in[67] & in2[67];
    assign P[180] = in[67] ^ in2[67];
    assign G[181] = in[66] & in2[66];
    assign P[181] = in[66] ^ in2[66];
    assign G[182] = in[65] & in2[65];
    assign P[182] = in[65] ^ in2[65];
    assign G[183] = in[64] & in2[64];
    assign P[183] = in[64] ^ in2[64];
    assign G[184] = in[63] & in2[63];
    assign P[184] = in[63] ^ in2[63];
    assign G[185] = in[62] & in2[62];
    assign P[185] = in[62] ^ in2[62];
    assign G[186] = in[61] & in2[61];
    assign P[186] = in[61] ^ in2[61];
    assign G[187] = in[60] & in2[60];
    assign P[187] = in[60] ^ in2[60];
    assign G[188] = in[59] & in2[59];
    assign P[188] = in[59] ^ in2[59];
    assign G[189] = in[58] & in2[58];
    assign P[189] = in[58] ^ in2[58];
    assign G[190] = in[57] & in2[57];
    assign P[190] = in[57] ^ in2[57];
    assign G[191] = in[56] & in2[56];
    assign P[191] = in[56] ^ in2[56];
    assign G[192] = in[55] & in2[55];
    assign P[192] = in[55] ^ in2[55];
    assign G[193] = in[54] & in2[54];
    assign P[193] = in[54] ^ in2[54];
    assign G[194] = in[53] & in2[53];
    assign P[194] = in[53] ^ in2[53];
    assign G[195] = in[52] & in2[52];
    assign P[195] = in[52] ^ in2[52];
    assign G[196] = in[51] & in2[51];
    assign P[196] = in[51] ^ in2[51];
    assign G[197] = in[50] & in2[50];
    assign P[197] = in[50] ^ in2[50];
    assign G[198] = in[49] & in2[49];
    assign P[198] = in[49] ^ in2[49];
    assign G[199] = in[48] & in2[48];
    assign P[199] = in[48] ^ in2[48];
    assign G[200] = in[47] & in2[47];
    assign P[200] = in[47] ^ in2[47];
    assign G[201] = in[46] & in2[46];
    assign P[201] = in[46] ^ in2[46];
    assign G[202] = in[45] & in2[45];
    assign P[202] = in[45] ^ in2[45];
    assign G[203] = in[44] & in2[44];
    assign P[203] = in[44] ^ in2[44];
    assign G[204] = in[43] & in2[43];
    assign P[204] = in[43] ^ in2[43];
    assign G[205] = in[42] & in2[42];
    assign P[205] = in[42] ^ in2[42];
    assign G[206] = in[41] & in2[41];
    assign P[206] = in[41] ^ in2[41];
    assign G[207] = in[40] & in2[40];
    assign P[207] = in[40] ^ in2[40];
    assign G[208] = in[39] & in2[39];
    assign P[208] = in[39] ^ in2[39];
    assign G[209] = in[38] & in2[38];
    assign P[209] = in[38] ^ in2[38];
    assign G[210] = in[37] & in2[37];
    assign P[210] = in[37] ^ in2[37];
    assign G[211] = in[36] & in2[36];
    assign P[211] = in[36] ^ in2[36];
    assign G[212] = in[35] & in2[35];
    assign P[212] = in[35] ^ in2[35];
    assign G[213] = in[34] & in2[34];
    assign P[213] = in[34] ^ in2[34];
    assign G[214] = in[33] & in2[33];
    assign P[214] = in[33] ^ in2[33];
    assign G[215] = in[32] & in2[32];
    assign P[215] = in[32] ^ in2[32];
    assign G[216] = in[31] & in2[31];
    assign P[216] = in[31] ^ in2[31];
    assign G[217] = in[30] & in2[30];
    assign P[217] = in[30] ^ in2[30];
    assign G[218] = in[29] & in2[29];
    assign P[218] = in[29] ^ in2[29];
    assign G[219] = in[28] & in2[28];
    assign P[219] = in[28] ^ in2[28];
    assign G[220] = in[27] & in2[27];
    assign P[220] = in[27] ^ in2[27];
    assign G[221] = in[26] & in2[26];
    assign P[221] = in[26] ^ in2[26];
    assign G[222] = in[25] & in2[25];
    assign P[222] = in[25] ^ in2[25];
    assign G[223] = in[24] & in2[24];
    assign P[223] = in[24] ^ in2[24];
    assign G[224] = in[23] & in2[23];
    assign P[224] = in[23] ^ in2[23];
    assign G[225] = in[22] & in2[22];
    assign P[225] = in[22] ^ in2[22];
    assign G[226] = in[21] & in2[21];
    assign P[226] = in[21] ^ in2[21];
    assign G[227] = in[20] & in2[20];
    assign P[227] = in[20] ^ in2[20];
    assign G[228] = in[19] & in2[19];
    assign P[228] = in[19] ^ in2[19];
    assign G[229] = in[18] & in2[18];
    assign P[229] = in[18] ^ in2[18];
    assign G[230] = in[17] & in2[17];
    assign P[230] = in[17] ^ in2[17];
    assign G[231] = in[16] & in2[16];
    assign P[231] = in[16] ^ in2[16];
    assign G[232] = in[15] & in2[15];
    assign P[232] = in[15] ^ in2[15];
    assign G[233] = in[14] & in2[14];
    assign P[233] = in[14] ^ in2[14];
    assign G[234] = in[13] & in2[13];
    assign P[234] = in[13] ^ in2[13];
    assign G[235] = in[12] & in2[12];
    assign P[235] = in[12] ^ in2[12];
    assign G[236] = in[11] & in2[11];
    assign P[236] = in[11] ^ in2[11];
    assign G[237] = in[10] & in2[10];
    assign P[237] = in[10] ^ in2[10];
    assign G[238] = in[9] & in2[9];
    assign P[238] = in[9] ^ in2[9];
    assign G[239] = in[8] & in2[8];
    assign P[239] = in[8] ^ in2[8];
    assign G[240] = in[7] & in2[7];
    assign P[240] = in[7] ^ in2[7];
    assign G[241] = in[6] & in2[6];
    assign P[241] = in[6] ^ in2[6];
    assign G[242] = in[5] & in2[5];
    assign P[242] = in[5] ^ in2[5];
    assign G[243] = in[4] & in2[4];
    assign P[243] = in[4] ^ in2[4];
    assign G[244] = in[3] & in2[3];
    assign P[244] = in[3] ^ in2[3];
    assign G[245] = in[2] & in2[2];
    assign P[245] = in[2] ^ in2[2];
    assign G[246] = in[1] & in2[1];
    assign P[246] = in[1] ^ in2[1];
    assign G[247] = in[0] & in2[0];
    assign P[247] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign C[247] = G[246] | (P[246] & C[246]);
    assign cout = G[247] | (P[247] & C[247]);
    assign sum = P ^ C;
endmodule

module CLA247(output [246:0] sum, output cout, input [246:0] in1, input [246:0] in2;

    wire[246:0] G;
    wire[246:0] C;
    wire[246:0] P;

    assign G[0] = in[246] & in2[246];
    assign P[0] = in[246] ^ in2[246];
    assign G[1] = in[245] & in2[245];
    assign P[1] = in[245] ^ in2[245];
    assign G[2] = in[244] & in2[244];
    assign P[2] = in[244] ^ in2[244];
    assign G[3] = in[243] & in2[243];
    assign P[3] = in[243] ^ in2[243];
    assign G[4] = in[242] & in2[242];
    assign P[4] = in[242] ^ in2[242];
    assign G[5] = in[241] & in2[241];
    assign P[5] = in[241] ^ in2[241];
    assign G[6] = in[240] & in2[240];
    assign P[6] = in[240] ^ in2[240];
    assign G[7] = in[239] & in2[239];
    assign P[7] = in[239] ^ in2[239];
    assign G[8] = in[238] & in2[238];
    assign P[8] = in[238] ^ in2[238];
    assign G[9] = in[237] & in2[237];
    assign P[9] = in[237] ^ in2[237];
    assign G[10] = in[236] & in2[236];
    assign P[10] = in[236] ^ in2[236];
    assign G[11] = in[235] & in2[235];
    assign P[11] = in[235] ^ in2[235];
    assign G[12] = in[234] & in2[234];
    assign P[12] = in[234] ^ in2[234];
    assign G[13] = in[233] & in2[233];
    assign P[13] = in[233] ^ in2[233];
    assign G[14] = in[232] & in2[232];
    assign P[14] = in[232] ^ in2[232];
    assign G[15] = in[231] & in2[231];
    assign P[15] = in[231] ^ in2[231];
    assign G[16] = in[230] & in2[230];
    assign P[16] = in[230] ^ in2[230];
    assign G[17] = in[229] & in2[229];
    assign P[17] = in[229] ^ in2[229];
    assign G[18] = in[228] & in2[228];
    assign P[18] = in[228] ^ in2[228];
    assign G[19] = in[227] & in2[227];
    assign P[19] = in[227] ^ in2[227];
    assign G[20] = in[226] & in2[226];
    assign P[20] = in[226] ^ in2[226];
    assign G[21] = in[225] & in2[225];
    assign P[21] = in[225] ^ in2[225];
    assign G[22] = in[224] & in2[224];
    assign P[22] = in[224] ^ in2[224];
    assign G[23] = in[223] & in2[223];
    assign P[23] = in[223] ^ in2[223];
    assign G[24] = in[222] & in2[222];
    assign P[24] = in[222] ^ in2[222];
    assign G[25] = in[221] & in2[221];
    assign P[25] = in[221] ^ in2[221];
    assign G[26] = in[220] & in2[220];
    assign P[26] = in[220] ^ in2[220];
    assign G[27] = in[219] & in2[219];
    assign P[27] = in[219] ^ in2[219];
    assign G[28] = in[218] & in2[218];
    assign P[28] = in[218] ^ in2[218];
    assign G[29] = in[217] & in2[217];
    assign P[29] = in[217] ^ in2[217];
    assign G[30] = in[216] & in2[216];
    assign P[30] = in[216] ^ in2[216];
    assign G[31] = in[215] & in2[215];
    assign P[31] = in[215] ^ in2[215];
    assign G[32] = in[214] & in2[214];
    assign P[32] = in[214] ^ in2[214];
    assign G[33] = in[213] & in2[213];
    assign P[33] = in[213] ^ in2[213];
    assign G[34] = in[212] & in2[212];
    assign P[34] = in[212] ^ in2[212];
    assign G[35] = in[211] & in2[211];
    assign P[35] = in[211] ^ in2[211];
    assign G[36] = in[210] & in2[210];
    assign P[36] = in[210] ^ in2[210];
    assign G[37] = in[209] & in2[209];
    assign P[37] = in[209] ^ in2[209];
    assign G[38] = in[208] & in2[208];
    assign P[38] = in[208] ^ in2[208];
    assign G[39] = in[207] & in2[207];
    assign P[39] = in[207] ^ in2[207];
    assign G[40] = in[206] & in2[206];
    assign P[40] = in[206] ^ in2[206];
    assign G[41] = in[205] & in2[205];
    assign P[41] = in[205] ^ in2[205];
    assign G[42] = in[204] & in2[204];
    assign P[42] = in[204] ^ in2[204];
    assign G[43] = in[203] & in2[203];
    assign P[43] = in[203] ^ in2[203];
    assign G[44] = in[202] & in2[202];
    assign P[44] = in[202] ^ in2[202];
    assign G[45] = in[201] & in2[201];
    assign P[45] = in[201] ^ in2[201];
    assign G[46] = in[200] & in2[200];
    assign P[46] = in[200] ^ in2[200];
    assign G[47] = in[199] & in2[199];
    assign P[47] = in[199] ^ in2[199];
    assign G[48] = in[198] & in2[198];
    assign P[48] = in[198] ^ in2[198];
    assign G[49] = in[197] & in2[197];
    assign P[49] = in[197] ^ in2[197];
    assign G[50] = in[196] & in2[196];
    assign P[50] = in[196] ^ in2[196];
    assign G[51] = in[195] & in2[195];
    assign P[51] = in[195] ^ in2[195];
    assign G[52] = in[194] & in2[194];
    assign P[52] = in[194] ^ in2[194];
    assign G[53] = in[193] & in2[193];
    assign P[53] = in[193] ^ in2[193];
    assign G[54] = in[192] & in2[192];
    assign P[54] = in[192] ^ in2[192];
    assign G[55] = in[191] & in2[191];
    assign P[55] = in[191] ^ in2[191];
    assign G[56] = in[190] & in2[190];
    assign P[56] = in[190] ^ in2[190];
    assign G[57] = in[189] & in2[189];
    assign P[57] = in[189] ^ in2[189];
    assign G[58] = in[188] & in2[188];
    assign P[58] = in[188] ^ in2[188];
    assign G[59] = in[187] & in2[187];
    assign P[59] = in[187] ^ in2[187];
    assign G[60] = in[186] & in2[186];
    assign P[60] = in[186] ^ in2[186];
    assign G[61] = in[185] & in2[185];
    assign P[61] = in[185] ^ in2[185];
    assign G[62] = in[184] & in2[184];
    assign P[62] = in[184] ^ in2[184];
    assign G[63] = in[183] & in2[183];
    assign P[63] = in[183] ^ in2[183];
    assign G[64] = in[182] & in2[182];
    assign P[64] = in[182] ^ in2[182];
    assign G[65] = in[181] & in2[181];
    assign P[65] = in[181] ^ in2[181];
    assign G[66] = in[180] & in2[180];
    assign P[66] = in[180] ^ in2[180];
    assign G[67] = in[179] & in2[179];
    assign P[67] = in[179] ^ in2[179];
    assign G[68] = in[178] & in2[178];
    assign P[68] = in[178] ^ in2[178];
    assign G[69] = in[177] & in2[177];
    assign P[69] = in[177] ^ in2[177];
    assign G[70] = in[176] & in2[176];
    assign P[70] = in[176] ^ in2[176];
    assign G[71] = in[175] & in2[175];
    assign P[71] = in[175] ^ in2[175];
    assign G[72] = in[174] & in2[174];
    assign P[72] = in[174] ^ in2[174];
    assign G[73] = in[173] & in2[173];
    assign P[73] = in[173] ^ in2[173];
    assign G[74] = in[172] & in2[172];
    assign P[74] = in[172] ^ in2[172];
    assign G[75] = in[171] & in2[171];
    assign P[75] = in[171] ^ in2[171];
    assign G[76] = in[170] & in2[170];
    assign P[76] = in[170] ^ in2[170];
    assign G[77] = in[169] & in2[169];
    assign P[77] = in[169] ^ in2[169];
    assign G[78] = in[168] & in2[168];
    assign P[78] = in[168] ^ in2[168];
    assign G[79] = in[167] & in2[167];
    assign P[79] = in[167] ^ in2[167];
    assign G[80] = in[166] & in2[166];
    assign P[80] = in[166] ^ in2[166];
    assign G[81] = in[165] & in2[165];
    assign P[81] = in[165] ^ in2[165];
    assign G[82] = in[164] & in2[164];
    assign P[82] = in[164] ^ in2[164];
    assign G[83] = in[163] & in2[163];
    assign P[83] = in[163] ^ in2[163];
    assign G[84] = in[162] & in2[162];
    assign P[84] = in[162] ^ in2[162];
    assign G[85] = in[161] & in2[161];
    assign P[85] = in[161] ^ in2[161];
    assign G[86] = in[160] & in2[160];
    assign P[86] = in[160] ^ in2[160];
    assign G[87] = in[159] & in2[159];
    assign P[87] = in[159] ^ in2[159];
    assign G[88] = in[158] & in2[158];
    assign P[88] = in[158] ^ in2[158];
    assign G[89] = in[157] & in2[157];
    assign P[89] = in[157] ^ in2[157];
    assign G[90] = in[156] & in2[156];
    assign P[90] = in[156] ^ in2[156];
    assign G[91] = in[155] & in2[155];
    assign P[91] = in[155] ^ in2[155];
    assign G[92] = in[154] & in2[154];
    assign P[92] = in[154] ^ in2[154];
    assign G[93] = in[153] & in2[153];
    assign P[93] = in[153] ^ in2[153];
    assign G[94] = in[152] & in2[152];
    assign P[94] = in[152] ^ in2[152];
    assign G[95] = in[151] & in2[151];
    assign P[95] = in[151] ^ in2[151];
    assign G[96] = in[150] & in2[150];
    assign P[96] = in[150] ^ in2[150];
    assign G[97] = in[149] & in2[149];
    assign P[97] = in[149] ^ in2[149];
    assign G[98] = in[148] & in2[148];
    assign P[98] = in[148] ^ in2[148];
    assign G[99] = in[147] & in2[147];
    assign P[99] = in[147] ^ in2[147];
    assign G[100] = in[146] & in2[146];
    assign P[100] = in[146] ^ in2[146];
    assign G[101] = in[145] & in2[145];
    assign P[101] = in[145] ^ in2[145];
    assign G[102] = in[144] & in2[144];
    assign P[102] = in[144] ^ in2[144];
    assign G[103] = in[143] & in2[143];
    assign P[103] = in[143] ^ in2[143];
    assign G[104] = in[142] & in2[142];
    assign P[104] = in[142] ^ in2[142];
    assign G[105] = in[141] & in2[141];
    assign P[105] = in[141] ^ in2[141];
    assign G[106] = in[140] & in2[140];
    assign P[106] = in[140] ^ in2[140];
    assign G[107] = in[139] & in2[139];
    assign P[107] = in[139] ^ in2[139];
    assign G[108] = in[138] & in2[138];
    assign P[108] = in[138] ^ in2[138];
    assign G[109] = in[137] & in2[137];
    assign P[109] = in[137] ^ in2[137];
    assign G[110] = in[136] & in2[136];
    assign P[110] = in[136] ^ in2[136];
    assign G[111] = in[135] & in2[135];
    assign P[111] = in[135] ^ in2[135];
    assign G[112] = in[134] & in2[134];
    assign P[112] = in[134] ^ in2[134];
    assign G[113] = in[133] & in2[133];
    assign P[113] = in[133] ^ in2[133];
    assign G[114] = in[132] & in2[132];
    assign P[114] = in[132] ^ in2[132];
    assign G[115] = in[131] & in2[131];
    assign P[115] = in[131] ^ in2[131];
    assign G[116] = in[130] & in2[130];
    assign P[116] = in[130] ^ in2[130];
    assign G[117] = in[129] & in2[129];
    assign P[117] = in[129] ^ in2[129];
    assign G[118] = in[128] & in2[128];
    assign P[118] = in[128] ^ in2[128];
    assign G[119] = in[127] & in2[127];
    assign P[119] = in[127] ^ in2[127];
    assign G[120] = in[126] & in2[126];
    assign P[120] = in[126] ^ in2[126];
    assign G[121] = in[125] & in2[125];
    assign P[121] = in[125] ^ in2[125];
    assign G[122] = in[124] & in2[124];
    assign P[122] = in[124] ^ in2[124];
    assign G[123] = in[123] & in2[123];
    assign P[123] = in[123] ^ in2[123];
    assign G[124] = in[122] & in2[122];
    assign P[124] = in[122] ^ in2[122];
    assign G[125] = in[121] & in2[121];
    assign P[125] = in[121] ^ in2[121];
    assign G[126] = in[120] & in2[120];
    assign P[126] = in[120] ^ in2[120];
    assign G[127] = in[119] & in2[119];
    assign P[127] = in[119] ^ in2[119];
    assign G[128] = in[118] & in2[118];
    assign P[128] = in[118] ^ in2[118];
    assign G[129] = in[117] & in2[117];
    assign P[129] = in[117] ^ in2[117];
    assign G[130] = in[116] & in2[116];
    assign P[130] = in[116] ^ in2[116];
    assign G[131] = in[115] & in2[115];
    assign P[131] = in[115] ^ in2[115];
    assign G[132] = in[114] & in2[114];
    assign P[132] = in[114] ^ in2[114];
    assign G[133] = in[113] & in2[113];
    assign P[133] = in[113] ^ in2[113];
    assign G[134] = in[112] & in2[112];
    assign P[134] = in[112] ^ in2[112];
    assign G[135] = in[111] & in2[111];
    assign P[135] = in[111] ^ in2[111];
    assign G[136] = in[110] & in2[110];
    assign P[136] = in[110] ^ in2[110];
    assign G[137] = in[109] & in2[109];
    assign P[137] = in[109] ^ in2[109];
    assign G[138] = in[108] & in2[108];
    assign P[138] = in[108] ^ in2[108];
    assign G[139] = in[107] & in2[107];
    assign P[139] = in[107] ^ in2[107];
    assign G[140] = in[106] & in2[106];
    assign P[140] = in[106] ^ in2[106];
    assign G[141] = in[105] & in2[105];
    assign P[141] = in[105] ^ in2[105];
    assign G[142] = in[104] & in2[104];
    assign P[142] = in[104] ^ in2[104];
    assign G[143] = in[103] & in2[103];
    assign P[143] = in[103] ^ in2[103];
    assign G[144] = in[102] & in2[102];
    assign P[144] = in[102] ^ in2[102];
    assign G[145] = in[101] & in2[101];
    assign P[145] = in[101] ^ in2[101];
    assign G[146] = in[100] & in2[100];
    assign P[146] = in[100] ^ in2[100];
    assign G[147] = in[99] & in2[99];
    assign P[147] = in[99] ^ in2[99];
    assign G[148] = in[98] & in2[98];
    assign P[148] = in[98] ^ in2[98];
    assign G[149] = in[97] & in2[97];
    assign P[149] = in[97] ^ in2[97];
    assign G[150] = in[96] & in2[96];
    assign P[150] = in[96] ^ in2[96];
    assign G[151] = in[95] & in2[95];
    assign P[151] = in[95] ^ in2[95];
    assign G[152] = in[94] & in2[94];
    assign P[152] = in[94] ^ in2[94];
    assign G[153] = in[93] & in2[93];
    assign P[153] = in[93] ^ in2[93];
    assign G[154] = in[92] & in2[92];
    assign P[154] = in[92] ^ in2[92];
    assign G[155] = in[91] & in2[91];
    assign P[155] = in[91] ^ in2[91];
    assign G[156] = in[90] & in2[90];
    assign P[156] = in[90] ^ in2[90];
    assign G[157] = in[89] & in2[89];
    assign P[157] = in[89] ^ in2[89];
    assign G[158] = in[88] & in2[88];
    assign P[158] = in[88] ^ in2[88];
    assign G[159] = in[87] & in2[87];
    assign P[159] = in[87] ^ in2[87];
    assign G[160] = in[86] & in2[86];
    assign P[160] = in[86] ^ in2[86];
    assign G[161] = in[85] & in2[85];
    assign P[161] = in[85] ^ in2[85];
    assign G[162] = in[84] & in2[84];
    assign P[162] = in[84] ^ in2[84];
    assign G[163] = in[83] & in2[83];
    assign P[163] = in[83] ^ in2[83];
    assign G[164] = in[82] & in2[82];
    assign P[164] = in[82] ^ in2[82];
    assign G[165] = in[81] & in2[81];
    assign P[165] = in[81] ^ in2[81];
    assign G[166] = in[80] & in2[80];
    assign P[166] = in[80] ^ in2[80];
    assign G[167] = in[79] & in2[79];
    assign P[167] = in[79] ^ in2[79];
    assign G[168] = in[78] & in2[78];
    assign P[168] = in[78] ^ in2[78];
    assign G[169] = in[77] & in2[77];
    assign P[169] = in[77] ^ in2[77];
    assign G[170] = in[76] & in2[76];
    assign P[170] = in[76] ^ in2[76];
    assign G[171] = in[75] & in2[75];
    assign P[171] = in[75] ^ in2[75];
    assign G[172] = in[74] & in2[74];
    assign P[172] = in[74] ^ in2[74];
    assign G[173] = in[73] & in2[73];
    assign P[173] = in[73] ^ in2[73];
    assign G[174] = in[72] & in2[72];
    assign P[174] = in[72] ^ in2[72];
    assign G[175] = in[71] & in2[71];
    assign P[175] = in[71] ^ in2[71];
    assign G[176] = in[70] & in2[70];
    assign P[176] = in[70] ^ in2[70];
    assign G[177] = in[69] & in2[69];
    assign P[177] = in[69] ^ in2[69];
    assign G[178] = in[68] & in2[68];
    assign P[178] = in[68] ^ in2[68];
    assign G[179] = in[67] & in2[67];
    assign P[179] = in[67] ^ in2[67];
    assign G[180] = in[66] & in2[66];
    assign P[180] = in[66] ^ in2[66];
    assign G[181] = in[65] & in2[65];
    assign P[181] = in[65] ^ in2[65];
    assign G[182] = in[64] & in2[64];
    assign P[182] = in[64] ^ in2[64];
    assign G[183] = in[63] & in2[63];
    assign P[183] = in[63] ^ in2[63];
    assign G[184] = in[62] & in2[62];
    assign P[184] = in[62] ^ in2[62];
    assign G[185] = in[61] & in2[61];
    assign P[185] = in[61] ^ in2[61];
    assign G[186] = in[60] & in2[60];
    assign P[186] = in[60] ^ in2[60];
    assign G[187] = in[59] & in2[59];
    assign P[187] = in[59] ^ in2[59];
    assign G[188] = in[58] & in2[58];
    assign P[188] = in[58] ^ in2[58];
    assign G[189] = in[57] & in2[57];
    assign P[189] = in[57] ^ in2[57];
    assign G[190] = in[56] & in2[56];
    assign P[190] = in[56] ^ in2[56];
    assign G[191] = in[55] & in2[55];
    assign P[191] = in[55] ^ in2[55];
    assign G[192] = in[54] & in2[54];
    assign P[192] = in[54] ^ in2[54];
    assign G[193] = in[53] & in2[53];
    assign P[193] = in[53] ^ in2[53];
    assign G[194] = in[52] & in2[52];
    assign P[194] = in[52] ^ in2[52];
    assign G[195] = in[51] & in2[51];
    assign P[195] = in[51] ^ in2[51];
    assign G[196] = in[50] & in2[50];
    assign P[196] = in[50] ^ in2[50];
    assign G[197] = in[49] & in2[49];
    assign P[197] = in[49] ^ in2[49];
    assign G[198] = in[48] & in2[48];
    assign P[198] = in[48] ^ in2[48];
    assign G[199] = in[47] & in2[47];
    assign P[199] = in[47] ^ in2[47];
    assign G[200] = in[46] & in2[46];
    assign P[200] = in[46] ^ in2[46];
    assign G[201] = in[45] & in2[45];
    assign P[201] = in[45] ^ in2[45];
    assign G[202] = in[44] & in2[44];
    assign P[202] = in[44] ^ in2[44];
    assign G[203] = in[43] & in2[43];
    assign P[203] = in[43] ^ in2[43];
    assign G[204] = in[42] & in2[42];
    assign P[204] = in[42] ^ in2[42];
    assign G[205] = in[41] & in2[41];
    assign P[205] = in[41] ^ in2[41];
    assign G[206] = in[40] & in2[40];
    assign P[206] = in[40] ^ in2[40];
    assign G[207] = in[39] & in2[39];
    assign P[207] = in[39] ^ in2[39];
    assign G[208] = in[38] & in2[38];
    assign P[208] = in[38] ^ in2[38];
    assign G[209] = in[37] & in2[37];
    assign P[209] = in[37] ^ in2[37];
    assign G[210] = in[36] & in2[36];
    assign P[210] = in[36] ^ in2[36];
    assign G[211] = in[35] & in2[35];
    assign P[211] = in[35] ^ in2[35];
    assign G[212] = in[34] & in2[34];
    assign P[212] = in[34] ^ in2[34];
    assign G[213] = in[33] & in2[33];
    assign P[213] = in[33] ^ in2[33];
    assign G[214] = in[32] & in2[32];
    assign P[214] = in[32] ^ in2[32];
    assign G[215] = in[31] & in2[31];
    assign P[215] = in[31] ^ in2[31];
    assign G[216] = in[30] & in2[30];
    assign P[216] = in[30] ^ in2[30];
    assign G[217] = in[29] & in2[29];
    assign P[217] = in[29] ^ in2[29];
    assign G[218] = in[28] & in2[28];
    assign P[218] = in[28] ^ in2[28];
    assign G[219] = in[27] & in2[27];
    assign P[219] = in[27] ^ in2[27];
    assign G[220] = in[26] & in2[26];
    assign P[220] = in[26] ^ in2[26];
    assign G[221] = in[25] & in2[25];
    assign P[221] = in[25] ^ in2[25];
    assign G[222] = in[24] & in2[24];
    assign P[222] = in[24] ^ in2[24];
    assign G[223] = in[23] & in2[23];
    assign P[223] = in[23] ^ in2[23];
    assign G[224] = in[22] & in2[22];
    assign P[224] = in[22] ^ in2[22];
    assign G[225] = in[21] & in2[21];
    assign P[225] = in[21] ^ in2[21];
    assign G[226] = in[20] & in2[20];
    assign P[226] = in[20] ^ in2[20];
    assign G[227] = in[19] & in2[19];
    assign P[227] = in[19] ^ in2[19];
    assign G[228] = in[18] & in2[18];
    assign P[228] = in[18] ^ in2[18];
    assign G[229] = in[17] & in2[17];
    assign P[229] = in[17] ^ in2[17];
    assign G[230] = in[16] & in2[16];
    assign P[230] = in[16] ^ in2[16];
    assign G[231] = in[15] & in2[15];
    assign P[231] = in[15] ^ in2[15];
    assign G[232] = in[14] & in2[14];
    assign P[232] = in[14] ^ in2[14];
    assign G[233] = in[13] & in2[13];
    assign P[233] = in[13] ^ in2[13];
    assign G[234] = in[12] & in2[12];
    assign P[234] = in[12] ^ in2[12];
    assign G[235] = in[11] & in2[11];
    assign P[235] = in[11] ^ in2[11];
    assign G[236] = in[10] & in2[10];
    assign P[236] = in[10] ^ in2[10];
    assign G[237] = in[9] & in2[9];
    assign P[237] = in[9] ^ in2[9];
    assign G[238] = in[8] & in2[8];
    assign P[238] = in[8] ^ in2[8];
    assign G[239] = in[7] & in2[7];
    assign P[239] = in[7] ^ in2[7];
    assign G[240] = in[6] & in2[6];
    assign P[240] = in[6] ^ in2[6];
    assign G[241] = in[5] & in2[5];
    assign P[241] = in[5] ^ in2[5];
    assign G[242] = in[4] & in2[4];
    assign P[242] = in[4] ^ in2[4];
    assign G[243] = in[3] & in2[3];
    assign P[243] = in[3] ^ in2[3];
    assign G[244] = in[2] & in2[2];
    assign P[244] = in[2] ^ in2[2];
    assign G[245] = in[1] & in2[1];
    assign P[245] = in[1] ^ in2[1];
    assign G[246] = in[0] & in2[0];
    assign P[246] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign C[246] = G[245] | (P[245] & C[245]);
    assign cout = G[246] | (P[246] & C[246]);
    assign sum = P ^ C;
endmodule

module CLA246(output [245:0] sum, output cout, input [245:0] in1, input [245:0] in2;

    wire[245:0] G;
    wire[245:0] C;
    wire[245:0] P;

    assign G[0] = in[245] & in2[245];
    assign P[0] = in[245] ^ in2[245];
    assign G[1] = in[244] & in2[244];
    assign P[1] = in[244] ^ in2[244];
    assign G[2] = in[243] & in2[243];
    assign P[2] = in[243] ^ in2[243];
    assign G[3] = in[242] & in2[242];
    assign P[3] = in[242] ^ in2[242];
    assign G[4] = in[241] & in2[241];
    assign P[4] = in[241] ^ in2[241];
    assign G[5] = in[240] & in2[240];
    assign P[5] = in[240] ^ in2[240];
    assign G[6] = in[239] & in2[239];
    assign P[6] = in[239] ^ in2[239];
    assign G[7] = in[238] & in2[238];
    assign P[7] = in[238] ^ in2[238];
    assign G[8] = in[237] & in2[237];
    assign P[8] = in[237] ^ in2[237];
    assign G[9] = in[236] & in2[236];
    assign P[9] = in[236] ^ in2[236];
    assign G[10] = in[235] & in2[235];
    assign P[10] = in[235] ^ in2[235];
    assign G[11] = in[234] & in2[234];
    assign P[11] = in[234] ^ in2[234];
    assign G[12] = in[233] & in2[233];
    assign P[12] = in[233] ^ in2[233];
    assign G[13] = in[232] & in2[232];
    assign P[13] = in[232] ^ in2[232];
    assign G[14] = in[231] & in2[231];
    assign P[14] = in[231] ^ in2[231];
    assign G[15] = in[230] & in2[230];
    assign P[15] = in[230] ^ in2[230];
    assign G[16] = in[229] & in2[229];
    assign P[16] = in[229] ^ in2[229];
    assign G[17] = in[228] & in2[228];
    assign P[17] = in[228] ^ in2[228];
    assign G[18] = in[227] & in2[227];
    assign P[18] = in[227] ^ in2[227];
    assign G[19] = in[226] & in2[226];
    assign P[19] = in[226] ^ in2[226];
    assign G[20] = in[225] & in2[225];
    assign P[20] = in[225] ^ in2[225];
    assign G[21] = in[224] & in2[224];
    assign P[21] = in[224] ^ in2[224];
    assign G[22] = in[223] & in2[223];
    assign P[22] = in[223] ^ in2[223];
    assign G[23] = in[222] & in2[222];
    assign P[23] = in[222] ^ in2[222];
    assign G[24] = in[221] & in2[221];
    assign P[24] = in[221] ^ in2[221];
    assign G[25] = in[220] & in2[220];
    assign P[25] = in[220] ^ in2[220];
    assign G[26] = in[219] & in2[219];
    assign P[26] = in[219] ^ in2[219];
    assign G[27] = in[218] & in2[218];
    assign P[27] = in[218] ^ in2[218];
    assign G[28] = in[217] & in2[217];
    assign P[28] = in[217] ^ in2[217];
    assign G[29] = in[216] & in2[216];
    assign P[29] = in[216] ^ in2[216];
    assign G[30] = in[215] & in2[215];
    assign P[30] = in[215] ^ in2[215];
    assign G[31] = in[214] & in2[214];
    assign P[31] = in[214] ^ in2[214];
    assign G[32] = in[213] & in2[213];
    assign P[32] = in[213] ^ in2[213];
    assign G[33] = in[212] & in2[212];
    assign P[33] = in[212] ^ in2[212];
    assign G[34] = in[211] & in2[211];
    assign P[34] = in[211] ^ in2[211];
    assign G[35] = in[210] & in2[210];
    assign P[35] = in[210] ^ in2[210];
    assign G[36] = in[209] & in2[209];
    assign P[36] = in[209] ^ in2[209];
    assign G[37] = in[208] & in2[208];
    assign P[37] = in[208] ^ in2[208];
    assign G[38] = in[207] & in2[207];
    assign P[38] = in[207] ^ in2[207];
    assign G[39] = in[206] & in2[206];
    assign P[39] = in[206] ^ in2[206];
    assign G[40] = in[205] & in2[205];
    assign P[40] = in[205] ^ in2[205];
    assign G[41] = in[204] & in2[204];
    assign P[41] = in[204] ^ in2[204];
    assign G[42] = in[203] & in2[203];
    assign P[42] = in[203] ^ in2[203];
    assign G[43] = in[202] & in2[202];
    assign P[43] = in[202] ^ in2[202];
    assign G[44] = in[201] & in2[201];
    assign P[44] = in[201] ^ in2[201];
    assign G[45] = in[200] & in2[200];
    assign P[45] = in[200] ^ in2[200];
    assign G[46] = in[199] & in2[199];
    assign P[46] = in[199] ^ in2[199];
    assign G[47] = in[198] & in2[198];
    assign P[47] = in[198] ^ in2[198];
    assign G[48] = in[197] & in2[197];
    assign P[48] = in[197] ^ in2[197];
    assign G[49] = in[196] & in2[196];
    assign P[49] = in[196] ^ in2[196];
    assign G[50] = in[195] & in2[195];
    assign P[50] = in[195] ^ in2[195];
    assign G[51] = in[194] & in2[194];
    assign P[51] = in[194] ^ in2[194];
    assign G[52] = in[193] & in2[193];
    assign P[52] = in[193] ^ in2[193];
    assign G[53] = in[192] & in2[192];
    assign P[53] = in[192] ^ in2[192];
    assign G[54] = in[191] & in2[191];
    assign P[54] = in[191] ^ in2[191];
    assign G[55] = in[190] & in2[190];
    assign P[55] = in[190] ^ in2[190];
    assign G[56] = in[189] & in2[189];
    assign P[56] = in[189] ^ in2[189];
    assign G[57] = in[188] & in2[188];
    assign P[57] = in[188] ^ in2[188];
    assign G[58] = in[187] & in2[187];
    assign P[58] = in[187] ^ in2[187];
    assign G[59] = in[186] & in2[186];
    assign P[59] = in[186] ^ in2[186];
    assign G[60] = in[185] & in2[185];
    assign P[60] = in[185] ^ in2[185];
    assign G[61] = in[184] & in2[184];
    assign P[61] = in[184] ^ in2[184];
    assign G[62] = in[183] & in2[183];
    assign P[62] = in[183] ^ in2[183];
    assign G[63] = in[182] & in2[182];
    assign P[63] = in[182] ^ in2[182];
    assign G[64] = in[181] & in2[181];
    assign P[64] = in[181] ^ in2[181];
    assign G[65] = in[180] & in2[180];
    assign P[65] = in[180] ^ in2[180];
    assign G[66] = in[179] & in2[179];
    assign P[66] = in[179] ^ in2[179];
    assign G[67] = in[178] & in2[178];
    assign P[67] = in[178] ^ in2[178];
    assign G[68] = in[177] & in2[177];
    assign P[68] = in[177] ^ in2[177];
    assign G[69] = in[176] & in2[176];
    assign P[69] = in[176] ^ in2[176];
    assign G[70] = in[175] & in2[175];
    assign P[70] = in[175] ^ in2[175];
    assign G[71] = in[174] & in2[174];
    assign P[71] = in[174] ^ in2[174];
    assign G[72] = in[173] & in2[173];
    assign P[72] = in[173] ^ in2[173];
    assign G[73] = in[172] & in2[172];
    assign P[73] = in[172] ^ in2[172];
    assign G[74] = in[171] & in2[171];
    assign P[74] = in[171] ^ in2[171];
    assign G[75] = in[170] & in2[170];
    assign P[75] = in[170] ^ in2[170];
    assign G[76] = in[169] & in2[169];
    assign P[76] = in[169] ^ in2[169];
    assign G[77] = in[168] & in2[168];
    assign P[77] = in[168] ^ in2[168];
    assign G[78] = in[167] & in2[167];
    assign P[78] = in[167] ^ in2[167];
    assign G[79] = in[166] & in2[166];
    assign P[79] = in[166] ^ in2[166];
    assign G[80] = in[165] & in2[165];
    assign P[80] = in[165] ^ in2[165];
    assign G[81] = in[164] & in2[164];
    assign P[81] = in[164] ^ in2[164];
    assign G[82] = in[163] & in2[163];
    assign P[82] = in[163] ^ in2[163];
    assign G[83] = in[162] & in2[162];
    assign P[83] = in[162] ^ in2[162];
    assign G[84] = in[161] & in2[161];
    assign P[84] = in[161] ^ in2[161];
    assign G[85] = in[160] & in2[160];
    assign P[85] = in[160] ^ in2[160];
    assign G[86] = in[159] & in2[159];
    assign P[86] = in[159] ^ in2[159];
    assign G[87] = in[158] & in2[158];
    assign P[87] = in[158] ^ in2[158];
    assign G[88] = in[157] & in2[157];
    assign P[88] = in[157] ^ in2[157];
    assign G[89] = in[156] & in2[156];
    assign P[89] = in[156] ^ in2[156];
    assign G[90] = in[155] & in2[155];
    assign P[90] = in[155] ^ in2[155];
    assign G[91] = in[154] & in2[154];
    assign P[91] = in[154] ^ in2[154];
    assign G[92] = in[153] & in2[153];
    assign P[92] = in[153] ^ in2[153];
    assign G[93] = in[152] & in2[152];
    assign P[93] = in[152] ^ in2[152];
    assign G[94] = in[151] & in2[151];
    assign P[94] = in[151] ^ in2[151];
    assign G[95] = in[150] & in2[150];
    assign P[95] = in[150] ^ in2[150];
    assign G[96] = in[149] & in2[149];
    assign P[96] = in[149] ^ in2[149];
    assign G[97] = in[148] & in2[148];
    assign P[97] = in[148] ^ in2[148];
    assign G[98] = in[147] & in2[147];
    assign P[98] = in[147] ^ in2[147];
    assign G[99] = in[146] & in2[146];
    assign P[99] = in[146] ^ in2[146];
    assign G[100] = in[145] & in2[145];
    assign P[100] = in[145] ^ in2[145];
    assign G[101] = in[144] & in2[144];
    assign P[101] = in[144] ^ in2[144];
    assign G[102] = in[143] & in2[143];
    assign P[102] = in[143] ^ in2[143];
    assign G[103] = in[142] & in2[142];
    assign P[103] = in[142] ^ in2[142];
    assign G[104] = in[141] & in2[141];
    assign P[104] = in[141] ^ in2[141];
    assign G[105] = in[140] & in2[140];
    assign P[105] = in[140] ^ in2[140];
    assign G[106] = in[139] & in2[139];
    assign P[106] = in[139] ^ in2[139];
    assign G[107] = in[138] & in2[138];
    assign P[107] = in[138] ^ in2[138];
    assign G[108] = in[137] & in2[137];
    assign P[108] = in[137] ^ in2[137];
    assign G[109] = in[136] & in2[136];
    assign P[109] = in[136] ^ in2[136];
    assign G[110] = in[135] & in2[135];
    assign P[110] = in[135] ^ in2[135];
    assign G[111] = in[134] & in2[134];
    assign P[111] = in[134] ^ in2[134];
    assign G[112] = in[133] & in2[133];
    assign P[112] = in[133] ^ in2[133];
    assign G[113] = in[132] & in2[132];
    assign P[113] = in[132] ^ in2[132];
    assign G[114] = in[131] & in2[131];
    assign P[114] = in[131] ^ in2[131];
    assign G[115] = in[130] & in2[130];
    assign P[115] = in[130] ^ in2[130];
    assign G[116] = in[129] & in2[129];
    assign P[116] = in[129] ^ in2[129];
    assign G[117] = in[128] & in2[128];
    assign P[117] = in[128] ^ in2[128];
    assign G[118] = in[127] & in2[127];
    assign P[118] = in[127] ^ in2[127];
    assign G[119] = in[126] & in2[126];
    assign P[119] = in[126] ^ in2[126];
    assign G[120] = in[125] & in2[125];
    assign P[120] = in[125] ^ in2[125];
    assign G[121] = in[124] & in2[124];
    assign P[121] = in[124] ^ in2[124];
    assign G[122] = in[123] & in2[123];
    assign P[122] = in[123] ^ in2[123];
    assign G[123] = in[122] & in2[122];
    assign P[123] = in[122] ^ in2[122];
    assign G[124] = in[121] & in2[121];
    assign P[124] = in[121] ^ in2[121];
    assign G[125] = in[120] & in2[120];
    assign P[125] = in[120] ^ in2[120];
    assign G[126] = in[119] & in2[119];
    assign P[126] = in[119] ^ in2[119];
    assign G[127] = in[118] & in2[118];
    assign P[127] = in[118] ^ in2[118];
    assign G[128] = in[117] & in2[117];
    assign P[128] = in[117] ^ in2[117];
    assign G[129] = in[116] & in2[116];
    assign P[129] = in[116] ^ in2[116];
    assign G[130] = in[115] & in2[115];
    assign P[130] = in[115] ^ in2[115];
    assign G[131] = in[114] & in2[114];
    assign P[131] = in[114] ^ in2[114];
    assign G[132] = in[113] & in2[113];
    assign P[132] = in[113] ^ in2[113];
    assign G[133] = in[112] & in2[112];
    assign P[133] = in[112] ^ in2[112];
    assign G[134] = in[111] & in2[111];
    assign P[134] = in[111] ^ in2[111];
    assign G[135] = in[110] & in2[110];
    assign P[135] = in[110] ^ in2[110];
    assign G[136] = in[109] & in2[109];
    assign P[136] = in[109] ^ in2[109];
    assign G[137] = in[108] & in2[108];
    assign P[137] = in[108] ^ in2[108];
    assign G[138] = in[107] & in2[107];
    assign P[138] = in[107] ^ in2[107];
    assign G[139] = in[106] & in2[106];
    assign P[139] = in[106] ^ in2[106];
    assign G[140] = in[105] & in2[105];
    assign P[140] = in[105] ^ in2[105];
    assign G[141] = in[104] & in2[104];
    assign P[141] = in[104] ^ in2[104];
    assign G[142] = in[103] & in2[103];
    assign P[142] = in[103] ^ in2[103];
    assign G[143] = in[102] & in2[102];
    assign P[143] = in[102] ^ in2[102];
    assign G[144] = in[101] & in2[101];
    assign P[144] = in[101] ^ in2[101];
    assign G[145] = in[100] & in2[100];
    assign P[145] = in[100] ^ in2[100];
    assign G[146] = in[99] & in2[99];
    assign P[146] = in[99] ^ in2[99];
    assign G[147] = in[98] & in2[98];
    assign P[147] = in[98] ^ in2[98];
    assign G[148] = in[97] & in2[97];
    assign P[148] = in[97] ^ in2[97];
    assign G[149] = in[96] & in2[96];
    assign P[149] = in[96] ^ in2[96];
    assign G[150] = in[95] & in2[95];
    assign P[150] = in[95] ^ in2[95];
    assign G[151] = in[94] & in2[94];
    assign P[151] = in[94] ^ in2[94];
    assign G[152] = in[93] & in2[93];
    assign P[152] = in[93] ^ in2[93];
    assign G[153] = in[92] & in2[92];
    assign P[153] = in[92] ^ in2[92];
    assign G[154] = in[91] & in2[91];
    assign P[154] = in[91] ^ in2[91];
    assign G[155] = in[90] & in2[90];
    assign P[155] = in[90] ^ in2[90];
    assign G[156] = in[89] & in2[89];
    assign P[156] = in[89] ^ in2[89];
    assign G[157] = in[88] & in2[88];
    assign P[157] = in[88] ^ in2[88];
    assign G[158] = in[87] & in2[87];
    assign P[158] = in[87] ^ in2[87];
    assign G[159] = in[86] & in2[86];
    assign P[159] = in[86] ^ in2[86];
    assign G[160] = in[85] & in2[85];
    assign P[160] = in[85] ^ in2[85];
    assign G[161] = in[84] & in2[84];
    assign P[161] = in[84] ^ in2[84];
    assign G[162] = in[83] & in2[83];
    assign P[162] = in[83] ^ in2[83];
    assign G[163] = in[82] & in2[82];
    assign P[163] = in[82] ^ in2[82];
    assign G[164] = in[81] & in2[81];
    assign P[164] = in[81] ^ in2[81];
    assign G[165] = in[80] & in2[80];
    assign P[165] = in[80] ^ in2[80];
    assign G[166] = in[79] & in2[79];
    assign P[166] = in[79] ^ in2[79];
    assign G[167] = in[78] & in2[78];
    assign P[167] = in[78] ^ in2[78];
    assign G[168] = in[77] & in2[77];
    assign P[168] = in[77] ^ in2[77];
    assign G[169] = in[76] & in2[76];
    assign P[169] = in[76] ^ in2[76];
    assign G[170] = in[75] & in2[75];
    assign P[170] = in[75] ^ in2[75];
    assign G[171] = in[74] & in2[74];
    assign P[171] = in[74] ^ in2[74];
    assign G[172] = in[73] & in2[73];
    assign P[172] = in[73] ^ in2[73];
    assign G[173] = in[72] & in2[72];
    assign P[173] = in[72] ^ in2[72];
    assign G[174] = in[71] & in2[71];
    assign P[174] = in[71] ^ in2[71];
    assign G[175] = in[70] & in2[70];
    assign P[175] = in[70] ^ in2[70];
    assign G[176] = in[69] & in2[69];
    assign P[176] = in[69] ^ in2[69];
    assign G[177] = in[68] & in2[68];
    assign P[177] = in[68] ^ in2[68];
    assign G[178] = in[67] & in2[67];
    assign P[178] = in[67] ^ in2[67];
    assign G[179] = in[66] & in2[66];
    assign P[179] = in[66] ^ in2[66];
    assign G[180] = in[65] & in2[65];
    assign P[180] = in[65] ^ in2[65];
    assign G[181] = in[64] & in2[64];
    assign P[181] = in[64] ^ in2[64];
    assign G[182] = in[63] & in2[63];
    assign P[182] = in[63] ^ in2[63];
    assign G[183] = in[62] & in2[62];
    assign P[183] = in[62] ^ in2[62];
    assign G[184] = in[61] & in2[61];
    assign P[184] = in[61] ^ in2[61];
    assign G[185] = in[60] & in2[60];
    assign P[185] = in[60] ^ in2[60];
    assign G[186] = in[59] & in2[59];
    assign P[186] = in[59] ^ in2[59];
    assign G[187] = in[58] & in2[58];
    assign P[187] = in[58] ^ in2[58];
    assign G[188] = in[57] & in2[57];
    assign P[188] = in[57] ^ in2[57];
    assign G[189] = in[56] & in2[56];
    assign P[189] = in[56] ^ in2[56];
    assign G[190] = in[55] & in2[55];
    assign P[190] = in[55] ^ in2[55];
    assign G[191] = in[54] & in2[54];
    assign P[191] = in[54] ^ in2[54];
    assign G[192] = in[53] & in2[53];
    assign P[192] = in[53] ^ in2[53];
    assign G[193] = in[52] & in2[52];
    assign P[193] = in[52] ^ in2[52];
    assign G[194] = in[51] & in2[51];
    assign P[194] = in[51] ^ in2[51];
    assign G[195] = in[50] & in2[50];
    assign P[195] = in[50] ^ in2[50];
    assign G[196] = in[49] & in2[49];
    assign P[196] = in[49] ^ in2[49];
    assign G[197] = in[48] & in2[48];
    assign P[197] = in[48] ^ in2[48];
    assign G[198] = in[47] & in2[47];
    assign P[198] = in[47] ^ in2[47];
    assign G[199] = in[46] & in2[46];
    assign P[199] = in[46] ^ in2[46];
    assign G[200] = in[45] & in2[45];
    assign P[200] = in[45] ^ in2[45];
    assign G[201] = in[44] & in2[44];
    assign P[201] = in[44] ^ in2[44];
    assign G[202] = in[43] & in2[43];
    assign P[202] = in[43] ^ in2[43];
    assign G[203] = in[42] & in2[42];
    assign P[203] = in[42] ^ in2[42];
    assign G[204] = in[41] & in2[41];
    assign P[204] = in[41] ^ in2[41];
    assign G[205] = in[40] & in2[40];
    assign P[205] = in[40] ^ in2[40];
    assign G[206] = in[39] & in2[39];
    assign P[206] = in[39] ^ in2[39];
    assign G[207] = in[38] & in2[38];
    assign P[207] = in[38] ^ in2[38];
    assign G[208] = in[37] & in2[37];
    assign P[208] = in[37] ^ in2[37];
    assign G[209] = in[36] & in2[36];
    assign P[209] = in[36] ^ in2[36];
    assign G[210] = in[35] & in2[35];
    assign P[210] = in[35] ^ in2[35];
    assign G[211] = in[34] & in2[34];
    assign P[211] = in[34] ^ in2[34];
    assign G[212] = in[33] & in2[33];
    assign P[212] = in[33] ^ in2[33];
    assign G[213] = in[32] & in2[32];
    assign P[213] = in[32] ^ in2[32];
    assign G[214] = in[31] & in2[31];
    assign P[214] = in[31] ^ in2[31];
    assign G[215] = in[30] & in2[30];
    assign P[215] = in[30] ^ in2[30];
    assign G[216] = in[29] & in2[29];
    assign P[216] = in[29] ^ in2[29];
    assign G[217] = in[28] & in2[28];
    assign P[217] = in[28] ^ in2[28];
    assign G[218] = in[27] & in2[27];
    assign P[218] = in[27] ^ in2[27];
    assign G[219] = in[26] & in2[26];
    assign P[219] = in[26] ^ in2[26];
    assign G[220] = in[25] & in2[25];
    assign P[220] = in[25] ^ in2[25];
    assign G[221] = in[24] & in2[24];
    assign P[221] = in[24] ^ in2[24];
    assign G[222] = in[23] & in2[23];
    assign P[222] = in[23] ^ in2[23];
    assign G[223] = in[22] & in2[22];
    assign P[223] = in[22] ^ in2[22];
    assign G[224] = in[21] & in2[21];
    assign P[224] = in[21] ^ in2[21];
    assign G[225] = in[20] & in2[20];
    assign P[225] = in[20] ^ in2[20];
    assign G[226] = in[19] & in2[19];
    assign P[226] = in[19] ^ in2[19];
    assign G[227] = in[18] & in2[18];
    assign P[227] = in[18] ^ in2[18];
    assign G[228] = in[17] & in2[17];
    assign P[228] = in[17] ^ in2[17];
    assign G[229] = in[16] & in2[16];
    assign P[229] = in[16] ^ in2[16];
    assign G[230] = in[15] & in2[15];
    assign P[230] = in[15] ^ in2[15];
    assign G[231] = in[14] & in2[14];
    assign P[231] = in[14] ^ in2[14];
    assign G[232] = in[13] & in2[13];
    assign P[232] = in[13] ^ in2[13];
    assign G[233] = in[12] & in2[12];
    assign P[233] = in[12] ^ in2[12];
    assign G[234] = in[11] & in2[11];
    assign P[234] = in[11] ^ in2[11];
    assign G[235] = in[10] & in2[10];
    assign P[235] = in[10] ^ in2[10];
    assign G[236] = in[9] & in2[9];
    assign P[236] = in[9] ^ in2[9];
    assign G[237] = in[8] & in2[8];
    assign P[237] = in[8] ^ in2[8];
    assign G[238] = in[7] & in2[7];
    assign P[238] = in[7] ^ in2[7];
    assign G[239] = in[6] & in2[6];
    assign P[239] = in[6] ^ in2[6];
    assign G[240] = in[5] & in2[5];
    assign P[240] = in[5] ^ in2[5];
    assign G[241] = in[4] & in2[4];
    assign P[241] = in[4] ^ in2[4];
    assign G[242] = in[3] & in2[3];
    assign P[242] = in[3] ^ in2[3];
    assign G[243] = in[2] & in2[2];
    assign P[243] = in[2] ^ in2[2];
    assign G[244] = in[1] & in2[1];
    assign P[244] = in[1] ^ in2[1];
    assign G[245] = in[0] & in2[0];
    assign P[245] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign C[245] = G[244] | (P[244] & C[244]);
    assign cout = G[245] | (P[245] & C[245]);
    assign sum = P ^ C;
endmodule

module CLA245(output [244:0] sum, output cout, input [244:0] in1, input [244:0] in2;

    wire[244:0] G;
    wire[244:0] C;
    wire[244:0] P;

    assign G[0] = in[244] & in2[244];
    assign P[0] = in[244] ^ in2[244];
    assign G[1] = in[243] & in2[243];
    assign P[1] = in[243] ^ in2[243];
    assign G[2] = in[242] & in2[242];
    assign P[2] = in[242] ^ in2[242];
    assign G[3] = in[241] & in2[241];
    assign P[3] = in[241] ^ in2[241];
    assign G[4] = in[240] & in2[240];
    assign P[4] = in[240] ^ in2[240];
    assign G[5] = in[239] & in2[239];
    assign P[5] = in[239] ^ in2[239];
    assign G[6] = in[238] & in2[238];
    assign P[6] = in[238] ^ in2[238];
    assign G[7] = in[237] & in2[237];
    assign P[7] = in[237] ^ in2[237];
    assign G[8] = in[236] & in2[236];
    assign P[8] = in[236] ^ in2[236];
    assign G[9] = in[235] & in2[235];
    assign P[9] = in[235] ^ in2[235];
    assign G[10] = in[234] & in2[234];
    assign P[10] = in[234] ^ in2[234];
    assign G[11] = in[233] & in2[233];
    assign P[11] = in[233] ^ in2[233];
    assign G[12] = in[232] & in2[232];
    assign P[12] = in[232] ^ in2[232];
    assign G[13] = in[231] & in2[231];
    assign P[13] = in[231] ^ in2[231];
    assign G[14] = in[230] & in2[230];
    assign P[14] = in[230] ^ in2[230];
    assign G[15] = in[229] & in2[229];
    assign P[15] = in[229] ^ in2[229];
    assign G[16] = in[228] & in2[228];
    assign P[16] = in[228] ^ in2[228];
    assign G[17] = in[227] & in2[227];
    assign P[17] = in[227] ^ in2[227];
    assign G[18] = in[226] & in2[226];
    assign P[18] = in[226] ^ in2[226];
    assign G[19] = in[225] & in2[225];
    assign P[19] = in[225] ^ in2[225];
    assign G[20] = in[224] & in2[224];
    assign P[20] = in[224] ^ in2[224];
    assign G[21] = in[223] & in2[223];
    assign P[21] = in[223] ^ in2[223];
    assign G[22] = in[222] & in2[222];
    assign P[22] = in[222] ^ in2[222];
    assign G[23] = in[221] & in2[221];
    assign P[23] = in[221] ^ in2[221];
    assign G[24] = in[220] & in2[220];
    assign P[24] = in[220] ^ in2[220];
    assign G[25] = in[219] & in2[219];
    assign P[25] = in[219] ^ in2[219];
    assign G[26] = in[218] & in2[218];
    assign P[26] = in[218] ^ in2[218];
    assign G[27] = in[217] & in2[217];
    assign P[27] = in[217] ^ in2[217];
    assign G[28] = in[216] & in2[216];
    assign P[28] = in[216] ^ in2[216];
    assign G[29] = in[215] & in2[215];
    assign P[29] = in[215] ^ in2[215];
    assign G[30] = in[214] & in2[214];
    assign P[30] = in[214] ^ in2[214];
    assign G[31] = in[213] & in2[213];
    assign P[31] = in[213] ^ in2[213];
    assign G[32] = in[212] & in2[212];
    assign P[32] = in[212] ^ in2[212];
    assign G[33] = in[211] & in2[211];
    assign P[33] = in[211] ^ in2[211];
    assign G[34] = in[210] & in2[210];
    assign P[34] = in[210] ^ in2[210];
    assign G[35] = in[209] & in2[209];
    assign P[35] = in[209] ^ in2[209];
    assign G[36] = in[208] & in2[208];
    assign P[36] = in[208] ^ in2[208];
    assign G[37] = in[207] & in2[207];
    assign P[37] = in[207] ^ in2[207];
    assign G[38] = in[206] & in2[206];
    assign P[38] = in[206] ^ in2[206];
    assign G[39] = in[205] & in2[205];
    assign P[39] = in[205] ^ in2[205];
    assign G[40] = in[204] & in2[204];
    assign P[40] = in[204] ^ in2[204];
    assign G[41] = in[203] & in2[203];
    assign P[41] = in[203] ^ in2[203];
    assign G[42] = in[202] & in2[202];
    assign P[42] = in[202] ^ in2[202];
    assign G[43] = in[201] & in2[201];
    assign P[43] = in[201] ^ in2[201];
    assign G[44] = in[200] & in2[200];
    assign P[44] = in[200] ^ in2[200];
    assign G[45] = in[199] & in2[199];
    assign P[45] = in[199] ^ in2[199];
    assign G[46] = in[198] & in2[198];
    assign P[46] = in[198] ^ in2[198];
    assign G[47] = in[197] & in2[197];
    assign P[47] = in[197] ^ in2[197];
    assign G[48] = in[196] & in2[196];
    assign P[48] = in[196] ^ in2[196];
    assign G[49] = in[195] & in2[195];
    assign P[49] = in[195] ^ in2[195];
    assign G[50] = in[194] & in2[194];
    assign P[50] = in[194] ^ in2[194];
    assign G[51] = in[193] & in2[193];
    assign P[51] = in[193] ^ in2[193];
    assign G[52] = in[192] & in2[192];
    assign P[52] = in[192] ^ in2[192];
    assign G[53] = in[191] & in2[191];
    assign P[53] = in[191] ^ in2[191];
    assign G[54] = in[190] & in2[190];
    assign P[54] = in[190] ^ in2[190];
    assign G[55] = in[189] & in2[189];
    assign P[55] = in[189] ^ in2[189];
    assign G[56] = in[188] & in2[188];
    assign P[56] = in[188] ^ in2[188];
    assign G[57] = in[187] & in2[187];
    assign P[57] = in[187] ^ in2[187];
    assign G[58] = in[186] & in2[186];
    assign P[58] = in[186] ^ in2[186];
    assign G[59] = in[185] & in2[185];
    assign P[59] = in[185] ^ in2[185];
    assign G[60] = in[184] & in2[184];
    assign P[60] = in[184] ^ in2[184];
    assign G[61] = in[183] & in2[183];
    assign P[61] = in[183] ^ in2[183];
    assign G[62] = in[182] & in2[182];
    assign P[62] = in[182] ^ in2[182];
    assign G[63] = in[181] & in2[181];
    assign P[63] = in[181] ^ in2[181];
    assign G[64] = in[180] & in2[180];
    assign P[64] = in[180] ^ in2[180];
    assign G[65] = in[179] & in2[179];
    assign P[65] = in[179] ^ in2[179];
    assign G[66] = in[178] & in2[178];
    assign P[66] = in[178] ^ in2[178];
    assign G[67] = in[177] & in2[177];
    assign P[67] = in[177] ^ in2[177];
    assign G[68] = in[176] & in2[176];
    assign P[68] = in[176] ^ in2[176];
    assign G[69] = in[175] & in2[175];
    assign P[69] = in[175] ^ in2[175];
    assign G[70] = in[174] & in2[174];
    assign P[70] = in[174] ^ in2[174];
    assign G[71] = in[173] & in2[173];
    assign P[71] = in[173] ^ in2[173];
    assign G[72] = in[172] & in2[172];
    assign P[72] = in[172] ^ in2[172];
    assign G[73] = in[171] & in2[171];
    assign P[73] = in[171] ^ in2[171];
    assign G[74] = in[170] & in2[170];
    assign P[74] = in[170] ^ in2[170];
    assign G[75] = in[169] & in2[169];
    assign P[75] = in[169] ^ in2[169];
    assign G[76] = in[168] & in2[168];
    assign P[76] = in[168] ^ in2[168];
    assign G[77] = in[167] & in2[167];
    assign P[77] = in[167] ^ in2[167];
    assign G[78] = in[166] & in2[166];
    assign P[78] = in[166] ^ in2[166];
    assign G[79] = in[165] & in2[165];
    assign P[79] = in[165] ^ in2[165];
    assign G[80] = in[164] & in2[164];
    assign P[80] = in[164] ^ in2[164];
    assign G[81] = in[163] & in2[163];
    assign P[81] = in[163] ^ in2[163];
    assign G[82] = in[162] & in2[162];
    assign P[82] = in[162] ^ in2[162];
    assign G[83] = in[161] & in2[161];
    assign P[83] = in[161] ^ in2[161];
    assign G[84] = in[160] & in2[160];
    assign P[84] = in[160] ^ in2[160];
    assign G[85] = in[159] & in2[159];
    assign P[85] = in[159] ^ in2[159];
    assign G[86] = in[158] & in2[158];
    assign P[86] = in[158] ^ in2[158];
    assign G[87] = in[157] & in2[157];
    assign P[87] = in[157] ^ in2[157];
    assign G[88] = in[156] & in2[156];
    assign P[88] = in[156] ^ in2[156];
    assign G[89] = in[155] & in2[155];
    assign P[89] = in[155] ^ in2[155];
    assign G[90] = in[154] & in2[154];
    assign P[90] = in[154] ^ in2[154];
    assign G[91] = in[153] & in2[153];
    assign P[91] = in[153] ^ in2[153];
    assign G[92] = in[152] & in2[152];
    assign P[92] = in[152] ^ in2[152];
    assign G[93] = in[151] & in2[151];
    assign P[93] = in[151] ^ in2[151];
    assign G[94] = in[150] & in2[150];
    assign P[94] = in[150] ^ in2[150];
    assign G[95] = in[149] & in2[149];
    assign P[95] = in[149] ^ in2[149];
    assign G[96] = in[148] & in2[148];
    assign P[96] = in[148] ^ in2[148];
    assign G[97] = in[147] & in2[147];
    assign P[97] = in[147] ^ in2[147];
    assign G[98] = in[146] & in2[146];
    assign P[98] = in[146] ^ in2[146];
    assign G[99] = in[145] & in2[145];
    assign P[99] = in[145] ^ in2[145];
    assign G[100] = in[144] & in2[144];
    assign P[100] = in[144] ^ in2[144];
    assign G[101] = in[143] & in2[143];
    assign P[101] = in[143] ^ in2[143];
    assign G[102] = in[142] & in2[142];
    assign P[102] = in[142] ^ in2[142];
    assign G[103] = in[141] & in2[141];
    assign P[103] = in[141] ^ in2[141];
    assign G[104] = in[140] & in2[140];
    assign P[104] = in[140] ^ in2[140];
    assign G[105] = in[139] & in2[139];
    assign P[105] = in[139] ^ in2[139];
    assign G[106] = in[138] & in2[138];
    assign P[106] = in[138] ^ in2[138];
    assign G[107] = in[137] & in2[137];
    assign P[107] = in[137] ^ in2[137];
    assign G[108] = in[136] & in2[136];
    assign P[108] = in[136] ^ in2[136];
    assign G[109] = in[135] & in2[135];
    assign P[109] = in[135] ^ in2[135];
    assign G[110] = in[134] & in2[134];
    assign P[110] = in[134] ^ in2[134];
    assign G[111] = in[133] & in2[133];
    assign P[111] = in[133] ^ in2[133];
    assign G[112] = in[132] & in2[132];
    assign P[112] = in[132] ^ in2[132];
    assign G[113] = in[131] & in2[131];
    assign P[113] = in[131] ^ in2[131];
    assign G[114] = in[130] & in2[130];
    assign P[114] = in[130] ^ in2[130];
    assign G[115] = in[129] & in2[129];
    assign P[115] = in[129] ^ in2[129];
    assign G[116] = in[128] & in2[128];
    assign P[116] = in[128] ^ in2[128];
    assign G[117] = in[127] & in2[127];
    assign P[117] = in[127] ^ in2[127];
    assign G[118] = in[126] & in2[126];
    assign P[118] = in[126] ^ in2[126];
    assign G[119] = in[125] & in2[125];
    assign P[119] = in[125] ^ in2[125];
    assign G[120] = in[124] & in2[124];
    assign P[120] = in[124] ^ in2[124];
    assign G[121] = in[123] & in2[123];
    assign P[121] = in[123] ^ in2[123];
    assign G[122] = in[122] & in2[122];
    assign P[122] = in[122] ^ in2[122];
    assign G[123] = in[121] & in2[121];
    assign P[123] = in[121] ^ in2[121];
    assign G[124] = in[120] & in2[120];
    assign P[124] = in[120] ^ in2[120];
    assign G[125] = in[119] & in2[119];
    assign P[125] = in[119] ^ in2[119];
    assign G[126] = in[118] & in2[118];
    assign P[126] = in[118] ^ in2[118];
    assign G[127] = in[117] & in2[117];
    assign P[127] = in[117] ^ in2[117];
    assign G[128] = in[116] & in2[116];
    assign P[128] = in[116] ^ in2[116];
    assign G[129] = in[115] & in2[115];
    assign P[129] = in[115] ^ in2[115];
    assign G[130] = in[114] & in2[114];
    assign P[130] = in[114] ^ in2[114];
    assign G[131] = in[113] & in2[113];
    assign P[131] = in[113] ^ in2[113];
    assign G[132] = in[112] & in2[112];
    assign P[132] = in[112] ^ in2[112];
    assign G[133] = in[111] & in2[111];
    assign P[133] = in[111] ^ in2[111];
    assign G[134] = in[110] & in2[110];
    assign P[134] = in[110] ^ in2[110];
    assign G[135] = in[109] & in2[109];
    assign P[135] = in[109] ^ in2[109];
    assign G[136] = in[108] & in2[108];
    assign P[136] = in[108] ^ in2[108];
    assign G[137] = in[107] & in2[107];
    assign P[137] = in[107] ^ in2[107];
    assign G[138] = in[106] & in2[106];
    assign P[138] = in[106] ^ in2[106];
    assign G[139] = in[105] & in2[105];
    assign P[139] = in[105] ^ in2[105];
    assign G[140] = in[104] & in2[104];
    assign P[140] = in[104] ^ in2[104];
    assign G[141] = in[103] & in2[103];
    assign P[141] = in[103] ^ in2[103];
    assign G[142] = in[102] & in2[102];
    assign P[142] = in[102] ^ in2[102];
    assign G[143] = in[101] & in2[101];
    assign P[143] = in[101] ^ in2[101];
    assign G[144] = in[100] & in2[100];
    assign P[144] = in[100] ^ in2[100];
    assign G[145] = in[99] & in2[99];
    assign P[145] = in[99] ^ in2[99];
    assign G[146] = in[98] & in2[98];
    assign P[146] = in[98] ^ in2[98];
    assign G[147] = in[97] & in2[97];
    assign P[147] = in[97] ^ in2[97];
    assign G[148] = in[96] & in2[96];
    assign P[148] = in[96] ^ in2[96];
    assign G[149] = in[95] & in2[95];
    assign P[149] = in[95] ^ in2[95];
    assign G[150] = in[94] & in2[94];
    assign P[150] = in[94] ^ in2[94];
    assign G[151] = in[93] & in2[93];
    assign P[151] = in[93] ^ in2[93];
    assign G[152] = in[92] & in2[92];
    assign P[152] = in[92] ^ in2[92];
    assign G[153] = in[91] & in2[91];
    assign P[153] = in[91] ^ in2[91];
    assign G[154] = in[90] & in2[90];
    assign P[154] = in[90] ^ in2[90];
    assign G[155] = in[89] & in2[89];
    assign P[155] = in[89] ^ in2[89];
    assign G[156] = in[88] & in2[88];
    assign P[156] = in[88] ^ in2[88];
    assign G[157] = in[87] & in2[87];
    assign P[157] = in[87] ^ in2[87];
    assign G[158] = in[86] & in2[86];
    assign P[158] = in[86] ^ in2[86];
    assign G[159] = in[85] & in2[85];
    assign P[159] = in[85] ^ in2[85];
    assign G[160] = in[84] & in2[84];
    assign P[160] = in[84] ^ in2[84];
    assign G[161] = in[83] & in2[83];
    assign P[161] = in[83] ^ in2[83];
    assign G[162] = in[82] & in2[82];
    assign P[162] = in[82] ^ in2[82];
    assign G[163] = in[81] & in2[81];
    assign P[163] = in[81] ^ in2[81];
    assign G[164] = in[80] & in2[80];
    assign P[164] = in[80] ^ in2[80];
    assign G[165] = in[79] & in2[79];
    assign P[165] = in[79] ^ in2[79];
    assign G[166] = in[78] & in2[78];
    assign P[166] = in[78] ^ in2[78];
    assign G[167] = in[77] & in2[77];
    assign P[167] = in[77] ^ in2[77];
    assign G[168] = in[76] & in2[76];
    assign P[168] = in[76] ^ in2[76];
    assign G[169] = in[75] & in2[75];
    assign P[169] = in[75] ^ in2[75];
    assign G[170] = in[74] & in2[74];
    assign P[170] = in[74] ^ in2[74];
    assign G[171] = in[73] & in2[73];
    assign P[171] = in[73] ^ in2[73];
    assign G[172] = in[72] & in2[72];
    assign P[172] = in[72] ^ in2[72];
    assign G[173] = in[71] & in2[71];
    assign P[173] = in[71] ^ in2[71];
    assign G[174] = in[70] & in2[70];
    assign P[174] = in[70] ^ in2[70];
    assign G[175] = in[69] & in2[69];
    assign P[175] = in[69] ^ in2[69];
    assign G[176] = in[68] & in2[68];
    assign P[176] = in[68] ^ in2[68];
    assign G[177] = in[67] & in2[67];
    assign P[177] = in[67] ^ in2[67];
    assign G[178] = in[66] & in2[66];
    assign P[178] = in[66] ^ in2[66];
    assign G[179] = in[65] & in2[65];
    assign P[179] = in[65] ^ in2[65];
    assign G[180] = in[64] & in2[64];
    assign P[180] = in[64] ^ in2[64];
    assign G[181] = in[63] & in2[63];
    assign P[181] = in[63] ^ in2[63];
    assign G[182] = in[62] & in2[62];
    assign P[182] = in[62] ^ in2[62];
    assign G[183] = in[61] & in2[61];
    assign P[183] = in[61] ^ in2[61];
    assign G[184] = in[60] & in2[60];
    assign P[184] = in[60] ^ in2[60];
    assign G[185] = in[59] & in2[59];
    assign P[185] = in[59] ^ in2[59];
    assign G[186] = in[58] & in2[58];
    assign P[186] = in[58] ^ in2[58];
    assign G[187] = in[57] & in2[57];
    assign P[187] = in[57] ^ in2[57];
    assign G[188] = in[56] & in2[56];
    assign P[188] = in[56] ^ in2[56];
    assign G[189] = in[55] & in2[55];
    assign P[189] = in[55] ^ in2[55];
    assign G[190] = in[54] & in2[54];
    assign P[190] = in[54] ^ in2[54];
    assign G[191] = in[53] & in2[53];
    assign P[191] = in[53] ^ in2[53];
    assign G[192] = in[52] & in2[52];
    assign P[192] = in[52] ^ in2[52];
    assign G[193] = in[51] & in2[51];
    assign P[193] = in[51] ^ in2[51];
    assign G[194] = in[50] & in2[50];
    assign P[194] = in[50] ^ in2[50];
    assign G[195] = in[49] & in2[49];
    assign P[195] = in[49] ^ in2[49];
    assign G[196] = in[48] & in2[48];
    assign P[196] = in[48] ^ in2[48];
    assign G[197] = in[47] & in2[47];
    assign P[197] = in[47] ^ in2[47];
    assign G[198] = in[46] & in2[46];
    assign P[198] = in[46] ^ in2[46];
    assign G[199] = in[45] & in2[45];
    assign P[199] = in[45] ^ in2[45];
    assign G[200] = in[44] & in2[44];
    assign P[200] = in[44] ^ in2[44];
    assign G[201] = in[43] & in2[43];
    assign P[201] = in[43] ^ in2[43];
    assign G[202] = in[42] & in2[42];
    assign P[202] = in[42] ^ in2[42];
    assign G[203] = in[41] & in2[41];
    assign P[203] = in[41] ^ in2[41];
    assign G[204] = in[40] & in2[40];
    assign P[204] = in[40] ^ in2[40];
    assign G[205] = in[39] & in2[39];
    assign P[205] = in[39] ^ in2[39];
    assign G[206] = in[38] & in2[38];
    assign P[206] = in[38] ^ in2[38];
    assign G[207] = in[37] & in2[37];
    assign P[207] = in[37] ^ in2[37];
    assign G[208] = in[36] & in2[36];
    assign P[208] = in[36] ^ in2[36];
    assign G[209] = in[35] & in2[35];
    assign P[209] = in[35] ^ in2[35];
    assign G[210] = in[34] & in2[34];
    assign P[210] = in[34] ^ in2[34];
    assign G[211] = in[33] & in2[33];
    assign P[211] = in[33] ^ in2[33];
    assign G[212] = in[32] & in2[32];
    assign P[212] = in[32] ^ in2[32];
    assign G[213] = in[31] & in2[31];
    assign P[213] = in[31] ^ in2[31];
    assign G[214] = in[30] & in2[30];
    assign P[214] = in[30] ^ in2[30];
    assign G[215] = in[29] & in2[29];
    assign P[215] = in[29] ^ in2[29];
    assign G[216] = in[28] & in2[28];
    assign P[216] = in[28] ^ in2[28];
    assign G[217] = in[27] & in2[27];
    assign P[217] = in[27] ^ in2[27];
    assign G[218] = in[26] & in2[26];
    assign P[218] = in[26] ^ in2[26];
    assign G[219] = in[25] & in2[25];
    assign P[219] = in[25] ^ in2[25];
    assign G[220] = in[24] & in2[24];
    assign P[220] = in[24] ^ in2[24];
    assign G[221] = in[23] & in2[23];
    assign P[221] = in[23] ^ in2[23];
    assign G[222] = in[22] & in2[22];
    assign P[222] = in[22] ^ in2[22];
    assign G[223] = in[21] & in2[21];
    assign P[223] = in[21] ^ in2[21];
    assign G[224] = in[20] & in2[20];
    assign P[224] = in[20] ^ in2[20];
    assign G[225] = in[19] & in2[19];
    assign P[225] = in[19] ^ in2[19];
    assign G[226] = in[18] & in2[18];
    assign P[226] = in[18] ^ in2[18];
    assign G[227] = in[17] & in2[17];
    assign P[227] = in[17] ^ in2[17];
    assign G[228] = in[16] & in2[16];
    assign P[228] = in[16] ^ in2[16];
    assign G[229] = in[15] & in2[15];
    assign P[229] = in[15] ^ in2[15];
    assign G[230] = in[14] & in2[14];
    assign P[230] = in[14] ^ in2[14];
    assign G[231] = in[13] & in2[13];
    assign P[231] = in[13] ^ in2[13];
    assign G[232] = in[12] & in2[12];
    assign P[232] = in[12] ^ in2[12];
    assign G[233] = in[11] & in2[11];
    assign P[233] = in[11] ^ in2[11];
    assign G[234] = in[10] & in2[10];
    assign P[234] = in[10] ^ in2[10];
    assign G[235] = in[9] & in2[9];
    assign P[235] = in[9] ^ in2[9];
    assign G[236] = in[8] & in2[8];
    assign P[236] = in[8] ^ in2[8];
    assign G[237] = in[7] & in2[7];
    assign P[237] = in[7] ^ in2[7];
    assign G[238] = in[6] & in2[6];
    assign P[238] = in[6] ^ in2[6];
    assign G[239] = in[5] & in2[5];
    assign P[239] = in[5] ^ in2[5];
    assign G[240] = in[4] & in2[4];
    assign P[240] = in[4] ^ in2[4];
    assign G[241] = in[3] & in2[3];
    assign P[241] = in[3] ^ in2[3];
    assign G[242] = in[2] & in2[2];
    assign P[242] = in[2] ^ in2[2];
    assign G[243] = in[1] & in2[1];
    assign P[243] = in[1] ^ in2[1];
    assign G[244] = in[0] & in2[0];
    assign P[244] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign C[244] = G[243] | (P[243] & C[243]);
    assign cout = G[244] | (P[244] & C[244]);
    assign sum = P ^ C;
endmodule

module CLA244(output [243:0] sum, output cout, input [243:0] in1, input [243:0] in2;

    wire[243:0] G;
    wire[243:0] C;
    wire[243:0] P;

    assign G[0] = in[243] & in2[243];
    assign P[0] = in[243] ^ in2[243];
    assign G[1] = in[242] & in2[242];
    assign P[1] = in[242] ^ in2[242];
    assign G[2] = in[241] & in2[241];
    assign P[2] = in[241] ^ in2[241];
    assign G[3] = in[240] & in2[240];
    assign P[3] = in[240] ^ in2[240];
    assign G[4] = in[239] & in2[239];
    assign P[4] = in[239] ^ in2[239];
    assign G[5] = in[238] & in2[238];
    assign P[5] = in[238] ^ in2[238];
    assign G[6] = in[237] & in2[237];
    assign P[6] = in[237] ^ in2[237];
    assign G[7] = in[236] & in2[236];
    assign P[7] = in[236] ^ in2[236];
    assign G[8] = in[235] & in2[235];
    assign P[8] = in[235] ^ in2[235];
    assign G[9] = in[234] & in2[234];
    assign P[9] = in[234] ^ in2[234];
    assign G[10] = in[233] & in2[233];
    assign P[10] = in[233] ^ in2[233];
    assign G[11] = in[232] & in2[232];
    assign P[11] = in[232] ^ in2[232];
    assign G[12] = in[231] & in2[231];
    assign P[12] = in[231] ^ in2[231];
    assign G[13] = in[230] & in2[230];
    assign P[13] = in[230] ^ in2[230];
    assign G[14] = in[229] & in2[229];
    assign P[14] = in[229] ^ in2[229];
    assign G[15] = in[228] & in2[228];
    assign P[15] = in[228] ^ in2[228];
    assign G[16] = in[227] & in2[227];
    assign P[16] = in[227] ^ in2[227];
    assign G[17] = in[226] & in2[226];
    assign P[17] = in[226] ^ in2[226];
    assign G[18] = in[225] & in2[225];
    assign P[18] = in[225] ^ in2[225];
    assign G[19] = in[224] & in2[224];
    assign P[19] = in[224] ^ in2[224];
    assign G[20] = in[223] & in2[223];
    assign P[20] = in[223] ^ in2[223];
    assign G[21] = in[222] & in2[222];
    assign P[21] = in[222] ^ in2[222];
    assign G[22] = in[221] & in2[221];
    assign P[22] = in[221] ^ in2[221];
    assign G[23] = in[220] & in2[220];
    assign P[23] = in[220] ^ in2[220];
    assign G[24] = in[219] & in2[219];
    assign P[24] = in[219] ^ in2[219];
    assign G[25] = in[218] & in2[218];
    assign P[25] = in[218] ^ in2[218];
    assign G[26] = in[217] & in2[217];
    assign P[26] = in[217] ^ in2[217];
    assign G[27] = in[216] & in2[216];
    assign P[27] = in[216] ^ in2[216];
    assign G[28] = in[215] & in2[215];
    assign P[28] = in[215] ^ in2[215];
    assign G[29] = in[214] & in2[214];
    assign P[29] = in[214] ^ in2[214];
    assign G[30] = in[213] & in2[213];
    assign P[30] = in[213] ^ in2[213];
    assign G[31] = in[212] & in2[212];
    assign P[31] = in[212] ^ in2[212];
    assign G[32] = in[211] & in2[211];
    assign P[32] = in[211] ^ in2[211];
    assign G[33] = in[210] & in2[210];
    assign P[33] = in[210] ^ in2[210];
    assign G[34] = in[209] & in2[209];
    assign P[34] = in[209] ^ in2[209];
    assign G[35] = in[208] & in2[208];
    assign P[35] = in[208] ^ in2[208];
    assign G[36] = in[207] & in2[207];
    assign P[36] = in[207] ^ in2[207];
    assign G[37] = in[206] & in2[206];
    assign P[37] = in[206] ^ in2[206];
    assign G[38] = in[205] & in2[205];
    assign P[38] = in[205] ^ in2[205];
    assign G[39] = in[204] & in2[204];
    assign P[39] = in[204] ^ in2[204];
    assign G[40] = in[203] & in2[203];
    assign P[40] = in[203] ^ in2[203];
    assign G[41] = in[202] & in2[202];
    assign P[41] = in[202] ^ in2[202];
    assign G[42] = in[201] & in2[201];
    assign P[42] = in[201] ^ in2[201];
    assign G[43] = in[200] & in2[200];
    assign P[43] = in[200] ^ in2[200];
    assign G[44] = in[199] & in2[199];
    assign P[44] = in[199] ^ in2[199];
    assign G[45] = in[198] & in2[198];
    assign P[45] = in[198] ^ in2[198];
    assign G[46] = in[197] & in2[197];
    assign P[46] = in[197] ^ in2[197];
    assign G[47] = in[196] & in2[196];
    assign P[47] = in[196] ^ in2[196];
    assign G[48] = in[195] & in2[195];
    assign P[48] = in[195] ^ in2[195];
    assign G[49] = in[194] & in2[194];
    assign P[49] = in[194] ^ in2[194];
    assign G[50] = in[193] & in2[193];
    assign P[50] = in[193] ^ in2[193];
    assign G[51] = in[192] & in2[192];
    assign P[51] = in[192] ^ in2[192];
    assign G[52] = in[191] & in2[191];
    assign P[52] = in[191] ^ in2[191];
    assign G[53] = in[190] & in2[190];
    assign P[53] = in[190] ^ in2[190];
    assign G[54] = in[189] & in2[189];
    assign P[54] = in[189] ^ in2[189];
    assign G[55] = in[188] & in2[188];
    assign P[55] = in[188] ^ in2[188];
    assign G[56] = in[187] & in2[187];
    assign P[56] = in[187] ^ in2[187];
    assign G[57] = in[186] & in2[186];
    assign P[57] = in[186] ^ in2[186];
    assign G[58] = in[185] & in2[185];
    assign P[58] = in[185] ^ in2[185];
    assign G[59] = in[184] & in2[184];
    assign P[59] = in[184] ^ in2[184];
    assign G[60] = in[183] & in2[183];
    assign P[60] = in[183] ^ in2[183];
    assign G[61] = in[182] & in2[182];
    assign P[61] = in[182] ^ in2[182];
    assign G[62] = in[181] & in2[181];
    assign P[62] = in[181] ^ in2[181];
    assign G[63] = in[180] & in2[180];
    assign P[63] = in[180] ^ in2[180];
    assign G[64] = in[179] & in2[179];
    assign P[64] = in[179] ^ in2[179];
    assign G[65] = in[178] & in2[178];
    assign P[65] = in[178] ^ in2[178];
    assign G[66] = in[177] & in2[177];
    assign P[66] = in[177] ^ in2[177];
    assign G[67] = in[176] & in2[176];
    assign P[67] = in[176] ^ in2[176];
    assign G[68] = in[175] & in2[175];
    assign P[68] = in[175] ^ in2[175];
    assign G[69] = in[174] & in2[174];
    assign P[69] = in[174] ^ in2[174];
    assign G[70] = in[173] & in2[173];
    assign P[70] = in[173] ^ in2[173];
    assign G[71] = in[172] & in2[172];
    assign P[71] = in[172] ^ in2[172];
    assign G[72] = in[171] & in2[171];
    assign P[72] = in[171] ^ in2[171];
    assign G[73] = in[170] & in2[170];
    assign P[73] = in[170] ^ in2[170];
    assign G[74] = in[169] & in2[169];
    assign P[74] = in[169] ^ in2[169];
    assign G[75] = in[168] & in2[168];
    assign P[75] = in[168] ^ in2[168];
    assign G[76] = in[167] & in2[167];
    assign P[76] = in[167] ^ in2[167];
    assign G[77] = in[166] & in2[166];
    assign P[77] = in[166] ^ in2[166];
    assign G[78] = in[165] & in2[165];
    assign P[78] = in[165] ^ in2[165];
    assign G[79] = in[164] & in2[164];
    assign P[79] = in[164] ^ in2[164];
    assign G[80] = in[163] & in2[163];
    assign P[80] = in[163] ^ in2[163];
    assign G[81] = in[162] & in2[162];
    assign P[81] = in[162] ^ in2[162];
    assign G[82] = in[161] & in2[161];
    assign P[82] = in[161] ^ in2[161];
    assign G[83] = in[160] & in2[160];
    assign P[83] = in[160] ^ in2[160];
    assign G[84] = in[159] & in2[159];
    assign P[84] = in[159] ^ in2[159];
    assign G[85] = in[158] & in2[158];
    assign P[85] = in[158] ^ in2[158];
    assign G[86] = in[157] & in2[157];
    assign P[86] = in[157] ^ in2[157];
    assign G[87] = in[156] & in2[156];
    assign P[87] = in[156] ^ in2[156];
    assign G[88] = in[155] & in2[155];
    assign P[88] = in[155] ^ in2[155];
    assign G[89] = in[154] & in2[154];
    assign P[89] = in[154] ^ in2[154];
    assign G[90] = in[153] & in2[153];
    assign P[90] = in[153] ^ in2[153];
    assign G[91] = in[152] & in2[152];
    assign P[91] = in[152] ^ in2[152];
    assign G[92] = in[151] & in2[151];
    assign P[92] = in[151] ^ in2[151];
    assign G[93] = in[150] & in2[150];
    assign P[93] = in[150] ^ in2[150];
    assign G[94] = in[149] & in2[149];
    assign P[94] = in[149] ^ in2[149];
    assign G[95] = in[148] & in2[148];
    assign P[95] = in[148] ^ in2[148];
    assign G[96] = in[147] & in2[147];
    assign P[96] = in[147] ^ in2[147];
    assign G[97] = in[146] & in2[146];
    assign P[97] = in[146] ^ in2[146];
    assign G[98] = in[145] & in2[145];
    assign P[98] = in[145] ^ in2[145];
    assign G[99] = in[144] & in2[144];
    assign P[99] = in[144] ^ in2[144];
    assign G[100] = in[143] & in2[143];
    assign P[100] = in[143] ^ in2[143];
    assign G[101] = in[142] & in2[142];
    assign P[101] = in[142] ^ in2[142];
    assign G[102] = in[141] & in2[141];
    assign P[102] = in[141] ^ in2[141];
    assign G[103] = in[140] & in2[140];
    assign P[103] = in[140] ^ in2[140];
    assign G[104] = in[139] & in2[139];
    assign P[104] = in[139] ^ in2[139];
    assign G[105] = in[138] & in2[138];
    assign P[105] = in[138] ^ in2[138];
    assign G[106] = in[137] & in2[137];
    assign P[106] = in[137] ^ in2[137];
    assign G[107] = in[136] & in2[136];
    assign P[107] = in[136] ^ in2[136];
    assign G[108] = in[135] & in2[135];
    assign P[108] = in[135] ^ in2[135];
    assign G[109] = in[134] & in2[134];
    assign P[109] = in[134] ^ in2[134];
    assign G[110] = in[133] & in2[133];
    assign P[110] = in[133] ^ in2[133];
    assign G[111] = in[132] & in2[132];
    assign P[111] = in[132] ^ in2[132];
    assign G[112] = in[131] & in2[131];
    assign P[112] = in[131] ^ in2[131];
    assign G[113] = in[130] & in2[130];
    assign P[113] = in[130] ^ in2[130];
    assign G[114] = in[129] & in2[129];
    assign P[114] = in[129] ^ in2[129];
    assign G[115] = in[128] & in2[128];
    assign P[115] = in[128] ^ in2[128];
    assign G[116] = in[127] & in2[127];
    assign P[116] = in[127] ^ in2[127];
    assign G[117] = in[126] & in2[126];
    assign P[117] = in[126] ^ in2[126];
    assign G[118] = in[125] & in2[125];
    assign P[118] = in[125] ^ in2[125];
    assign G[119] = in[124] & in2[124];
    assign P[119] = in[124] ^ in2[124];
    assign G[120] = in[123] & in2[123];
    assign P[120] = in[123] ^ in2[123];
    assign G[121] = in[122] & in2[122];
    assign P[121] = in[122] ^ in2[122];
    assign G[122] = in[121] & in2[121];
    assign P[122] = in[121] ^ in2[121];
    assign G[123] = in[120] & in2[120];
    assign P[123] = in[120] ^ in2[120];
    assign G[124] = in[119] & in2[119];
    assign P[124] = in[119] ^ in2[119];
    assign G[125] = in[118] & in2[118];
    assign P[125] = in[118] ^ in2[118];
    assign G[126] = in[117] & in2[117];
    assign P[126] = in[117] ^ in2[117];
    assign G[127] = in[116] & in2[116];
    assign P[127] = in[116] ^ in2[116];
    assign G[128] = in[115] & in2[115];
    assign P[128] = in[115] ^ in2[115];
    assign G[129] = in[114] & in2[114];
    assign P[129] = in[114] ^ in2[114];
    assign G[130] = in[113] & in2[113];
    assign P[130] = in[113] ^ in2[113];
    assign G[131] = in[112] & in2[112];
    assign P[131] = in[112] ^ in2[112];
    assign G[132] = in[111] & in2[111];
    assign P[132] = in[111] ^ in2[111];
    assign G[133] = in[110] & in2[110];
    assign P[133] = in[110] ^ in2[110];
    assign G[134] = in[109] & in2[109];
    assign P[134] = in[109] ^ in2[109];
    assign G[135] = in[108] & in2[108];
    assign P[135] = in[108] ^ in2[108];
    assign G[136] = in[107] & in2[107];
    assign P[136] = in[107] ^ in2[107];
    assign G[137] = in[106] & in2[106];
    assign P[137] = in[106] ^ in2[106];
    assign G[138] = in[105] & in2[105];
    assign P[138] = in[105] ^ in2[105];
    assign G[139] = in[104] & in2[104];
    assign P[139] = in[104] ^ in2[104];
    assign G[140] = in[103] & in2[103];
    assign P[140] = in[103] ^ in2[103];
    assign G[141] = in[102] & in2[102];
    assign P[141] = in[102] ^ in2[102];
    assign G[142] = in[101] & in2[101];
    assign P[142] = in[101] ^ in2[101];
    assign G[143] = in[100] & in2[100];
    assign P[143] = in[100] ^ in2[100];
    assign G[144] = in[99] & in2[99];
    assign P[144] = in[99] ^ in2[99];
    assign G[145] = in[98] & in2[98];
    assign P[145] = in[98] ^ in2[98];
    assign G[146] = in[97] & in2[97];
    assign P[146] = in[97] ^ in2[97];
    assign G[147] = in[96] & in2[96];
    assign P[147] = in[96] ^ in2[96];
    assign G[148] = in[95] & in2[95];
    assign P[148] = in[95] ^ in2[95];
    assign G[149] = in[94] & in2[94];
    assign P[149] = in[94] ^ in2[94];
    assign G[150] = in[93] & in2[93];
    assign P[150] = in[93] ^ in2[93];
    assign G[151] = in[92] & in2[92];
    assign P[151] = in[92] ^ in2[92];
    assign G[152] = in[91] & in2[91];
    assign P[152] = in[91] ^ in2[91];
    assign G[153] = in[90] & in2[90];
    assign P[153] = in[90] ^ in2[90];
    assign G[154] = in[89] & in2[89];
    assign P[154] = in[89] ^ in2[89];
    assign G[155] = in[88] & in2[88];
    assign P[155] = in[88] ^ in2[88];
    assign G[156] = in[87] & in2[87];
    assign P[156] = in[87] ^ in2[87];
    assign G[157] = in[86] & in2[86];
    assign P[157] = in[86] ^ in2[86];
    assign G[158] = in[85] & in2[85];
    assign P[158] = in[85] ^ in2[85];
    assign G[159] = in[84] & in2[84];
    assign P[159] = in[84] ^ in2[84];
    assign G[160] = in[83] & in2[83];
    assign P[160] = in[83] ^ in2[83];
    assign G[161] = in[82] & in2[82];
    assign P[161] = in[82] ^ in2[82];
    assign G[162] = in[81] & in2[81];
    assign P[162] = in[81] ^ in2[81];
    assign G[163] = in[80] & in2[80];
    assign P[163] = in[80] ^ in2[80];
    assign G[164] = in[79] & in2[79];
    assign P[164] = in[79] ^ in2[79];
    assign G[165] = in[78] & in2[78];
    assign P[165] = in[78] ^ in2[78];
    assign G[166] = in[77] & in2[77];
    assign P[166] = in[77] ^ in2[77];
    assign G[167] = in[76] & in2[76];
    assign P[167] = in[76] ^ in2[76];
    assign G[168] = in[75] & in2[75];
    assign P[168] = in[75] ^ in2[75];
    assign G[169] = in[74] & in2[74];
    assign P[169] = in[74] ^ in2[74];
    assign G[170] = in[73] & in2[73];
    assign P[170] = in[73] ^ in2[73];
    assign G[171] = in[72] & in2[72];
    assign P[171] = in[72] ^ in2[72];
    assign G[172] = in[71] & in2[71];
    assign P[172] = in[71] ^ in2[71];
    assign G[173] = in[70] & in2[70];
    assign P[173] = in[70] ^ in2[70];
    assign G[174] = in[69] & in2[69];
    assign P[174] = in[69] ^ in2[69];
    assign G[175] = in[68] & in2[68];
    assign P[175] = in[68] ^ in2[68];
    assign G[176] = in[67] & in2[67];
    assign P[176] = in[67] ^ in2[67];
    assign G[177] = in[66] & in2[66];
    assign P[177] = in[66] ^ in2[66];
    assign G[178] = in[65] & in2[65];
    assign P[178] = in[65] ^ in2[65];
    assign G[179] = in[64] & in2[64];
    assign P[179] = in[64] ^ in2[64];
    assign G[180] = in[63] & in2[63];
    assign P[180] = in[63] ^ in2[63];
    assign G[181] = in[62] & in2[62];
    assign P[181] = in[62] ^ in2[62];
    assign G[182] = in[61] & in2[61];
    assign P[182] = in[61] ^ in2[61];
    assign G[183] = in[60] & in2[60];
    assign P[183] = in[60] ^ in2[60];
    assign G[184] = in[59] & in2[59];
    assign P[184] = in[59] ^ in2[59];
    assign G[185] = in[58] & in2[58];
    assign P[185] = in[58] ^ in2[58];
    assign G[186] = in[57] & in2[57];
    assign P[186] = in[57] ^ in2[57];
    assign G[187] = in[56] & in2[56];
    assign P[187] = in[56] ^ in2[56];
    assign G[188] = in[55] & in2[55];
    assign P[188] = in[55] ^ in2[55];
    assign G[189] = in[54] & in2[54];
    assign P[189] = in[54] ^ in2[54];
    assign G[190] = in[53] & in2[53];
    assign P[190] = in[53] ^ in2[53];
    assign G[191] = in[52] & in2[52];
    assign P[191] = in[52] ^ in2[52];
    assign G[192] = in[51] & in2[51];
    assign P[192] = in[51] ^ in2[51];
    assign G[193] = in[50] & in2[50];
    assign P[193] = in[50] ^ in2[50];
    assign G[194] = in[49] & in2[49];
    assign P[194] = in[49] ^ in2[49];
    assign G[195] = in[48] & in2[48];
    assign P[195] = in[48] ^ in2[48];
    assign G[196] = in[47] & in2[47];
    assign P[196] = in[47] ^ in2[47];
    assign G[197] = in[46] & in2[46];
    assign P[197] = in[46] ^ in2[46];
    assign G[198] = in[45] & in2[45];
    assign P[198] = in[45] ^ in2[45];
    assign G[199] = in[44] & in2[44];
    assign P[199] = in[44] ^ in2[44];
    assign G[200] = in[43] & in2[43];
    assign P[200] = in[43] ^ in2[43];
    assign G[201] = in[42] & in2[42];
    assign P[201] = in[42] ^ in2[42];
    assign G[202] = in[41] & in2[41];
    assign P[202] = in[41] ^ in2[41];
    assign G[203] = in[40] & in2[40];
    assign P[203] = in[40] ^ in2[40];
    assign G[204] = in[39] & in2[39];
    assign P[204] = in[39] ^ in2[39];
    assign G[205] = in[38] & in2[38];
    assign P[205] = in[38] ^ in2[38];
    assign G[206] = in[37] & in2[37];
    assign P[206] = in[37] ^ in2[37];
    assign G[207] = in[36] & in2[36];
    assign P[207] = in[36] ^ in2[36];
    assign G[208] = in[35] & in2[35];
    assign P[208] = in[35] ^ in2[35];
    assign G[209] = in[34] & in2[34];
    assign P[209] = in[34] ^ in2[34];
    assign G[210] = in[33] & in2[33];
    assign P[210] = in[33] ^ in2[33];
    assign G[211] = in[32] & in2[32];
    assign P[211] = in[32] ^ in2[32];
    assign G[212] = in[31] & in2[31];
    assign P[212] = in[31] ^ in2[31];
    assign G[213] = in[30] & in2[30];
    assign P[213] = in[30] ^ in2[30];
    assign G[214] = in[29] & in2[29];
    assign P[214] = in[29] ^ in2[29];
    assign G[215] = in[28] & in2[28];
    assign P[215] = in[28] ^ in2[28];
    assign G[216] = in[27] & in2[27];
    assign P[216] = in[27] ^ in2[27];
    assign G[217] = in[26] & in2[26];
    assign P[217] = in[26] ^ in2[26];
    assign G[218] = in[25] & in2[25];
    assign P[218] = in[25] ^ in2[25];
    assign G[219] = in[24] & in2[24];
    assign P[219] = in[24] ^ in2[24];
    assign G[220] = in[23] & in2[23];
    assign P[220] = in[23] ^ in2[23];
    assign G[221] = in[22] & in2[22];
    assign P[221] = in[22] ^ in2[22];
    assign G[222] = in[21] & in2[21];
    assign P[222] = in[21] ^ in2[21];
    assign G[223] = in[20] & in2[20];
    assign P[223] = in[20] ^ in2[20];
    assign G[224] = in[19] & in2[19];
    assign P[224] = in[19] ^ in2[19];
    assign G[225] = in[18] & in2[18];
    assign P[225] = in[18] ^ in2[18];
    assign G[226] = in[17] & in2[17];
    assign P[226] = in[17] ^ in2[17];
    assign G[227] = in[16] & in2[16];
    assign P[227] = in[16] ^ in2[16];
    assign G[228] = in[15] & in2[15];
    assign P[228] = in[15] ^ in2[15];
    assign G[229] = in[14] & in2[14];
    assign P[229] = in[14] ^ in2[14];
    assign G[230] = in[13] & in2[13];
    assign P[230] = in[13] ^ in2[13];
    assign G[231] = in[12] & in2[12];
    assign P[231] = in[12] ^ in2[12];
    assign G[232] = in[11] & in2[11];
    assign P[232] = in[11] ^ in2[11];
    assign G[233] = in[10] & in2[10];
    assign P[233] = in[10] ^ in2[10];
    assign G[234] = in[9] & in2[9];
    assign P[234] = in[9] ^ in2[9];
    assign G[235] = in[8] & in2[8];
    assign P[235] = in[8] ^ in2[8];
    assign G[236] = in[7] & in2[7];
    assign P[236] = in[7] ^ in2[7];
    assign G[237] = in[6] & in2[6];
    assign P[237] = in[6] ^ in2[6];
    assign G[238] = in[5] & in2[5];
    assign P[238] = in[5] ^ in2[5];
    assign G[239] = in[4] & in2[4];
    assign P[239] = in[4] ^ in2[4];
    assign G[240] = in[3] & in2[3];
    assign P[240] = in[3] ^ in2[3];
    assign G[241] = in[2] & in2[2];
    assign P[241] = in[2] ^ in2[2];
    assign G[242] = in[1] & in2[1];
    assign P[242] = in[1] ^ in2[1];
    assign G[243] = in[0] & in2[0];
    assign P[243] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign C[243] = G[242] | (P[242] & C[242]);
    assign cout = G[243] | (P[243] & C[243]);
    assign sum = P ^ C;
endmodule

module CLA243(output [242:0] sum, output cout, input [242:0] in1, input [242:0] in2;

    wire[242:0] G;
    wire[242:0] C;
    wire[242:0] P;

    assign G[0] = in[242] & in2[242];
    assign P[0] = in[242] ^ in2[242];
    assign G[1] = in[241] & in2[241];
    assign P[1] = in[241] ^ in2[241];
    assign G[2] = in[240] & in2[240];
    assign P[2] = in[240] ^ in2[240];
    assign G[3] = in[239] & in2[239];
    assign P[3] = in[239] ^ in2[239];
    assign G[4] = in[238] & in2[238];
    assign P[4] = in[238] ^ in2[238];
    assign G[5] = in[237] & in2[237];
    assign P[5] = in[237] ^ in2[237];
    assign G[6] = in[236] & in2[236];
    assign P[6] = in[236] ^ in2[236];
    assign G[7] = in[235] & in2[235];
    assign P[7] = in[235] ^ in2[235];
    assign G[8] = in[234] & in2[234];
    assign P[8] = in[234] ^ in2[234];
    assign G[9] = in[233] & in2[233];
    assign P[9] = in[233] ^ in2[233];
    assign G[10] = in[232] & in2[232];
    assign P[10] = in[232] ^ in2[232];
    assign G[11] = in[231] & in2[231];
    assign P[11] = in[231] ^ in2[231];
    assign G[12] = in[230] & in2[230];
    assign P[12] = in[230] ^ in2[230];
    assign G[13] = in[229] & in2[229];
    assign P[13] = in[229] ^ in2[229];
    assign G[14] = in[228] & in2[228];
    assign P[14] = in[228] ^ in2[228];
    assign G[15] = in[227] & in2[227];
    assign P[15] = in[227] ^ in2[227];
    assign G[16] = in[226] & in2[226];
    assign P[16] = in[226] ^ in2[226];
    assign G[17] = in[225] & in2[225];
    assign P[17] = in[225] ^ in2[225];
    assign G[18] = in[224] & in2[224];
    assign P[18] = in[224] ^ in2[224];
    assign G[19] = in[223] & in2[223];
    assign P[19] = in[223] ^ in2[223];
    assign G[20] = in[222] & in2[222];
    assign P[20] = in[222] ^ in2[222];
    assign G[21] = in[221] & in2[221];
    assign P[21] = in[221] ^ in2[221];
    assign G[22] = in[220] & in2[220];
    assign P[22] = in[220] ^ in2[220];
    assign G[23] = in[219] & in2[219];
    assign P[23] = in[219] ^ in2[219];
    assign G[24] = in[218] & in2[218];
    assign P[24] = in[218] ^ in2[218];
    assign G[25] = in[217] & in2[217];
    assign P[25] = in[217] ^ in2[217];
    assign G[26] = in[216] & in2[216];
    assign P[26] = in[216] ^ in2[216];
    assign G[27] = in[215] & in2[215];
    assign P[27] = in[215] ^ in2[215];
    assign G[28] = in[214] & in2[214];
    assign P[28] = in[214] ^ in2[214];
    assign G[29] = in[213] & in2[213];
    assign P[29] = in[213] ^ in2[213];
    assign G[30] = in[212] & in2[212];
    assign P[30] = in[212] ^ in2[212];
    assign G[31] = in[211] & in2[211];
    assign P[31] = in[211] ^ in2[211];
    assign G[32] = in[210] & in2[210];
    assign P[32] = in[210] ^ in2[210];
    assign G[33] = in[209] & in2[209];
    assign P[33] = in[209] ^ in2[209];
    assign G[34] = in[208] & in2[208];
    assign P[34] = in[208] ^ in2[208];
    assign G[35] = in[207] & in2[207];
    assign P[35] = in[207] ^ in2[207];
    assign G[36] = in[206] & in2[206];
    assign P[36] = in[206] ^ in2[206];
    assign G[37] = in[205] & in2[205];
    assign P[37] = in[205] ^ in2[205];
    assign G[38] = in[204] & in2[204];
    assign P[38] = in[204] ^ in2[204];
    assign G[39] = in[203] & in2[203];
    assign P[39] = in[203] ^ in2[203];
    assign G[40] = in[202] & in2[202];
    assign P[40] = in[202] ^ in2[202];
    assign G[41] = in[201] & in2[201];
    assign P[41] = in[201] ^ in2[201];
    assign G[42] = in[200] & in2[200];
    assign P[42] = in[200] ^ in2[200];
    assign G[43] = in[199] & in2[199];
    assign P[43] = in[199] ^ in2[199];
    assign G[44] = in[198] & in2[198];
    assign P[44] = in[198] ^ in2[198];
    assign G[45] = in[197] & in2[197];
    assign P[45] = in[197] ^ in2[197];
    assign G[46] = in[196] & in2[196];
    assign P[46] = in[196] ^ in2[196];
    assign G[47] = in[195] & in2[195];
    assign P[47] = in[195] ^ in2[195];
    assign G[48] = in[194] & in2[194];
    assign P[48] = in[194] ^ in2[194];
    assign G[49] = in[193] & in2[193];
    assign P[49] = in[193] ^ in2[193];
    assign G[50] = in[192] & in2[192];
    assign P[50] = in[192] ^ in2[192];
    assign G[51] = in[191] & in2[191];
    assign P[51] = in[191] ^ in2[191];
    assign G[52] = in[190] & in2[190];
    assign P[52] = in[190] ^ in2[190];
    assign G[53] = in[189] & in2[189];
    assign P[53] = in[189] ^ in2[189];
    assign G[54] = in[188] & in2[188];
    assign P[54] = in[188] ^ in2[188];
    assign G[55] = in[187] & in2[187];
    assign P[55] = in[187] ^ in2[187];
    assign G[56] = in[186] & in2[186];
    assign P[56] = in[186] ^ in2[186];
    assign G[57] = in[185] & in2[185];
    assign P[57] = in[185] ^ in2[185];
    assign G[58] = in[184] & in2[184];
    assign P[58] = in[184] ^ in2[184];
    assign G[59] = in[183] & in2[183];
    assign P[59] = in[183] ^ in2[183];
    assign G[60] = in[182] & in2[182];
    assign P[60] = in[182] ^ in2[182];
    assign G[61] = in[181] & in2[181];
    assign P[61] = in[181] ^ in2[181];
    assign G[62] = in[180] & in2[180];
    assign P[62] = in[180] ^ in2[180];
    assign G[63] = in[179] & in2[179];
    assign P[63] = in[179] ^ in2[179];
    assign G[64] = in[178] & in2[178];
    assign P[64] = in[178] ^ in2[178];
    assign G[65] = in[177] & in2[177];
    assign P[65] = in[177] ^ in2[177];
    assign G[66] = in[176] & in2[176];
    assign P[66] = in[176] ^ in2[176];
    assign G[67] = in[175] & in2[175];
    assign P[67] = in[175] ^ in2[175];
    assign G[68] = in[174] & in2[174];
    assign P[68] = in[174] ^ in2[174];
    assign G[69] = in[173] & in2[173];
    assign P[69] = in[173] ^ in2[173];
    assign G[70] = in[172] & in2[172];
    assign P[70] = in[172] ^ in2[172];
    assign G[71] = in[171] & in2[171];
    assign P[71] = in[171] ^ in2[171];
    assign G[72] = in[170] & in2[170];
    assign P[72] = in[170] ^ in2[170];
    assign G[73] = in[169] & in2[169];
    assign P[73] = in[169] ^ in2[169];
    assign G[74] = in[168] & in2[168];
    assign P[74] = in[168] ^ in2[168];
    assign G[75] = in[167] & in2[167];
    assign P[75] = in[167] ^ in2[167];
    assign G[76] = in[166] & in2[166];
    assign P[76] = in[166] ^ in2[166];
    assign G[77] = in[165] & in2[165];
    assign P[77] = in[165] ^ in2[165];
    assign G[78] = in[164] & in2[164];
    assign P[78] = in[164] ^ in2[164];
    assign G[79] = in[163] & in2[163];
    assign P[79] = in[163] ^ in2[163];
    assign G[80] = in[162] & in2[162];
    assign P[80] = in[162] ^ in2[162];
    assign G[81] = in[161] & in2[161];
    assign P[81] = in[161] ^ in2[161];
    assign G[82] = in[160] & in2[160];
    assign P[82] = in[160] ^ in2[160];
    assign G[83] = in[159] & in2[159];
    assign P[83] = in[159] ^ in2[159];
    assign G[84] = in[158] & in2[158];
    assign P[84] = in[158] ^ in2[158];
    assign G[85] = in[157] & in2[157];
    assign P[85] = in[157] ^ in2[157];
    assign G[86] = in[156] & in2[156];
    assign P[86] = in[156] ^ in2[156];
    assign G[87] = in[155] & in2[155];
    assign P[87] = in[155] ^ in2[155];
    assign G[88] = in[154] & in2[154];
    assign P[88] = in[154] ^ in2[154];
    assign G[89] = in[153] & in2[153];
    assign P[89] = in[153] ^ in2[153];
    assign G[90] = in[152] & in2[152];
    assign P[90] = in[152] ^ in2[152];
    assign G[91] = in[151] & in2[151];
    assign P[91] = in[151] ^ in2[151];
    assign G[92] = in[150] & in2[150];
    assign P[92] = in[150] ^ in2[150];
    assign G[93] = in[149] & in2[149];
    assign P[93] = in[149] ^ in2[149];
    assign G[94] = in[148] & in2[148];
    assign P[94] = in[148] ^ in2[148];
    assign G[95] = in[147] & in2[147];
    assign P[95] = in[147] ^ in2[147];
    assign G[96] = in[146] & in2[146];
    assign P[96] = in[146] ^ in2[146];
    assign G[97] = in[145] & in2[145];
    assign P[97] = in[145] ^ in2[145];
    assign G[98] = in[144] & in2[144];
    assign P[98] = in[144] ^ in2[144];
    assign G[99] = in[143] & in2[143];
    assign P[99] = in[143] ^ in2[143];
    assign G[100] = in[142] & in2[142];
    assign P[100] = in[142] ^ in2[142];
    assign G[101] = in[141] & in2[141];
    assign P[101] = in[141] ^ in2[141];
    assign G[102] = in[140] & in2[140];
    assign P[102] = in[140] ^ in2[140];
    assign G[103] = in[139] & in2[139];
    assign P[103] = in[139] ^ in2[139];
    assign G[104] = in[138] & in2[138];
    assign P[104] = in[138] ^ in2[138];
    assign G[105] = in[137] & in2[137];
    assign P[105] = in[137] ^ in2[137];
    assign G[106] = in[136] & in2[136];
    assign P[106] = in[136] ^ in2[136];
    assign G[107] = in[135] & in2[135];
    assign P[107] = in[135] ^ in2[135];
    assign G[108] = in[134] & in2[134];
    assign P[108] = in[134] ^ in2[134];
    assign G[109] = in[133] & in2[133];
    assign P[109] = in[133] ^ in2[133];
    assign G[110] = in[132] & in2[132];
    assign P[110] = in[132] ^ in2[132];
    assign G[111] = in[131] & in2[131];
    assign P[111] = in[131] ^ in2[131];
    assign G[112] = in[130] & in2[130];
    assign P[112] = in[130] ^ in2[130];
    assign G[113] = in[129] & in2[129];
    assign P[113] = in[129] ^ in2[129];
    assign G[114] = in[128] & in2[128];
    assign P[114] = in[128] ^ in2[128];
    assign G[115] = in[127] & in2[127];
    assign P[115] = in[127] ^ in2[127];
    assign G[116] = in[126] & in2[126];
    assign P[116] = in[126] ^ in2[126];
    assign G[117] = in[125] & in2[125];
    assign P[117] = in[125] ^ in2[125];
    assign G[118] = in[124] & in2[124];
    assign P[118] = in[124] ^ in2[124];
    assign G[119] = in[123] & in2[123];
    assign P[119] = in[123] ^ in2[123];
    assign G[120] = in[122] & in2[122];
    assign P[120] = in[122] ^ in2[122];
    assign G[121] = in[121] & in2[121];
    assign P[121] = in[121] ^ in2[121];
    assign G[122] = in[120] & in2[120];
    assign P[122] = in[120] ^ in2[120];
    assign G[123] = in[119] & in2[119];
    assign P[123] = in[119] ^ in2[119];
    assign G[124] = in[118] & in2[118];
    assign P[124] = in[118] ^ in2[118];
    assign G[125] = in[117] & in2[117];
    assign P[125] = in[117] ^ in2[117];
    assign G[126] = in[116] & in2[116];
    assign P[126] = in[116] ^ in2[116];
    assign G[127] = in[115] & in2[115];
    assign P[127] = in[115] ^ in2[115];
    assign G[128] = in[114] & in2[114];
    assign P[128] = in[114] ^ in2[114];
    assign G[129] = in[113] & in2[113];
    assign P[129] = in[113] ^ in2[113];
    assign G[130] = in[112] & in2[112];
    assign P[130] = in[112] ^ in2[112];
    assign G[131] = in[111] & in2[111];
    assign P[131] = in[111] ^ in2[111];
    assign G[132] = in[110] & in2[110];
    assign P[132] = in[110] ^ in2[110];
    assign G[133] = in[109] & in2[109];
    assign P[133] = in[109] ^ in2[109];
    assign G[134] = in[108] & in2[108];
    assign P[134] = in[108] ^ in2[108];
    assign G[135] = in[107] & in2[107];
    assign P[135] = in[107] ^ in2[107];
    assign G[136] = in[106] & in2[106];
    assign P[136] = in[106] ^ in2[106];
    assign G[137] = in[105] & in2[105];
    assign P[137] = in[105] ^ in2[105];
    assign G[138] = in[104] & in2[104];
    assign P[138] = in[104] ^ in2[104];
    assign G[139] = in[103] & in2[103];
    assign P[139] = in[103] ^ in2[103];
    assign G[140] = in[102] & in2[102];
    assign P[140] = in[102] ^ in2[102];
    assign G[141] = in[101] & in2[101];
    assign P[141] = in[101] ^ in2[101];
    assign G[142] = in[100] & in2[100];
    assign P[142] = in[100] ^ in2[100];
    assign G[143] = in[99] & in2[99];
    assign P[143] = in[99] ^ in2[99];
    assign G[144] = in[98] & in2[98];
    assign P[144] = in[98] ^ in2[98];
    assign G[145] = in[97] & in2[97];
    assign P[145] = in[97] ^ in2[97];
    assign G[146] = in[96] & in2[96];
    assign P[146] = in[96] ^ in2[96];
    assign G[147] = in[95] & in2[95];
    assign P[147] = in[95] ^ in2[95];
    assign G[148] = in[94] & in2[94];
    assign P[148] = in[94] ^ in2[94];
    assign G[149] = in[93] & in2[93];
    assign P[149] = in[93] ^ in2[93];
    assign G[150] = in[92] & in2[92];
    assign P[150] = in[92] ^ in2[92];
    assign G[151] = in[91] & in2[91];
    assign P[151] = in[91] ^ in2[91];
    assign G[152] = in[90] & in2[90];
    assign P[152] = in[90] ^ in2[90];
    assign G[153] = in[89] & in2[89];
    assign P[153] = in[89] ^ in2[89];
    assign G[154] = in[88] & in2[88];
    assign P[154] = in[88] ^ in2[88];
    assign G[155] = in[87] & in2[87];
    assign P[155] = in[87] ^ in2[87];
    assign G[156] = in[86] & in2[86];
    assign P[156] = in[86] ^ in2[86];
    assign G[157] = in[85] & in2[85];
    assign P[157] = in[85] ^ in2[85];
    assign G[158] = in[84] & in2[84];
    assign P[158] = in[84] ^ in2[84];
    assign G[159] = in[83] & in2[83];
    assign P[159] = in[83] ^ in2[83];
    assign G[160] = in[82] & in2[82];
    assign P[160] = in[82] ^ in2[82];
    assign G[161] = in[81] & in2[81];
    assign P[161] = in[81] ^ in2[81];
    assign G[162] = in[80] & in2[80];
    assign P[162] = in[80] ^ in2[80];
    assign G[163] = in[79] & in2[79];
    assign P[163] = in[79] ^ in2[79];
    assign G[164] = in[78] & in2[78];
    assign P[164] = in[78] ^ in2[78];
    assign G[165] = in[77] & in2[77];
    assign P[165] = in[77] ^ in2[77];
    assign G[166] = in[76] & in2[76];
    assign P[166] = in[76] ^ in2[76];
    assign G[167] = in[75] & in2[75];
    assign P[167] = in[75] ^ in2[75];
    assign G[168] = in[74] & in2[74];
    assign P[168] = in[74] ^ in2[74];
    assign G[169] = in[73] & in2[73];
    assign P[169] = in[73] ^ in2[73];
    assign G[170] = in[72] & in2[72];
    assign P[170] = in[72] ^ in2[72];
    assign G[171] = in[71] & in2[71];
    assign P[171] = in[71] ^ in2[71];
    assign G[172] = in[70] & in2[70];
    assign P[172] = in[70] ^ in2[70];
    assign G[173] = in[69] & in2[69];
    assign P[173] = in[69] ^ in2[69];
    assign G[174] = in[68] & in2[68];
    assign P[174] = in[68] ^ in2[68];
    assign G[175] = in[67] & in2[67];
    assign P[175] = in[67] ^ in2[67];
    assign G[176] = in[66] & in2[66];
    assign P[176] = in[66] ^ in2[66];
    assign G[177] = in[65] & in2[65];
    assign P[177] = in[65] ^ in2[65];
    assign G[178] = in[64] & in2[64];
    assign P[178] = in[64] ^ in2[64];
    assign G[179] = in[63] & in2[63];
    assign P[179] = in[63] ^ in2[63];
    assign G[180] = in[62] & in2[62];
    assign P[180] = in[62] ^ in2[62];
    assign G[181] = in[61] & in2[61];
    assign P[181] = in[61] ^ in2[61];
    assign G[182] = in[60] & in2[60];
    assign P[182] = in[60] ^ in2[60];
    assign G[183] = in[59] & in2[59];
    assign P[183] = in[59] ^ in2[59];
    assign G[184] = in[58] & in2[58];
    assign P[184] = in[58] ^ in2[58];
    assign G[185] = in[57] & in2[57];
    assign P[185] = in[57] ^ in2[57];
    assign G[186] = in[56] & in2[56];
    assign P[186] = in[56] ^ in2[56];
    assign G[187] = in[55] & in2[55];
    assign P[187] = in[55] ^ in2[55];
    assign G[188] = in[54] & in2[54];
    assign P[188] = in[54] ^ in2[54];
    assign G[189] = in[53] & in2[53];
    assign P[189] = in[53] ^ in2[53];
    assign G[190] = in[52] & in2[52];
    assign P[190] = in[52] ^ in2[52];
    assign G[191] = in[51] & in2[51];
    assign P[191] = in[51] ^ in2[51];
    assign G[192] = in[50] & in2[50];
    assign P[192] = in[50] ^ in2[50];
    assign G[193] = in[49] & in2[49];
    assign P[193] = in[49] ^ in2[49];
    assign G[194] = in[48] & in2[48];
    assign P[194] = in[48] ^ in2[48];
    assign G[195] = in[47] & in2[47];
    assign P[195] = in[47] ^ in2[47];
    assign G[196] = in[46] & in2[46];
    assign P[196] = in[46] ^ in2[46];
    assign G[197] = in[45] & in2[45];
    assign P[197] = in[45] ^ in2[45];
    assign G[198] = in[44] & in2[44];
    assign P[198] = in[44] ^ in2[44];
    assign G[199] = in[43] & in2[43];
    assign P[199] = in[43] ^ in2[43];
    assign G[200] = in[42] & in2[42];
    assign P[200] = in[42] ^ in2[42];
    assign G[201] = in[41] & in2[41];
    assign P[201] = in[41] ^ in2[41];
    assign G[202] = in[40] & in2[40];
    assign P[202] = in[40] ^ in2[40];
    assign G[203] = in[39] & in2[39];
    assign P[203] = in[39] ^ in2[39];
    assign G[204] = in[38] & in2[38];
    assign P[204] = in[38] ^ in2[38];
    assign G[205] = in[37] & in2[37];
    assign P[205] = in[37] ^ in2[37];
    assign G[206] = in[36] & in2[36];
    assign P[206] = in[36] ^ in2[36];
    assign G[207] = in[35] & in2[35];
    assign P[207] = in[35] ^ in2[35];
    assign G[208] = in[34] & in2[34];
    assign P[208] = in[34] ^ in2[34];
    assign G[209] = in[33] & in2[33];
    assign P[209] = in[33] ^ in2[33];
    assign G[210] = in[32] & in2[32];
    assign P[210] = in[32] ^ in2[32];
    assign G[211] = in[31] & in2[31];
    assign P[211] = in[31] ^ in2[31];
    assign G[212] = in[30] & in2[30];
    assign P[212] = in[30] ^ in2[30];
    assign G[213] = in[29] & in2[29];
    assign P[213] = in[29] ^ in2[29];
    assign G[214] = in[28] & in2[28];
    assign P[214] = in[28] ^ in2[28];
    assign G[215] = in[27] & in2[27];
    assign P[215] = in[27] ^ in2[27];
    assign G[216] = in[26] & in2[26];
    assign P[216] = in[26] ^ in2[26];
    assign G[217] = in[25] & in2[25];
    assign P[217] = in[25] ^ in2[25];
    assign G[218] = in[24] & in2[24];
    assign P[218] = in[24] ^ in2[24];
    assign G[219] = in[23] & in2[23];
    assign P[219] = in[23] ^ in2[23];
    assign G[220] = in[22] & in2[22];
    assign P[220] = in[22] ^ in2[22];
    assign G[221] = in[21] & in2[21];
    assign P[221] = in[21] ^ in2[21];
    assign G[222] = in[20] & in2[20];
    assign P[222] = in[20] ^ in2[20];
    assign G[223] = in[19] & in2[19];
    assign P[223] = in[19] ^ in2[19];
    assign G[224] = in[18] & in2[18];
    assign P[224] = in[18] ^ in2[18];
    assign G[225] = in[17] & in2[17];
    assign P[225] = in[17] ^ in2[17];
    assign G[226] = in[16] & in2[16];
    assign P[226] = in[16] ^ in2[16];
    assign G[227] = in[15] & in2[15];
    assign P[227] = in[15] ^ in2[15];
    assign G[228] = in[14] & in2[14];
    assign P[228] = in[14] ^ in2[14];
    assign G[229] = in[13] & in2[13];
    assign P[229] = in[13] ^ in2[13];
    assign G[230] = in[12] & in2[12];
    assign P[230] = in[12] ^ in2[12];
    assign G[231] = in[11] & in2[11];
    assign P[231] = in[11] ^ in2[11];
    assign G[232] = in[10] & in2[10];
    assign P[232] = in[10] ^ in2[10];
    assign G[233] = in[9] & in2[9];
    assign P[233] = in[9] ^ in2[9];
    assign G[234] = in[8] & in2[8];
    assign P[234] = in[8] ^ in2[8];
    assign G[235] = in[7] & in2[7];
    assign P[235] = in[7] ^ in2[7];
    assign G[236] = in[6] & in2[6];
    assign P[236] = in[6] ^ in2[6];
    assign G[237] = in[5] & in2[5];
    assign P[237] = in[5] ^ in2[5];
    assign G[238] = in[4] & in2[4];
    assign P[238] = in[4] ^ in2[4];
    assign G[239] = in[3] & in2[3];
    assign P[239] = in[3] ^ in2[3];
    assign G[240] = in[2] & in2[2];
    assign P[240] = in[2] ^ in2[2];
    assign G[241] = in[1] & in2[1];
    assign P[241] = in[1] ^ in2[1];
    assign G[242] = in[0] & in2[0];
    assign P[242] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign C[242] = G[241] | (P[241] & C[241]);
    assign cout = G[242] | (P[242] & C[242]);
    assign sum = P ^ C;
endmodule

module CLA242(output [241:0] sum, output cout, input [241:0] in1, input [241:0] in2;

    wire[241:0] G;
    wire[241:0] C;
    wire[241:0] P;

    assign G[0] = in[241] & in2[241];
    assign P[0] = in[241] ^ in2[241];
    assign G[1] = in[240] & in2[240];
    assign P[1] = in[240] ^ in2[240];
    assign G[2] = in[239] & in2[239];
    assign P[2] = in[239] ^ in2[239];
    assign G[3] = in[238] & in2[238];
    assign P[3] = in[238] ^ in2[238];
    assign G[4] = in[237] & in2[237];
    assign P[4] = in[237] ^ in2[237];
    assign G[5] = in[236] & in2[236];
    assign P[5] = in[236] ^ in2[236];
    assign G[6] = in[235] & in2[235];
    assign P[6] = in[235] ^ in2[235];
    assign G[7] = in[234] & in2[234];
    assign P[7] = in[234] ^ in2[234];
    assign G[8] = in[233] & in2[233];
    assign P[8] = in[233] ^ in2[233];
    assign G[9] = in[232] & in2[232];
    assign P[9] = in[232] ^ in2[232];
    assign G[10] = in[231] & in2[231];
    assign P[10] = in[231] ^ in2[231];
    assign G[11] = in[230] & in2[230];
    assign P[11] = in[230] ^ in2[230];
    assign G[12] = in[229] & in2[229];
    assign P[12] = in[229] ^ in2[229];
    assign G[13] = in[228] & in2[228];
    assign P[13] = in[228] ^ in2[228];
    assign G[14] = in[227] & in2[227];
    assign P[14] = in[227] ^ in2[227];
    assign G[15] = in[226] & in2[226];
    assign P[15] = in[226] ^ in2[226];
    assign G[16] = in[225] & in2[225];
    assign P[16] = in[225] ^ in2[225];
    assign G[17] = in[224] & in2[224];
    assign P[17] = in[224] ^ in2[224];
    assign G[18] = in[223] & in2[223];
    assign P[18] = in[223] ^ in2[223];
    assign G[19] = in[222] & in2[222];
    assign P[19] = in[222] ^ in2[222];
    assign G[20] = in[221] & in2[221];
    assign P[20] = in[221] ^ in2[221];
    assign G[21] = in[220] & in2[220];
    assign P[21] = in[220] ^ in2[220];
    assign G[22] = in[219] & in2[219];
    assign P[22] = in[219] ^ in2[219];
    assign G[23] = in[218] & in2[218];
    assign P[23] = in[218] ^ in2[218];
    assign G[24] = in[217] & in2[217];
    assign P[24] = in[217] ^ in2[217];
    assign G[25] = in[216] & in2[216];
    assign P[25] = in[216] ^ in2[216];
    assign G[26] = in[215] & in2[215];
    assign P[26] = in[215] ^ in2[215];
    assign G[27] = in[214] & in2[214];
    assign P[27] = in[214] ^ in2[214];
    assign G[28] = in[213] & in2[213];
    assign P[28] = in[213] ^ in2[213];
    assign G[29] = in[212] & in2[212];
    assign P[29] = in[212] ^ in2[212];
    assign G[30] = in[211] & in2[211];
    assign P[30] = in[211] ^ in2[211];
    assign G[31] = in[210] & in2[210];
    assign P[31] = in[210] ^ in2[210];
    assign G[32] = in[209] & in2[209];
    assign P[32] = in[209] ^ in2[209];
    assign G[33] = in[208] & in2[208];
    assign P[33] = in[208] ^ in2[208];
    assign G[34] = in[207] & in2[207];
    assign P[34] = in[207] ^ in2[207];
    assign G[35] = in[206] & in2[206];
    assign P[35] = in[206] ^ in2[206];
    assign G[36] = in[205] & in2[205];
    assign P[36] = in[205] ^ in2[205];
    assign G[37] = in[204] & in2[204];
    assign P[37] = in[204] ^ in2[204];
    assign G[38] = in[203] & in2[203];
    assign P[38] = in[203] ^ in2[203];
    assign G[39] = in[202] & in2[202];
    assign P[39] = in[202] ^ in2[202];
    assign G[40] = in[201] & in2[201];
    assign P[40] = in[201] ^ in2[201];
    assign G[41] = in[200] & in2[200];
    assign P[41] = in[200] ^ in2[200];
    assign G[42] = in[199] & in2[199];
    assign P[42] = in[199] ^ in2[199];
    assign G[43] = in[198] & in2[198];
    assign P[43] = in[198] ^ in2[198];
    assign G[44] = in[197] & in2[197];
    assign P[44] = in[197] ^ in2[197];
    assign G[45] = in[196] & in2[196];
    assign P[45] = in[196] ^ in2[196];
    assign G[46] = in[195] & in2[195];
    assign P[46] = in[195] ^ in2[195];
    assign G[47] = in[194] & in2[194];
    assign P[47] = in[194] ^ in2[194];
    assign G[48] = in[193] & in2[193];
    assign P[48] = in[193] ^ in2[193];
    assign G[49] = in[192] & in2[192];
    assign P[49] = in[192] ^ in2[192];
    assign G[50] = in[191] & in2[191];
    assign P[50] = in[191] ^ in2[191];
    assign G[51] = in[190] & in2[190];
    assign P[51] = in[190] ^ in2[190];
    assign G[52] = in[189] & in2[189];
    assign P[52] = in[189] ^ in2[189];
    assign G[53] = in[188] & in2[188];
    assign P[53] = in[188] ^ in2[188];
    assign G[54] = in[187] & in2[187];
    assign P[54] = in[187] ^ in2[187];
    assign G[55] = in[186] & in2[186];
    assign P[55] = in[186] ^ in2[186];
    assign G[56] = in[185] & in2[185];
    assign P[56] = in[185] ^ in2[185];
    assign G[57] = in[184] & in2[184];
    assign P[57] = in[184] ^ in2[184];
    assign G[58] = in[183] & in2[183];
    assign P[58] = in[183] ^ in2[183];
    assign G[59] = in[182] & in2[182];
    assign P[59] = in[182] ^ in2[182];
    assign G[60] = in[181] & in2[181];
    assign P[60] = in[181] ^ in2[181];
    assign G[61] = in[180] & in2[180];
    assign P[61] = in[180] ^ in2[180];
    assign G[62] = in[179] & in2[179];
    assign P[62] = in[179] ^ in2[179];
    assign G[63] = in[178] & in2[178];
    assign P[63] = in[178] ^ in2[178];
    assign G[64] = in[177] & in2[177];
    assign P[64] = in[177] ^ in2[177];
    assign G[65] = in[176] & in2[176];
    assign P[65] = in[176] ^ in2[176];
    assign G[66] = in[175] & in2[175];
    assign P[66] = in[175] ^ in2[175];
    assign G[67] = in[174] & in2[174];
    assign P[67] = in[174] ^ in2[174];
    assign G[68] = in[173] & in2[173];
    assign P[68] = in[173] ^ in2[173];
    assign G[69] = in[172] & in2[172];
    assign P[69] = in[172] ^ in2[172];
    assign G[70] = in[171] & in2[171];
    assign P[70] = in[171] ^ in2[171];
    assign G[71] = in[170] & in2[170];
    assign P[71] = in[170] ^ in2[170];
    assign G[72] = in[169] & in2[169];
    assign P[72] = in[169] ^ in2[169];
    assign G[73] = in[168] & in2[168];
    assign P[73] = in[168] ^ in2[168];
    assign G[74] = in[167] & in2[167];
    assign P[74] = in[167] ^ in2[167];
    assign G[75] = in[166] & in2[166];
    assign P[75] = in[166] ^ in2[166];
    assign G[76] = in[165] & in2[165];
    assign P[76] = in[165] ^ in2[165];
    assign G[77] = in[164] & in2[164];
    assign P[77] = in[164] ^ in2[164];
    assign G[78] = in[163] & in2[163];
    assign P[78] = in[163] ^ in2[163];
    assign G[79] = in[162] & in2[162];
    assign P[79] = in[162] ^ in2[162];
    assign G[80] = in[161] & in2[161];
    assign P[80] = in[161] ^ in2[161];
    assign G[81] = in[160] & in2[160];
    assign P[81] = in[160] ^ in2[160];
    assign G[82] = in[159] & in2[159];
    assign P[82] = in[159] ^ in2[159];
    assign G[83] = in[158] & in2[158];
    assign P[83] = in[158] ^ in2[158];
    assign G[84] = in[157] & in2[157];
    assign P[84] = in[157] ^ in2[157];
    assign G[85] = in[156] & in2[156];
    assign P[85] = in[156] ^ in2[156];
    assign G[86] = in[155] & in2[155];
    assign P[86] = in[155] ^ in2[155];
    assign G[87] = in[154] & in2[154];
    assign P[87] = in[154] ^ in2[154];
    assign G[88] = in[153] & in2[153];
    assign P[88] = in[153] ^ in2[153];
    assign G[89] = in[152] & in2[152];
    assign P[89] = in[152] ^ in2[152];
    assign G[90] = in[151] & in2[151];
    assign P[90] = in[151] ^ in2[151];
    assign G[91] = in[150] & in2[150];
    assign P[91] = in[150] ^ in2[150];
    assign G[92] = in[149] & in2[149];
    assign P[92] = in[149] ^ in2[149];
    assign G[93] = in[148] & in2[148];
    assign P[93] = in[148] ^ in2[148];
    assign G[94] = in[147] & in2[147];
    assign P[94] = in[147] ^ in2[147];
    assign G[95] = in[146] & in2[146];
    assign P[95] = in[146] ^ in2[146];
    assign G[96] = in[145] & in2[145];
    assign P[96] = in[145] ^ in2[145];
    assign G[97] = in[144] & in2[144];
    assign P[97] = in[144] ^ in2[144];
    assign G[98] = in[143] & in2[143];
    assign P[98] = in[143] ^ in2[143];
    assign G[99] = in[142] & in2[142];
    assign P[99] = in[142] ^ in2[142];
    assign G[100] = in[141] & in2[141];
    assign P[100] = in[141] ^ in2[141];
    assign G[101] = in[140] & in2[140];
    assign P[101] = in[140] ^ in2[140];
    assign G[102] = in[139] & in2[139];
    assign P[102] = in[139] ^ in2[139];
    assign G[103] = in[138] & in2[138];
    assign P[103] = in[138] ^ in2[138];
    assign G[104] = in[137] & in2[137];
    assign P[104] = in[137] ^ in2[137];
    assign G[105] = in[136] & in2[136];
    assign P[105] = in[136] ^ in2[136];
    assign G[106] = in[135] & in2[135];
    assign P[106] = in[135] ^ in2[135];
    assign G[107] = in[134] & in2[134];
    assign P[107] = in[134] ^ in2[134];
    assign G[108] = in[133] & in2[133];
    assign P[108] = in[133] ^ in2[133];
    assign G[109] = in[132] & in2[132];
    assign P[109] = in[132] ^ in2[132];
    assign G[110] = in[131] & in2[131];
    assign P[110] = in[131] ^ in2[131];
    assign G[111] = in[130] & in2[130];
    assign P[111] = in[130] ^ in2[130];
    assign G[112] = in[129] & in2[129];
    assign P[112] = in[129] ^ in2[129];
    assign G[113] = in[128] & in2[128];
    assign P[113] = in[128] ^ in2[128];
    assign G[114] = in[127] & in2[127];
    assign P[114] = in[127] ^ in2[127];
    assign G[115] = in[126] & in2[126];
    assign P[115] = in[126] ^ in2[126];
    assign G[116] = in[125] & in2[125];
    assign P[116] = in[125] ^ in2[125];
    assign G[117] = in[124] & in2[124];
    assign P[117] = in[124] ^ in2[124];
    assign G[118] = in[123] & in2[123];
    assign P[118] = in[123] ^ in2[123];
    assign G[119] = in[122] & in2[122];
    assign P[119] = in[122] ^ in2[122];
    assign G[120] = in[121] & in2[121];
    assign P[120] = in[121] ^ in2[121];
    assign G[121] = in[120] & in2[120];
    assign P[121] = in[120] ^ in2[120];
    assign G[122] = in[119] & in2[119];
    assign P[122] = in[119] ^ in2[119];
    assign G[123] = in[118] & in2[118];
    assign P[123] = in[118] ^ in2[118];
    assign G[124] = in[117] & in2[117];
    assign P[124] = in[117] ^ in2[117];
    assign G[125] = in[116] & in2[116];
    assign P[125] = in[116] ^ in2[116];
    assign G[126] = in[115] & in2[115];
    assign P[126] = in[115] ^ in2[115];
    assign G[127] = in[114] & in2[114];
    assign P[127] = in[114] ^ in2[114];
    assign G[128] = in[113] & in2[113];
    assign P[128] = in[113] ^ in2[113];
    assign G[129] = in[112] & in2[112];
    assign P[129] = in[112] ^ in2[112];
    assign G[130] = in[111] & in2[111];
    assign P[130] = in[111] ^ in2[111];
    assign G[131] = in[110] & in2[110];
    assign P[131] = in[110] ^ in2[110];
    assign G[132] = in[109] & in2[109];
    assign P[132] = in[109] ^ in2[109];
    assign G[133] = in[108] & in2[108];
    assign P[133] = in[108] ^ in2[108];
    assign G[134] = in[107] & in2[107];
    assign P[134] = in[107] ^ in2[107];
    assign G[135] = in[106] & in2[106];
    assign P[135] = in[106] ^ in2[106];
    assign G[136] = in[105] & in2[105];
    assign P[136] = in[105] ^ in2[105];
    assign G[137] = in[104] & in2[104];
    assign P[137] = in[104] ^ in2[104];
    assign G[138] = in[103] & in2[103];
    assign P[138] = in[103] ^ in2[103];
    assign G[139] = in[102] & in2[102];
    assign P[139] = in[102] ^ in2[102];
    assign G[140] = in[101] & in2[101];
    assign P[140] = in[101] ^ in2[101];
    assign G[141] = in[100] & in2[100];
    assign P[141] = in[100] ^ in2[100];
    assign G[142] = in[99] & in2[99];
    assign P[142] = in[99] ^ in2[99];
    assign G[143] = in[98] & in2[98];
    assign P[143] = in[98] ^ in2[98];
    assign G[144] = in[97] & in2[97];
    assign P[144] = in[97] ^ in2[97];
    assign G[145] = in[96] & in2[96];
    assign P[145] = in[96] ^ in2[96];
    assign G[146] = in[95] & in2[95];
    assign P[146] = in[95] ^ in2[95];
    assign G[147] = in[94] & in2[94];
    assign P[147] = in[94] ^ in2[94];
    assign G[148] = in[93] & in2[93];
    assign P[148] = in[93] ^ in2[93];
    assign G[149] = in[92] & in2[92];
    assign P[149] = in[92] ^ in2[92];
    assign G[150] = in[91] & in2[91];
    assign P[150] = in[91] ^ in2[91];
    assign G[151] = in[90] & in2[90];
    assign P[151] = in[90] ^ in2[90];
    assign G[152] = in[89] & in2[89];
    assign P[152] = in[89] ^ in2[89];
    assign G[153] = in[88] & in2[88];
    assign P[153] = in[88] ^ in2[88];
    assign G[154] = in[87] & in2[87];
    assign P[154] = in[87] ^ in2[87];
    assign G[155] = in[86] & in2[86];
    assign P[155] = in[86] ^ in2[86];
    assign G[156] = in[85] & in2[85];
    assign P[156] = in[85] ^ in2[85];
    assign G[157] = in[84] & in2[84];
    assign P[157] = in[84] ^ in2[84];
    assign G[158] = in[83] & in2[83];
    assign P[158] = in[83] ^ in2[83];
    assign G[159] = in[82] & in2[82];
    assign P[159] = in[82] ^ in2[82];
    assign G[160] = in[81] & in2[81];
    assign P[160] = in[81] ^ in2[81];
    assign G[161] = in[80] & in2[80];
    assign P[161] = in[80] ^ in2[80];
    assign G[162] = in[79] & in2[79];
    assign P[162] = in[79] ^ in2[79];
    assign G[163] = in[78] & in2[78];
    assign P[163] = in[78] ^ in2[78];
    assign G[164] = in[77] & in2[77];
    assign P[164] = in[77] ^ in2[77];
    assign G[165] = in[76] & in2[76];
    assign P[165] = in[76] ^ in2[76];
    assign G[166] = in[75] & in2[75];
    assign P[166] = in[75] ^ in2[75];
    assign G[167] = in[74] & in2[74];
    assign P[167] = in[74] ^ in2[74];
    assign G[168] = in[73] & in2[73];
    assign P[168] = in[73] ^ in2[73];
    assign G[169] = in[72] & in2[72];
    assign P[169] = in[72] ^ in2[72];
    assign G[170] = in[71] & in2[71];
    assign P[170] = in[71] ^ in2[71];
    assign G[171] = in[70] & in2[70];
    assign P[171] = in[70] ^ in2[70];
    assign G[172] = in[69] & in2[69];
    assign P[172] = in[69] ^ in2[69];
    assign G[173] = in[68] & in2[68];
    assign P[173] = in[68] ^ in2[68];
    assign G[174] = in[67] & in2[67];
    assign P[174] = in[67] ^ in2[67];
    assign G[175] = in[66] & in2[66];
    assign P[175] = in[66] ^ in2[66];
    assign G[176] = in[65] & in2[65];
    assign P[176] = in[65] ^ in2[65];
    assign G[177] = in[64] & in2[64];
    assign P[177] = in[64] ^ in2[64];
    assign G[178] = in[63] & in2[63];
    assign P[178] = in[63] ^ in2[63];
    assign G[179] = in[62] & in2[62];
    assign P[179] = in[62] ^ in2[62];
    assign G[180] = in[61] & in2[61];
    assign P[180] = in[61] ^ in2[61];
    assign G[181] = in[60] & in2[60];
    assign P[181] = in[60] ^ in2[60];
    assign G[182] = in[59] & in2[59];
    assign P[182] = in[59] ^ in2[59];
    assign G[183] = in[58] & in2[58];
    assign P[183] = in[58] ^ in2[58];
    assign G[184] = in[57] & in2[57];
    assign P[184] = in[57] ^ in2[57];
    assign G[185] = in[56] & in2[56];
    assign P[185] = in[56] ^ in2[56];
    assign G[186] = in[55] & in2[55];
    assign P[186] = in[55] ^ in2[55];
    assign G[187] = in[54] & in2[54];
    assign P[187] = in[54] ^ in2[54];
    assign G[188] = in[53] & in2[53];
    assign P[188] = in[53] ^ in2[53];
    assign G[189] = in[52] & in2[52];
    assign P[189] = in[52] ^ in2[52];
    assign G[190] = in[51] & in2[51];
    assign P[190] = in[51] ^ in2[51];
    assign G[191] = in[50] & in2[50];
    assign P[191] = in[50] ^ in2[50];
    assign G[192] = in[49] & in2[49];
    assign P[192] = in[49] ^ in2[49];
    assign G[193] = in[48] & in2[48];
    assign P[193] = in[48] ^ in2[48];
    assign G[194] = in[47] & in2[47];
    assign P[194] = in[47] ^ in2[47];
    assign G[195] = in[46] & in2[46];
    assign P[195] = in[46] ^ in2[46];
    assign G[196] = in[45] & in2[45];
    assign P[196] = in[45] ^ in2[45];
    assign G[197] = in[44] & in2[44];
    assign P[197] = in[44] ^ in2[44];
    assign G[198] = in[43] & in2[43];
    assign P[198] = in[43] ^ in2[43];
    assign G[199] = in[42] & in2[42];
    assign P[199] = in[42] ^ in2[42];
    assign G[200] = in[41] & in2[41];
    assign P[200] = in[41] ^ in2[41];
    assign G[201] = in[40] & in2[40];
    assign P[201] = in[40] ^ in2[40];
    assign G[202] = in[39] & in2[39];
    assign P[202] = in[39] ^ in2[39];
    assign G[203] = in[38] & in2[38];
    assign P[203] = in[38] ^ in2[38];
    assign G[204] = in[37] & in2[37];
    assign P[204] = in[37] ^ in2[37];
    assign G[205] = in[36] & in2[36];
    assign P[205] = in[36] ^ in2[36];
    assign G[206] = in[35] & in2[35];
    assign P[206] = in[35] ^ in2[35];
    assign G[207] = in[34] & in2[34];
    assign P[207] = in[34] ^ in2[34];
    assign G[208] = in[33] & in2[33];
    assign P[208] = in[33] ^ in2[33];
    assign G[209] = in[32] & in2[32];
    assign P[209] = in[32] ^ in2[32];
    assign G[210] = in[31] & in2[31];
    assign P[210] = in[31] ^ in2[31];
    assign G[211] = in[30] & in2[30];
    assign P[211] = in[30] ^ in2[30];
    assign G[212] = in[29] & in2[29];
    assign P[212] = in[29] ^ in2[29];
    assign G[213] = in[28] & in2[28];
    assign P[213] = in[28] ^ in2[28];
    assign G[214] = in[27] & in2[27];
    assign P[214] = in[27] ^ in2[27];
    assign G[215] = in[26] & in2[26];
    assign P[215] = in[26] ^ in2[26];
    assign G[216] = in[25] & in2[25];
    assign P[216] = in[25] ^ in2[25];
    assign G[217] = in[24] & in2[24];
    assign P[217] = in[24] ^ in2[24];
    assign G[218] = in[23] & in2[23];
    assign P[218] = in[23] ^ in2[23];
    assign G[219] = in[22] & in2[22];
    assign P[219] = in[22] ^ in2[22];
    assign G[220] = in[21] & in2[21];
    assign P[220] = in[21] ^ in2[21];
    assign G[221] = in[20] & in2[20];
    assign P[221] = in[20] ^ in2[20];
    assign G[222] = in[19] & in2[19];
    assign P[222] = in[19] ^ in2[19];
    assign G[223] = in[18] & in2[18];
    assign P[223] = in[18] ^ in2[18];
    assign G[224] = in[17] & in2[17];
    assign P[224] = in[17] ^ in2[17];
    assign G[225] = in[16] & in2[16];
    assign P[225] = in[16] ^ in2[16];
    assign G[226] = in[15] & in2[15];
    assign P[226] = in[15] ^ in2[15];
    assign G[227] = in[14] & in2[14];
    assign P[227] = in[14] ^ in2[14];
    assign G[228] = in[13] & in2[13];
    assign P[228] = in[13] ^ in2[13];
    assign G[229] = in[12] & in2[12];
    assign P[229] = in[12] ^ in2[12];
    assign G[230] = in[11] & in2[11];
    assign P[230] = in[11] ^ in2[11];
    assign G[231] = in[10] & in2[10];
    assign P[231] = in[10] ^ in2[10];
    assign G[232] = in[9] & in2[9];
    assign P[232] = in[9] ^ in2[9];
    assign G[233] = in[8] & in2[8];
    assign P[233] = in[8] ^ in2[8];
    assign G[234] = in[7] & in2[7];
    assign P[234] = in[7] ^ in2[7];
    assign G[235] = in[6] & in2[6];
    assign P[235] = in[6] ^ in2[6];
    assign G[236] = in[5] & in2[5];
    assign P[236] = in[5] ^ in2[5];
    assign G[237] = in[4] & in2[4];
    assign P[237] = in[4] ^ in2[4];
    assign G[238] = in[3] & in2[3];
    assign P[238] = in[3] ^ in2[3];
    assign G[239] = in[2] & in2[2];
    assign P[239] = in[2] ^ in2[2];
    assign G[240] = in[1] & in2[1];
    assign P[240] = in[1] ^ in2[1];
    assign G[241] = in[0] & in2[0];
    assign P[241] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign C[241] = G[240] | (P[240] & C[240]);
    assign cout = G[241] | (P[241] & C[241]);
    assign sum = P ^ C;
endmodule

module CLA241(output [240:0] sum, output cout, input [240:0] in1, input [240:0] in2;

    wire[240:0] G;
    wire[240:0] C;
    wire[240:0] P;

    assign G[0] = in[240] & in2[240];
    assign P[0] = in[240] ^ in2[240];
    assign G[1] = in[239] & in2[239];
    assign P[1] = in[239] ^ in2[239];
    assign G[2] = in[238] & in2[238];
    assign P[2] = in[238] ^ in2[238];
    assign G[3] = in[237] & in2[237];
    assign P[3] = in[237] ^ in2[237];
    assign G[4] = in[236] & in2[236];
    assign P[4] = in[236] ^ in2[236];
    assign G[5] = in[235] & in2[235];
    assign P[5] = in[235] ^ in2[235];
    assign G[6] = in[234] & in2[234];
    assign P[6] = in[234] ^ in2[234];
    assign G[7] = in[233] & in2[233];
    assign P[7] = in[233] ^ in2[233];
    assign G[8] = in[232] & in2[232];
    assign P[8] = in[232] ^ in2[232];
    assign G[9] = in[231] & in2[231];
    assign P[9] = in[231] ^ in2[231];
    assign G[10] = in[230] & in2[230];
    assign P[10] = in[230] ^ in2[230];
    assign G[11] = in[229] & in2[229];
    assign P[11] = in[229] ^ in2[229];
    assign G[12] = in[228] & in2[228];
    assign P[12] = in[228] ^ in2[228];
    assign G[13] = in[227] & in2[227];
    assign P[13] = in[227] ^ in2[227];
    assign G[14] = in[226] & in2[226];
    assign P[14] = in[226] ^ in2[226];
    assign G[15] = in[225] & in2[225];
    assign P[15] = in[225] ^ in2[225];
    assign G[16] = in[224] & in2[224];
    assign P[16] = in[224] ^ in2[224];
    assign G[17] = in[223] & in2[223];
    assign P[17] = in[223] ^ in2[223];
    assign G[18] = in[222] & in2[222];
    assign P[18] = in[222] ^ in2[222];
    assign G[19] = in[221] & in2[221];
    assign P[19] = in[221] ^ in2[221];
    assign G[20] = in[220] & in2[220];
    assign P[20] = in[220] ^ in2[220];
    assign G[21] = in[219] & in2[219];
    assign P[21] = in[219] ^ in2[219];
    assign G[22] = in[218] & in2[218];
    assign P[22] = in[218] ^ in2[218];
    assign G[23] = in[217] & in2[217];
    assign P[23] = in[217] ^ in2[217];
    assign G[24] = in[216] & in2[216];
    assign P[24] = in[216] ^ in2[216];
    assign G[25] = in[215] & in2[215];
    assign P[25] = in[215] ^ in2[215];
    assign G[26] = in[214] & in2[214];
    assign P[26] = in[214] ^ in2[214];
    assign G[27] = in[213] & in2[213];
    assign P[27] = in[213] ^ in2[213];
    assign G[28] = in[212] & in2[212];
    assign P[28] = in[212] ^ in2[212];
    assign G[29] = in[211] & in2[211];
    assign P[29] = in[211] ^ in2[211];
    assign G[30] = in[210] & in2[210];
    assign P[30] = in[210] ^ in2[210];
    assign G[31] = in[209] & in2[209];
    assign P[31] = in[209] ^ in2[209];
    assign G[32] = in[208] & in2[208];
    assign P[32] = in[208] ^ in2[208];
    assign G[33] = in[207] & in2[207];
    assign P[33] = in[207] ^ in2[207];
    assign G[34] = in[206] & in2[206];
    assign P[34] = in[206] ^ in2[206];
    assign G[35] = in[205] & in2[205];
    assign P[35] = in[205] ^ in2[205];
    assign G[36] = in[204] & in2[204];
    assign P[36] = in[204] ^ in2[204];
    assign G[37] = in[203] & in2[203];
    assign P[37] = in[203] ^ in2[203];
    assign G[38] = in[202] & in2[202];
    assign P[38] = in[202] ^ in2[202];
    assign G[39] = in[201] & in2[201];
    assign P[39] = in[201] ^ in2[201];
    assign G[40] = in[200] & in2[200];
    assign P[40] = in[200] ^ in2[200];
    assign G[41] = in[199] & in2[199];
    assign P[41] = in[199] ^ in2[199];
    assign G[42] = in[198] & in2[198];
    assign P[42] = in[198] ^ in2[198];
    assign G[43] = in[197] & in2[197];
    assign P[43] = in[197] ^ in2[197];
    assign G[44] = in[196] & in2[196];
    assign P[44] = in[196] ^ in2[196];
    assign G[45] = in[195] & in2[195];
    assign P[45] = in[195] ^ in2[195];
    assign G[46] = in[194] & in2[194];
    assign P[46] = in[194] ^ in2[194];
    assign G[47] = in[193] & in2[193];
    assign P[47] = in[193] ^ in2[193];
    assign G[48] = in[192] & in2[192];
    assign P[48] = in[192] ^ in2[192];
    assign G[49] = in[191] & in2[191];
    assign P[49] = in[191] ^ in2[191];
    assign G[50] = in[190] & in2[190];
    assign P[50] = in[190] ^ in2[190];
    assign G[51] = in[189] & in2[189];
    assign P[51] = in[189] ^ in2[189];
    assign G[52] = in[188] & in2[188];
    assign P[52] = in[188] ^ in2[188];
    assign G[53] = in[187] & in2[187];
    assign P[53] = in[187] ^ in2[187];
    assign G[54] = in[186] & in2[186];
    assign P[54] = in[186] ^ in2[186];
    assign G[55] = in[185] & in2[185];
    assign P[55] = in[185] ^ in2[185];
    assign G[56] = in[184] & in2[184];
    assign P[56] = in[184] ^ in2[184];
    assign G[57] = in[183] & in2[183];
    assign P[57] = in[183] ^ in2[183];
    assign G[58] = in[182] & in2[182];
    assign P[58] = in[182] ^ in2[182];
    assign G[59] = in[181] & in2[181];
    assign P[59] = in[181] ^ in2[181];
    assign G[60] = in[180] & in2[180];
    assign P[60] = in[180] ^ in2[180];
    assign G[61] = in[179] & in2[179];
    assign P[61] = in[179] ^ in2[179];
    assign G[62] = in[178] & in2[178];
    assign P[62] = in[178] ^ in2[178];
    assign G[63] = in[177] & in2[177];
    assign P[63] = in[177] ^ in2[177];
    assign G[64] = in[176] & in2[176];
    assign P[64] = in[176] ^ in2[176];
    assign G[65] = in[175] & in2[175];
    assign P[65] = in[175] ^ in2[175];
    assign G[66] = in[174] & in2[174];
    assign P[66] = in[174] ^ in2[174];
    assign G[67] = in[173] & in2[173];
    assign P[67] = in[173] ^ in2[173];
    assign G[68] = in[172] & in2[172];
    assign P[68] = in[172] ^ in2[172];
    assign G[69] = in[171] & in2[171];
    assign P[69] = in[171] ^ in2[171];
    assign G[70] = in[170] & in2[170];
    assign P[70] = in[170] ^ in2[170];
    assign G[71] = in[169] & in2[169];
    assign P[71] = in[169] ^ in2[169];
    assign G[72] = in[168] & in2[168];
    assign P[72] = in[168] ^ in2[168];
    assign G[73] = in[167] & in2[167];
    assign P[73] = in[167] ^ in2[167];
    assign G[74] = in[166] & in2[166];
    assign P[74] = in[166] ^ in2[166];
    assign G[75] = in[165] & in2[165];
    assign P[75] = in[165] ^ in2[165];
    assign G[76] = in[164] & in2[164];
    assign P[76] = in[164] ^ in2[164];
    assign G[77] = in[163] & in2[163];
    assign P[77] = in[163] ^ in2[163];
    assign G[78] = in[162] & in2[162];
    assign P[78] = in[162] ^ in2[162];
    assign G[79] = in[161] & in2[161];
    assign P[79] = in[161] ^ in2[161];
    assign G[80] = in[160] & in2[160];
    assign P[80] = in[160] ^ in2[160];
    assign G[81] = in[159] & in2[159];
    assign P[81] = in[159] ^ in2[159];
    assign G[82] = in[158] & in2[158];
    assign P[82] = in[158] ^ in2[158];
    assign G[83] = in[157] & in2[157];
    assign P[83] = in[157] ^ in2[157];
    assign G[84] = in[156] & in2[156];
    assign P[84] = in[156] ^ in2[156];
    assign G[85] = in[155] & in2[155];
    assign P[85] = in[155] ^ in2[155];
    assign G[86] = in[154] & in2[154];
    assign P[86] = in[154] ^ in2[154];
    assign G[87] = in[153] & in2[153];
    assign P[87] = in[153] ^ in2[153];
    assign G[88] = in[152] & in2[152];
    assign P[88] = in[152] ^ in2[152];
    assign G[89] = in[151] & in2[151];
    assign P[89] = in[151] ^ in2[151];
    assign G[90] = in[150] & in2[150];
    assign P[90] = in[150] ^ in2[150];
    assign G[91] = in[149] & in2[149];
    assign P[91] = in[149] ^ in2[149];
    assign G[92] = in[148] & in2[148];
    assign P[92] = in[148] ^ in2[148];
    assign G[93] = in[147] & in2[147];
    assign P[93] = in[147] ^ in2[147];
    assign G[94] = in[146] & in2[146];
    assign P[94] = in[146] ^ in2[146];
    assign G[95] = in[145] & in2[145];
    assign P[95] = in[145] ^ in2[145];
    assign G[96] = in[144] & in2[144];
    assign P[96] = in[144] ^ in2[144];
    assign G[97] = in[143] & in2[143];
    assign P[97] = in[143] ^ in2[143];
    assign G[98] = in[142] & in2[142];
    assign P[98] = in[142] ^ in2[142];
    assign G[99] = in[141] & in2[141];
    assign P[99] = in[141] ^ in2[141];
    assign G[100] = in[140] & in2[140];
    assign P[100] = in[140] ^ in2[140];
    assign G[101] = in[139] & in2[139];
    assign P[101] = in[139] ^ in2[139];
    assign G[102] = in[138] & in2[138];
    assign P[102] = in[138] ^ in2[138];
    assign G[103] = in[137] & in2[137];
    assign P[103] = in[137] ^ in2[137];
    assign G[104] = in[136] & in2[136];
    assign P[104] = in[136] ^ in2[136];
    assign G[105] = in[135] & in2[135];
    assign P[105] = in[135] ^ in2[135];
    assign G[106] = in[134] & in2[134];
    assign P[106] = in[134] ^ in2[134];
    assign G[107] = in[133] & in2[133];
    assign P[107] = in[133] ^ in2[133];
    assign G[108] = in[132] & in2[132];
    assign P[108] = in[132] ^ in2[132];
    assign G[109] = in[131] & in2[131];
    assign P[109] = in[131] ^ in2[131];
    assign G[110] = in[130] & in2[130];
    assign P[110] = in[130] ^ in2[130];
    assign G[111] = in[129] & in2[129];
    assign P[111] = in[129] ^ in2[129];
    assign G[112] = in[128] & in2[128];
    assign P[112] = in[128] ^ in2[128];
    assign G[113] = in[127] & in2[127];
    assign P[113] = in[127] ^ in2[127];
    assign G[114] = in[126] & in2[126];
    assign P[114] = in[126] ^ in2[126];
    assign G[115] = in[125] & in2[125];
    assign P[115] = in[125] ^ in2[125];
    assign G[116] = in[124] & in2[124];
    assign P[116] = in[124] ^ in2[124];
    assign G[117] = in[123] & in2[123];
    assign P[117] = in[123] ^ in2[123];
    assign G[118] = in[122] & in2[122];
    assign P[118] = in[122] ^ in2[122];
    assign G[119] = in[121] & in2[121];
    assign P[119] = in[121] ^ in2[121];
    assign G[120] = in[120] & in2[120];
    assign P[120] = in[120] ^ in2[120];
    assign G[121] = in[119] & in2[119];
    assign P[121] = in[119] ^ in2[119];
    assign G[122] = in[118] & in2[118];
    assign P[122] = in[118] ^ in2[118];
    assign G[123] = in[117] & in2[117];
    assign P[123] = in[117] ^ in2[117];
    assign G[124] = in[116] & in2[116];
    assign P[124] = in[116] ^ in2[116];
    assign G[125] = in[115] & in2[115];
    assign P[125] = in[115] ^ in2[115];
    assign G[126] = in[114] & in2[114];
    assign P[126] = in[114] ^ in2[114];
    assign G[127] = in[113] & in2[113];
    assign P[127] = in[113] ^ in2[113];
    assign G[128] = in[112] & in2[112];
    assign P[128] = in[112] ^ in2[112];
    assign G[129] = in[111] & in2[111];
    assign P[129] = in[111] ^ in2[111];
    assign G[130] = in[110] & in2[110];
    assign P[130] = in[110] ^ in2[110];
    assign G[131] = in[109] & in2[109];
    assign P[131] = in[109] ^ in2[109];
    assign G[132] = in[108] & in2[108];
    assign P[132] = in[108] ^ in2[108];
    assign G[133] = in[107] & in2[107];
    assign P[133] = in[107] ^ in2[107];
    assign G[134] = in[106] & in2[106];
    assign P[134] = in[106] ^ in2[106];
    assign G[135] = in[105] & in2[105];
    assign P[135] = in[105] ^ in2[105];
    assign G[136] = in[104] & in2[104];
    assign P[136] = in[104] ^ in2[104];
    assign G[137] = in[103] & in2[103];
    assign P[137] = in[103] ^ in2[103];
    assign G[138] = in[102] & in2[102];
    assign P[138] = in[102] ^ in2[102];
    assign G[139] = in[101] & in2[101];
    assign P[139] = in[101] ^ in2[101];
    assign G[140] = in[100] & in2[100];
    assign P[140] = in[100] ^ in2[100];
    assign G[141] = in[99] & in2[99];
    assign P[141] = in[99] ^ in2[99];
    assign G[142] = in[98] & in2[98];
    assign P[142] = in[98] ^ in2[98];
    assign G[143] = in[97] & in2[97];
    assign P[143] = in[97] ^ in2[97];
    assign G[144] = in[96] & in2[96];
    assign P[144] = in[96] ^ in2[96];
    assign G[145] = in[95] & in2[95];
    assign P[145] = in[95] ^ in2[95];
    assign G[146] = in[94] & in2[94];
    assign P[146] = in[94] ^ in2[94];
    assign G[147] = in[93] & in2[93];
    assign P[147] = in[93] ^ in2[93];
    assign G[148] = in[92] & in2[92];
    assign P[148] = in[92] ^ in2[92];
    assign G[149] = in[91] & in2[91];
    assign P[149] = in[91] ^ in2[91];
    assign G[150] = in[90] & in2[90];
    assign P[150] = in[90] ^ in2[90];
    assign G[151] = in[89] & in2[89];
    assign P[151] = in[89] ^ in2[89];
    assign G[152] = in[88] & in2[88];
    assign P[152] = in[88] ^ in2[88];
    assign G[153] = in[87] & in2[87];
    assign P[153] = in[87] ^ in2[87];
    assign G[154] = in[86] & in2[86];
    assign P[154] = in[86] ^ in2[86];
    assign G[155] = in[85] & in2[85];
    assign P[155] = in[85] ^ in2[85];
    assign G[156] = in[84] & in2[84];
    assign P[156] = in[84] ^ in2[84];
    assign G[157] = in[83] & in2[83];
    assign P[157] = in[83] ^ in2[83];
    assign G[158] = in[82] & in2[82];
    assign P[158] = in[82] ^ in2[82];
    assign G[159] = in[81] & in2[81];
    assign P[159] = in[81] ^ in2[81];
    assign G[160] = in[80] & in2[80];
    assign P[160] = in[80] ^ in2[80];
    assign G[161] = in[79] & in2[79];
    assign P[161] = in[79] ^ in2[79];
    assign G[162] = in[78] & in2[78];
    assign P[162] = in[78] ^ in2[78];
    assign G[163] = in[77] & in2[77];
    assign P[163] = in[77] ^ in2[77];
    assign G[164] = in[76] & in2[76];
    assign P[164] = in[76] ^ in2[76];
    assign G[165] = in[75] & in2[75];
    assign P[165] = in[75] ^ in2[75];
    assign G[166] = in[74] & in2[74];
    assign P[166] = in[74] ^ in2[74];
    assign G[167] = in[73] & in2[73];
    assign P[167] = in[73] ^ in2[73];
    assign G[168] = in[72] & in2[72];
    assign P[168] = in[72] ^ in2[72];
    assign G[169] = in[71] & in2[71];
    assign P[169] = in[71] ^ in2[71];
    assign G[170] = in[70] & in2[70];
    assign P[170] = in[70] ^ in2[70];
    assign G[171] = in[69] & in2[69];
    assign P[171] = in[69] ^ in2[69];
    assign G[172] = in[68] & in2[68];
    assign P[172] = in[68] ^ in2[68];
    assign G[173] = in[67] & in2[67];
    assign P[173] = in[67] ^ in2[67];
    assign G[174] = in[66] & in2[66];
    assign P[174] = in[66] ^ in2[66];
    assign G[175] = in[65] & in2[65];
    assign P[175] = in[65] ^ in2[65];
    assign G[176] = in[64] & in2[64];
    assign P[176] = in[64] ^ in2[64];
    assign G[177] = in[63] & in2[63];
    assign P[177] = in[63] ^ in2[63];
    assign G[178] = in[62] & in2[62];
    assign P[178] = in[62] ^ in2[62];
    assign G[179] = in[61] & in2[61];
    assign P[179] = in[61] ^ in2[61];
    assign G[180] = in[60] & in2[60];
    assign P[180] = in[60] ^ in2[60];
    assign G[181] = in[59] & in2[59];
    assign P[181] = in[59] ^ in2[59];
    assign G[182] = in[58] & in2[58];
    assign P[182] = in[58] ^ in2[58];
    assign G[183] = in[57] & in2[57];
    assign P[183] = in[57] ^ in2[57];
    assign G[184] = in[56] & in2[56];
    assign P[184] = in[56] ^ in2[56];
    assign G[185] = in[55] & in2[55];
    assign P[185] = in[55] ^ in2[55];
    assign G[186] = in[54] & in2[54];
    assign P[186] = in[54] ^ in2[54];
    assign G[187] = in[53] & in2[53];
    assign P[187] = in[53] ^ in2[53];
    assign G[188] = in[52] & in2[52];
    assign P[188] = in[52] ^ in2[52];
    assign G[189] = in[51] & in2[51];
    assign P[189] = in[51] ^ in2[51];
    assign G[190] = in[50] & in2[50];
    assign P[190] = in[50] ^ in2[50];
    assign G[191] = in[49] & in2[49];
    assign P[191] = in[49] ^ in2[49];
    assign G[192] = in[48] & in2[48];
    assign P[192] = in[48] ^ in2[48];
    assign G[193] = in[47] & in2[47];
    assign P[193] = in[47] ^ in2[47];
    assign G[194] = in[46] & in2[46];
    assign P[194] = in[46] ^ in2[46];
    assign G[195] = in[45] & in2[45];
    assign P[195] = in[45] ^ in2[45];
    assign G[196] = in[44] & in2[44];
    assign P[196] = in[44] ^ in2[44];
    assign G[197] = in[43] & in2[43];
    assign P[197] = in[43] ^ in2[43];
    assign G[198] = in[42] & in2[42];
    assign P[198] = in[42] ^ in2[42];
    assign G[199] = in[41] & in2[41];
    assign P[199] = in[41] ^ in2[41];
    assign G[200] = in[40] & in2[40];
    assign P[200] = in[40] ^ in2[40];
    assign G[201] = in[39] & in2[39];
    assign P[201] = in[39] ^ in2[39];
    assign G[202] = in[38] & in2[38];
    assign P[202] = in[38] ^ in2[38];
    assign G[203] = in[37] & in2[37];
    assign P[203] = in[37] ^ in2[37];
    assign G[204] = in[36] & in2[36];
    assign P[204] = in[36] ^ in2[36];
    assign G[205] = in[35] & in2[35];
    assign P[205] = in[35] ^ in2[35];
    assign G[206] = in[34] & in2[34];
    assign P[206] = in[34] ^ in2[34];
    assign G[207] = in[33] & in2[33];
    assign P[207] = in[33] ^ in2[33];
    assign G[208] = in[32] & in2[32];
    assign P[208] = in[32] ^ in2[32];
    assign G[209] = in[31] & in2[31];
    assign P[209] = in[31] ^ in2[31];
    assign G[210] = in[30] & in2[30];
    assign P[210] = in[30] ^ in2[30];
    assign G[211] = in[29] & in2[29];
    assign P[211] = in[29] ^ in2[29];
    assign G[212] = in[28] & in2[28];
    assign P[212] = in[28] ^ in2[28];
    assign G[213] = in[27] & in2[27];
    assign P[213] = in[27] ^ in2[27];
    assign G[214] = in[26] & in2[26];
    assign P[214] = in[26] ^ in2[26];
    assign G[215] = in[25] & in2[25];
    assign P[215] = in[25] ^ in2[25];
    assign G[216] = in[24] & in2[24];
    assign P[216] = in[24] ^ in2[24];
    assign G[217] = in[23] & in2[23];
    assign P[217] = in[23] ^ in2[23];
    assign G[218] = in[22] & in2[22];
    assign P[218] = in[22] ^ in2[22];
    assign G[219] = in[21] & in2[21];
    assign P[219] = in[21] ^ in2[21];
    assign G[220] = in[20] & in2[20];
    assign P[220] = in[20] ^ in2[20];
    assign G[221] = in[19] & in2[19];
    assign P[221] = in[19] ^ in2[19];
    assign G[222] = in[18] & in2[18];
    assign P[222] = in[18] ^ in2[18];
    assign G[223] = in[17] & in2[17];
    assign P[223] = in[17] ^ in2[17];
    assign G[224] = in[16] & in2[16];
    assign P[224] = in[16] ^ in2[16];
    assign G[225] = in[15] & in2[15];
    assign P[225] = in[15] ^ in2[15];
    assign G[226] = in[14] & in2[14];
    assign P[226] = in[14] ^ in2[14];
    assign G[227] = in[13] & in2[13];
    assign P[227] = in[13] ^ in2[13];
    assign G[228] = in[12] & in2[12];
    assign P[228] = in[12] ^ in2[12];
    assign G[229] = in[11] & in2[11];
    assign P[229] = in[11] ^ in2[11];
    assign G[230] = in[10] & in2[10];
    assign P[230] = in[10] ^ in2[10];
    assign G[231] = in[9] & in2[9];
    assign P[231] = in[9] ^ in2[9];
    assign G[232] = in[8] & in2[8];
    assign P[232] = in[8] ^ in2[8];
    assign G[233] = in[7] & in2[7];
    assign P[233] = in[7] ^ in2[7];
    assign G[234] = in[6] & in2[6];
    assign P[234] = in[6] ^ in2[6];
    assign G[235] = in[5] & in2[5];
    assign P[235] = in[5] ^ in2[5];
    assign G[236] = in[4] & in2[4];
    assign P[236] = in[4] ^ in2[4];
    assign G[237] = in[3] & in2[3];
    assign P[237] = in[3] ^ in2[3];
    assign G[238] = in[2] & in2[2];
    assign P[238] = in[2] ^ in2[2];
    assign G[239] = in[1] & in2[1];
    assign P[239] = in[1] ^ in2[1];
    assign G[240] = in[0] & in2[0];
    assign P[240] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign C[240] = G[239] | (P[239] & C[239]);
    assign cout = G[240] | (P[240] & C[240]);
    assign sum = P ^ C;
endmodule

module CLA240(output [239:0] sum, output cout, input [239:0] in1, input [239:0] in2;

    wire[239:0] G;
    wire[239:0] C;
    wire[239:0] P;

    assign G[0] = in[239] & in2[239];
    assign P[0] = in[239] ^ in2[239];
    assign G[1] = in[238] & in2[238];
    assign P[1] = in[238] ^ in2[238];
    assign G[2] = in[237] & in2[237];
    assign P[2] = in[237] ^ in2[237];
    assign G[3] = in[236] & in2[236];
    assign P[3] = in[236] ^ in2[236];
    assign G[4] = in[235] & in2[235];
    assign P[4] = in[235] ^ in2[235];
    assign G[5] = in[234] & in2[234];
    assign P[5] = in[234] ^ in2[234];
    assign G[6] = in[233] & in2[233];
    assign P[6] = in[233] ^ in2[233];
    assign G[7] = in[232] & in2[232];
    assign P[7] = in[232] ^ in2[232];
    assign G[8] = in[231] & in2[231];
    assign P[8] = in[231] ^ in2[231];
    assign G[9] = in[230] & in2[230];
    assign P[9] = in[230] ^ in2[230];
    assign G[10] = in[229] & in2[229];
    assign P[10] = in[229] ^ in2[229];
    assign G[11] = in[228] & in2[228];
    assign P[11] = in[228] ^ in2[228];
    assign G[12] = in[227] & in2[227];
    assign P[12] = in[227] ^ in2[227];
    assign G[13] = in[226] & in2[226];
    assign P[13] = in[226] ^ in2[226];
    assign G[14] = in[225] & in2[225];
    assign P[14] = in[225] ^ in2[225];
    assign G[15] = in[224] & in2[224];
    assign P[15] = in[224] ^ in2[224];
    assign G[16] = in[223] & in2[223];
    assign P[16] = in[223] ^ in2[223];
    assign G[17] = in[222] & in2[222];
    assign P[17] = in[222] ^ in2[222];
    assign G[18] = in[221] & in2[221];
    assign P[18] = in[221] ^ in2[221];
    assign G[19] = in[220] & in2[220];
    assign P[19] = in[220] ^ in2[220];
    assign G[20] = in[219] & in2[219];
    assign P[20] = in[219] ^ in2[219];
    assign G[21] = in[218] & in2[218];
    assign P[21] = in[218] ^ in2[218];
    assign G[22] = in[217] & in2[217];
    assign P[22] = in[217] ^ in2[217];
    assign G[23] = in[216] & in2[216];
    assign P[23] = in[216] ^ in2[216];
    assign G[24] = in[215] & in2[215];
    assign P[24] = in[215] ^ in2[215];
    assign G[25] = in[214] & in2[214];
    assign P[25] = in[214] ^ in2[214];
    assign G[26] = in[213] & in2[213];
    assign P[26] = in[213] ^ in2[213];
    assign G[27] = in[212] & in2[212];
    assign P[27] = in[212] ^ in2[212];
    assign G[28] = in[211] & in2[211];
    assign P[28] = in[211] ^ in2[211];
    assign G[29] = in[210] & in2[210];
    assign P[29] = in[210] ^ in2[210];
    assign G[30] = in[209] & in2[209];
    assign P[30] = in[209] ^ in2[209];
    assign G[31] = in[208] & in2[208];
    assign P[31] = in[208] ^ in2[208];
    assign G[32] = in[207] & in2[207];
    assign P[32] = in[207] ^ in2[207];
    assign G[33] = in[206] & in2[206];
    assign P[33] = in[206] ^ in2[206];
    assign G[34] = in[205] & in2[205];
    assign P[34] = in[205] ^ in2[205];
    assign G[35] = in[204] & in2[204];
    assign P[35] = in[204] ^ in2[204];
    assign G[36] = in[203] & in2[203];
    assign P[36] = in[203] ^ in2[203];
    assign G[37] = in[202] & in2[202];
    assign P[37] = in[202] ^ in2[202];
    assign G[38] = in[201] & in2[201];
    assign P[38] = in[201] ^ in2[201];
    assign G[39] = in[200] & in2[200];
    assign P[39] = in[200] ^ in2[200];
    assign G[40] = in[199] & in2[199];
    assign P[40] = in[199] ^ in2[199];
    assign G[41] = in[198] & in2[198];
    assign P[41] = in[198] ^ in2[198];
    assign G[42] = in[197] & in2[197];
    assign P[42] = in[197] ^ in2[197];
    assign G[43] = in[196] & in2[196];
    assign P[43] = in[196] ^ in2[196];
    assign G[44] = in[195] & in2[195];
    assign P[44] = in[195] ^ in2[195];
    assign G[45] = in[194] & in2[194];
    assign P[45] = in[194] ^ in2[194];
    assign G[46] = in[193] & in2[193];
    assign P[46] = in[193] ^ in2[193];
    assign G[47] = in[192] & in2[192];
    assign P[47] = in[192] ^ in2[192];
    assign G[48] = in[191] & in2[191];
    assign P[48] = in[191] ^ in2[191];
    assign G[49] = in[190] & in2[190];
    assign P[49] = in[190] ^ in2[190];
    assign G[50] = in[189] & in2[189];
    assign P[50] = in[189] ^ in2[189];
    assign G[51] = in[188] & in2[188];
    assign P[51] = in[188] ^ in2[188];
    assign G[52] = in[187] & in2[187];
    assign P[52] = in[187] ^ in2[187];
    assign G[53] = in[186] & in2[186];
    assign P[53] = in[186] ^ in2[186];
    assign G[54] = in[185] & in2[185];
    assign P[54] = in[185] ^ in2[185];
    assign G[55] = in[184] & in2[184];
    assign P[55] = in[184] ^ in2[184];
    assign G[56] = in[183] & in2[183];
    assign P[56] = in[183] ^ in2[183];
    assign G[57] = in[182] & in2[182];
    assign P[57] = in[182] ^ in2[182];
    assign G[58] = in[181] & in2[181];
    assign P[58] = in[181] ^ in2[181];
    assign G[59] = in[180] & in2[180];
    assign P[59] = in[180] ^ in2[180];
    assign G[60] = in[179] & in2[179];
    assign P[60] = in[179] ^ in2[179];
    assign G[61] = in[178] & in2[178];
    assign P[61] = in[178] ^ in2[178];
    assign G[62] = in[177] & in2[177];
    assign P[62] = in[177] ^ in2[177];
    assign G[63] = in[176] & in2[176];
    assign P[63] = in[176] ^ in2[176];
    assign G[64] = in[175] & in2[175];
    assign P[64] = in[175] ^ in2[175];
    assign G[65] = in[174] & in2[174];
    assign P[65] = in[174] ^ in2[174];
    assign G[66] = in[173] & in2[173];
    assign P[66] = in[173] ^ in2[173];
    assign G[67] = in[172] & in2[172];
    assign P[67] = in[172] ^ in2[172];
    assign G[68] = in[171] & in2[171];
    assign P[68] = in[171] ^ in2[171];
    assign G[69] = in[170] & in2[170];
    assign P[69] = in[170] ^ in2[170];
    assign G[70] = in[169] & in2[169];
    assign P[70] = in[169] ^ in2[169];
    assign G[71] = in[168] & in2[168];
    assign P[71] = in[168] ^ in2[168];
    assign G[72] = in[167] & in2[167];
    assign P[72] = in[167] ^ in2[167];
    assign G[73] = in[166] & in2[166];
    assign P[73] = in[166] ^ in2[166];
    assign G[74] = in[165] & in2[165];
    assign P[74] = in[165] ^ in2[165];
    assign G[75] = in[164] & in2[164];
    assign P[75] = in[164] ^ in2[164];
    assign G[76] = in[163] & in2[163];
    assign P[76] = in[163] ^ in2[163];
    assign G[77] = in[162] & in2[162];
    assign P[77] = in[162] ^ in2[162];
    assign G[78] = in[161] & in2[161];
    assign P[78] = in[161] ^ in2[161];
    assign G[79] = in[160] & in2[160];
    assign P[79] = in[160] ^ in2[160];
    assign G[80] = in[159] & in2[159];
    assign P[80] = in[159] ^ in2[159];
    assign G[81] = in[158] & in2[158];
    assign P[81] = in[158] ^ in2[158];
    assign G[82] = in[157] & in2[157];
    assign P[82] = in[157] ^ in2[157];
    assign G[83] = in[156] & in2[156];
    assign P[83] = in[156] ^ in2[156];
    assign G[84] = in[155] & in2[155];
    assign P[84] = in[155] ^ in2[155];
    assign G[85] = in[154] & in2[154];
    assign P[85] = in[154] ^ in2[154];
    assign G[86] = in[153] & in2[153];
    assign P[86] = in[153] ^ in2[153];
    assign G[87] = in[152] & in2[152];
    assign P[87] = in[152] ^ in2[152];
    assign G[88] = in[151] & in2[151];
    assign P[88] = in[151] ^ in2[151];
    assign G[89] = in[150] & in2[150];
    assign P[89] = in[150] ^ in2[150];
    assign G[90] = in[149] & in2[149];
    assign P[90] = in[149] ^ in2[149];
    assign G[91] = in[148] & in2[148];
    assign P[91] = in[148] ^ in2[148];
    assign G[92] = in[147] & in2[147];
    assign P[92] = in[147] ^ in2[147];
    assign G[93] = in[146] & in2[146];
    assign P[93] = in[146] ^ in2[146];
    assign G[94] = in[145] & in2[145];
    assign P[94] = in[145] ^ in2[145];
    assign G[95] = in[144] & in2[144];
    assign P[95] = in[144] ^ in2[144];
    assign G[96] = in[143] & in2[143];
    assign P[96] = in[143] ^ in2[143];
    assign G[97] = in[142] & in2[142];
    assign P[97] = in[142] ^ in2[142];
    assign G[98] = in[141] & in2[141];
    assign P[98] = in[141] ^ in2[141];
    assign G[99] = in[140] & in2[140];
    assign P[99] = in[140] ^ in2[140];
    assign G[100] = in[139] & in2[139];
    assign P[100] = in[139] ^ in2[139];
    assign G[101] = in[138] & in2[138];
    assign P[101] = in[138] ^ in2[138];
    assign G[102] = in[137] & in2[137];
    assign P[102] = in[137] ^ in2[137];
    assign G[103] = in[136] & in2[136];
    assign P[103] = in[136] ^ in2[136];
    assign G[104] = in[135] & in2[135];
    assign P[104] = in[135] ^ in2[135];
    assign G[105] = in[134] & in2[134];
    assign P[105] = in[134] ^ in2[134];
    assign G[106] = in[133] & in2[133];
    assign P[106] = in[133] ^ in2[133];
    assign G[107] = in[132] & in2[132];
    assign P[107] = in[132] ^ in2[132];
    assign G[108] = in[131] & in2[131];
    assign P[108] = in[131] ^ in2[131];
    assign G[109] = in[130] & in2[130];
    assign P[109] = in[130] ^ in2[130];
    assign G[110] = in[129] & in2[129];
    assign P[110] = in[129] ^ in2[129];
    assign G[111] = in[128] & in2[128];
    assign P[111] = in[128] ^ in2[128];
    assign G[112] = in[127] & in2[127];
    assign P[112] = in[127] ^ in2[127];
    assign G[113] = in[126] & in2[126];
    assign P[113] = in[126] ^ in2[126];
    assign G[114] = in[125] & in2[125];
    assign P[114] = in[125] ^ in2[125];
    assign G[115] = in[124] & in2[124];
    assign P[115] = in[124] ^ in2[124];
    assign G[116] = in[123] & in2[123];
    assign P[116] = in[123] ^ in2[123];
    assign G[117] = in[122] & in2[122];
    assign P[117] = in[122] ^ in2[122];
    assign G[118] = in[121] & in2[121];
    assign P[118] = in[121] ^ in2[121];
    assign G[119] = in[120] & in2[120];
    assign P[119] = in[120] ^ in2[120];
    assign G[120] = in[119] & in2[119];
    assign P[120] = in[119] ^ in2[119];
    assign G[121] = in[118] & in2[118];
    assign P[121] = in[118] ^ in2[118];
    assign G[122] = in[117] & in2[117];
    assign P[122] = in[117] ^ in2[117];
    assign G[123] = in[116] & in2[116];
    assign P[123] = in[116] ^ in2[116];
    assign G[124] = in[115] & in2[115];
    assign P[124] = in[115] ^ in2[115];
    assign G[125] = in[114] & in2[114];
    assign P[125] = in[114] ^ in2[114];
    assign G[126] = in[113] & in2[113];
    assign P[126] = in[113] ^ in2[113];
    assign G[127] = in[112] & in2[112];
    assign P[127] = in[112] ^ in2[112];
    assign G[128] = in[111] & in2[111];
    assign P[128] = in[111] ^ in2[111];
    assign G[129] = in[110] & in2[110];
    assign P[129] = in[110] ^ in2[110];
    assign G[130] = in[109] & in2[109];
    assign P[130] = in[109] ^ in2[109];
    assign G[131] = in[108] & in2[108];
    assign P[131] = in[108] ^ in2[108];
    assign G[132] = in[107] & in2[107];
    assign P[132] = in[107] ^ in2[107];
    assign G[133] = in[106] & in2[106];
    assign P[133] = in[106] ^ in2[106];
    assign G[134] = in[105] & in2[105];
    assign P[134] = in[105] ^ in2[105];
    assign G[135] = in[104] & in2[104];
    assign P[135] = in[104] ^ in2[104];
    assign G[136] = in[103] & in2[103];
    assign P[136] = in[103] ^ in2[103];
    assign G[137] = in[102] & in2[102];
    assign P[137] = in[102] ^ in2[102];
    assign G[138] = in[101] & in2[101];
    assign P[138] = in[101] ^ in2[101];
    assign G[139] = in[100] & in2[100];
    assign P[139] = in[100] ^ in2[100];
    assign G[140] = in[99] & in2[99];
    assign P[140] = in[99] ^ in2[99];
    assign G[141] = in[98] & in2[98];
    assign P[141] = in[98] ^ in2[98];
    assign G[142] = in[97] & in2[97];
    assign P[142] = in[97] ^ in2[97];
    assign G[143] = in[96] & in2[96];
    assign P[143] = in[96] ^ in2[96];
    assign G[144] = in[95] & in2[95];
    assign P[144] = in[95] ^ in2[95];
    assign G[145] = in[94] & in2[94];
    assign P[145] = in[94] ^ in2[94];
    assign G[146] = in[93] & in2[93];
    assign P[146] = in[93] ^ in2[93];
    assign G[147] = in[92] & in2[92];
    assign P[147] = in[92] ^ in2[92];
    assign G[148] = in[91] & in2[91];
    assign P[148] = in[91] ^ in2[91];
    assign G[149] = in[90] & in2[90];
    assign P[149] = in[90] ^ in2[90];
    assign G[150] = in[89] & in2[89];
    assign P[150] = in[89] ^ in2[89];
    assign G[151] = in[88] & in2[88];
    assign P[151] = in[88] ^ in2[88];
    assign G[152] = in[87] & in2[87];
    assign P[152] = in[87] ^ in2[87];
    assign G[153] = in[86] & in2[86];
    assign P[153] = in[86] ^ in2[86];
    assign G[154] = in[85] & in2[85];
    assign P[154] = in[85] ^ in2[85];
    assign G[155] = in[84] & in2[84];
    assign P[155] = in[84] ^ in2[84];
    assign G[156] = in[83] & in2[83];
    assign P[156] = in[83] ^ in2[83];
    assign G[157] = in[82] & in2[82];
    assign P[157] = in[82] ^ in2[82];
    assign G[158] = in[81] & in2[81];
    assign P[158] = in[81] ^ in2[81];
    assign G[159] = in[80] & in2[80];
    assign P[159] = in[80] ^ in2[80];
    assign G[160] = in[79] & in2[79];
    assign P[160] = in[79] ^ in2[79];
    assign G[161] = in[78] & in2[78];
    assign P[161] = in[78] ^ in2[78];
    assign G[162] = in[77] & in2[77];
    assign P[162] = in[77] ^ in2[77];
    assign G[163] = in[76] & in2[76];
    assign P[163] = in[76] ^ in2[76];
    assign G[164] = in[75] & in2[75];
    assign P[164] = in[75] ^ in2[75];
    assign G[165] = in[74] & in2[74];
    assign P[165] = in[74] ^ in2[74];
    assign G[166] = in[73] & in2[73];
    assign P[166] = in[73] ^ in2[73];
    assign G[167] = in[72] & in2[72];
    assign P[167] = in[72] ^ in2[72];
    assign G[168] = in[71] & in2[71];
    assign P[168] = in[71] ^ in2[71];
    assign G[169] = in[70] & in2[70];
    assign P[169] = in[70] ^ in2[70];
    assign G[170] = in[69] & in2[69];
    assign P[170] = in[69] ^ in2[69];
    assign G[171] = in[68] & in2[68];
    assign P[171] = in[68] ^ in2[68];
    assign G[172] = in[67] & in2[67];
    assign P[172] = in[67] ^ in2[67];
    assign G[173] = in[66] & in2[66];
    assign P[173] = in[66] ^ in2[66];
    assign G[174] = in[65] & in2[65];
    assign P[174] = in[65] ^ in2[65];
    assign G[175] = in[64] & in2[64];
    assign P[175] = in[64] ^ in2[64];
    assign G[176] = in[63] & in2[63];
    assign P[176] = in[63] ^ in2[63];
    assign G[177] = in[62] & in2[62];
    assign P[177] = in[62] ^ in2[62];
    assign G[178] = in[61] & in2[61];
    assign P[178] = in[61] ^ in2[61];
    assign G[179] = in[60] & in2[60];
    assign P[179] = in[60] ^ in2[60];
    assign G[180] = in[59] & in2[59];
    assign P[180] = in[59] ^ in2[59];
    assign G[181] = in[58] & in2[58];
    assign P[181] = in[58] ^ in2[58];
    assign G[182] = in[57] & in2[57];
    assign P[182] = in[57] ^ in2[57];
    assign G[183] = in[56] & in2[56];
    assign P[183] = in[56] ^ in2[56];
    assign G[184] = in[55] & in2[55];
    assign P[184] = in[55] ^ in2[55];
    assign G[185] = in[54] & in2[54];
    assign P[185] = in[54] ^ in2[54];
    assign G[186] = in[53] & in2[53];
    assign P[186] = in[53] ^ in2[53];
    assign G[187] = in[52] & in2[52];
    assign P[187] = in[52] ^ in2[52];
    assign G[188] = in[51] & in2[51];
    assign P[188] = in[51] ^ in2[51];
    assign G[189] = in[50] & in2[50];
    assign P[189] = in[50] ^ in2[50];
    assign G[190] = in[49] & in2[49];
    assign P[190] = in[49] ^ in2[49];
    assign G[191] = in[48] & in2[48];
    assign P[191] = in[48] ^ in2[48];
    assign G[192] = in[47] & in2[47];
    assign P[192] = in[47] ^ in2[47];
    assign G[193] = in[46] & in2[46];
    assign P[193] = in[46] ^ in2[46];
    assign G[194] = in[45] & in2[45];
    assign P[194] = in[45] ^ in2[45];
    assign G[195] = in[44] & in2[44];
    assign P[195] = in[44] ^ in2[44];
    assign G[196] = in[43] & in2[43];
    assign P[196] = in[43] ^ in2[43];
    assign G[197] = in[42] & in2[42];
    assign P[197] = in[42] ^ in2[42];
    assign G[198] = in[41] & in2[41];
    assign P[198] = in[41] ^ in2[41];
    assign G[199] = in[40] & in2[40];
    assign P[199] = in[40] ^ in2[40];
    assign G[200] = in[39] & in2[39];
    assign P[200] = in[39] ^ in2[39];
    assign G[201] = in[38] & in2[38];
    assign P[201] = in[38] ^ in2[38];
    assign G[202] = in[37] & in2[37];
    assign P[202] = in[37] ^ in2[37];
    assign G[203] = in[36] & in2[36];
    assign P[203] = in[36] ^ in2[36];
    assign G[204] = in[35] & in2[35];
    assign P[204] = in[35] ^ in2[35];
    assign G[205] = in[34] & in2[34];
    assign P[205] = in[34] ^ in2[34];
    assign G[206] = in[33] & in2[33];
    assign P[206] = in[33] ^ in2[33];
    assign G[207] = in[32] & in2[32];
    assign P[207] = in[32] ^ in2[32];
    assign G[208] = in[31] & in2[31];
    assign P[208] = in[31] ^ in2[31];
    assign G[209] = in[30] & in2[30];
    assign P[209] = in[30] ^ in2[30];
    assign G[210] = in[29] & in2[29];
    assign P[210] = in[29] ^ in2[29];
    assign G[211] = in[28] & in2[28];
    assign P[211] = in[28] ^ in2[28];
    assign G[212] = in[27] & in2[27];
    assign P[212] = in[27] ^ in2[27];
    assign G[213] = in[26] & in2[26];
    assign P[213] = in[26] ^ in2[26];
    assign G[214] = in[25] & in2[25];
    assign P[214] = in[25] ^ in2[25];
    assign G[215] = in[24] & in2[24];
    assign P[215] = in[24] ^ in2[24];
    assign G[216] = in[23] & in2[23];
    assign P[216] = in[23] ^ in2[23];
    assign G[217] = in[22] & in2[22];
    assign P[217] = in[22] ^ in2[22];
    assign G[218] = in[21] & in2[21];
    assign P[218] = in[21] ^ in2[21];
    assign G[219] = in[20] & in2[20];
    assign P[219] = in[20] ^ in2[20];
    assign G[220] = in[19] & in2[19];
    assign P[220] = in[19] ^ in2[19];
    assign G[221] = in[18] & in2[18];
    assign P[221] = in[18] ^ in2[18];
    assign G[222] = in[17] & in2[17];
    assign P[222] = in[17] ^ in2[17];
    assign G[223] = in[16] & in2[16];
    assign P[223] = in[16] ^ in2[16];
    assign G[224] = in[15] & in2[15];
    assign P[224] = in[15] ^ in2[15];
    assign G[225] = in[14] & in2[14];
    assign P[225] = in[14] ^ in2[14];
    assign G[226] = in[13] & in2[13];
    assign P[226] = in[13] ^ in2[13];
    assign G[227] = in[12] & in2[12];
    assign P[227] = in[12] ^ in2[12];
    assign G[228] = in[11] & in2[11];
    assign P[228] = in[11] ^ in2[11];
    assign G[229] = in[10] & in2[10];
    assign P[229] = in[10] ^ in2[10];
    assign G[230] = in[9] & in2[9];
    assign P[230] = in[9] ^ in2[9];
    assign G[231] = in[8] & in2[8];
    assign P[231] = in[8] ^ in2[8];
    assign G[232] = in[7] & in2[7];
    assign P[232] = in[7] ^ in2[7];
    assign G[233] = in[6] & in2[6];
    assign P[233] = in[6] ^ in2[6];
    assign G[234] = in[5] & in2[5];
    assign P[234] = in[5] ^ in2[5];
    assign G[235] = in[4] & in2[4];
    assign P[235] = in[4] ^ in2[4];
    assign G[236] = in[3] & in2[3];
    assign P[236] = in[3] ^ in2[3];
    assign G[237] = in[2] & in2[2];
    assign P[237] = in[2] ^ in2[2];
    assign G[238] = in[1] & in2[1];
    assign P[238] = in[1] ^ in2[1];
    assign G[239] = in[0] & in2[0];
    assign P[239] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign C[239] = G[238] | (P[238] & C[238]);
    assign cout = G[239] | (P[239] & C[239]);
    assign sum = P ^ C;
endmodule

module CLA239(output [238:0] sum, output cout, input [238:0] in1, input [238:0] in2;

    wire[238:0] G;
    wire[238:0] C;
    wire[238:0] P;

    assign G[0] = in[238] & in2[238];
    assign P[0] = in[238] ^ in2[238];
    assign G[1] = in[237] & in2[237];
    assign P[1] = in[237] ^ in2[237];
    assign G[2] = in[236] & in2[236];
    assign P[2] = in[236] ^ in2[236];
    assign G[3] = in[235] & in2[235];
    assign P[3] = in[235] ^ in2[235];
    assign G[4] = in[234] & in2[234];
    assign P[4] = in[234] ^ in2[234];
    assign G[5] = in[233] & in2[233];
    assign P[5] = in[233] ^ in2[233];
    assign G[6] = in[232] & in2[232];
    assign P[6] = in[232] ^ in2[232];
    assign G[7] = in[231] & in2[231];
    assign P[7] = in[231] ^ in2[231];
    assign G[8] = in[230] & in2[230];
    assign P[8] = in[230] ^ in2[230];
    assign G[9] = in[229] & in2[229];
    assign P[9] = in[229] ^ in2[229];
    assign G[10] = in[228] & in2[228];
    assign P[10] = in[228] ^ in2[228];
    assign G[11] = in[227] & in2[227];
    assign P[11] = in[227] ^ in2[227];
    assign G[12] = in[226] & in2[226];
    assign P[12] = in[226] ^ in2[226];
    assign G[13] = in[225] & in2[225];
    assign P[13] = in[225] ^ in2[225];
    assign G[14] = in[224] & in2[224];
    assign P[14] = in[224] ^ in2[224];
    assign G[15] = in[223] & in2[223];
    assign P[15] = in[223] ^ in2[223];
    assign G[16] = in[222] & in2[222];
    assign P[16] = in[222] ^ in2[222];
    assign G[17] = in[221] & in2[221];
    assign P[17] = in[221] ^ in2[221];
    assign G[18] = in[220] & in2[220];
    assign P[18] = in[220] ^ in2[220];
    assign G[19] = in[219] & in2[219];
    assign P[19] = in[219] ^ in2[219];
    assign G[20] = in[218] & in2[218];
    assign P[20] = in[218] ^ in2[218];
    assign G[21] = in[217] & in2[217];
    assign P[21] = in[217] ^ in2[217];
    assign G[22] = in[216] & in2[216];
    assign P[22] = in[216] ^ in2[216];
    assign G[23] = in[215] & in2[215];
    assign P[23] = in[215] ^ in2[215];
    assign G[24] = in[214] & in2[214];
    assign P[24] = in[214] ^ in2[214];
    assign G[25] = in[213] & in2[213];
    assign P[25] = in[213] ^ in2[213];
    assign G[26] = in[212] & in2[212];
    assign P[26] = in[212] ^ in2[212];
    assign G[27] = in[211] & in2[211];
    assign P[27] = in[211] ^ in2[211];
    assign G[28] = in[210] & in2[210];
    assign P[28] = in[210] ^ in2[210];
    assign G[29] = in[209] & in2[209];
    assign P[29] = in[209] ^ in2[209];
    assign G[30] = in[208] & in2[208];
    assign P[30] = in[208] ^ in2[208];
    assign G[31] = in[207] & in2[207];
    assign P[31] = in[207] ^ in2[207];
    assign G[32] = in[206] & in2[206];
    assign P[32] = in[206] ^ in2[206];
    assign G[33] = in[205] & in2[205];
    assign P[33] = in[205] ^ in2[205];
    assign G[34] = in[204] & in2[204];
    assign P[34] = in[204] ^ in2[204];
    assign G[35] = in[203] & in2[203];
    assign P[35] = in[203] ^ in2[203];
    assign G[36] = in[202] & in2[202];
    assign P[36] = in[202] ^ in2[202];
    assign G[37] = in[201] & in2[201];
    assign P[37] = in[201] ^ in2[201];
    assign G[38] = in[200] & in2[200];
    assign P[38] = in[200] ^ in2[200];
    assign G[39] = in[199] & in2[199];
    assign P[39] = in[199] ^ in2[199];
    assign G[40] = in[198] & in2[198];
    assign P[40] = in[198] ^ in2[198];
    assign G[41] = in[197] & in2[197];
    assign P[41] = in[197] ^ in2[197];
    assign G[42] = in[196] & in2[196];
    assign P[42] = in[196] ^ in2[196];
    assign G[43] = in[195] & in2[195];
    assign P[43] = in[195] ^ in2[195];
    assign G[44] = in[194] & in2[194];
    assign P[44] = in[194] ^ in2[194];
    assign G[45] = in[193] & in2[193];
    assign P[45] = in[193] ^ in2[193];
    assign G[46] = in[192] & in2[192];
    assign P[46] = in[192] ^ in2[192];
    assign G[47] = in[191] & in2[191];
    assign P[47] = in[191] ^ in2[191];
    assign G[48] = in[190] & in2[190];
    assign P[48] = in[190] ^ in2[190];
    assign G[49] = in[189] & in2[189];
    assign P[49] = in[189] ^ in2[189];
    assign G[50] = in[188] & in2[188];
    assign P[50] = in[188] ^ in2[188];
    assign G[51] = in[187] & in2[187];
    assign P[51] = in[187] ^ in2[187];
    assign G[52] = in[186] & in2[186];
    assign P[52] = in[186] ^ in2[186];
    assign G[53] = in[185] & in2[185];
    assign P[53] = in[185] ^ in2[185];
    assign G[54] = in[184] & in2[184];
    assign P[54] = in[184] ^ in2[184];
    assign G[55] = in[183] & in2[183];
    assign P[55] = in[183] ^ in2[183];
    assign G[56] = in[182] & in2[182];
    assign P[56] = in[182] ^ in2[182];
    assign G[57] = in[181] & in2[181];
    assign P[57] = in[181] ^ in2[181];
    assign G[58] = in[180] & in2[180];
    assign P[58] = in[180] ^ in2[180];
    assign G[59] = in[179] & in2[179];
    assign P[59] = in[179] ^ in2[179];
    assign G[60] = in[178] & in2[178];
    assign P[60] = in[178] ^ in2[178];
    assign G[61] = in[177] & in2[177];
    assign P[61] = in[177] ^ in2[177];
    assign G[62] = in[176] & in2[176];
    assign P[62] = in[176] ^ in2[176];
    assign G[63] = in[175] & in2[175];
    assign P[63] = in[175] ^ in2[175];
    assign G[64] = in[174] & in2[174];
    assign P[64] = in[174] ^ in2[174];
    assign G[65] = in[173] & in2[173];
    assign P[65] = in[173] ^ in2[173];
    assign G[66] = in[172] & in2[172];
    assign P[66] = in[172] ^ in2[172];
    assign G[67] = in[171] & in2[171];
    assign P[67] = in[171] ^ in2[171];
    assign G[68] = in[170] & in2[170];
    assign P[68] = in[170] ^ in2[170];
    assign G[69] = in[169] & in2[169];
    assign P[69] = in[169] ^ in2[169];
    assign G[70] = in[168] & in2[168];
    assign P[70] = in[168] ^ in2[168];
    assign G[71] = in[167] & in2[167];
    assign P[71] = in[167] ^ in2[167];
    assign G[72] = in[166] & in2[166];
    assign P[72] = in[166] ^ in2[166];
    assign G[73] = in[165] & in2[165];
    assign P[73] = in[165] ^ in2[165];
    assign G[74] = in[164] & in2[164];
    assign P[74] = in[164] ^ in2[164];
    assign G[75] = in[163] & in2[163];
    assign P[75] = in[163] ^ in2[163];
    assign G[76] = in[162] & in2[162];
    assign P[76] = in[162] ^ in2[162];
    assign G[77] = in[161] & in2[161];
    assign P[77] = in[161] ^ in2[161];
    assign G[78] = in[160] & in2[160];
    assign P[78] = in[160] ^ in2[160];
    assign G[79] = in[159] & in2[159];
    assign P[79] = in[159] ^ in2[159];
    assign G[80] = in[158] & in2[158];
    assign P[80] = in[158] ^ in2[158];
    assign G[81] = in[157] & in2[157];
    assign P[81] = in[157] ^ in2[157];
    assign G[82] = in[156] & in2[156];
    assign P[82] = in[156] ^ in2[156];
    assign G[83] = in[155] & in2[155];
    assign P[83] = in[155] ^ in2[155];
    assign G[84] = in[154] & in2[154];
    assign P[84] = in[154] ^ in2[154];
    assign G[85] = in[153] & in2[153];
    assign P[85] = in[153] ^ in2[153];
    assign G[86] = in[152] & in2[152];
    assign P[86] = in[152] ^ in2[152];
    assign G[87] = in[151] & in2[151];
    assign P[87] = in[151] ^ in2[151];
    assign G[88] = in[150] & in2[150];
    assign P[88] = in[150] ^ in2[150];
    assign G[89] = in[149] & in2[149];
    assign P[89] = in[149] ^ in2[149];
    assign G[90] = in[148] & in2[148];
    assign P[90] = in[148] ^ in2[148];
    assign G[91] = in[147] & in2[147];
    assign P[91] = in[147] ^ in2[147];
    assign G[92] = in[146] & in2[146];
    assign P[92] = in[146] ^ in2[146];
    assign G[93] = in[145] & in2[145];
    assign P[93] = in[145] ^ in2[145];
    assign G[94] = in[144] & in2[144];
    assign P[94] = in[144] ^ in2[144];
    assign G[95] = in[143] & in2[143];
    assign P[95] = in[143] ^ in2[143];
    assign G[96] = in[142] & in2[142];
    assign P[96] = in[142] ^ in2[142];
    assign G[97] = in[141] & in2[141];
    assign P[97] = in[141] ^ in2[141];
    assign G[98] = in[140] & in2[140];
    assign P[98] = in[140] ^ in2[140];
    assign G[99] = in[139] & in2[139];
    assign P[99] = in[139] ^ in2[139];
    assign G[100] = in[138] & in2[138];
    assign P[100] = in[138] ^ in2[138];
    assign G[101] = in[137] & in2[137];
    assign P[101] = in[137] ^ in2[137];
    assign G[102] = in[136] & in2[136];
    assign P[102] = in[136] ^ in2[136];
    assign G[103] = in[135] & in2[135];
    assign P[103] = in[135] ^ in2[135];
    assign G[104] = in[134] & in2[134];
    assign P[104] = in[134] ^ in2[134];
    assign G[105] = in[133] & in2[133];
    assign P[105] = in[133] ^ in2[133];
    assign G[106] = in[132] & in2[132];
    assign P[106] = in[132] ^ in2[132];
    assign G[107] = in[131] & in2[131];
    assign P[107] = in[131] ^ in2[131];
    assign G[108] = in[130] & in2[130];
    assign P[108] = in[130] ^ in2[130];
    assign G[109] = in[129] & in2[129];
    assign P[109] = in[129] ^ in2[129];
    assign G[110] = in[128] & in2[128];
    assign P[110] = in[128] ^ in2[128];
    assign G[111] = in[127] & in2[127];
    assign P[111] = in[127] ^ in2[127];
    assign G[112] = in[126] & in2[126];
    assign P[112] = in[126] ^ in2[126];
    assign G[113] = in[125] & in2[125];
    assign P[113] = in[125] ^ in2[125];
    assign G[114] = in[124] & in2[124];
    assign P[114] = in[124] ^ in2[124];
    assign G[115] = in[123] & in2[123];
    assign P[115] = in[123] ^ in2[123];
    assign G[116] = in[122] & in2[122];
    assign P[116] = in[122] ^ in2[122];
    assign G[117] = in[121] & in2[121];
    assign P[117] = in[121] ^ in2[121];
    assign G[118] = in[120] & in2[120];
    assign P[118] = in[120] ^ in2[120];
    assign G[119] = in[119] & in2[119];
    assign P[119] = in[119] ^ in2[119];
    assign G[120] = in[118] & in2[118];
    assign P[120] = in[118] ^ in2[118];
    assign G[121] = in[117] & in2[117];
    assign P[121] = in[117] ^ in2[117];
    assign G[122] = in[116] & in2[116];
    assign P[122] = in[116] ^ in2[116];
    assign G[123] = in[115] & in2[115];
    assign P[123] = in[115] ^ in2[115];
    assign G[124] = in[114] & in2[114];
    assign P[124] = in[114] ^ in2[114];
    assign G[125] = in[113] & in2[113];
    assign P[125] = in[113] ^ in2[113];
    assign G[126] = in[112] & in2[112];
    assign P[126] = in[112] ^ in2[112];
    assign G[127] = in[111] & in2[111];
    assign P[127] = in[111] ^ in2[111];
    assign G[128] = in[110] & in2[110];
    assign P[128] = in[110] ^ in2[110];
    assign G[129] = in[109] & in2[109];
    assign P[129] = in[109] ^ in2[109];
    assign G[130] = in[108] & in2[108];
    assign P[130] = in[108] ^ in2[108];
    assign G[131] = in[107] & in2[107];
    assign P[131] = in[107] ^ in2[107];
    assign G[132] = in[106] & in2[106];
    assign P[132] = in[106] ^ in2[106];
    assign G[133] = in[105] & in2[105];
    assign P[133] = in[105] ^ in2[105];
    assign G[134] = in[104] & in2[104];
    assign P[134] = in[104] ^ in2[104];
    assign G[135] = in[103] & in2[103];
    assign P[135] = in[103] ^ in2[103];
    assign G[136] = in[102] & in2[102];
    assign P[136] = in[102] ^ in2[102];
    assign G[137] = in[101] & in2[101];
    assign P[137] = in[101] ^ in2[101];
    assign G[138] = in[100] & in2[100];
    assign P[138] = in[100] ^ in2[100];
    assign G[139] = in[99] & in2[99];
    assign P[139] = in[99] ^ in2[99];
    assign G[140] = in[98] & in2[98];
    assign P[140] = in[98] ^ in2[98];
    assign G[141] = in[97] & in2[97];
    assign P[141] = in[97] ^ in2[97];
    assign G[142] = in[96] & in2[96];
    assign P[142] = in[96] ^ in2[96];
    assign G[143] = in[95] & in2[95];
    assign P[143] = in[95] ^ in2[95];
    assign G[144] = in[94] & in2[94];
    assign P[144] = in[94] ^ in2[94];
    assign G[145] = in[93] & in2[93];
    assign P[145] = in[93] ^ in2[93];
    assign G[146] = in[92] & in2[92];
    assign P[146] = in[92] ^ in2[92];
    assign G[147] = in[91] & in2[91];
    assign P[147] = in[91] ^ in2[91];
    assign G[148] = in[90] & in2[90];
    assign P[148] = in[90] ^ in2[90];
    assign G[149] = in[89] & in2[89];
    assign P[149] = in[89] ^ in2[89];
    assign G[150] = in[88] & in2[88];
    assign P[150] = in[88] ^ in2[88];
    assign G[151] = in[87] & in2[87];
    assign P[151] = in[87] ^ in2[87];
    assign G[152] = in[86] & in2[86];
    assign P[152] = in[86] ^ in2[86];
    assign G[153] = in[85] & in2[85];
    assign P[153] = in[85] ^ in2[85];
    assign G[154] = in[84] & in2[84];
    assign P[154] = in[84] ^ in2[84];
    assign G[155] = in[83] & in2[83];
    assign P[155] = in[83] ^ in2[83];
    assign G[156] = in[82] & in2[82];
    assign P[156] = in[82] ^ in2[82];
    assign G[157] = in[81] & in2[81];
    assign P[157] = in[81] ^ in2[81];
    assign G[158] = in[80] & in2[80];
    assign P[158] = in[80] ^ in2[80];
    assign G[159] = in[79] & in2[79];
    assign P[159] = in[79] ^ in2[79];
    assign G[160] = in[78] & in2[78];
    assign P[160] = in[78] ^ in2[78];
    assign G[161] = in[77] & in2[77];
    assign P[161] = in[77] ^ in2[77];
    assign G[162] = in[76] & in2[76];
    assign P[162] = in[76] ^ in2[76];
    assign G[163] = in[75] & in2[75];
    assign P[163] = in[75] ^ in2[75];
    assign G[164] = in[74] & in2[74];
    assign P[164] = in[74] ^ in2[74];
    assign G[165] = in[73] & in2[73];
    assign P[165] = in[73] ^ in2[73];
    assign G[166] = in[72] & in2[72];
    assign P[166] = in[72] ^ in2[72];
    assign G[167] = in[71] & in2[71];
    assign P[167] = in[71] ^ in2[71];
    assign G[168] = in[70] & in2[70];
    assign P[168] = in[70] ^ in2[70];
    assign G[169] = in[69] & in2[69];
    assign P[169] = in[69] ^ in2[69];
    assign G[170] = in[68] & in2[68];
    assign P[170] = in[68] ^ in2[68];
    assign G[171] = in[67] & in2[67];
    assign P[171] = in[67] ^ in2[67];
    assign G[172] = in[66] & in2[66];
    assign P[172] = in[66] ^ in2[66];
    assign G[173] = in[65] & in2[65];
    assign P[173] = in[65] ^ in2[65];
    assign G[174] = in[64] & in2[64];
    assign P[174] = in[64] ^ in2[64];
    assign G[175] = in[63] & in2[63];
    assign P[175] = in[63] ^ in2[63];
    assign G[176] = in[62] & in2[62];
    assign P[176] = in[62] ^ in2[62];
    assign G[177] = in[61] & in2[61];
    assign P[177] = in[61] ^ in2[61];
    assign G[178] = in[60] & in2[60];
    assign P[178] = in[60] ^ in2[60];
    assign G[179] = in[59] & in2[59];
    assign P[179] = in[59] ^ in2[59];
    assign G[180] = in[58] & in2[58];
    assign P[180] = in[58] ^ in2[58];
    assign G[181] = in[57] & in2[57];
    assign P[181] = in[57] ^ in2[57];
    assign G[182] = in[56] & in2[56];
    assign P[182] = in[56] ^ in2[56];
    assign G[183] = in[55] & in2[55];
    assign P[183] = in[55] ^ in2[55];
    assign G[184] = in[54] & in2[54];
    assign P[184] = in[54] ^ in2[54];
    assign G[185] = in[53] & in2[53];
    assign P[185] = in[53] ^ in2[53];
    assign G[186] = in[52] & in2[52];
    assign P[186] = in[52] ^ in2[52];
    assign G[187] = in[51] & in2[51];
    assign P[187] = in[51] ^ in2[51];
    assign G[188] = in[50] & in2[50];
    assign P[188] = in[50] ^ in2[50];
    assign G[189] = in[49] & in2[49];
    assign P[189] = in[49] ^ in2[49];
    assign G[190] = in[48] & in2[48];
    assign P[190] = in[48] ^ in2[48];
    assign G[191] = in[47] & in2[47];
    assign P[191] = in[47] ^ in2[47];
    assign G[192] = in[46] & in2[46];
    assign P[192] = in[46] ^ in2[46];
    assign G[193] = in[45] & in2[45];
    assign P[193] = in[45] ^ in2[45];
    assign G[194] = in[44] & in2[44];
    assign P[194] = in[44] ^ in2[44];
    assign G[195] = in[43] & in2[43];
    assign P[195] = in[43] ^ in2[43];
    assign G[196] = in[42] & in2[42];
    assign P[196] = in[42] ^ in2[42];
    assign G[197] = in[41] & in2[41];
    assign P[197] = in[41] ^ in2[41];
    assign G[198] = in[40] & in2[40];
    assign P[198] = in[40] ^ in2[40];
    assign G[199] = in[39] & in2[39];
    assign P[199] = in[39] ^ in2[39];
    assign G[200] = in[38] & in2[38];
    assign P[200] = in[38] ^ in2[38];
    assign G[201] = in[37] & in2[37];
    assign P[201] = in[37] ^ in2[37];
    assign G[202] = in[36] & in2[36];
    assign P[202] = in[36] ^ in2[36];
    assign G[203] = in[35] & in2[35];
    assign P[203] = in[35] ^ in2[35];
    assign G[204] = in[34] & in2[34];
    assign P[204] = in[34] ^ in2[34];
    assign G[205] = in[33] & in2[33];
    assign P[205] = in[33] ^ in2[33];
    assign G[206] = in[32] & in2[32];
    assign P[206] = in[32] ^ in2[32];
    assign G[207] = in[31] & in2[31];
    assign P[207] = in[31] ^ in2[31];
    assign G[208] = in[30] & in2[30];
    assign P[208] = in[30] ^ in2[30];
    assign G[209] = in[29] & in2[29];
    assign P[209] = in[29] ^ in2[29];
    assign G[210] = in[28] & in2[28];
    assign P[210] = in[28] ^ in2[28];
    assign G[211] = in[27] & in2[27];
    assign P[211] = in[27] ^ in2[27];
    assign G[212] = in[26] & in2[26];
    assign P[212] = in[26] ^ in2[26];
    assign G[213] = in[25] & in2[25];
    assign P[213] = in[25] ^ in2[25];
    assign G[214] = in[24] & in2[24];
    assign P[214] = in[24] ^ in2[24];
    assign G[215] = in[23] & in2[23];
    assign P[215] = in[23] ^ in2[23];
    assign G[216] = in[22] & in2[22];
    assign P[216] = in[22] ^ in2[22];
    assign G[217] = in[21] & in2[21];
    assign P[217] = in[21] ^ in2[21];
    assign G[218] = in[20] & in2[20];
    assign P[218] = in[20] ^ in2[20];
    assign G[219] = in[19] & in2[19];
    assign P[219] = in[19] ^ in2[19];
    assign G[220] = in[18] & in2[18];
    assign P[220] = in[18] ^ in2[18];
    assign G[221] = in[17] & in2[17];
    assign P[221] = in[17] ^ in2[17];
    assign G[222] = in[16] & in2[16];
    assign P[222] = in[16] ^ in2[16];
    assign G[223] = in[15] & in2[15];
    assign P[223] = in[15] ^ in2[15];
    assign G[224] = in[14] & in2[14];
    assign P[224] = in[14] ^ in2[14];
    assign G[225] = in[13] & in2[13];
    assign P[225] = in[13] ^ in2[13];
    assign G[226] = in[12] & in2[12];
    assign P[226] = in[12] ^ in2[12];
    assign G[227] = in[11] & in2[11];
    assign P[227] = in[11] ^ in2[11];
    assign G[228] = in[10] & in2[10];
    assign P[228] = in[10] ^ in2[10];
    assign G[229] = in[9] & in2[9];
    assign P[229] = in[9] ^ in2[9];
    assign G[230] = in[8] & in2[8];
    assign P[230] = in[8] ^ in2[8];
    assign G[231] = in[7] & in2[7];
    assign P[231] = in[7] ^ in2[7];
    assign G[232] = in[6] & in2[6];
    assign P[232] = in[6] ^ in2[6];
    assign G[233] = in[5] & in2[5];
    assign P[233] = in[5] ^ in2[5];
    assign G[234] = in[4] & in2[4];
    assign P[234] = in[4] ^ in2[4];
    assign G[235] = in[3] & in2[3];
    assign P[235] = in[3] ^ in2[3];
    assign G[236] = in[2] & in2[2];
    assign P[236] = in[2] ^ in2[2];
    assign G[237] = in[1] & in2[1];
    assign P[237] = in[1] ^ in2[1];
    assign G[238] = in[0] & in2[0];
    assign P[238] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign C[238] = G[237] | (P[237] & C[237]);
    assign cout = G[238] | (P[238] & C[238]);
    assign sum = P ^ C;
endmodule

module CLA238(output [237:0] sum, output cout, input [237:0] in1, input [237:0] in2;

    wire[237:0] G;
    wire[237:0] C;
    wire[237:0] P;

    assign G[0] = in[237] & in2[237];
    assign P[0] = in[237] ^ in2[237];
    assign G[1] = in[236] & in2[236];
    assign P[1] = in[236] ^ in2[236];
    assign G[2] = in[235] & in2[235];
    assign P[2] = in[235] ^ in2[235];
    assign G[3] = in[234] & in2[234];
    assign P[3] = in[234] ^ in2[234];
    assign G[4] = in[233] & in2[233];
    assign P[4] = in[233] ^ in2[233];
    assign G[5] = in[232] & in2[232];
    assign P[5] = in[232] ^ in2[232];
    assign G[6] = in[231] & in2[231];
    assign P[6] = in[231] ^ in2[231];
    assign G[7] = in[230] & in2[230];
    assign P[7] = in[230] ^ in2[230];
    assign G[8] = in[229] & in2[229];
    assign P[8] = in[229] ^ in2[229];
    assign G[9] = in[228] & in2[228];
    assign P[9] = in[228] ^ in2[228];
    assign G[10] = in[227] & in2[227];
    assign P[10] = in[227] ^ in2[227];
    assign G[11] = in[226] & in2[226];
    assign P[11] = in[226] ^ in2[226];
    assign G[12] = in[225] & in2[225];
    assign P[12] = in[225] ^ in2[225];
    assign G[13] = in[224] & in2[224];
    assign P[13] = in[224] ^ in2[224];
    assign G[14] = in[223] & in2[223];
    assign P[14] = in[223] ^ in2[223];
    assign G[15] = in[222] & in2[222];
    assign P[15] = in[222] ^ in2[222];
    assign G[16] = in[221] & in2[221];
    assign P[16] = in[221] ^ in2[221];
    assign G[17] = in[220] & in2[220];
    assign P[17] = in[220] ^ in2[220];
    assign G[18] = in[219] & in2[219];
    assign P[18] = in[219] ^ in2[219];
    assign G[19] = in[218] & in2[218];
    assign P[19] = in[218] ^ in2[218];
    assign G[20] = in[217] & in2[217];
    assign P[20] = in[217] ^ in2[217];
    assign G[21] = in[216] & in2[216];
    assign P[21] = in[216] ^ in2[216];
    assign G[22] = in[215] & in2[215];
    assign P[22] = in[215] ^ in2[215];
    assign G[23] = in[214] & in2[214];
    assign P[23] = in[214] ^ in2[214];
    assign G[24] = in[213] & in2[213];
    assign P[24] = in[213] ^ in2[213];
    assign G[25] = in[212] & in2[212];
    assign P[25] = in[212] ^ in2[212];
    assign G[26] = in[211] & in2[211];
    assign P[26] = in[211] ^ in2[211];
    assign G[27] = in[210] & in2[210];
    assign P[27] = in[210] ^ in2[210];
    assign G[28] = in[209] & in2[209];
    assign P[28] = in[209] ^ in2[209];
    assign G[29] = in[208] & in2[208];
    assign P[29] = in[208] ^ in2[208];
    assign G[30] = in[207] & in2[207];
    assign P[30] = in[207] ^ in2[207];
    assign G[31] = in[206] & in2[206];
    assign P[31] = in[206] ^ in2[206];
    assign G[32] = in[205] & in2[205];
    assign P[32] = in[205] ^ in2[205];
    assign G[33] = in[204] & in2[204];
    assign P[33] = in[204] ^ in2[204];
    assign G[34] = in[203] & in2[203];
    assign P[34] = in[203] ^ in2[203];
    assign G[35] = in[202] & in2[202];
    assign P[35] = in[202] ^ in2[202];
    assign G[36] = in[201] & in2[201];
    assign P[36] = in[201] ^ in2[201];
    assign G[37] = in[200] & in2[200];
    assign P[37] = in[200] ^ in2[200];
    assign G[38] = in[199] & in2[199];
    assign P[38] = in[199] ^ in2[199];
    assign G[39] = in[198] & in2[198];
    assign P[39] = in[198] ^ in2[198];
    assign G[40] = in[197] & in2[197];
    assign P[40] = in[197] ^ in2[197];
    assign G[41] = in[196] & in2[196];
    assign P[41] = in[196] ^ in2[196];
    assign G[42] = in[195] & in2[195];
    assign P[42] = in[195] ^ in2[195];
    assign G[43] = in[194] & in2[194];
    assign P[43] = in[194] ^ in2[194];
    assign G[44] = in[193] & in2[193];
    assign P[44] = in[193] ^ in2[193];
    assign G[45] = in[192] & in2[192];
    assign P[45] = in[192] ^ in2[192];
    assign G[46] = in[191] & in2[191];
    assign P[46] = in[191] ^ in2[191];
    assign G[47] = in[190] & in2[190];
    assign P[47] = in[190] ^ in2[190];
    assign G[48] = in[189] & in2[189];
    assign P[48] = in[189] ^ in2[189];
    assign G[49] = in[188] & in2[188];
    assign P[49] = in[188] ^ in2[188];
    assign G[50] = in[187] & in2[187];
    assign P[50] = in[187] ^ in2[187];
    assign G[51] = in[186] & in2[186];
    assign P[51] = in[186] ^ in2[186];
    assign G[52] = in[185] & in2[185];
    assign P[52] = in[185] ^ in2[185];
    assign G[53] = in[184] & in2[184];
    assign P[53] = in[184] ^ in2[184];
    assign G[54] = in[183] & in2[183];
    assign P[54] = in[183] ^ in2[183];
    assign G[55] = in[182] & in2[182];
    assign P[55] = in[182] ^ in2[182];
    assign G[56] = in[181] & in2[181];
    assign P[56] = in[181] ^ in2[181];
    assign G[57] = in[180] & in2[180];
    assign P[57] = in[180] ^ in2[180];
    assign G[58] = in[179] & in2[179];
    assign P[58] = in[179] ^ in2[179];
    assign G[59] = in[178] & in2[178];
    assign P[59] = in[178] ^ in2[178];
    assign G[60] = in[177] & in2[177];
    assign P[60] = in[177] ^ in2[177];
    assign G[61] = in[176] & in2[176];
    assign P[61] = in[176] ^ in2[176];
    assign G[62] = in[175] & in2[175];
    assign P[62] = in[175] ^ in2[175];
    assign G[63] = in[174] & in2[174];
    assign P[63] = in[174] ^ in2[174];
    assign G[64] = in[173] & in2[173];
    assign P[64] = in[173] ^ in2[173];
    assign G[65] = in[172] & in2[172];
    assign P[65] = in[172] ^ in2[172];
    assign G[66] = in[171] & in2[171];
    assign P[66] = in[171] ^ in2[171];
    assign G[67] = in[170] & in2[170];
    assign P[67] = in[170] ^ in2[170];
    assign G[68] = in[169] & in2[169];
    assign P[68] = in[169] ^ in2[169];
    assign G[69] = in[168] & in2[168];
    assign P[69] = in[168] ^ in2[168];
    assign G[70] = in[167] & in2[167];
    assign P[70] = in[167] ^ in2[167];
    assign G[71] = in[166] & in2[166];
    assign P[71] = in[166] ^ in2[166];
    assign G[72] = in[165] & in2[165];
    assign P[72] = in[165] ^ in2[165];
    assign G[73] = in[164] & in2[164];
    assign P[73] = in[164] ^ in2[164];
    assign G[74] = in[163] & in2[163];
    assign P[74] = in[163] ^ in2[163];
    assign G[75] = in[162] & in2[162];
    assign P[75] = in[162] ^ in2[162];
    assign G[76] = in[161] & in2[161];
    assign P[76] = in[161] ^ in2[161];
    assign G[77] = in[160] & in2[160];
    assign P[77] = in[160] ^ in2[160];
    assign G[78] = in[159] & in2[159];
    assign P[78] = in[159] ^ in2[159];
    assign G[79] = in[158] & in2[158];
    assign P[79] = in[158] ^ in2[158];
    assign G[80] = in[157] & in2[157];
    assign P[80] = in[157] ^ in2[157];
    assign G[81] = in[156] & in2[156];
    assign P[81] = in[156] ^ in2[156];
    assign G[82] = in[155] & in2[155];
    assign P[82] = in[155] ^ in2[155];
    assign G[83] = in[154] & in2[154];
    assign P[83] = in[154] ^ in2[154];
    assign G[84] = in[153] & in2[153];
    assign P[84] = in[153] ^ in2[153];
    assign G[85] = in[152] & in2[152];
    assign P[85] = in[152] ^ in2[152];
    assign G[86] = in[151] & in2[151];
    assign P[86] = in[151] ^ in2[151];
    assign G[87] = in[150] & in2[150];
    assign P[87] = in[150] ^ in2[150];
    assign G[88] = in[149] & in2[149];
    assign P[88] = in[149] ^ in2[149];
    assign G[89] = in[148] & in2[148];
    assign P[89] = in[148] ^ in2[148];
    assign G[90] = in[147] & in2[147];
    assign P[90] = in[147] ^ in2[147];
    assign G[91] = in[146] & in2[146];
    assign P[91] = in[146] ^ in2[146];
    assign G[92] = in[145] & in2[145];
    assign P[92] = in[145] ^ in2[145];
    assign G[93] = in[144] & in2[144];
    assign P[93] = in[144] ^ in2[144];
    assign G[94] = in[143] & in2[143];
    assign P[94] = in[143] ^ in2[143];
    assign G[95] = in[142] & in2[142];
    assign P[95] = in[142] ^ in2[142];
    assign G[96] = in[141] & in2[141];
    assign P[96] = in[141] ^ in2[141];
    assign G[97] = in[140] & in2[140];
    assign P[97] = in[140] ^ in2[140];
    assign G[98] = in[139] & in2[139];
    assign P[98] = in[139] ^ in2[139];
    assign G[99] = in[138] & in2[138];
    assign P[99] = in[138] ^ in2[138];
    assign G[100] = in[137] & in2[137];
    assign P[100] = in[137] ^ in2[137];
    assign G[101] = in[136] & in2[136];
    assign P[101] = in[136] ^ in2[136];
    assign G[102] = in[135] & in2[135];
    assign P[102] = in[135] ^ in2[135];
    assign G[103] = in[134] & in2[134];
    assign P[103] = in[134] ^ in2[134];
    assign G[104] = in[133] & in2[133];
    assign P[104] = in[133] ^ in2[133];
    assign G[105] = in[132] & in2[132];
    assign P[105] = in[132] ^ in2[132];
    assign G[106] = in[131] & in2[131];
    assign P[106] = in[131] ^ in2[131];
    assign G[107] = in[130] & in2[130];
    assign P[107] = in[130] ^ in2[130];
    assign G[108] = in[129] & in2[129];
    assign P[108] = in[129] ^ in2[129];
    assign G[109] = in[128] & in2[128];
    assign P[109] = in[128] ^ in2[128];
    assign G[110] = in[127] & in2[127];
    assign P[110] = in[127] ^ in2[127];
    assign G[111] = in[126] & in2[126];
    assign P[111] = in[126] ^ in2[126];
    assign G[112] = in[125] & in2[125];
    assign P[112] = in[125] ^ in2[125];
    assign G[113] = in[124] & in2[124];
    assign P[113] = in[124] ^ in2[124];
    assign G[114] = in[123] & in2[123];
    assign P[114] = in[123] ^ in2[123];
    assign G[115] = in[122] & in2[122];
    assign P[115] = in[122] ^ in2[122];
    assign G[116] = in[121] & in2[121];
    assign P[116] = in[121] ^ in2[121];
    assign G[117] = in[120] & in2[120];
    assign P[117] = in[120] ^ in2[120];
    assign G[118] = in[119] & in2[119];
    assign P[118] = in[119] ^ in2[119];
    assign G[119] = in[118] & in2[118];
    assign P[119] = in[118] ^ in2[118];
    assign G[120] = in[117] & in2[117];
    assign P[120] = in[117] ^ in2[117];
    assign G[121] = in[116] & in2[116];
    assign P[121] = in[116] ^ in2[116];
    assign G[122] = in[115] & in2[115];
    assign P[122] = in[115] ^ in2[115];
    assign G[123] = in[114] & in2[114];
    assign P[123] = in[114] ^ in2[114];
    assign G[124] = in[113] & in2[113];
    assign P[124] = in[113] ^ in2[113];
    assign G[125] = in[112] & in2[112];
    assign P[125] = in[112] ^ in2[112];
    assign G[126] = in[111] & in2[111];
    assign P[126] = in[111] ^ in2[111];
    assign G[127] = in[110] & in2[110];
    assign P[127] = in[110] ^ in2[110];
    assign G[128] = in[109] & in2[109];
    assign P[128] = in[109] ^ in2[109];
    assign G[129] = in[108] & in2[108];
    assign P[129] = in[108] ^ in2[108];
    assign G[130] = in[107] & in2[107];
    assign P[130] = in[107] ^ in2[107];
    assign G[131] = in[106] & in2[106];
    assign P[131] = in[106] ^ in2[106];
    assign G[132] = in[105] & in2[105];
    assign P[132] = in[105] ^ in2[105];
    assign G[133] = in[104] & in2[104];
    assign P[133] = in[104] ^ in2[104];
    assign G[134] = in[103] & in2[103];
    assign P[134] = in[103] ^ in2[103];
    assign G[135] = in[102] & in2[102];
    assign P[135] = in[102] ^ in2[102];
    assign G[136] = in[101] & in2[101];
    assign P[136] = in[101] ^ in2[101];
    assign G[137] = in[100] & in2[100];
    assign P[137] = in[100] ^ in2[100];
    assign G[138] = in[99] & in2[99];
    assign P[138] = in[99] ^ in2[99];
    assign G[139] = in[98] & in2[98];
    assign P[139] = in[98] ^ in2[98];
    assign G[140] = in[97] & in2[97];
    assign P[140] = in[97] ^ in2[97];
    assign G[141] = in[96] & in2[96];
    assign P[141] = in[96] ^ in2[96];
    assign G[142] = in[95] & in2[95];
    assign P[142] = in[95] ^ in2[95];
    assign G[143] = in[94] & in2[94];
    assign P[143] = in[94] ^ in2[94];
    assign G[144] = in[93] & in2[93];
    assign P[144] = in[93] ^ in2[93];
    assign G[145] = in[92] & in2[92];
    assign P[145] = in[92] ^ in2[92];
    assign G[146] = in[91] & in2[91];
    assign P[146] = in[91] ^ in2[91];
    assign G[147] = in[90] & in2[90];
    assign P[147] = in[90] ^ in2[90];
    assign G[148] = in[89] & in2[89];
    assign P[148] = in[89] ^ in2[89];
    assign G[149] = in[88] & in2[88];
    assign P[149] = in[88] ^ in2[88];
    assign G[150] = in[87] & in2[87];
    assign P[150] = in[87] ^ in2[87];
    assign G[151] = in[86] & in2[86];
    assign P[151] = in[86] ^ in2[86];
    assign G[152] = in[85] & in2[85];
    assign P[152] = in[85] ^ in2[85];
    assign G[153] = in[84] & in2[84];
    assign P[153] = in[84] ^ in2[84];
    assign G[154] = in[83] & in2[83];
    assign P[154] = in[83] ^ in2[83];
    assign G[155] = in[82] & in2[82];
    assign P[155] = in[82] ^ in2[82];
    assign G[156] = in[81] & in2[81];
    assign P[156] = in[81] ^ in2[81];
    assign G[157] = in[80] & in2[80];
    assign P[157] = in[80] ^ in2[80];
    assign G[158] = in[79] & in2[79];
    assign P[158] = in[79] ^ in2[79];
    assign G[159] = in[78] & in2[78];
    assign P[159] = in[78] ^ in2[78];
    assign G[160] = in[77] & in2[77];
    assign P[160] = in[77] ^ in2[77];
    assign G[161] = in[76] & in2[76];
    assign P[161] = in[76] ^ in2[76];
    assign G[162] = in[75] & in2[75];
    assign P[162] = in[75] ^ in2[75];
    assign G[163] = in[74] & in2[74];
    assign P[163] = in[74] ^ in2[74];
    assign G[164] = in[73] & in2[73];
    assign P[164] = in[73] ^ in2[73];
    assign G[165] = in[72] & in2[72];
    assign P[165] = in[72] ^ in2[72];
    assign G[166] = in[71] & in2[71];
    assign P[166] = in[71] ^ in2[71];
    assign G[167] = in[70] & in2[70];
    assign P[167] = in[70] ^ in2[70];
    assign G[168] = in[69] & in2[69];
    assign P[168] = in[69] ^ in2[69];
    assign G[169] = in[68] & in2[68];
    assign P[169] = in[68] ^ in2[68];
    assign G[170] = in[67] & in2[67];
    assign P[170] = in[67] ^ in2[67];
    assign G[171] = in[66] & in2[66];
    assign P[171] = in[66] ^ in2[66];
    assign G[172] = in[65] & in2[65];
    assign P[172] = in[65] ^ in2[65];
    assign G[173] = in[64] & in2[64];
    assign P[173] = in[64] ^ in2[64];
    assign G[174] = in[63] & in2[63];
    assign P[174] = in[63] ^ in2[63];
    assign G[175] = in[62] & in2[62];
    assign P[175] = in[62] ^ in2[62];
    assign G[176] = in[61] & in2[61];
    assign P[176] = in[61] ^ in2[61];
    assign G[177] = in[60] & in2[60];
    assign P[177] = in[60] ^ in2[60];
    assign G[178] = in[59] & in2[59];
    assign P[178] = in[59] ^ in2[59];
    assign G[179] = in[58] & in2[58];
    assign P[179] = in[58] ^ in2[58];
    assign G[180] = in[57] & in2[57];
    assign P[180] = in[57] ^ in2[57];
    assign G[181] = in[56] & in2[56];
    assign P[181] = in[56] ^ in2[56];
    assign G[182] = in[55] & in2[55];
    assign P[182] = in[55] ^ in2[55];
    assign G[183] = in[54] & in2[54];
    assign P[183] = in[54] ^ in2[54];
    assign G[184] = in[53] & in2[53];
    assign P[184] = in[53] ^ in2[53];
    assign G[185] = in[52] & in2[52];
    assign P[185] = in[52] ^ in2[52];
    assign G[186] = in[51] & in2[51];
    assign P[186] = in[51] ^ in2[51];
    assign G[187] = in[50] & in2[50];
    assign P[187] = in[50] ^ in2[50];
    assign G[188] = in[49] & in2[49];
    assign P[188] = in[49] ^ in2[49];
    assign G[189] = in[48] & in2[48];
    assign P[189] = in[48] ^ in2[48];
    assign G[190] = in[47] & in2[47];
    assign P[190] = in[47] ^ in2[47];
    assign G[191] = in[46] & in2[46];
    assign P[191] = in[46] ^ in2[46];
    assign G[192] = in[45] & in2[45];
    assign P[192] = in[45] ^ in2[45];
    assign G[193] = in[44] & in2[44];
    assign P[193] = in[44] ^ in2[44];
    assign G[194] = in[43] & in2[43];
    assign P[194] = in[43] ^ in2[43];
    assign G[195] = in[42] & in2[42];
    assign P[195] = in[42] ^ in2[42];
    assign G[196] = in[41] & in2[41];
    assign P[196] = in[41] ^ in2[41];
    assign G[197] = in[40] & in2[40];
    assign P[197] = in[40] ^ in2[40];
    assign G[198] = in[39] & in2[39];
    assign P[198] = in[39] ^ in2[39];
    assign G[199] = in[38] & in2[38];
    assign P[199] = in[38] ^ in2[38];
    assign G[200] = in[37] & in2[37];
    assign P[200] = in[37] ^ in2[37];
    assign G[201] = in[36] & in2[36];
    assign P[201] = in[36] ^ in2[36];
    assign G[202] = in[35] & in2[35];
    assign P[202] = in[35] ^ in2[35];
    assign G[203] = in[34] & in2[34];
    assign P[203] = in[34] ^ in2[34];
    assign G[204] = in[33] & in2[33];
    assign P[204] = in[33] ^ in2[33];
    assign G[205] = in[32] & in2[32];
    assign P[205] = in[32] ^ in2[32];
    assign G[206] = in[31] & in2[31];
    assign P[206] = in[31] ^ in2[31];
    assign G[207] = in[30] & in2[30];
    assign P[207] = in[30] ^ in2[30];
    assign G[208] = in[29] & in2[29];
    assign P[208] = in[29] ^ in2[29];
    assign G[209] = in[28] & in2[28];
    assign P[209] = in[28] ^ in2[28];
    assign G[210] = in[27] & in2[27];
    assign P[210] = in[27] ^ in2[27];
    assign G[211] = in[26] & in2[26];
    assign P[211] = in[26] ^ in2[26];
    assign G[212] = in[25] & in2[25];
    assign P[212] = in[25] ^ in2[25];
    assign G[213] = in[24] & in2[24];
    assign P[213] = in[24] ^ in2[24];
    assign G[214] = in[23] & in2[23];
    assign P[214] = in[23] ^ in2[23];
    assign G[215] = in[22] & in2[22];
    assign P[215] = in[22] ^ in2[22];
    assign G[216] = in[21] & in2[21];
    assign P[216] = in[21] ^ in2[21];
    assign G[217] = in[20] & in2[20];
    assign P[217] = in[20] ^ in2[20];
    assign G[218] = in[19] & in2[19];
    assign P[218] = in[19] ^ in2[19];
    assign G[219] = in[18] & in2[18];
    assign P[219] = in[18] ^ in2[18];
    assign G[220] = in[17] & in2[17];
    assign P[220] = in[17] ^ in2[17];
    assign G[221] = in[16] & in2[16];
    assign P[221] = in[16] ^ in2[16];
    assign G[222] = in[15] & in2[15];
    assign P[222] = in[15] ^ in2[15];
    assign G[223] = in[14] & in2[14];
    assign P[223] = in[14] ^ in2[14];
    assign G[224] = in[13] & in2[13];
    assign P[224] = in[13] ^ in2[13];
    assign G[225] = in[12] & in2[12];
    assign P[225] = in[12] ^ in2[12];
    assign G[226] = in[11] & in2[11];
    assign P[226] = in[11] ^ in2[11];
    assign G[227] = in[10] & in2[10];
    assign P[227] = in[10] ^ in2[10];
    assign G[228] = in[9] & in2[9];
    assign P[228] = in[9] ^ in2[9];
    assign G[229] = in[8] & in2[8];
    assign P[229] = in[8] ^ in2[8];
    assign G[230] = in[7] & in2[7];
    assign P[230] = in[7] ^ in2[7];
    assign G[231] = in[6] & in2[6];
    assign P[231] = in[6] ^ in2[6];
    assign G[232] = in[5] & in2[5];
    assign P[232] = in[5] ^ in2[5];
    assign G[233] = in[4] & in2[4];
    assign P[233] = in[4] ^ in2[4];
    assign G[234] = in[3] & in2[3];
    assign P[234] = in[3] ^ in2[3];
    assign G[235] = in[2] & in2[2];
    assign P[235] = in[2] ^ in2[2];
    assign G[236] = in[1] & in2[1];
    assign P[236] = in[1] ^ in2[1];
    assign G[237] = in[0] & in2[0];
    assign P[237] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign C[237] = G[236] | (P[236] & C[236]);
    assign cout = G[237] | (P[237] & C[237]);
    assign sum = P ^ C;
endmodule

module CLA237(output [236:0] sum, output cout, input [236:0] in1, input [236:0] in2;

    wire[236:0] G;
    wire[236:0] C;
    wire[236:0] P;

    assign G[0] = in[236] & in2[236];
    assign P[0] = in[236] ^ in2[236];
    assign G[1] = in[235] & in2[235];
    assign P[1] = in[235] ^ in2[235];
    assign G[2] = in[234] & in2[234];
    assign P[2] = in[234] ^ in2[234];
    assign G[3] = in[233] & in2[233];
    assign P[3] = in[233] ^ in2[233];
    assign G[4] = in[232] & in2[232];
    assign P[4] = in[232] ^ in2[232];
    assign G[5] = in[231] & in2[231];
    assign P[5] = in[231] ^ in2[231];
    assign G[6] = in[230] & in2[230];
    assign P[6] = in[230] ^ in2[230];
    assign G[7] = in[229] & in2[229];
    assign P[7] = in[229] ^ in2[229];
    assign G[8] = in[228] & in2[228];
    assign P[8] = in[228] ^ in2[228];
    assign G[9] = in[227] & in2[227];
    assign P[9] = in[227] ^ in2[227];
    assign G[10] = in[226] & in2[226];
    assign P[10] = in[226] ^ in2[226];
    assign G[11] = in[225] & in2[225];
    assign P[11] = in[225] ^ in2[225];
    assign G[12] = in[224] & in2[224];
    assign P[12] = in[224] ^ in2[224];
    assign G[13] = in[223] & in2[223];
    assign P[13] = in[223] ^ in2[223];
    assign G[14] = in[222] & in2[222];
    assign P[14] = in[222] ^ in2[222];
    assign G[15] = in[221] & in2[221];
    assign P[15] = in[221] ^ in2[221];
    assign G[16] = in[220] & in2[220];
    assign P[16] = in[220] ^ in2[220];
    assign G[17] = in[219] & in2[219];
    assign P[17] = in[219] ^ in2[219];
    assign G[18] = in[218] & in2[218];
    assign P[18] = in[218] ^ in2[218];
    assign G[19] = in[217] & in2[217];
    assign P[19] = in[217] ^ in2[217];
    assign G[20] = in[216] & in2[216];
    assign P[20] = in[216] ^ in2[216];
    assign G[21] = in[215] & in2[215];
    assign P[21] = in[215] ^ in2[215];
    assign G[22] = in[214] & in2[214];
    assign P[22] = in[214] ^ in2[214];
    assign G[23] = in[213] & in2[213];
    assign P[23] = in[213] ^ in2[213];
    assign G[24] = in[212] & in2[212];
    assign P[24] = in[212] ^ in2[212];
    assign G[25] = in[211] & in2[211];
    assign P[25] = in[211] ^ in2[211];
    assign G[26] = in[210] & in2[210];
    assign P[26] = in[210] ^ in2[210];
    assign G[27] = in[209] & in2[209];
    assign P[27] = in[209] ^ in2[209];
    assign G[28] = in[208] & in2[208];
    assign P[28] = in[208] ^ in2[208];
    assign G[29] = in[207] & in2[207];
    assign P[29] = in[207] ^ in2[207];
    assign G[30] = in[206] & in2[206];
    assign P[30] = in[206] ^ in2[206];
    assign G[31] = in[205] & in2[205];
    assign P[31] = in[205] ^ in2[205];
    assign G[32] = in[204] & in2[204];
    assign P[32] = in[204] ^ in2[204];
    assign G[33] = in[203] & in2[203];
    assign P[33] = in[203] ^ in2[203];
    assign G[34] = in[202] & in2[202];
    assign P[34] = in[202] ^ in2[202];
    assign G[35] = in[201] & in2[201];
    assign P[35] = in[201] ^ in2[201];
    assign G[36] = in[200] & in2[200];
    assign P[36] = in[200] ^ in2[200];
    assign G[37] = in[199] & in2[199];
    assign P[37] = in[199] ^ in2[199];
    assign G[38] = in[198] & in2[198];
    assign P[38] = in[198] ^ in2[198];
    assign G[39] = in[197] & in2[197];
    assign P[39] = in[197] ^ in2[197];
    assign G[40] = in[196] & in2[196];
    assign P[40] = in[196] ^ in2[196];
    assign G[41] = in[195] & in2[195];
    assign P[41] = in[195] ^ in2[195];
    assign G[42] = in[194] & in2[194];
    assign P[42] = in[194] ^ in2[194];
    assign G[43] = in[193] & in2[193];
    assign P[43] = in[193] ^ in2[193];
    assign G[44] = in[192] & in2[192];
    assign P[44] = in[192] ^ in2[192];
    assign G[45] = in[191] & in2[191];
    assign P[45] = in[191] ^ in2[191];
    assign G[46] = in[190] & in2[190];
    assign P[46] = in[190] ^ in2[190];
    assign G[47] = in[189] & in2[189];
    assign P[47] = in[189] ^ in2[189];
    assign G[48] = in[188] & in2[188];
    assign P[48] = in[188] ^ in2[188];
    assign G[49] = in[187] & in2[187];
    assign P[49] = in[187] ^ in2[187];
    assign G[50] = in[186] & in2[186];
    assign P[50] = in[186] ^ in2[186];
    assign G[51] = in[185] & in2[185];
    assign P[51] = in[185] ^ in2[185];
    assign G[52] = in[184] & in2[184];
    assign P[52] = in[184] ^ in2[184];
    assign G[53] = in[183] & in2[183];
    assign P[53] = in[183] ^ in2[183];
    assign G[54] = in[182] & in2[182];
    assign P[54] = in[182] ^ in2[182];
    assign G[55] = in[181] & in2[181];
    assign P[55] = in[181] ^ in2[181];
    assign G[56] = in[180] & in2[180];
    assign P[56] = in[180] ^ in2[180];
    assign G[57] = in[179] & in2[179];
    assign P[57] = in[179] ^ in2[179];
    assign G[58] = in[178] & in2[178];
    assign P[58] = in[178] ^ in2[178];
    assign G[59] = in[177] & in2[177];
    assign P[59] = in[177] ^ in2[177];
    assign G[60] = in[176] & in2[176];
    assign P[60] = in[176] ^ in2[176];
    assign G[61] = in[175] & in2[175];
    assign P[61] = in[175] ^ in2[175];
    assign G[62] = in[174] & in2[174];
    assign P[62] = in[174] ^ in2[174];
    assign G[63] = in[173] & in2[173];
    assign P[63] = in[173] ^ in2[173];
    assign G[64] = in[172] & in2[172];
    assign P[64] = in[172] ^ in2[172];
    assign G[65] = in[171] & in2[171];
    assign P[65] = in[171] ^ in2[171];
    assign G[66] = in[170] & in2[170];
    assign P[66] = in[170] ^ in2[170];
    assign G[67] = in[169] & in2[169];
    assign P[67] = in[169] ^ in2[169];
    assign G[68] = in[168] & in2[168];
    assign P[68] = in[168] ^ in2[168];
    assign G[69] = in[167] & in2[167];
    assign P[69] = in[167] ^ in2[167];
    assign G[70] = in[166] & in2[166];
    assign P[70] = in[166] ^ in2[166];
    assign G[71] = in[165] & in2[165];
    assign P[71] = in[165] ^ in2[165];
    assign G[72] = in[164] & in2[164];
    assign P[72] = in[164] ^ in2[164];
    assign G[73] = in[163] & in2[163];
    assign P[73] = in[163] ^ in2[163];
    assign G[74] = in[162] & in2[162];
    assign P[74] = in[162] ^ in2[162];
    assign G[75] = in[161] & in2[161];
    assign P[75] = in[161] ^ in2[161];
    assign G[76] = in[160] & in2[160];
    assign P[76] = in[160] ^ in2[160];
    assign G[77] = in[159] & in2[159];
    assign P[77] = in[159] ^ in2[159];
    assign G[78] = in[158] & in2[158];
    assign P[78] = in[158] ^ in2[158];
    assign G[79] = in[157] & in2[157];
    assign P[79] = in[157] ^ in2[157];
    assign G[80] = in[156] & in2[156];
    assign P[80] = in[156] ^ in2[156];
    assign G[81] = in[155] & in2[155];
    assign P[81] = in[155] ^ in2[155];
    assign G[82] = in[154] & in2[154];
    assign P[82] = in[154] ^ in2[154];
    assign G[83] = in[153] & in2[153];
    assign P[83] = in[153] ^ in2[153];
    assign G[84] = in[152] & in2[152];
    assign P[84] = in[152] ^ in2[152];
    assign G[85] = in[151] & in2[151];
    assign P[85] = in[151] ^ in2[151];
    assign G[86] = in[150] & in2[150];
    assign P[86] = in[150] ^ in2[150];
    assign G[87] = in[149] & in2[149];
    assign P[87] = in[149] ^ in2[149];
    assign G[88] = in[148] & in2[148];
    assign P[88] = in[148] ^ in2[148];
    assign G[89] = in[147] & in2[147];
    assign P[89] = in[147] ^ in2[147];
    assign G[90] = in[146] & in2[146];
    assign P[90] = in[146] ^ in2[146];
    assign G[91] = in[145] & in2[145];
    assign P[91] = in[145] ^ in2[145];
    assign G[92] = in[144] & in2[144];
    assign P[92] = in[144] ^ in2[144];
    assign G[93] = in[143] & in2[143];
    assign P[93] = in[143] ^ in2[143];
    assign G[94] = in[142] & in2[142];
    assign P[94] = in[142] ^ in2[142];
    assign G[95] = in[141] & in2[141];
    assign P[95] = in[141] ^ in2[141];
    assign G[96] = in[140] & in2[140];
    assign P[96] = in[140] ^ in2[140];
    assign G[97] = in[139] & in2[139];
    assign P[97] = in[139] ^ in2[139];
    assign G[98] = in[138] & in2[138];
    assign P[98] = in[138] ^ in2[138];
    assign G[99] = in[137] & in2[137];
    assign P[99] = in[137] ^ in2[137];
    assign G[100] = in[136] & in2[136];
    assign P[100] = in[136] ^ in2[136];
    assign G[101] = in[135] & in2[135];
    assign P[101] = in[135] ^ in2[135];
    assign G[102] = in[134] & in2[134];
    assign P[102] = in[134] ^ in2[134];
    assign G[103] = in[133] & in2[133];
    assign P[103] = in[133] ^ in2[133];
    assign G[104] = in[132] & in2[132];
    assign P[104] = in[132] ^ in2[132];
    assign G[105] = in[131] & in2[131];
    assign P[105] = in[131] ^ in2[131];
    assign G[106] = in[130] & in2[130];
    assign P[106] = in[130] ^ in2[130];
    assign G[107] = in[129] & in2[129];
    assign P[107] = in[129] ^ in2[129];
    assign G[108] = in[128] & in2[128];
    assign P[108] = in[128] ^ in2[128];
    assign G[109] = in[127] & in2[127];
    assign P[109] = in[127] ^ in2[127];
    assign G[110] = in[126] & in2[126];
    assign P[110] = in[126] ^ in2[126];
    assign G[111] = in[125] & in2[125];
    assign P[111] = in[125] ^ in2[125];
    assign G[112] = in[124] & in2[124];
    assign P[112] = in[124] ^ in2[124];
    assign G[113] = in[123] & in2[123];
    assign P[113] = in[123] ^ in2[123];
    assign G[114] = in[122] & in2[122];
    assign P[114] = in[122] ^ in2[122];
    assign G[115] = in[121] & in2[121];
    assign P[115] = in[121] ^ in2[121];
    assign G[116] = in[120] & in2[120];
    assign P[116] = in[120] ^ in2[120];
    assign G[117] = in[119] & in2[119];
    assign P[117] = in[119] ^ in2[119];
    assign G[118] = in[118] & in2[118];
    assign P[118] = in[118] ^ in2[118];
    assign G[119] = in[117] & in2[117];
    assign P[119] = in[117] ^ in2[117];
    assign G[120] = in[116] & in2[116];
    assign P[120] = in[116] ^ in2[116];
    assign G[121] = in[115] & in2[115];
    assign P[121] = in[115] ^ in2[115];
    assign G[122] = in[114] & in2[114];
    assign P[122] = in[114] ^ in2[114];
    assign G[123] = in[113] & in2[113];
    assign P[123] = in[113] ^ in2[113];
    assign G[124] = in[112] & in2[112];
    assign P[124] = in[112] ^ in2[112];
    assign G[125] = in[111] & in2[111];
    assign P[125] = in[111] ^ in2[111];
    assign G[126] = in[110] & in2[110];
    assign P[126] = in[110] ^ in2[110];
    assign G[127] = in[109] & in2[109];
    assign P[127] = in[109] ^ in2[109];
    assign G[128] = in[108] & in2[108];
    assign P[128] = in[108] ^ in2[108];
    assign G[129] = in[107] & in2[107];
    assign P[129] = in[107] ^ in2[107];
    assign G[130] = in[106] & in2[106];
    assign P[130] = in[106] ^ in2[106];
    assign G[131] = in[105] & in2[105];
    assign P[131] = in[105] ^ in2[105];
    assign G[132] = in[104] & in2[104];
    assign P[132] = in[104] ^ in2[104];
    assign G[133] = in[103] & in2[103];
    assign P[133] = in[103] ^ in2[103];
    assign G[134] = in[102] & in2[102];
    assign P[134] = in[102] ^ in2[102];
    assign G[135] = in[101] & in2[101];
    assign P[135] = in[101] ^ in2[101];
    assign G[136] = in[100] & in2[100];
    assign P[136] = in[100] ^ in2[100];
    assign G[137] = in[99] & in2[99];
    assign P[137] = in[99] ^ in2[99];
    assign G[138] = in[98] & in2[98];
    assign P[138] = in[98] ^ in2[98];
    assign G[139] = in[97] & in2[97];
    assign P[139] = in[97] ^ in2[97];
    assign G[140] = in[96] & in2[96];
    assign P[140] = in[96] ^ in2[96];
    assign G[141] = in[95] & in2[95];
    assign P[141] = in[95] ^ in2[95];
    assign G[142] = in[94] & in2[94];
    assign P[142] = in[94] ^ in2[94];
    assign G[143] = in[93] & in2[93];
    assign P[143] = in[93] ^ in2[93];
    assign G[144] = in[92] & in2[92];
    assign P[144] = in[92] ^ in2[92];
    assign G[145] = in[91] & in2[91];
    assign P[145] = in[91] ^ in2[91];
    assign G[146] = in[90] & in2[90];
    assign P[146] = in[90] ^ in2[90];
    assign G[147] = in[89] & in2[89];
    assign P[147] = in[89] ^ in2[89];
    assign G[148] = in[88] & in2[88];
    assign P[148] = in[88] ^ in2[88];
    assign G[149] = in[87] & in2[87];
    assign P[149] = in[87] ^ in2[87];
    assign G[150] = in[86] & in2[86];
    assign P[150] = in[86] ^ in2[86];
    assign G[151] = in[85] & in2[85];
    assign P[151] = in[85] ^ in2[85];
    assign G[152] = in[84] & in2[84];
    assign P[152] = in[84] ^ in2[84];
    assign G[153] = in[83] & in2[83];
    assign P[153] = in[83] ^ in2[83];
    assign G[154] = in[82] & in2[82];
    assign P[154] = in[82] ^ in2[82];
    assign G[155] = in[81] & in2[81];
    assign P[155] = in[81] ^ in2[81];
    assign G[156] = in[80] & in2[80];
    assign P[156] = in[80] ^ in2[80];
    assign G[157] = in[79] & in2[79];
    assign P[157] = in[79] ^ in2[79];
    assign G[158] = in[78] & in2[78];
    assign P[158] = in[78] ^ in2[78];
    assign G[159] = in[77] & in2[77];
    assign P[159] = in[77] ^ in2[77];
    assign G[160] = in[76] & in2[76];
    assign P[160] = in[76] ^ in2[76];
    assign G[161] = in[75] & in2[75];
    assign P[161] = in[75] ^ in2[75];
    assign G[162] = in[74] & in2[74];
    assign P[162] = in[74] ^ in2[74];
    assign G[163] = in[73] & in2[73];
    assign P[163] = in[73] ^ in2[73];
    assign G[164] = in[72] & in2[72];
    assign P[164] = in[72] ^ in2[72];
    assign G[165] = in[71] & in2[71];
    assign P[165] = in[71] ^ in2[71];
    assign G[166] = in[70] & in2[70];
    assign P[166] = in[70] ^ in2[70];
    assign G[167] = in[69] & in2[69];
    assign P[167] = in[69] ^ in2[69];
    assign G[168] = in[68] & in2[68];
    assign P[168] = in[68] ^ in2[68];
    assign G[169] = in[67] & in2[67];
    assign P[169] = in[67] ^ in2[67];
    assign G[170] = in[66] & in2[66];
    assign P[170] = in[66] ^ in2[66];
    assign G[171] = in[65] & in2[65];
    assign P[171] = in[65] ^ in2[65];
    assign G[172] = in[64] & in2[64];
    assign P[172] = in[64] ^ in2[64];
    assign G[173] = in[63] & in2[63];
    assign P[173] = in[63] ^ in2[63];
    assign G[174] = in[62] & in2[62];
    assign P[174] = in[62] ^ in2[62];
    assign G[175] = in[61] & in2[61];
    assign P[175] = in[61] ^ in2[61];
    assign G[176] = in[60] & in2[60];
    assign P[176] = in[60] ^ in2[60];
    assign G[177] = in[59] & in2[59];
    assign P[177] = in[59] ^ in2[59];
    assign G[178] = in[58] & in2[58];
    assign P[178] = in[58] ^ in2[58];
    assign G[179] = in[57] & in2[57];
    assign P[179] = in[57] ^ in2[57];
    assign G[180] = in[56] & in2[56];
    assign P[180] = in[56] ^ in2[56];
    assign G[181] = in[55] & in2[55];
    assign P[181] = in[55] ^ in2[55];
    assign G[182] = in[54] & in2[54];
    assign P[182] = in[54] ^ in2[54];
    assign G[183] = in[53] & in2[53];
    assign P[183] = in[53] ^ in2[53];
    assign G[184] = in[52] & in2[52];
    assign P[184] = in[52] ^ in2[52];
    assign G[185] = in[51] & in2[51];
    assign P[185] = in[51] ^ in2[51];
    assign G[186] = in[50] & in2[50];
    assign P[186] = in[50] ^ in2[50];
    assign G[187] = in[49] & in2[49];
    assign P[187] = in[49] ^ in2[49];
    assign G[188] = in[48] & in2[48];
    assign P[188] = in[48] ^ in2[48];
    assign G[189] = in[47] & in2[47];
    assign P[189] = in[47] ^ in2[47];
    assign G[190] = in[46] & in2[46];
    assign P[190] = in[46] ^ in2[46];
    assign G[191] = in[45] & in2[45];
    assign P[191] = in[45] ^ in2[45];
    assign G[192] = in[44] & in2[44];
    assign P[192] = in[44] ^ in2[44];
    assign G[193] = in[43] & in2[43];
    assign P[193] = in[43] ^ in2[43];
    assign G[194] = in[42] & in2[42];
    assign P[194] = in[42] ^ in2[42];
    assign G[195] = in[41] & in2[41];
    assign P[195] = in[41] ^ in2[41];
    assign G[196] = in[40] & in2[40];
    assign P[196] = in[40] ^ in2[40];
    assign G[197] = in[39] & in2[39];
    assign P[197] = in[39] ^ in2[39];
    assign G[198] = in[38] & in2[38];
    assign P[198] = in[38] ^ in2[38];
    assign G[199] = in[37] & in2[37];
    assign P[199] = in[37] ^ in2[37];
    assign G[200] = in[36] & in2[36];
    assign P[200] = in[36] ^ in2[36];
    assign G[201] = in[35] & in2[35];
    assign P[201] = in[35] ^ in2[35];
    assign G[202] = in[34] & in2[34];
    assign P[202] = in[34] ^ in2[34];
    assign G[203] = in[33] & in2[33];
    assign P[203] = in[33] ^ in2[33];
    assign G[204] = in[32] & in2[32];
    assign P[204] = in[32] ^ in2[32];
    assign G[205] = in[31] & in2[31];
    assign P[205] = in[31] ^ in2[31];
    assign G[206] = in[30] & in2[30];
    assign P[206] = in[30] ^ in2[30];
    assign G[207] = in[29] & in2[29];
    assign P[207] = in[29] ^ in2[29];
    assign G[208] = in[28] & in2[28];
    assign P[208] = in[28] ^ in2[28];
    assign G[209] = in[27] & in2[27];
    assign P[209] = in[27] ^ in2[27];
    assign G[210] = in[26] & in2[26];
    assign P[210] = in[26] ^ in2[26];
    assign G[211] = in[25] & in2[25];
    assign P[211] = in[25] ^ in2[25];
    assign G[212] = in[24] & in2[24];
    assign P[212] = in[24] ^ in2[24];
    assign G[213] = in[23] & in2[23];
    assign P[213] = in[23] ^ in2[23];
    assign G[214] = in[22] & in2[22];
    assign P[214] = in[22] ^ in2[22];
    assign G[215] = in[21] & in2[21];
    assign P[215] = in[21] ^ in2[21];
    assign G[216] = in[20] & in2[20];
    assign P[216] = in[20] ^ in2[20];
    assign G[217] = in[19] & in2[19];
    assign P[217] = in[19] ^ in2[19];
    assign G[218] = in[18] & in2[18];
    assign P[218] = in[18] ^ in2[18];
    assign G[219] = in[17] & in2[17];
    assign P[219] = in[17] ^ in2[17];
    assign G[220] = in[16] & in2[16];
    assign P[220] = in[16] ^ in2[16];
    assign G[221] = in[15] & in2[15];
    assign P[221] = in[15] ^ in2[15];
    assign G[222] = in[14] & in2[14];
    assign P[222] = in[14] ^ in2[14];
    assign G[223] = in[13] & in2[13];
    assign P[223] = in[13] ^ in2[13];
    assign G[224] = in[12] & in2[12];
    assign P[224] = in[12] ^ in2[12];
    assign G[225] = in[11] & in2[11];
    assign P[225] = in[11] ^ in2[11];
    assign G[226] = in[10] & in2[10];
    assign P[226] = in[10] ^ in2[10];
    assign G[227] = in[9] & in2[9];
    assign P[227] = in[9] ^ in2[9];
    assign G[228] = in[8] & in2[8];
    assign P[228] = in[8] ^ in2[8];
    assign G[229] = in[7] & in2[7];
    assign P[229] = in[7] ^ in2[7];
    assign G[230] = in[6] & in2[6];
    assign P[230] = in[6] ^ in2[6];
    assign G[231] = in[5] & in2[5];
    assign P[231] = in[5] ^ in2[5];
    assign G[232] = in[4] & in2[4];
    assign P[232] = in[4] ^ in2[4];
    assign G[233] = in[3] & in2[3];
    assign P[233] = in[3] ^ in2[3];
    assign G[234] = in[2] & in2[2];
    assign P[234] = in[2] ^ in2[2];
    assign G[235] = in[1] & in2[1];
    assign P[235] = in[1] ^ in2[1];
    assign G[236] = in[0] & in2[0];
    assign P[236] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign C[236] = G[235] | (P[235] & C[235]);
    assign cout = G[236] | (P[236] & C[236]);
    assign sum = P ^ C;
endmodule

module CLA236(output [235:0] sum, output cout, input [235:0] in1, input [235:0] in2;

    wire[235:0] G;
    wire[235:0] C;
    wire[235:0] P;

    assign G[0] = in[235] & in2[235];
    assign P[0] = in[235] ^ in2[235];
    assign G[1] = in[234] & in2[234];
    assign P[1] = in[234] ^ in2[234];
    assign G[2] = in[233] & in2[233];
    assign P[2] = in[233] ^ in2[233];
    assign G[3] = in[232] & in2[232];
    assign P[3] = in[232] ^ in2[232];
    assign G[4] = in[231] & in2[231];
    assign P[4] = in[231] ^ in2[231];
    assign G[5] = in[230] & in2[230];
    assign P[5] = in[230] ^ in2[230];
    assign G[6] = in[229] & in2[229];
    assign P[6] = in[229] ^ in2[229];
    assign G[7] = in[228] & in2[228];
    assign P[7] = in[228] ^ in2[228];
    assign G[8] = in[227] & in2[227];
    assign P[8] = in[227] ^ in2[227];
    assign G[9] = in[226] & in2[226];
    assign P[9] = in[226] ^ in2[226];
    assign G[10] = in[225] & in2[225];
    assign P[10] = in[225] ^ in2[225];
    assign G[11] = in[224] & in2[224];
    assign P[11] = in[224] ^ in2[224];
    assign G[12] = in[223] & in2[223];
    assign P[12] = in[223] ^ in2[223];
    assign G[13] = in[222] & in2[222];
    assign P[13] = in[222] ^ in2[222];
    assign G[14] = in[221] & in2[221];
    assign P[14] = in[221] ^ in2[221];
    assign G[15] = in[220] & in2[220];
    assign P[15] = in[220] ^ in2[220];
    assign G[16] = in[219] & in2[219];
    assign P[16] = in[219] ^ in2[219];
    assign G[17] = in[218] & in2[218];
    assign P[17] = in[218] ^ in2[218];
    assign G[18] = in[217] & in2[217];
    assign P[18] = in[217] ^ in2[217];
    assign G[19] = in[216] & in2[216];
    assign P[19] = in[216] ^ in2[216];
    assign G[20] = in[215] & in2[215];
    assign P[20] = in[215] ^ in2[215];
    assign G[21] = in[214] & in2[214];
    assign P[21] = in[214] ^ in2[214];
    assign G[22] = in[213] & in2[213];
    assign P[22] = in[213] ^ in2[213];
    assign G[23] = in[212] & in2[212];
    assign P[23] = in[212] ^ in2[212];
    assign G[24] = in[211] & in2[211];
    assign P[24] = in[211] ^ in2[211];
    assign G[25] = in[210] & in2[210];
    assign P[25] = in[210] ^ in2[210];
    assign G[26] = in[209] & in2[209];
    assign P[26] = in[209] ^ in2[209];
    assign G[27] = in[208] & in2[208];
    assign P[27] = in[208] ^ in2[208];
    assign G[28] = in[207] & in2[207];
    assign P[28] = in[207] ^ in2[207];
    assign G[29] = in[206] & in2[206];
    assign P[29] = in[206] ^ in2[206];
    assign G[30] = in[205] & in2[205];
    assign P[30] = in[205] ^ in2[205];
    assign G[31] = in[204] & in2[204];
    assign P[31] = in[204] ^ in2[204];
    assign G[32] = in[203] & in2[203];
    assign P[32] = in[203] ^ in2[203];
    assign G[33] = in[202] & in2[202];
    assign P[33] = in[202] ^ in2[202];
    assign G[34] = in[201] & in2[201];
    assign P[34] = in[201] ^ in2[201];
    assign G[35] = in[200] & in2[200];
    assign P[35] = in[200] ^ in2[200];
    assign G[36] = in[199] & in2[199];
    assign P[36] = in[199] ^ in2[199];
    assign G[37] = in[198] & in2[198];
    assign P[37] = in[198] ^ in2[198];
    assign G[38] = in[197] & in2[197];
    assign P[38] = in[197] ^ in2[197];
    assign G[39] = in[196] & in2[196];
    assign P[39] = in[196] ^ in2[196];
    assign G[40] = in[195] & in2[195];
    assign P[40] = in[195] ^ in2[195];
    assign G[41] = in[194] & in2[194];
    assign P[41] = in[194] ^ in2[194];
    assign G[42] = in[193] & in2[193];
    assign P[42] = in[193] ^ in2[193];
    assign G[43] = in[192] & in2[192];
    assign P[43] = in[192] ^ in2[192];
    assign G[44] = in[191] & in2[191];
    assign P[44] = in[191] ^ in2[191];
    assign G[45] = in[190] & in2[190];
    assign P[45] = in[190] ^ in2[190];
    assign G[46] = in[189] & in2[189];
    assign P[46] = in[189] ^ in2[189];
    assign G[47] = in[188] & in2[188];
    assign P[47] = in[188] ^ in2[188];
    assign G[48] = in[187] & in2[187];
    assign P[48] = in[187] ^ in2[187];
    assign G[49] = in[186] & in2[186];
    assign P[49] = in[186] ^ in2[186];
    assign G[50] = in[185] & in2[185];
    assign P[50] = in[185] ^ in2[185];
    assign G[51] = in[184] & in2[184];
    assign P[51] = in[184] ^ in2[184];
    assign G[52] = in[183] & in2[183];
    assign P[52] = in[183] ^ in2[183];
    assign G[53] = in[182] & in2[182];
    assign P[53] = in[182] ^ in2[182];
    assign G[54] = in[181] & in2[181];
    assign P[54] = in[181] ^ in2[181];
    assign G[55] = in[180] & in2[180];
    assign P[55] = in[180] ^ in2[180];
    assign G[56] = in[179] & in2[179];
    assign P[56] = in[179] ^ in2[179];
    assign G[57] = in[178] & in2[178];
    assign P[57] = in[178] ^ in2[178];
    assign G[58] = in[177] & in2[177];
    assign P[58] = in[177] ^ in2[177];
    assign G[59] = in[176] & in2[176];
    assign P[59] = in[176] ^ in2[176];
    assign G[60] = in[175] & in2[175];
    assign P[60] = in[175] ^ in2[175];
    assign G[61] = in[174] & in2[174];
    assign P[61] = in[174] ^ in2[174];
    assign G[62] = in[173] & in2[173];
    assign P[62] = in[173] ^ in2[173];
    assign G[63] = in[172] & in2[172];
    assign P[63] = in[172] ^ in2[172];
    assign G[64] = in[171] & in2[171];
    assign P[64] = in[171] ^ in2[171];
    assign G[65] = in[170] & in2[170];
    assign P[65] = in[170] ^ in2[170];
    assign G[66] = in[169] & in2[169];
    assign P[66] = in[169] ^ in2[169];
    assign G[67] = in[168] & in2[168];
    assign P[67] = in[168] ^ in2[168];
    assign G[68] = in[167] & in2[167];
    assign P[68] = in[167] ^ in2[167];
    assign G[69] = in[166] & in2[166];
    assign P[69] = in[166] ^ in2[166];
    assign G[70] = in[165] & in2[165];
    assign P[70] = in[165] ^ in2[165];
    assign G[71] = in[164] & in2[164];
    assign P[71] = in[164] ^ in2[164];
    assign G[72] = in[163] & in2[163];
    assign P[72] = in[163] ^ in2[163];
    assign G[73] = in[162] & in2[162];
    assign P[73] = in[162] ^ in2[162];
    assign G[74] = in[161] & in2[161];
    assign P[74] = in[161] ^ in2[161];
    assign G[75] = in[160] & in2[160];
    assign P[75] = in[160] ^ in2[160];
    assign G[76] = in[159] & in2[159];
    assign P[76] = in[159] ^ in2[159];
    assign G[77] = in[158] & in2[158];
    assign P[77] = in[158] ^ in2[158];
    assign G[78] = in[157] & in2[157];
    assign P[78] = in[157] ^ in2[157];
    assign G[79] = in[156] & in2[156];
    assign P[79] = in[156] ^ in2[156];
    assign G[80] = in[155] & in2[155];
    assign P[80] = in[155] ^ in2[155];
    assign G[81] = in[154] & in2[154];
    assign P[81] = in[154] ^ in2[154];
    assign G[82] = in[153] & in2[153];
    assign P[82] = in[153] ^ in2[153];
    assign G[83] = in[152] & in2[152];
    assign P[83] = in[152] ^ in2[152];
    assign G[84] = in[151] & in2[151];
    assign P[84] = in[151] ^ in2[151];
    assign G[85] = in[150] & in2[150];
    assign P[85] = in[150] ^ in2[150];
    assign G[86] = in[149] & in2[149];
    assign P[86] = in[149] ^ in2[149];
    assign G[87] = in[148] & in2[148];
    assign P[87] = in[148] ^ in2[148];
    assign G[88] = in[147] & in2[147];
    assign P[88] = in[147] ^ in2[147];
    assign G[89] = in[146] & in2[146];
    assign P[89] = in[146] ^ in2[146];
    assign G[90] = in[145] & in2[145];
    assign P[90] = in[145] ^ in2[145];
    assign G[91] = in[144] & in2[144];
    assign P[91] = in[144] ^ in2[144];
    assign G[92] = in[143] & in2[143];
    assign P[92] = in[143] ^ in2[143];
    assign G[93] = in[142] & in2[142];
    assign P[93] = in[142] ^ in2[142];
    assign G[94] = in[141] & in2[141];
    assign P[94] = in[141] ^ in2[141];
    assign G[95] = in[140] & in2[140];
    assign P[95] = in[140] ^ in2[140];
    assign G[96] = in[139] & in2[139];
    assign P[96] = in[139] ^ in2[139];
    assign G[97] = in[138] & in2[138];
    assign P[97] = in[138] ^ in2[138];
    assign G[98] = in[137] & in2[137];
    assign P[98] = in[137] ^ in2[137];
    assign G[99] = in[136] & in2[136];
    assign P[99] = in[136] ^ in2[136];
    assign G[100] = in[135] & in2[135];
    assign P[100] = in[135] ^ in2[135];
    assign G[101] = in[134] & in2[134];
    assign P[101] = in[134] ^ in2[134];
    assign G[102] = in[133] & in2[133];
    assign P[102] = in[133] ^ in2[133];
    assign G[103] = in[132] & in2[132];
    assign P[103] = in[132] ^ in2[132];
    assign G[104] = in[131] & in2[131];
    assign P[104] = in[131] ^ in2[131];
    assign G[105] = in[130] & in2[130];
    assign P[105] = in[130] ^ in2[130];
    assign G[106] = in[129] & in2[129];
    assign P[106] = in[129] ^ in2[129];
    assign G[107] = in[128] & in2[128];
    assign P[107] = in[128] ^ in2[128];
    assign G[108] = in[127] & in2[127];
    assign P[108] = in[127] ^ in2[127];
    assign G[109] = in[126] & in2[126];
    assign P[109] = in[126] ^ in2[126];
    assign G[110] = in[125] & in2[125];
    assign P[110] = in[125] ^ in2[125];
    assign G[111] = in[124] & in2[124];
    assign P[111] = in[124] ^ in2[124];
    assign G[112] = in[123] & in2[123];
    assign P[112] = in[123] ^ in2[123];
    assign G[113] = in[122] & in2[122];
    assign P[113] = in[122] ^ in2[122];
    assign G[114] = in[121] & in2[121];
    assign P[114] = in[121] ^ in2[121];
    assign G[115] = in[120] & in2[120];
    assign P[115] = in[120] ^ in2[120];
    assign G[116] = in[119] & in2[119];
    assign P[116] = in[119] ^ in2[119];
    assign G[117] = in[118] & in2[118];
    assign P[117] = in[118] ^ in2[118];
    assign G[118] = in[117] & in2[117];
    assign P[118] = in[117] ^ in2[117];
    assign G[119] = in[116] & in2[116];
    assign P[119] = in[116] ^ in2[116];
    assign G[120] = in[115] & in2[115];
    assign P[120] = in[115] ^ in2[115];
    assign G[121] = in[114] & in2[114];
    assign P[121] = in[114] ^ in2[114];
    assign G[122] = in[113] & in2[113];
    assign P[122] = in[113] ^ in2[113];
    assign G[123] = in[112] & in2[112];
    assign P[123] = in[112] ^ in2[112];
    assign G[124] = in[111] & in2[111];
    assign P[124] = in[111] ^ in2[111];
    assign G[125] = in[110] & in2[110];
    assign P[125] = in[110] ^ in2[110];
    assign G[126] = in[109] & in2[109];
    assign P[126] = in[109] ^ in2[109];
    assign G[127] = in[108] & in2[108];
    assign P[127] = in[108] ^ in2[108];
    assign G[128] = in[107] & in2[107];
    assign P[128] = in[107] ^ in2[107];
    assign G[129] = in[106] & in2[106];
    assign P[129] = in[106] ^ in2[106];
    assign G[130] = in[105] & in2[105];
    assign P[130] = in[105] ^ in2[105];
    assign G[131] = in[104] & in2[104];
    assign P[131] = in[104] ^ in2[104];
    assign G[132] = in[103] & in2[103];
    assign P[132] = in[103] ^ in2[103];
    assign G[133] = in[102] & in2[102];
    assign P[133] = in[102] ^ in2[102];
    assign G[134] = in[101] & in2[101];
    assign P[134] = in[101] ^ in2[101];
    assign G[135] = in[100] & in2[100];
    assign P[135] = in[100] ^ in2[100];
    assign G[136] = in[99] & in2[99];
    assign P[136] = in[99] ^ in2[99];
    assign G[137] = in[98] & in2[98];
    assign P[137] = in[98] ^ in2[98];
    assign G[138] = in[97] & in2[97];
    assign P[138] = in[97] ^ in2[97];
    assign G[139] = in[96] & in2[96];
    assign P[139] = in[96] ^ in2[96];
    assign G[140] = in[95] & in2[95];
    assign P[140] = in[95] ^ in2[95];
    assign G[141] = in[94] & in2[94];
    assign P[141] = in[94] ^ in2[94];
    assign G[142] = in[93] & in2[93];
    assign P[142] = in[93] ^ in2[93];
    assign G[143] = in[92] & in2[92];
    assign P[143] = in[92] ^ in2[92];
    assign G[144] = in[91] & in2[91];
    assign P[144] = in[91] ^ in2[91];
    assign G[145] = in[90] & in2[90];
    assign P[145] = in[90] ^ in2[90];
    assign G[146] = in[89] & in2[89];
    assign P[146] = in[89] ^ in2[89];
    assign G[147] = in[88] & in2[88];
    assign P[147] = in[88] ^ in2[88];
    assign G[148] = in[87] & in2[87];
    assign P[148] = in[87] ^ in2[87];
    assign G[149] = in[86] & in2[86];
    assign P[149] = in[86] ^ in2[86];
    assign G[150] = in[85] & in2[85];
    assign P[150] = in[85] ^ in2[85];
    assign G[151] = in[84] & in2[84];
    assign P[151] = in[84] ^ in2[84];
    assign G[152] = in[83] & in2[83];
    assign P[152] = in[83] ^ in2[83];
    assign G[153] = in[82] & in2[82];
    assign P[153] = in[82] ^ in2[82];
    assign G[154] = in[81] & in2[81];
    assign P[154] = in[81] ^ in2[81];
    assign G[155] = in[80] & in2[80];
    assign P[155] = in[80] ^ in2[80];
    assign G[156] = in[79] & in2[79];
    assign P[156] = in[79] ^ in2[79];
    assign G[157] = in[78] & in2[78];
    assign P[157] = in[78] ^ in2[78];
    assign G[158] = in[77] & in2[77];
    assign P[158] = in[77] ^ in2[77];
    assign G[159] = in[76] & in2[76];
    assign P[159] = in[76] ^ in2[76];
    assign G[160] = in[75] & in2[75];
    assign P[160] = in[75] ^ in2[75];
    assign G[161] = in[74] & in2[74];
    assign P[161] = in[74] ^ in2[74];
    assign G[162] = in[73] & in2[73];
    assign P[162] = in[73] ^ in2[73];
    assign G[163] = in[72] & in2[72];
    assign P[163] = in[72] ^ in2[72];
    assign G[164] = in[71] & in2[71];
    assign P[164] = in[71] ^ in2[71];
    assign G[165] = in[70] & in2[70];
    assign P[165] = in[70] ^ in2[70];
    assign G[166] = in[69] & in2[69];
    assign P[166] = in[69] ^ in2[69];
    assign G[167] = in[68] & in2[68];
    assign P[167] = in[68] ^ in2[68];
    assign G[168] = in[67] & in2[67];
    assign P[168] = in[67] ^ in2[67];
    assign G[169] = in[66] & in2[66];
    assign P[169] = in[66] ^ in2[66];
    assign G[170] = in[65] & in2[65];
    assign P[170] = in[65] ^ in2[65];
    assign G[171] = in[64] & in2[64];
    assign P[171] = in[64] ^ in2[64];
    assign G[172] = in[63] & in2[63];
    assign P[172] = in[63] ^ in2[63];
    assign G[173] = in[62] & in2[62];
    assign P[173] = in[62] ^ in2[62];
    assign G[174] = in[61] & in2[61];
    assign P[174] = in[61] ^ in2[61];
    assign G[175] = in[60] & in2[60];
    assign P[175] = in[60] ^ in2[60];
    assign G[176] = in[59] & in2[59];
    assign P[176] = in[59] ^ in2[59];
    assign G[177] = in[58] & in2[58];
    assign P[177] = in[58] ^ in2[58];
    assign G[178] = in[57] & in2[57];
    assign P[178] = in[57] ^ in2[57];
    assign G[179] = in[56] & in2[56];
    assign P[179] = in[56] ^ in2[56];
    assign G[180] = in[55] & in2[55];
    assign P[180] = in[55] ^ in2[55];
    assign G[181] = in[54] & in2[54];
    assign P[181] = in[54] ^ in2[54];
    assign G[182] = in[53] & in2[53];
    assign P[182] = in[53] ^ in2[53];
    assign G[183] = in[52] & in2[52];
    assign P[183] = in[52] ^ in2[52];
    assign G[184] = in[51] & in2[51];
    assign P[184] = in[51] ^ in2[51];
    assign G[185] = in[50] & in2[50];
    assign P[185] = in[50] ^ in2[50];
    assign G[186] = in[49] & in2[49];
    assign P[186] = in[49] ^ in2[49];
    assign G[187] = in[48] & in2[48];
    assign P[187] = in[48] ^ in2[48];
    assign G[188] = in[47] & in2[47];
    assign P[188] = in[47] ^ in2[47];
    assign G[189] = in[46] & in2[46];
    assign P[189] = in[46] ^ in2[46];
    assign G[190] = in[45] & in2[45];
    assign P[190] = in[45] ^ in2[45];
    assign G[191] = in[44] & in2[44];
    assign P[191] = in[44] ^ in2[44];
    assign G[192] = in[43] & in2[43];
    assign P[192] = in[43] ^ in2[43];
    assign G[193] = in[42] & in2[42];
    assign P[193] = in[42] ^ in2[42];
    assign G[194] = in[41] & in2[41];
    assign P[194] = in[41] ^ in2[41];
    assign G[195] = in[40] & in2[40];
    assign P[195] = in[40] ^ in2[40];
    assign G[196] = in[39] & in2[39];
    assign P[196] = in[39] ^ in2[39];
    assign G[197] = in[38] & in2[38];
    assign P[197] = in[38] ^ in2[38];
    assign G[198] = in[37] & in2[37];
    assign P[198] = in[37] ^ in2[37];
    assign G[199] = in[36] & in2[36];
    assign P[199] = in[36] ^ in2[36];
    assign G[200] = in[35] & in2[35];
    assign P[200] = in[35] ^ in2[35];
    assign G[201] = in[34] & in2[34];
    assign P[201] = in[34] ^ in2[34];
    assign G[202] = in[33] & in2[33];
    assign P[202] = in[33] ^ in2[33];
    assign G[203] = in[32] & in2[32];
    assign P[203] = in[32] ^ in2[32];
    assign G[204] = in[31] & in2[31];
    assign P[204] = in[31] ^ in2[31];
    assign G[205] = in[30] & in2[30];
    assign P[205] = in[30] ^ in2[30];
    assign G[206] = in[29] & in2[29];
    assign P[206] = in[29] ^ in2[29];
    assign G[207] = in[28] & in2[28];
    assign P[207] = in[28] ^ in2[28];
    assign G[208] = in[27] & in2[27];
    assign P[208] = in[27] ^ in2[27];
    assign G[209] = in[26] & in2[26];
    assign P[209] = in[26] ^ in2[26];
    assign G[210] = in[25] & in2[25];
    assign P[210] = in[25] ^ in2[25];
    assign G[211] = in[24] & in2[24];
    assign P[211] = in[24] ^ in2[24];
    assign G[212] = in[23] & in2[23];
    assign P[212] = in[23] ^ in2[23];
    assign G[213] = in[22] & in2[22];
    assign P[213] = in[22] ^ in2[22];
    assign G[214] = in[21] & in2[21];
    assign P[214] = in[21] ^ in2[21];
    assign G[215] = in[20] & in2[20];
    assign P[215] = in[20] ^ in2[20];
    assign G[216] = in[19] & in2[19];
    assign P[216] = in[19] ^ in2[19];
    assign G[217] = in[18] & in2[18];
    assign P[217] = in[18] ^ in2[18];
    assign G[218] = in[17] & in2[17];
    assign P[218] = in[17] ^ in2[17];
    assign G[219] = in[16] & in2[16];
    assign P[219] = in[16] ^ in2[16];
    assign G[220] = in[15] & in2[15];
    assign P[220] = in[15] ^ in2[15];
    assign G[221] = in[14] & in2[14];
    assign P[221] = in[14] ^ in2[14];
    assign G[222] = in[13] & in2[13];
    assign P[222] = in[13] ^ in2[13];
    assign G[223] = in[12] & in2[12];
    assign P[223] = in[12] ^ in2[12];
    assign G[224] = in[11] & in2[11];
    assign P[224] = in[11] ^ in2[11];
    assign G[225] = in[10] & in2[10];
    assign P[225] = in[10] ^ in2[10];
    assign G[226] = in[9] & in2[9];
    assign P[226] = in[9] ^ in2[9];
    assign G[227] = in[8] & in2[8];
    assign P[227] = in[8] ^ in2[8];
    assign G[228] = in[7] & in2[7];
    assign P[228] = in[7] ^ in2[7];
    assign G[229] = in[6] & in2[6];
    assign P[229] = in[6] ^ in2[6];
    assign G[230] = in[5] & in2[5];
    assign P[230] = in[5] ^ in2[5];
    assign G[231] = in[4] & in2[4];
    assign P[231] = in[4] ^ in2[4];
    assign G[232] = in[3] & in2[3];
    assign P[232] = in[3] ^ in2[3];
    assign G[233] = in[2] & in2[2];
    assign P[233] = in[2] ^ in2[2];
    assign G[234] = in[1] & in2[1];
    assign P[234] = in[1] ^ in2[1];
    assign G[235] = in[0] & in2[0];
    assign P[235] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign C[235] = G[234] | (P[234] & C[234]);
    assign cout = G[235] | (P[235] & C[235]);
    assign sum = P ^ C;
endmodule

module CLA235(output [234:0] sum, output cout, input [234:0] in1, input [234:0] in2;

    wire[234:0] G;
    wire[234:0] C;
    wire[234:0] P;

    assign G[0] = in[234] & in2[234];
    assign P[0] = in[234] ^ in2[234];
    assign G[1] = in[233] & in2[233];
    assign P[1] = in[233] ^ in2[233];
    assign G[2] = in[232] & in2[232];
    assign P[2] = in[232] ^ in2[232];
    assign G[3] = in[231] & in2[231];
    assign P[3] = in[231] ^ in2[231];
    assign G[4] = in[230] & in2[230];
    assign P[4] = in[230] ^ in2[230];
    assign G[5] = in[229] & in2[229];
    assign P[5] = in[229] ^ in2[229];
    assign G[6] = in[228] & in2[228];
    assign P[6] = in[228] ^ in2[228];
    assign G[7] = in[227] & in2[227];
    assign P[7] = in[227] ^ in2[227];
    assign G[8] = in[226] & in2[226];
    assign P[8] = in[226] ^ in2[226];
    assign G[9] = in[225] & in2[225];
    assign P[9] = in[225] ^ in2[225];
    assign G[10] = in[224] & in2[224];
    assign P[10] = in[224] ^ in2[224];
    assign G[11] = in[223] & in2[223];
    assign P[11] = in[223] ^ in2[223];
    assign G[12] = in[222] & in2[222];
    assign P[12] = in[222] ^ in2[222];
    assign G[13] = in[221] & in2[221];
    assign P[13] = in[221] ^ in2[221];
    assign G[14] = in[220] & in2[220];
    assign P[14] = in[220] ^ in2[220];
    assign G[15] = in[219] & in2[219];
    assign P[15] = in[219] ^ in2[219];
    assign G[16] = in[218] & in2[218];
    assign P[16] = in[218] ^ in2[218];
    assign G[17] = in[217] & in2[217];
    assign P[17] = in[217] ^ in2[217];
    assign G[18] = in[216] & in2[216];
    assign P[18] = in[216] ^ in2[216];
    assign G[19] = in[215] & in2[215];
    assign P[19] = in[215] ^ in2[215];
    assign G[20] = in[214] & in2[214];
    assign P[20] = in[214] ^ in2[214];
    assign G[21] = in[213] & in2[213];
    assign P[21] = in[213] ^ in2[213];
    assign G[22] = in[212] & in2[212];
    assign P[22] = in[212] ^ in2[212];
    assign G[23] = in[211] & in2[211];
    assign P[23] = in[211] ^ in2[211];
    assign G[24] = in[210] & in2[210];
    assign P[24] = in[210] ^ in2[210];
    assign G[25] = in[209] & in2[209];
    assign P[25] = in[209] ^ in2[209];
    assign G[26] = in[208] & in2[208];
    assign P[26] = in[208] ^ in2[208];
    assign G[27] = in[207] & in2[207];
    assign P[27] = in[207] ^ in2[207];
    assign G[28] = in[206] & in2[206];
    assign P[28] = in[206] ^ in2[206];
    assign G[29] = in[205] & in2[205];
    assign P[29] = in[205] ^ in2[205];
    assign G[30] = in[204] & in2[204];
    assign P[30] = in[204] ^ in2[204];
    assign G[31] = in[203] & in2[203];
    assign P[31] = in[203] ^ in2[203];
    assign G[32] = in[202] & in2[202];
    assign P[32] = in[202] ^ in2[202];
    assign G[33] = in[201] & in2[201];
    assign P[33] = in[201] ^ in2[201];
    assign G[34] = in[200] & in2[200];
    assign P[34] = in[200] ^ in2[200];
    assign G[35] = in[199] & in2[199];
    assign P[35] = in[199] ^ in2[199];
    assign G[36] = in[198] & in2[198];
    assign P[36] = in[198] ^ in2[198];
    assign G[37] = in[197] & in2[197];
    assign P[37] = in[197] ^ in2[197];
    assign G[38] = in[196] & in2[196];
    assign P[38] = in[196] ^ in2[196];
    assign G[39] = in[195] & in2[195];
    assign P[39] = in[195] ^ in2[195];
    assign G[40] = in[194] & in2[194];
    assign P[40] = in[194] ^ in2[194];
    assign G[41] = in[193] & in2[193];
    assign P[41] = in[193] ^ in2[193];
    assign G[42] = in[192] & in2[192];
    assign P[42] = in[192] ^ in2[192];
    assign G[43] = in[191] & in2[191];
    assign P[43] = in[191] ^ in2[191];
    assign G[44] = in[190] & in2[190];
    assign P[44] = in[190] ^ in2[190];
    assign G[45] = in[189] & in2[189];
    assign P[45] = in[189] ^ in2[189];
    assign G[46] = in[188] & in2[188];
    assign P[46] = in[188] ^ in2[188];
    assign G[47] = in[187] & in2[187];
    assign P[47] = in[187] ^ in2[187];
    assign G[48] = in[186] & in2[186];
    assign P[48] = in[186] ^ in2[186];
    assign G[49] = in[185] & in2[185];
    assign P[49] = in[185] ^ in2[185];
    assign G[50] = in[184] & in2[184];
    assign P[50] = in[184] ^ in2[184];
    assign G[51] = in[183] & in2[183];
    assign P[51] = in[183] ^ in2[183];
    assign G[52] = in[182] & in2[182];
    assign P[52] = in[182] ^ in2[182];
    assign G[53] = in[181] & in2[181];
    assign P[53] = in[181] ^ in2[181];
    assign G[54] = in[180] & in2[180];
    assign P[54] = in[180] ^ in2[180];
    assign G[55] = in[179] & in2[179];
    assign P[55] = in[179] ^ in2[179];
    assign G[56] = in[178] & in2[178];
    assign P[56] = in[178] ^ in2[178];
    assign G[57] = in[177] & in2[177];
    assign P[57] = in[177] ^ in2[177];
    assign G[58] = in[176] & in2[176];
    assign P[58] = in[176] ^ in2[176];
    assign G[59] = in[175] & in2[175];
    assign P[59] = in[175] ^ in2[175];
    assign G[60] = in[174] & in2[174];
    assign P[60] = in[174] ^ in2[174];
    assign G[61] = in[173] & in2[173];
    assign P[61] = in[173] ^ in2[173];
    assign G[62] = in[172] & in2[172];
    assign P[62] = in[172] ^ in2[172];
    assign G[63] = in[171] & in2[171];
    assign P[63] = in[171] ^ in2[171];
    assign G[64] = in[170] & in2[170];
    assign P[64] = in[170] ^ in2[170];
    assign G[65] = in[169] & in2[169];
    assign P[65] = in[169] ^ in2[169];
    assign G[66] = in[168] & in2[168];
    assign P[66] = in[168] ^ in2[168];
    assign G[67] = in[167] & in2[167];
    assign P[67] = in[167] ^ in2[167];
    assign G[68] = in[166] & in2[166];
    assign P[68] = in[166] ^ in2[166];
    assign G[69] = in[165] & in2[165];
    assign P[69] = in[165] ^ in2[165];
    assign G[70] = in[164] & in2[164];
    assign P[70] = in[164] ^ in2[164];
    assign G[71] = in[163] & in2[163];
    assign P[71] = in[163] ^ in2[163];
    assign G[72] = in[162] & in2[162];
    assign P[72] = in[162] ^ in2[162];
    assign G[73] = in[161] & in2[161];
    assign P[73] = in[161] ^ in2[161];
    assign G[74] = in[160] & in2[160];
    assign P[74] = in[160] ^ in2[160];
    assign G[75] = in[159] & in2[159];
    assign P[75] = in[159] ^ in2[159];
    assign G[76] = in[158] & in2[158];
    assign P[76] = in[158] ^ in2[158];
    assign G[77] = in[157] & in2[157];
    assign P[77] = in[157] ^ in2[157];
    assign G[78] = in[156] & in2[156];
    assign P[78] = in[156] ^ in2[156];
    assign G[79] = in[155] & in2[155];
    assign P[79] = in[155] ^ in2[155];
    assign G[80] = in[154] & in2[154];
    assign P[80] = in[154] ^ in2[154];
    assign G[81] = in[153] & in2[153];
    assign P[81] = in[153] ^ in2[153];
    assign G[82] = in[152] & in2[152];
    assign P[82] = in[152] ^ in2[152];
    assign G[83] = in[151] & in2[151];
    assign P[83] = in[151] ^ in2[151];
    assign G[84] = in[150] & in2[150];
    assign P[84] = in[150] ^ in2[150];
    assign G[85] = in[149] & in2[149];
    assign P[85] = in[149] ^ in2[149];
    assign G[86] = in[148] & in2[148];
    assign P[86] = in[148] ^ in2[148];
    assign G[87] = in[147] & in2[147];
    assign P[87] = in[147] ^ in2[147];
    assign G[88] = in[146] & in2[146];
    assign P[88] = in[146] ^ in2[146];
    assign G[89] = in[145] & in2[145];
    assign P[89] = in[145] ^ in2[145];
    assign G[90] = in[144] & in2[144];
    assign P[90] = in[144] ^ in2[144];
    assign G[91] = in[143] & in2[143];
    assign P[91] = in[143] ^ in2[143];
    assign G[92] = in[142] & in2[142];
    assign P[92] = in[142] ^ in2[142];
    assign G[93] = in[141] & in2[141];
    assign P[93] = in[141] ^ in2[141];
    assign G[94] = in[140] & in2[140];
    assign P[94] = in[140] ^ in2[140];
    assign G[95] = in[139] & in2[139];
    assign P[95] = in[139] ^ in2[139];
    assign G[96] = in[138] & in2[138];
    assign P[96] = in[138] ^ in2[138];
    assign G[97] = in[137] & in2[137];
    assign P[97] = in[137] ^ in2[137];
    assign G[98] = in[136] & in2[136];
    assign P[98] = in[136] ^ in2[136];
    assign G[99] = in[135] & in2[135];
    assign P[99] = in[135] ^ in2[135];
    assign G[100] = in[134] & in2[134];
    assign P[100] = in[134] ^ in2[134];
    assign G[101] = in[133] & in2[133];
    assign P[101] = in[133] ^ in2[133];
    assign G[102] = in[132] & in2[132];
    assign P[102] = in[132] ^ in2[132];
    assign G[103] = in[131] & in2[131];
    assign P[103] = in[131] ^ in2[131];
    assign G[104] = in[130] & in2[130];
    assign P[104] = in[130] ^ in2[130];
    assign G[105] = in[129] & in2[129];
    assign P[105] = in[129] ^ in2[129];
    assign G[106] = in[128] & in2[128];
    assign P[106] = in[128] ^ in2[128];
    assign G[107] = in[127] & in2[127];
    assign P[107] = in[127] ^ in2[127];
    assign G[108] = in[126] & in2[126];
    assign P[108] = in[126] ^ in2[126];
    assign G[109] = in[125] & in2[125];
    assign P[109] = in[125] ^ in2[125];
    assign G[110] = in[124] & in2[124];
    assign P[110] = in[124] ^ in2[124];
    assign G[111] = in[123] & in2[123];
    assign P[111] = in[123] ^ in2[123];
    assign G[112] = in[122] & in2[122];
    assign P[112] = in[122] ^ in2[122];
    assign G[113] = in[121] & in2[121];
    assign P[113] = in[121] ^ in2[121];
    assign G[114] = in[120] & in2[120];
    assign P[114] = in[120] ^ in2[120];
    assign G[115] = in[119] & in2[119];
    assign P[115] = in[119] ^ in2[119];
    assign G[116] = in[118] & in2[118];
    assign P[116] = in[118] ^ in2[118];
    assign G[117] = in[117] & in2[117];
    assign P[117] = in[117] ^ in2[117];
    assign G[118] = in[116] & in2[116];
    assign P[118] = in[116] ^ in2[116];
    assign G[119] = in[115] & in2[115];
    assign P[119] = in[115] ^ in2[115];
    assign G[120] = in[114] & in2[114];
    assign P[120] = in[114] ^ in2[114];
    assign G[121] = in[113] & in2[113];
    assign P[121] = in[113] ^ in2[113];
    assign G[122] = in[112] & in2[112];
    assign P[122] = in[112] ^ in2[112];
    assign G[123] = in[111] & in2[111];
    assign P[123] = in[111] ^ in2[111];
    assign G[124] = in[110] & in2[110];
    assign P[124] = in[110] ^ in2[110];
    assign G[125] = in[109] & in2[109];
    assign P[125] = in[109] ^ in2[109];
    assign G[126] = in[108] & in2[108];
    assign P[126] = in[108] ^ in2[108];
    assign G[127] = in[107] & in2[107];
    assign P[127] = in[107] ^ in2[107];
    assign G[128] = in[106] & in2[106];
    assign P[128] = in[106] ^ in2[106];
    assign G[129] = in[105] & in2[105];
    assign P[129] = in[105] ^ in2[105];
    assign G[130] = in[104] & in2[104];
    assign P[130] = in[104] ^ in2[104];
    assign G[131] = in[103] & in2[103];
    assign P[131] = in[103] ^ in2[103];
    assign G[132] = in[102] & in2[102];
    assign P[132] = in[102] ^ in2[102];
    assign G[133] = in[101] & in2[101];
    assign P[133] = in[101] ^ in2[101];
    assign G[134] = in[100] & in2[100];
    assign P[134] = in[100] ^ in2[100];
    assign G[135] = in[99] & in2[99];
    assign P[135] = in[99] ^ in2[99];
    assign G[136] = in[98] & in2[98];
    assign P[136] = in[98] ^ in2[98];
    assign G[137] = in[97] & in2[97];
    assign P[137] = in[97] ^ in2[97];
    assign G[138] = in[96] & in2[96];
    assign P[138] = in[96] ^ in2[96];
    assign G[139] = in[95] & in2[95];
    assign P[139] = in[95] ^ in2[95];
    assign G[140] = in[94] & in2[94];
    assign P[140] = in[94] ^ in2[94];
    assign G[141] = in[93] & in2[93];
    assign P[141] = in[93] ^ in2[93];
    assign G[142] = in[92] & in2[92];
    assign P[142] = in[92] ^ in2[92];
    assign G[143] = in[91] & in2[91];
    assign P[143] = in[91] ^ in2[91];
    assign G[144] = in[90] & in2[90];
    assign P[144] = in[90] ^ in2[90];
    assign G[145] = in[89] & in2[89];
    assign P[145] = in[89] ^ in2[89];
    assign G[146] = in[88] & in2[88];
    assign P[146] = in[88] ^ in2[88];
    assign G[147] = in[87] & in2[87];
    assign P[147] = in[87] ^ in2[87];
    assign G[148] = in[86] & in2[86];
    assign P[148] = in[86] ^ in2[86];
    assign G[149] = in[85] & in2[85];
    assign P[149] = in[85] ^ in2[85];
    assign G[150] = in[84] & in2[84];
    assign P[150] = in[84] ^ in2[84];
    assign G[151] = in[83] & in2[83];
    assign P[151] = in[83] ^ in2[83];
    assign G[152] = in[82] & in2[82];
    assign P[152] = in[82] ^ in2[82];
    assign G[153] = in[81] & in2[81];
    assign P[153] = in[81] ^ in2[81];
    assign G[154] = in[80] & in2[80];
    assign P[154] = in[80] ^ in2[80];
    assign G[155] = in[79] & in2[79];
    assign P[155] = in[79] ^ in2[79];
    assign G[156] = in[78] & in2[78];
    assign P[156] = in[78] ^ in2[78];
    assign G[157] = in[77] & in2[77];
    assign P[157] = in[77] ^ in2[77];
    assign G[158] = in[76] & in2[76];
    assign P[158] = in[76] ^ in2[76];
    assign G[159] = in[75] & in2[75];
    assign P[159] = in[75] ^ in2[75];
    assign G[160] = in[74] & in2[74];
    assign P[160] = in[74] ^ in2[74];
    assign G[161] = in[73] & in2[73];
    assign P[161] = in[73] ^ in2[73];
    assign G[162] = in[72] & in2[72];
    assign P[162] = in[72] ^ in2[72];
    assign G[163] = in[71] & in2[71];
    assign P[163] = in[71] ^ in2[71];
    assign G[164] = in[70] & in2[70];
    assign P[164] = in[70] ^ in2[70];
    assign G[165] = in[69] & in2[69];
    assign P[165] = in[69] ^ in2[69];
    assign G[166] = in[68] & in2[68];
    assign P[166] = in[68] ^ in2[68];
    assign G[167] = in[67] & in2[67];
    assign P[167] = in[67] ^ in2[67];
    assign G[168] = in[66] & in2[66];
    assign P[168] = in[66] ^ in2[66];
    assign G[169] = in[65] & in2[65];
    assign P[169] = in[65] ^ in2[65];
    assign G[170] = in[64] & in2[64];
    assign P[170] = in[64] ^ in2[64];
    assign G[171] = in[63] & in2[63];
    assign P[171] = in[63] ^ in2[63];
    assign G[172] = in[62] & in2[62];
    assign P[172] = in[62] ^ in2[62];
    assign G[173] = in[61] & in2[61];
    assign P[173] = in[61] ^ in2[61];
    assign G[174] = in[60] & in2[60];
    assign P[174] = in[60] ^ in2[60];
    assign G[175] = in[59] & in2[59];
    assign P[175] = in[59] ^ in2[59];
    assign G[176] = in[58] & in2[58];
    assign P[176] = in[58] ^ in2[58];
    assign G[177] = in[57] & in2[57];
    assign P[177] = in[57] ^ in2[57];
    assign G[178] = in[56] & in2[56];
    assign P[178] = in[56] ^ in2[56];
    assign G[179] = in[55] & in2[55];
    assign P[179] = in[55] ^ in2[55];
    assign G[180] = in[54] & in2[54];
    assign P[180] = in[54] ^ in2[54];
    assign G[181] = in[53] & in2[53];
    assign P[181] = in[53] ^ in2[53];
    assign G[182] = in[52] & in2[52];
    assign P[182] = in[52] ^ in2[52];
    assign G[183] = in[51] & in2[51];
    assign P[183] = in[51] ^ in2[51];
    assign G[184] = in[50] & in2[50];
    assign P[184] = in[50] ^ in2[50];
    assign G[185] = in[49] & in2[49];
    assign P[185] = in[49] ^ in2[49];
    assign G[186] = in[48] & in2[48];
    assign P[186] = in[48] ^ in2[48];
    assign G[187] = in[47] & in2[47];
    assign P[187] = in[47] ^ in2[47];
    assign G[188] = in[46] & in2[46];
    assign P[188] = in[46] ^ in2[46];
    assign G[189] = in[45] & in2[45];
    assign P[189] = in[45] ^ in2[45];
    assign G[190] = in[44] & in2[44];
    assign P[190] = in[44] ^ in2[44];
    assign G[191] = in[43] & in2[43];
    assign P[191] = in[43] ^ in2[43];
    assign G[192] = in[42] & in2[42];
    assign P[192] = in[42] ^ in2[42];
    assign G[193] = in[41] & in2[41];
    assign P[193] = in[41] ^ in2[41];
    assign G[194] = in[40] & in2[40];
    assign P[194] = in[40] ^ in2[40];
    assign G[195] = in[39] & in2[39];
    assign P[195] = in[39] ^ in2[39];
    assign G[196] = in[38] & in2[38];
    assign P[196] = in[38] ^ in2[38];
    assign G[197] = in[37] & in2[37];
    assign P[197] = in[37] ^ in2[37];
    assign G[198] = in[36] & in2[36];
    assign P[198] = in[36] ^ in2[36];
    assign G[199] = in[35] & in2[35];
    assign P[199] = in[35] ^ in2[35];
    assign G[200] = in[34] & in2[34];
    assign P[200] = in[34] ^ in2[34];
    assign G[201] = in[33] & in2[33];
    assign P[201] = in[33] ^ in2[33];
    assign G[202] = in[32] & in2[32];
    assign P[202] = in[32] ^ in2[32];
    assign G[203] = in[31] & in2[31];
    assign P[203] = in[31] ^ in2[31];
    assign G[204] = in[30] & in2[30];
    assign P[204] = in[30] ^ in2[30];
    assign G[205] = in[29] & in2[29];
    assign P[205] = in[29] ^ in2[29];
    assign G[206] = in[28] & in2[28];
    assign P[206] = in[28] ^ in2[28];
    assign G[207] = in[27] & in2[27];
    assign P[207] = in[27] ^ in2[27];
    assign G[208] = in[26] & in2[26];
    assign P[208] = in[26] ^ in2[26];
    assign G[209] = in[25] & in2[25];
    assign P[209] = in[25] ^ in2[25];
    assign G[210] = in[24] & in2[24];
    assign P[210] = in[24] ^ in2[24];
    assign G[211] = in[23] & in2[23];
    assign P[211] = in[23] ^ in2[23];
    assign G[212] = in[22] & in2[22];
    assign P[212] = in[22] ^ in2[22];
    assign G[213] = in[21] & in2[21];
    assign P[213] = in[21] ^ in2[21];
    assign G[214] = in[20] & in2[20];
    assign P[214] = in[20] ^ in2[20];
    assign G[215] = in[19] & in2[19];
    assign P[215] = in[19] ^ in2[19];
    assign G[216] = in[18] & in2[18];
    assign P[216] = in[18] ^ in2[18];
    assign G[217] = in[17] & in2[17];
    assign P[217] = in[17] ^ in2[17];
    assign G[218] = in[16] & in2[16];
    assign P[218] = in[16] ^ in2[16];
    assign G[219] = in[15] & in2[15];
    assign P[219] = in[15] ^ in2[15];
    assign G[220] = in[14] & in2[14];
    assign P[220] = in[14] ^ in2[14];
    assign G[221] = in[13] & in2[13];
    assign P[221] = in[13] ^ in2[13];
    assign G[222] = in[12] & in2[12];
    assign P[222] = in[12] ^ in2[12];
    assign G[223] = in[11] & in2[11];
    assign P[223] = in[11] ^ in2[11];
    assign G[224] = in[10] & in2[10];
    assign P[224] = in[10] ^ in2[10];
    assign G[225] = in[9] & in2[9];
    assign P[225] = in[9] ^ in2[9];
    assign G[226] = in[8] & in2[8];
    assign P[226] = in[8] ^ in2[8];
    assign G[227] = in[7] & in2[7];
    assign P[227] = in[7] ^ in2[7];
    assign G[228] = in[6] & in2[6];
    assign P[228] = in[6] ^ in2[6];
    assign G[229] = in[5] & in2[5];
    assign P[229] = in[5] ^ in2[5];
    assign G[230] = in[4] & in2[4];
    assign P[230] = in[4] ^ in2[4];
    assign G[231] = in[3] & in2[3];
    assign P[231] = in[3] ^ in2[3];
    assign G[232] = in[2] & in2[2];
    assign P[232] = in[2] ^ in2[2];
    assign G[233] = in[1] & in2[1];
    assign P[233] = in[1] ^ in2[1];
    assign G[234] = in[0] & in2[0];
    assign P[234] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign C[234] = G[233] | (P[233] & C[233]);
    assign cout = G[234] | (P[234] & C[234]);
    assign sum = P ^ C;
endmodule

module CLA234(output [233:0] sum, output cout, input [233:0] in1, input [233:0] in2;

    wire[233:0] G;
    wire[233:0] C;
    wire[233:0] P;

    assign G[0] = in[233] & in2[233];
    assign P[0] = in[233] ^ in2[233];
    assign G[1] = in[232] & in2[232];
    assign P[1] = in[232] ^ in2[232];
    assign G[2] = in[231] & in2[231];
    assign P[2] = in[231] ^ in2[231];
    assign G[3] = in[230] & in2[230];
    assign P[3] = in[230] ^ in2[230];
    assign G[4] = in[229] & in2[229];
    assign P[4] = in[229] ^ in2[229];
    assign G[5] = in[228] & in2[228];
    assign P[5] = in[228] ^ in2[228];
    assign G[6] = in[227] & in2[227];
    assign P[6] = in[227] ^ in2[227];
    assign G[7] = in[226] & in2[226];
    assign P[7] = in[226] ^ in2[226];
    assign G[8] = in[225] & in2[225];
    assign P[8] = in[225] ^ in2[225];
    assign G[9] = in[224] & in2[224];
    assign P[9] = in[224] ^ in2[224];
    assign G[10] = in[223] & in2[223];
    assign P[10] = in[223] ^ in2[223];
    assign G[11] = in[222] & in2[222];
    assign P[11] = in[222] ^ in2[222];
    assign G[12] = in[221] & in2[221];
    assign P[12] = in[221] ^ in2[221];
    assign G[13] = in[220] & in2[220];
    assign P[13] = in[220] ^ in2[220];
    assign G[14] = in[219] & in2[219];
    assign P[14] = in[219] ^ in2[219];
    assign G[15] = in[218] & in2[218];
    assign P[15] = in[218] ^ in2[218];
    assign G[16] = in[217] & in2[217];
    assign P[16] = in[217] ^ in2[217];
    assign G[17] = in[216] & in2[216];
    assign P[17] = in[216] ^ in2[216];
    assign G[18] = in[215] & in2[215];
    assign P[18] = in[215] ^ in2[215];
    assign G[19] = in[214] & in2[214];
    assign P[19] = in[214] ^ in2[214];
    assign G[20] = in[213] & in2[213];
    assign P[20] = in[213] ^ in2[213];
    assign G[21] = in[212] & in2[212];
    assign P[21] = in[212] ^ in2[212];
    assign G[22] = in[211] & in2[211];
    assign P[22] = in[211] ^ in2[211];
    assign G[23] = in[210] & in2[210];
    assign P[23] = in[210] ^ in2[210];
    assign G[24] = in[209] & in2[209];
    assign P[24] = in[209] ^ in2[209];
    assign G[25] = in[208] & in2[208];
    assign P[25] = in[208] ^ in2[208];
    assign G[26] = in[207] & in2[207];
    assign P[26] = in[207] ^ in2[207];
    assign G[27] = in[206] & in2[206];
    assign P[27] = in[206] ^ in2[206];
    assign G[28] = in[205] & in2[205];
    assign P[28] = in[205] ^ in2[205];
    assign G[29] = in[204] & in2[204];
    assign P[29] = in[204] ^ in2[204];
    assign G[30] = in[203] & in2[203];
    assign P[30] = in[203] ^ in2[203];
    assign G[31] = in[202] & in2[202];
    assign P[31] = in[202] ^ in2[202];
    assign G[32] = in[201] & in2[201];
    assign P[32] = in[201] ^ in2[201];
    assign G[33] = in[200] & in2[200];
    assign P[33] = in[200] ^ in2[200];
    assign G[34] = in[199] & in2[199];
    assign P[34] = in[199] ^ in2[199];
    assign G[35] = in[198] & in2[198];
    assign P[35] = in[198] ^ in2[198];
    assign G[36] = in[197] & in2[197];
    assign P[36] = in[197] ^ in2[197];
    assign G[37] = in[196] & in2[196];
    assign P[37] = in[196] ^ in2[196];
    assign G[38] = in[195] & in2[195];
    assign P[38] = in[195] ^ in2[195];
    assign G[39] = in[194] & in2[194];
    assign P[39] = in[194] ^ in2[194];
    assign G[40] = in[193] & in2[193];
    assign P[40] = in[193] ^ in2[193];
    assign G[41] = in[192] & in2[192];
    assign P[41] = in[192] ^ in2[192];
    assign G[42] = in[191] & in2[191];
    assign P[42] = in[191] ^ in2[191];
    assign G[43] = in[190] & in2[190];
    assign P[43] = in[190] ^ in2[190];
    assign G[44] = in[189] & in2[189];
    assign P[44] = in[189] ^ in2[189];
    assign G[45] = in[188] & in2[188];
    assign P[45] = in[188] ^ in2[188];
    assign G[46] = in[187] & in2[187];
    assign P[46] = in[187] ^ in2[187];
    assign G[47] = in[186] & in2[186];
    assign P[47] = in[186] ^ in2[186];
    assign G[48] = in[185] & in2[185];
    assign P[48] = in[185] ^ in2[185];
    assign G[49] = in[184] & in2[184];
    assign P[49] = in[184] ^ in2[184];
    assign G[50] = in[183] & in2[183];
    assign P[50] = in[183] ^ in2[183];
    assign G[51] = in[182] & in2[182];
    assign P[51] = in[182] ^ in2[182];
    assign G[52] = in[181] & in2[181];
    assign P[52] = in[181] ^ in2[181];
    assign G[53] = in[180] & in2[180];
    assign P[53] = in[180] ^ in2[180];
    assign G[54] = in[179] & in2[179];
    assign P[54] = in[179] ^ in2[179];
    assign G[55] = in[178] & in2[178];
    assign P[55] = in[178] ^ in2[178];
    assign G[56] = in[177] & in2[177];
    assign P[56] = in[177] ^ in2[177];
    assign G[57] = in[176] & in2[176];
    assign P[57] = in[176] ^ in2[176];
    assign G[58] = in[175] & in2[175];
    assign P[58] = in[175] ^ in2[175];
    assign G[59] = in[174] & in2[174];
    assign P[59] = in[174] ^ in2[174];
    assign G[60] = in[173] & in2[173];
    assign P[60] = in[173] ^ in2[173];
    assign G[61] = in[172] & in2[172];
    assign P[61] = in[172] ^ in2[172];
    assign G[62] = in[171] & in2[171];
    assign P[62] = in[171] ^ in2[171];
    assign G[63] = in[170] & in2[170];
    assign P[63] = in[170] ^ in2[170];
    assign G[64] = in[169] & in2[169];
    assign P[64] = in[169] ^ in2[169];
    assign G[65] = in[168] & in2[168];
    assign P[65] = in[168] ^ in2[168];
    assign G[66] = in[167] & in2[167];
    assign P[66] = in[167] ^ in2[167];
    assign G[67] = in[166] & in2[166];
    assign P[67] = in[166] ^ in2[166];
    assign G[68] = in[165] & in2[165];
    assign P[68] = in[165] ^ in2[165];
    assign G[69] = in[164] & in2[164];
    assign P[69] = in[164] ^ in2[164];
    assign G[70] = in[163] & in2[163];
    assign P[70] = in[163] ^ in2[163];
    assign G[71] = in[162] & in2[162];
    assign P[71] = in[162] ^ in2[162];
    assign G[72] = in[161] & in2[161];
    assign P[72] = in[161] ^ in2[161];
    assign G[73] = in[160] & in2[160];
    assign P[73] = in[160] ^ in2[160];
    assign G[74] = in[159] & in2[159];
    assign P[74] = in[159] ^ in2[159];
    assign G[75] = in[158] & in2[158];
    assign P[75] = in[158] ^ in2[158];
    assign G[76] = in[157] & in2[157];
    assign P[76] = in[157] ^ in2[157];
    assign G[77] = in[156] & in2[156];
    assign P[77] = in[156] ^ in2[156];
    assign G[78] = in[155] & in2[155];
    assign P[78] = in[155] ^ in2[155];
    assign G[79] = in[154] & in2[154];
    assign P[79] = in[154] ^ in2[154];
    assign G[80] = in[153] & in2[153];
    assign P[80] = in[153] ^ in2[153];
    assign G[81] = in[152] & in2[152];
    assign P[81] = in[152] ^ in2[152];
    assign G[82] = in[151] & in2[151];
    assign P[82] = in[151] ^ in2[151];
    assign G[83] = in[150] & in2[150];
    assign P[83] = in[150] ^ in2[150];
    assign G[84] = in[149] & in2[149];
    assign P[84] = in[149] ^ in2[149];
    assign G[85] = in[148] & in2[148];
    assign P[85] = in[148] ^ in2[148];
    assign G[86] = in[147] & in2[147];
    assign P[86] = in[147] ^ in2[147];
    assign G[87] = in[146] & in2[146];
    assign P[87] = in[146] ^ in2[146];
    assign G[88] = in[145] & in2[145];
    assign P[88] = in[145] ^ in2[145];
    assign G[89] = in[144] & in2[144];
    assign P[89] = in[144] ^ in2[144];
    assign G[90] = in[143] & in2[143];
    assign P[90] = in[143] ^ in2[143];
    assign G[91] = in[142] & in2[142];
    assign P[91] = in[142] ^ in2[142];
    assign G[92] = in[141] & in2[141];
    assign P[92] = in[141] ^ in2[141];
    assign G[93] = in[140] & in2[140];
    assign P[93] = in[140] ^ in2[140];
    assign G[94] = in[139] & in2[139];
    assign P[94] = in[139] ^ in2[139];
    assign G[95] = in[138] & in2[138];
    assign P[95] = in[138] ^ in2[138];
    assign G[96] = in[137] & in2[137];
    assign P[96] = in[137] ^ in2[137];
    assign G[97] = in[136] & in2[136];
    assign P[97] = in[136] ^ in2[136];
    assign G[98] = in[135] & in2[135];
    assign P[98] = in[135] ^ in2[135];
    assign G[99] = in[134] & in2[134];
    assign P[99] = in[134] ^ in2[134];
    assign G[100] = in[133] & in2[133];
    assign P[100] = in[133] ^ in2[133];
    assign G[101] = in[132] & in2[132];
    assign P[101] = in[132] ^ in2[132];
    assign G[102] = in[131] & in2[131];
    assign P[102] = in[131] ^ in2[131];
    assign G[103] = in[130] & in2[130];
    assign P[103] = in[130] ^ in2[130];
    assign G[104] = in[129] & in2[129];
    assign P[104] = in[129] ^ in2[129];
    assign G[105] = in[128] & in2[128];
    assign P[105] = in[128] ^ in2[128];
    assign G[106] = in[127] & in2[127];
    assign P[106] = in[127] ^ in2[127];
    assign G[107] = in[126] & in2[126];
    assign P[107] = in[126] ^ in2[126];
    assign G[108] = in[125] & in2[125];
    assign P[108] = in[125] ^ in2[125];
    assign G[109] = in[124] & in2[124];
    assign P[109] = in[124] ^ in2[124];
    assign G[110] = in[123] & in2[123];
    assign P[110] = in[123] ^ in2[123];
    assign G[111] = in[122] & in2[122];
    assign P[111] = in[122] ^ in2[122];
    assign G[112] = in[121] & in2[121];
    assign P[112] = in[121] ^ in2[121];
    assign G[113] = in[120] & in2[120];
    assign P[113] = in[120] ^ in2[120];
    assign G[114] = in[119] & in2[119];
    assign P[114] = in[119] ^ in2[119];
    assign G[115] = in[118] & in2[118];
    assign P[115] = in[118] ^ in2[118];
    assign G[116] = in[117] & in2[117];
    assign P[116] = in[117] ^ in2[117];
    assign G[117] = in[116] & in2[116];
    assign P[117] = in[116] ^ in2[116];
    assign G[118] = in[115] & in2[115];
    assign P[118] = in[115] ^ in2[115];
    assign G[119] = in[114] & in2[114];
    assign P[119] = in[114] ^ in2[114];
    assign G[120] = in[113] & in2[113];
    assign P[120] = in[113] ^ in2[113];
    assign G[121] = in[112] & in2[112];
    assign P[121] = in[112] ^ in2[112];
    assign G[122] = in[111] & in2[111];
    assign P[122] = in[111] ^ in2[111];
    assign G[123] = in[110] & in2[110];
    assign P[123] = in[110] ^ in2[110];
    assign G[124] = in[109] & in2[109];
    assign P[124] = in[109] ^ in2[109];
    assign G[125] = in[108] & in2[108];
    assign P[125] = in[108] ^ in2[108];
    assign G[126] = in[107] & in2[107];
    assign P[126] = in[107] ^ in2[107];
    assign G[127] = in[106] & in2[106];
    assign P[127] = in[106] ^ in2[106];
    assign G[128] = in[105] & in2[105];
    assign P[128] = in[105] ^ in2[105];
    assign G[129] = in[104] & in2[104];
    assign P[129] = in[104] ^ in2[104];
    assign G[130] = in[103] & in2[103];
    assign P[130] = in[103] ^ in2[103];
    assign G[131] = in[102] & in2[102];
    assign P[131] = in[102] ^ in2[102];
    assign G[132] = in[101] & in2[101];
    assign P[132] = in[101] ^ in2[101];
    assign G[133] = in[100] & in2[100];
    assign P[133] = in[100] ^ in2[100];
    assign G[134] = in[99] & in2[99];
    assign P[134] = in[99] ^ in2[99];
    assign G[135] = in[98] & in2[98];
    assign P[135] = in[98] ^ in2[98];
    assign G[136] = in[97] & in2[97];
    assign P[136] = in[97] ^ in2[97];
    assign G[137] = in[96] & in2[96];
    assign P[137] = in[96] ^ in2[96];
    assign G[138] = in[95] & in2[95];
    assign P[138] = in[95] ^ in2[95];
    assign G[139] = in[94] & in2[94];
    assign P[139] = in[94] ^ in2[94];
    assign G[140] = in[93] & in2[93];
    assign P[140] = in[93] ^ in2[93];
    assign G[141] = in[92] & in2[92];
    assign P[141] = in[92] ^ in2[92];
    assign G[142] = in[91] & in2[91];
    assign P[142] = in[91] ^ in2[91];
    assign G[143] = in[90] & in2[90];
    assign P[143] = in[90] ^ in2[90];
    assign G[144] = in[89] & in2[89];
    assign P[144] = in[89] ^ in2[89];
    assign G[145] = in[88] & in2[88];
    assign P[145] = in[88] ^ in2[88];
    assign G[146] = in[87] & in2[87];
    assign P[146] = in[87] ^ in2[87];
    assign G[147] = in[86] & in2[86];
    assign P[147] = in[86] ^ in2[86];
    assign G[148] = in[85] & in2[85];
    assign P[148] = in[85] ^ in2[85];
    assign G[149] = in[84] & in2[84];
    assign P[149] = in[84] ^ in2[84];
    assign G[150] = in[83] & in2[83];
    assign P[150] = in[83] ^ in2[83];
    assign G[151] = in[82] & in2[82];
    assign P[151] = in[82] ^ in2[82];
    assign G[152] = in[81] & in2[81];
    assign P[152] = in[81] ^ in2[81];
    assign G[153] = in[80] & in2[80];
    assign P[153] = in[80] ^ in2[80];
    assign G[154] = in[79] & in2[79];
    assign P[154] = in[79] ^ in2[79];
    assign G[155] = in[78] & in2[78];
    assign P[155] = in[78] ^ in2[78];
    assign G[156] = in[77] & in2[77];
    assign P[156] = in[77] ^ in2[77];
    assign G[157] = in[76] & in2[76];
    assign P[157] = in[76] ^ in2[76];
    assign G[158] = in[75] & in2[75];
    assign P[158] = in[75] ^ in2[75];
    assign G[159] = in[74] & in2[74];
    assign P[159] = in[74] ^ in2[74];
    assign G[160] = in[73] & in2[73];
    assign P[160] = in[73] ^ in2[73];
    assign G[161] = in[72] & in2[72];
    assign P[161] = in[72] ^ in2[72];
    assign G[162] = in[71] & in2[71];
    assign P[162] = in[71] ^ in2[71];
    assign G[163] = in[70] & in2[70];
    assign P[163] = in[70] ^ in2[70];
    assign G[164] = in[69] & in2[69];
    assign P[164] = in[69] ^ in2[69];
    assign G[165] = in[68] & in2[68];
    assign P[165] = in[68] ^ in2[68];
    assign G[166] = in[67] & in2[67];
    assign P[166] = in[67] ^ in2[67];
    assign G[167] = in[66] & in2[66];
    assign P[167] = in[66] ^ in2[66];
    assign G[168] = in[65] & in2[65];
    assign P[168] = in[65] ^ in2[65];
    assign G[169] = in[64] & in2[64];
    assign P[169] = in[64] ^ in2[64];
    assign G[170] = in[63] & in2[63];
    assign P[170] = in[63] ^ in2[63];
    assign G[171] = in[62] & in2[62];
    assign P[171] = in[62] ^ in2[62];
    assign G[172] = in[61] & in2[61];
    assign P[172] = in[61] ^ in2[61];
    assign G[173] = in[60] & in2[60];
    assign P[173] = in[60] ^ in2[60];
    assign G[174] = in[59] & in2[59];
    assign P[174] = in[59] ^ in2[59];
    assign G[175] = in[58] & in2[58];
    assign P[175] = in[58] ^ in2[58];
    assign G[176] = in[57] & in2[57];
    assign P[176] = in[57] ^ in2[57];
    assign G[177] = in[56] & in2[56];
    assign P[177] = in[56] ^ in2[56];
    assign G[178] = in[55] & in2[55];
    assign P[178] = in[55] ^ in2[55];
    assign G[179] = in[54] & in2[54];
    assign P[179] = in[54] ^ in2[54];
    assign G[180] = in[53] & in2[53];
    assign P[180] = in[53] ^ in2[53];
    assign G[181] = in[52] & in2[52];
    assign P[181] = in[52] ^ in2[52];
    assign G[182] = in[51] & in2[51];
    assign P[182] = in[51] ^ in2[51];
    assign G[183] = in[50] & in2[50];
    assign P[183] = in[50] ^ in2[50];
    assign G[184] = in[49] & in2[49];
    assign P[184] = in[49] ^ in2[49];
    assign G[185] = in[48] & in2[48];
    assign P[185] = in[48] ^ in2[48];
    assign G[186] = in[47] & in2[47];
    assign P[186] = in[47] ^ in2[47];
    assign G[187] = in[46] & in2[46];
    assign P[187] = in[46] ^ in2[46];
    assign G[188] = in[45] & in2[45];
    assign P[188] = in[45] ^ in2[45];
    assign G[189] = in[44] & in2[44];
    assign P[189] = in[44] ^ in2[44];
    assign G[190] = in[43] & in2[43];
    assign P[190] = in[43] ^ in2[43];
    assign G[191] = in[42] & in2[42];
    assign P[191] = in[42] ^ in2[42];
    assign G[192] = in[41] & in2[41];
    assign P[192] = in[41] ^ in2[41];
    assign G[193] = in[40] & in2[40];
    assign P[193] = in[40] ^ in2[40];
    assign G[194] = in[39] & in2[39];
    assign P[194] = in[39] ^ in2[39];
    assign G[195] = in[38] & in2[38];
    assign P[195] = in[38] ^ in2[38];
    assign G[196] = in[37] & in2[37];
    assign P[196] = in[37] ^ in2[37];
    assign G[197] = in[36] & in2[36];
    assign P[197] = in[36] ^ in2[36];
    assign G[198] = in[35] & in2[35];
    assign P[198] = in[35] ^ in2[35];
    assign G[199] = in[34] & in2[34];
    assign P[199] = in[34] ^ in2[34];
    assign G[200] = in[33] & in2[33];
    assign P[200] = in[33] ^ in2[33];
    assign G[201] = in[32] & in2[32];
    assign P[201] = in[32] ^ in2[32];
    assign G[202] = in[31] & in2[31];
    assign P[202] = in[31] ^ in2[31];
    assign G[203] = in[30] & in2[30];
    assign P[203] = in[30] ^ in2[30];
    assign G[204] = in[29] & in2[29];
    assign P[204] = in[29] ^ in2[29];
    assign G[205] = in[28] & in2[28];
    assign P[205] = in[28] ^ in2[28];
    assign G[206] = in[27] & in2[27];
    assign P[206] = in[27] ^ in2[27];
    assign G[207] = in[26] & in2[26];
    assign P[207] = in[26] ^ in2[26];
    assign G[208] = in[25] & in2[25];
    assign P[208] = in[25] ^ in2[25];
    assign G[209] = in[24] & in2[24];
    assign P[209] = in[24] ^ in2[24];
    assign G[210] = in[23] & in2[23];
    assign P[210] = in[23] ^ in2[23];
    assign G[211] = in[22] & in2[22];
    assign P[211] = in[22] ^ in2[22];
    assign G[212] = in[21] & in2[21];
    assign P[212] = in[21] ^ in2[21];
    assign G[213] = in[20] & in2[20];
    assign P[213] = in[20] ^ in2[20];
    assign G[214] = in[19] & in2[19];
    assign P[214] = in[19] ^ in2[19];
    assign G[215] = in[18] & in2[18];
    assign P[215] = in[18] ^ in2[18];
    assign G[216] = in[17] & in2[17];
    assign P[216] = in[17] ^ in2[17];
    assign G[217] = in[16] & in2[16];
    assign P[217] = in[16] ^ in2[16];
    assign G[218] = in[15] & in2[15];
    assign P[218] = in[15] ^ in2[15];
    assign G[219] = in[14] & in2[14];
    assign P[219] = in[14] ^ in2[14];
    assign G[220] = in[13] & in2[13];
    assign P[220] = in[13] ^ in2[13];
    assign G[221] = in[12] & in2[12];
    assign P[221] = in[12] ^ in2[12];
    assign G[222] = in[11] & in2[11];
    assign P[222] = in[11] ^ in2[11];
    assign G[223] = in[10] & in2[10];
    assign P[223] = in[10] ^ in2[10];
    assign G[224] = in[9] & in2[9];
    assign P[224] = in[9] ^ in2[9];
    assign G[225] = in[8] & in2[8];
    assign P[225] = in[8] ^ in2[8];
    assign G[226] = in[7] & in2[7];
    assign P[226] = in[7] ^ in2[7];
    assign G[227] = in[6] & in2[6];
    assign P[227] = in[6] ^ in2[6];
    assign G[228] = in[5] & in2[5];
    assign P[228] = in[5] ^ in2[5];
    assign G[229] = in[4] & in2[4];
    assign P[229] = in[4] ^ in2[4];
    assign G[230] = in[3] & in2[3];
    assign P[230] = in[3] ^ in2[3];
    assign G[231] = in[2] & in2[2];
    assign P[231] = in[2] ^ in2[2];
    assign G[232] = in[1] & in2[1];
    assign P[232] = in[1] ^ in2[1];
    assign G[233] = in[0] & in2[0];
    assign P[233] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign C[233] = G[232] | (P[232] & C[232]);
    assign cout = G[233] | (P[233] & C[233]);
    assign sum = P ^ C;
endmodule

module CLA233(output [232:0] sum, output cout, input [232:0] in1, input [232:0] in2;

    wire[232:0] G;
    wire[232:0] C;
    wire[232:0] P;

    assign G[0] = in[232] & in2[232];
    assign P[0] = in[232] ^ in2[232];
    assign G[1] = in[231] & in2[231];
    assign P[1] = in[231] ^ in2[231];
    assign G[2] = in[230] & in2[230];
    assign P[2] = in[230] ^ in2[230];
    assign G[3] = in[229] & in2[229];
    assign P[3] = in[229] ^ in2[229];
    assign G[4] = in[228] & in2[228];
    assign P[4] = in[228] ^ in2[228];
    assign G[5] = in[227] & in2[227];
    assign P[5] = in[227] ^ in2[227];
    assign G[6] = in[226] & in2[226];
    assign P[6] = in[226] ^ in2[226];
    assign G[7] = in[225] & in2[225];
    assign P[7] = in[225] ^ in2[225];
    assign G[8] = in[224] & in2[224];
    assign P[8] = in[224] ^ in2[224];
    assign G[9] = in[223] & in2[223];
    assign P[9] = in[223] ^ in2[223];
    assign G[10] = in[222] & in2[222];
    assign P[10] = in[222] ^ in2[222];
    assign G[11] = in[221] & in2[221];
    assign P[11] = in[221] ^ in2[221];
    assign G[12] = in[220] & in2[220];
    assign P[12] = in[220] ^ in2[220];
    assign G[13] = in[219] & in2[219];
    assign P[13] = in[219] ^ in2[219];
    assign G[14] = in[218] & in2[218];
    assign P[14] = in[218] ^ in2[218];
    assign G[15] = in[217] & in2[217];
    assign P[15] = in[217] ^ in2[217];
    assign G[16] = in[216] & in2[216];
    assign P[16] = in[216] ^ in2[216];
    assign G[17] = in[215] & in2[215];
    assign P[17] = in[215] ^ in2[215];
    assign G[18] = in[214] & in2[214];
    assign P[18] = in[214] ^ in2[214];
    assign G[19] = in[213] & in2[213];
    assign P[19] = in[213] ^ in2[213];
    assign G[20] = in[212] & in2[212];
    assign P[20] = in[212] ^ in2[212];
    assign G[21] = in[211] & in2[211];
    assign P[21] = in[211] ^ in2[211];
    assign G[22] = in[210] & in2[210];
    assign P[22] = in[210] ^ in2[210];
    assign G[23] = in[209] & in2[209];
    assign P[23] = in[209] ^ in2[209];
    assign G[24] = in[208] & in2[208];
    assign P[24] = in[208] ^ in2[208];
    assign G[25] = in[207] & in2[207];
    assign P[25] = in[207] ^ in2[207];
    assign G[26] = in[206] & in2[206];
    assign P[26] = in[206] ^ in2[206];
    assign G[27] = in[205] & in2[205];
    assign P[27] = in[205] ^ in2[205];
    assign G[28] = in[204] & in2[204];
    assign P[28] = in[204] ^ in2[204];
    assign G[29] = in[203] & in2[203];
    assign P[29] = in[203] ^ in2[203];
    assign G[30] = in[202] & in2[202];
    assign P[30] = in[202] ^ in2[202];
    assign G[31] = in[201] & in2[201];
    assign P[31] = in[201] ^ in2[201];
    assign G[32] = in[200] & in2[200];
    assign P[32] = in[200] ^ in2[200];
    assign G[33] = in[199] & in2[199];
    assign P[33] = in[199] ^ in2[199];
    assign G[34] = in[198] & in2[198];
    assign P[34] = in[198] ^ in2[198];
    assign G[35] = in[197] & in2[197];
    assign P[35] = in[197] ^ in2[197];
    assign G[36] = in[196] & in2[196];
    assign P[36] = in[196] ^ in2[196];
    assign G[37] = in[195] & in2[195];
    assign P[37] = in[195] ^ in2[195];
    assign G[38] = in[194] & in2[194];
    assign P[38] = in[194] ^ in2[194];
    assign G[39] = in[193] & in2[193];
    assign P[39] = in[193] ^ in2[193];
    assign G[40] = in[192] & in2[192];
    assign P[40] = in[192] ^ in2[192];
    assign G[41] = in[191] & in2[191];
    assign P[41] = in[191] ^ in2[191];
    assign G[42] = in[190] & in2[190];
    assign P[42] = in[190] ^ in2[190];
    assign G[43] = in[189] & in2[189];
    assign P[43] = in[189] ^ in2[189];
    assign G[44] = in[188] & in2[188];
    assign P[44] = in[188] ^ in2[188];
    assign G[45] = in[187] & in2[187];
    assign P[45] = in[187] ^ in2[187];
    assign G[46] = in[186] & in2[186];
    assign P[46] = in[186] ^ in2[186];
    assign G[47] = in[185] & in2[185];
    assign P[47] = in[185] ^ in2[185];
    assign G[48] = in[184] & in2[184];
    assign P[48] = in[184] ^ in2[184];
    assign G[49] = in[183] & in2[183];
    assign P[49] = in[183] ^ in2[183];
    assign G[50] = in[182] & in2[182];
    assign P[50] = in[182] ^ in2[182];
    assign G[51] = in[181] & in2[181];
    assign P[51] = in[181] ^ in2[181];
    assign G[52] = in[180] & in2[180];
    assign P[52] = in[180] ^ in2[180];
    assign G[53] = in[179] & in2[179];
    assign P[53] = in[179] ^ in2[179];
    assign G[54] = in[178] & in2[178];
    assign P[54] = in[178] ^ in2[178];
    assign G[55] = in[177] & in2[177];
    assign P[55] = in[177] ^ in2[177];
    assign G[56] = in[176] & in2[176];
    assign P[56] = in[176] ^ in2[176];
    assign G[57] = in[175] & in2[175];
    assign P[57] = in[175] ^ in2[175];
    assign G[58] = in[174] & in2[174];
    assign P[58] = in[174] ^ in2[174];
    assign G[59] = in[173] & in2[173];
    assign P[59] = in[173] ^ in2[173];
    assign G[60] = in[172] & in2[172];
    assign P[60] = in[172] ^ in2[172];
    assign G[61] = in[171] & in2[171];
    assign P[61] = in[171] ^ in2[171];
    assign G[62] = in[170] & in2[170];
    assign P[62] = in[170] ^ in2[170];
    assign G[63] = in[169] & in2[169];
    assign P[63] = in[169] ^ in2[169];
    assign G[64] = in[168] & in2[168];
    assign P[64] = in[168] ^ in2[168];
    assign G[65] = in[167] & in2[167];
    assign P[65] = in[167] ^ in2[167];
    assign G[66] = in[166] & in2[166];
    assign P[66] = in[166] ^ in2[166];
    assign G[67] = in[165] & in2[165];
    assign P[67] = in[165] ^ in2[165];
    assign G[68] = in[164] & in2[164];
    assign P[68] = in[164] ^ in2[164];
    assign G[69] = in[163] & in2[163];
    assign P[69] = in[163] ^ in2[163];
    assign G[70] = in[162] & in2[162];
    assign P[70] = in[162] ^ in2[162];
    assign G[71] = in[161] & in2[161];
    assign P[71] = in[161] ^ in2[161];
    assign G[72] = in[160] & in2[160];
    assign P[72] = in[160] ^ in2[160];
    assign G[73] = in[159] & in2[159];
    assign P[73] = in[159] ^ in2[159];
    assign G[74] = in[158] & in2[158];
    assign P[74] = in[158] ^ in2[158];
    assign G[75] = in[157] & in2[157];
    assign P[75] = in[157] ^ in2[157];
    assign G[76] = in[156] & in2[156];
    assign P[76] = in[156] ^ in2[156];
    assign G[77] = in[155] & in2[155];
    assign P[77] = in[155] ^ in2[155];
    assign G[78] = in[154] & in2[154];
    assign P[78] = in[154] ^ in2[154];
    assign G[79] = in[153] & in2[153];
    assign P[79] = in[153] ^ in2[153];
    assign G[80] = in[152] & in2[152];
    assign P[80] = in[152] ^ in2[152];
    assign G[81] = in[151] & in2[151];
    assign P[81] = in[151] ^ in2[151];
    assign G[82] = in[150] & in2[150];
    assign P[82] = in[150] ^ in2[150];
    assign G[83] = in[149] & in2[149];
    assign P[83] = in[149] ^ in2[149];
    assign G[84] = in[148] & in2[148];
    assign P[84] = in[148] ^ in2[148];
    assign G[85] = in[147] & in2[147];
    assign P[85] = in[147] ^ in2[147];
    assign G[86] = in[146] & in2[146];
    assign P[86] = in[146] ^ in2[146];
    assign G[87] = in[145] & in2[145];
    assign P[87] = in[145] ^ in2[145];
    assign G[88] = in[144] & in2[144];
    assign P[88] = in[144] ^ in2[144];
    assign G[89] = in[143] & in2[143];
    assign P[89] = in[143] ^ in2[143];
    assign G[90] = in[142] & in2[142];
    assign P[90] = in[142] ^ in2[142];
    assign G[91] = in[141] & in2[141];
    assign P[91] = in[141] ^ in2[141];
    assign G[92] = in[140] & in2[140];
    assign P[92] = in[140] ^ in2[140];
    assign G[93] = in[139] & in2[139];
    assign P[93] = in[139] ^ in2[139];
    assign G[94] = in[138] & in2[138];
    assign P[94] = in[138] ^ in2[138];
    assign G[95] = in[137] & in2[137];
    assign P[95] = in[137] ^ in2[137];
    assign G[96] = in[136] & in2[136];
    assign P[96] = in[136] ^ in2[136];
    assign G[97] = in[135] & in2[135];
    assign P[97] = in[135] ^ in2[135];
    assign G[98] = in[134] & in2[134];
    assign P[98] = in[134] ^ in2[134];
    assign G[99] = in[133] & in2[133];
    assign P[99] = in[133] ^ in2[133];
    assign G[100] = in[132] & in2[132];
    assign P[100] = in[132] ^ in2[132];
    assign G[101] = in[131] & in2[131];
    assign P[101] = in[131] ^ in2[131];
    assign G[102] = in[130] & in2[130];
    assign P[102] = in[130] ^ in2[130];
    assign G[103] = in[129] & in2[129];
    assign P[103] = in[129] ^ in2[129];
    assign G[104] = in[128] & in2[128];
    assign P[104] = in[128] ^ in2[128];
    assign G[105] = in[127] & in2[127];
    assign P[105] = in[127] ^ in2[127];
    assign G[106] = in[126] & in2[126];
    assign P[106] = in[126] ^ in2[126];
    assign G[107] = in[125] & in2[125];
    assign P[107] = in[125] ^ in2[125];
    assign G[108] = in[124] & in2[124];
    assign P[108] = in[124] ^ in2[124];
    assign G[109] = in[123] & in2[123];
    assign P[109] = in[123] ^ in2[123];
    assign G[110] = in[122] & in2[122];
    assign P[110] = in[122] ^ in2[122];
    assign G[111] = in[121] & in2[121];
    assign P[111] = in[121] ^ in2[121];
    assign G[112] = in[120] & in2[120];
    assign P[112] = in[120] ^ in2[120];
    assign G[113] = in[119] & in2[119];
    assign P[113] = in[119] ^ in2[119];
    assign G[114] = in[118] & in2[118];
    assign P[114] = in[118] ^ in2[118];
    assign G[115] = in[117] & in2[117];
    assign P[115] = in[117] ^ in2[117];
    assign G[116] = in[116] & in2[116];
    assign P[116] = in[116] ^ in2[116];
    assign G[117] = in[115] & in2[115];
    assign P[117] = in[115] ^ in2[115];
    assign G[118] = in[114] & in2[114];
    assign P[118] = in[114] ^ in2[114];
    assign G[119] = in[113] & in2[113];
    assign P[119] = in[113] ^ in2[113];
    assign G[120] = in[112] & in2[112];
    assign P[120] = in[112] ^ in2[112];
    assign G[121] = in[111] & in2[111];
    assign P[121] = in[111] ^ in2[111];
    assign G[122] = in[110] & in2[110];
    assign P[122] = in[110] ^ in2[110];
    assign G[123] = in[109] & in2[109];
    assign P[123] = in[109] ^ in2[109];
    assign G[124] = in[108] & in2[108];
    assign P[124] = in[108] ^ in2[108];
    assign G[125] = in[107] & in2[107];
    assign P[125] = in[107] ^ in2[107];
    assign G[126] = in[106] & in2[106];
    assign P[126] = in[106] ^ in2[106];
    assign G[127] = in[105] & in2[105];
    assign P[127] = in[105] ^ in2[105];
    assign G[128] = in[104] & in2[104];
    assign P[128] = in[104] ^ in2[104];
    assign G[129] = in[103] & in2[103];
    assign P[129] = in[103] ^ in2[103];
    assign G[130] = in[102] & in2[102];
    assign P[130] = in[102] ^ in2[102];
    assign G[131] = in[101] & in2[101];
    assign P[131] = in[101] ^ in2[101];
    assign G[132] = in[100] & in2[100];
    assign P[132] = in[100] ^ in2[100];
    assign G[133] = in[99] & in2[99];
    assign P[133] = in[99] ^ in2[99];
    assign G[134] = in[98] & in2[98];
    assign P[134] = in[98] ^ in2[98];
    assign G[135] = in[97] & in2[97];
    assign P[135] = in[97] ^ in2[97];
    assign G[136] = in[96] & in2[96];
    assign P[136] = in[96] ^ in2[96];
    assign G[137] = in[95] & in2[95];
    assign P[137] = in[95] ^ in2[95];
    assign G[138] = in[94] & in2[94];
    assign P[138] = in[94] ^ in2[94];
    assign G[139] = in[93] & in2[93];
    assign P[139] = in[93] ^ in2[93];
    assign G[140] = in[92] & in2[92];
    assign P[140] = in[92] ^ in2[92];
    assign G[141] = in[91] & in2[91];
    assign P[141] = in[91] ^ in2[91];
    assign G[142] = in[90] & in2[90];
    assign P[142] = in[90] ^ in2[90];
    assign G[143] = in[89] & in2[89];
    assign P[143] = in[89] ^ in2[89];
    assign G[144] = in[88] & in2[88];
    assign P[144] = in[88] ^ in2[88];
    assign G[145] = in[87] & in2[87];
    assign P[145] = in[87] ^ in2[87];
    assign G[146] = in[86] & in2[86];
    assign P[146] = in[86] ^ in2[86];
    assign G[147] = in[85] & in2[85];
    assign P[147] = in[85] ^ in2[85];
    assign G[148] = in[84] & in2[84];
    assign P[148] = in[84] ^ in2[84];
    assign G[149] = in[83] & in2[83];
    assign P[149] = in[83] ^ in2[83];
    assign G[150] = in[82] & in2[82];
    assign P[150] = in[82] ^ in2[82];
    assign G[151] = in[81] & in2[81];
    assign P[151] = in[81] ^ in2[81];
    assign G[152] = in[80] & in2[80];
    assign P[152] = in[80] ^ in2[80];
    assign G[153] = in[79] & in2[79];
    assign P[153] = in[79] ^ in2[79];
    assign G[154] = in[78] & in2[78];
    assign P[154] = in[78] ^ in2[78];
    assign G[155] = in[77] & in2[77];
    assign P[155] = in[77] ^ in2[77];
    assign G[156] = in[76] & in2[76];
    assign P[156] = in[76] ^ in2[76];
    assign G[157] = in[75] & in2[75];
    assign P[157] = in[75] ^ in2[75];
    assign G[158] = in[74] & in2[74];
    assign P[158] = in[74] ^ in2[74];
    assign G[159] = in[73] & in2[73];
    assign P[159] = in[73] ^ in2[73];
    assign G[160] = in[72] & in2[72];
    assign P[160] = in[72] ^ in2[72];
    assign G[161] = in[71] & in2[71];
    assign P[161] = in[71] ^ in2[71];
    assign G[162] = in[70] & in2[70];
    assign P[162] = in[70] ^ in2[70];
    assign G[163] = in[69] & in2[69];
    assign P[163] = in[69] ^ in2[69];
    assign G[164] = in[68] & in2[68];
    assign P[164] = in[68] ^ in2[68];
    assign G[165] = in[67] & in2[67];
    assign P[165] = in[67] ^ in2[67];
    assign G[166] = in[66] & in2[66];
    assign P[166] = in[66] ^ in2[66];
    assign G[167] = in[65] & in2[65];
    assign P[167] = in[65] ^ in2[65];
    assign G[168] = in[64] & in2[64];
    assign P[168] = in[64] ^ in2[64];
    assign G[169] = in[63] & in2[63];
    assign P[169] = in[63] ^ in2[63];
    assign G[170] = in[62] & in2[62];
    assign P[170] = in[62] ^ in2[62];
    assign G[171] = in[61] & in2[61];
    assign P[171] = in[61] ^ in2[61];
    assign G[172] = in[60] & in2[60];
    assign P[172] = in[60] ^ in2[60];
    assign G[173] = in[59] & in2[59];
    assign P[173] = in[59] ^ in2[59];
    assign G[174] = in[58] & in2[58];
    assign P[174] = in[58] ^ in2[58];
    assign G[175] = in[57] & in2[57];
    assign P[175] = in[57] ^ in2[57];
    assign G[176] = in[56] & in2[56];
    assign P[176] = in[56] ^ in2[56];
    assign G[177] = in[55] & in2[55];
    assign P[177] = in[55] ^ in2[55];
    assign G[178] = in[54] & in2[54];
    assign P[178] = in[54] ^ in2[54];
    assign G[179] = in[53] & in2[53];
    assign P[179] = in[53] ^ in2[53];
    assign G[180] = in[52] & in2[52];
    assign P[180] = in[52] ^ in2[52];
    assign G[181] = in[51] & in2[51];
    assign P[181] = in[51] ^ in2[51];
    assign G[182] = in[50] & in2[50];
    assign P[182] = in[50] ^ in2[50];
    assign G[183] = in[49] & in2[49];
    assign P[183] = in[49] ^ in2[49];
    assign G[184] = in[48] & in2[48];
    assign P[184] = in[48] ^ in2[48];
    assign G[185] = in[47] & in2[47];
    assign P[185] = in[47] ^ in2[47];
    assign G[186] = in[46] & in2[46];
    assign P[186] = in[46] ^ in2[46];
    assign G[187] = in[45] & in2[45];
    assign P[187] = in[45] ^ in2[45];
    assign G[188] = in[44] & in2[44];
    assign P[188] = in[44] ^ in2[44];
    assign G[189] = in[43] & in2[43];
    assign P[189] = in[43] ^ in2[43];
    assign G[190] = in[42] & in2[42];
    assign P[190] = in[42] ^ in2[42];
    assign G[191] = in[41] & in2[41];
    assign P[191] = in[41] ^ in2[41];
    assign G[192] = in[40] & in2[40];
    assign P[192] = in[40] ^ in2[40];
    assign G[193] = in[39] & in2[39];
    assign P[193] = in[39] ^ in2[39];
    assign G[194] = in[38] & in2[38];
    assign P[194] = in[38] ^ in2[38];
    assign G[195] = in[37] & in2[37];
    assign P[195] = in[37] ^ in2[37];
    assign G[196] = in[36] & in2[36];
    assign P[196] = in[36] ^ in2[36];
    assign G[197] = in[35] & in2[35];
    assign P[197] = in[35] ^ in2[35];
    assign G[198] = in[34] & in2[34];
    assign P[198] = in[34] ^ in2[34];
    assign G[199] = in[33] & in2[33];
    assign P[199] = in[33] ^ in2[33];
    assign G[200] = in[32] & in2[32];
    assign P[200] = in[32] ^ in2[32];
    assign G[201] = in[31] & in2[31];
    assign P[201] = in[31] ^ in2[31];
    assign G[202] = in[30] & in2[30];
    assign P[202] = in[30] ^ in2[30];
    assign G[203] = in[29] & in2[29];
    assign P[203] = in[29] ^ in2[29];
    assign G[204] = in[28] & in2[28];
    assign P[204] = in[28] ^ in2[28];
    assign G[205] = in[27] & in2[27];
    assign P[205] = in[27] ^ in2[27];
    assign G[206] = in[26] & in2[26];
    assign P[206] = in[26] ^ in2[26];
    assign G[207] = in[25] & in2[25];
    assign P[207] = in[25] ^ in2[25];
    assign G[208] = in[24] & in2[24];
    assign P[208] = in[24] ^ in2[24];
    assign G[209] = in[23] & in2[23];
    assign P[209] = in[23] ^ in2[23];
    assign G[210] = in[22] & in2[22];
    assign P[210] = in[22] ^ in2[22];
    assign G[211] = in[21] & in2[21];
    assign P[211] = in[21] ^ in2[21];
    assign G[212] = in[20] & in2[20];
    assign P[212] = in[20] ^ in2[20];
    assign G[213] = in[19] & in2[19];
    assign P[213] = in[19] ^ in2[19];
    assign G[214] = in[18] & in2[18];
    assign P[214] = in[18] ^ in2[18];
    assign G[215] = in[17] & in2[17];
    assign P[215] = in[17] ^ in2[17];
    assign G[216] = in[16] & in2[16];
    assign P[216] = in[16] ^ in2[16];
    assign G[217] = in[15] & in2[15];
    assign P[217] = in[15] ^ in2[15];
    assign G[218] = in[14] & in2[14];
    assign P[218] = in[14] ^ in2[14];
    assign G[219] = in[13] & in2[13];
    assign P[219] = in[13] ^ in2[13];
    assign G[220] = in[12] & in2[12];
    assign P[220] = in[12] ^ in2[12];
    assign G[221] = in[11] & in2[11];
    assign P[221] = in[11] ^ in2[11];
    assign G[222] = in[10] & in2[10];
    assign P[222] = in[10] ^ in2[10];
    assign G[223] = in[9] & in2[9];
    assign P[223] = in[9] ^ in2[9];
    assign G[224] = in[8] & in2[8];
    assign P[224] = in[8] ^ in2[8];
    assign G[225] = in[7] & in2[7];
    assign P[225] = in[7] ^ in2[7];
    assign G[226] = in[6] & in2[6];
    assign P[226] = in[6] ^ in2[6];
    assign G[227] = in[5] & in2[5];
    assign P[227] = in[5] ^ in2[5];
    assign G[228] = in[4] & in2[4];
    assign P[228] = in[4] ^ in2[4];
    assign G[229] = in[3] & in2[3];
    assign P[229] = in[3] ^ in2[3];
    assign G[230] = in[2] & in2[2];
    assign P[230] = in[2] ^ in2[2];
    assign G[231] = in[1] & in2[1];
    assign P[231] = in[1] ^ in2[1];
    assign G[232] = in[0] & in2[0];
    assign P[232] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign C[232] = G[231] | (P[231] & C[231]);
    assign cout = G[232] | (P[232] & C[232]);
    assign sum = P ^ C;
endmodule

module CLA232(output [231:0] sum, output cout, input [231:0] in1, input [231:0] in2;

    wire[231:0] G;
    wire[231:0] C;
    wire[231:0] P;

    assign G[0] = in[231] & in2[231];
    assign P[0] = in[231] ^ in2[231];
    assign G[1] = in[230] & in2[230];
    assign P[1] = in[230] ^ in2[230];
    assign G[2] = in[229] & in2[229];
    assign P[2] = in[229] ^ in2[229];
    assign G[3] = in[228] & in2[228];
    assign P[3] = in[228] ^ in2[228];
    assign G[4] = in[227] & in2[227];
    assign P[4] = in[227] ^ in2[227];
    assign G[5] = in[226] & in2[226];
    assign P[5] = in[226] ^ in2[226];
    assign G[6] = in[225] & in2[225];
    assign P[6] = in[225] ^ in2[225];
    assign G[7] = in[224] & in2[224];
    assign P[7] = in[224] ^ in2[224];
    assign G[8] = in[223] & in2[223];
    assign P[8] = in[223] ^ in2[223];
    assign G[9] = in[222] & in2[222];
    assign P[9] = in[222] ^ in2[222];
    assign G[10] = in[221] & in2[221];
    assign P[10] = in[221] ^ in2[221];
    assign G[11] = in[220] & in2[220];
    assign P[11] = in[220] ^ in2[220];
    assign G[12] = in[219] & in2[219];
    assign P[12] = in[219] ^ in2[219];
    assign G[13] = in[218] & in2[218];
    assign P[13] = in[218] ^ in2[218];
    assign G[14] = in[217] & in2[217];
    assign P[14] = in[217] ^ in2[217];
    assign G[15] = in[216] & in2[216];
    assign P[15] = in[216] ^ in2[216];
    assign G[16] = in[215] & in2[215];
    assign P[16] = in[215] ^ in2[215];
    assign G[17] = in[214] & in2[214];
    assign P[17] = in[214] ^ in2[214];
    assign G[18] = in[213] & in2[213];
    assign P[18] = in[213] ^ in2[213];
    assign G[19] = in[212] & in2[212];
    assign P[19] = in[212] ^ in2[212];
    assign G[20] = in[211] & in2[211];
    assign P[20] = in[211] ^ in2[211];
    assign G[21] = in[210] & in2[210];
    assign P[21] = in[210] ^ in2[210];
    assign G[22] = in[209] & in2[209];
    assign P[22] = in[209] ^ in2[209];
    assign G[23] = in[208] & in2[208];
    assign P[23] = in[208] ^ in2[208];
    assign G[24] = in[207] & in2[207];
    assign P[24] = in[207] ^ in2[207];
    assign G[25] = in[206] & in2[206];
    assign P[25] = in[206] ^ in2[206];
    assign G[26] = in[205] & in2[205];
    assign P[26] = in[205] ^ in2[205];
    assign G[27] = in[204] & in2[204];
    assign P[27] = in[204] ^ in2[204];
    assign G[28] = in[203] & in2[203];
    assign P[28] = in[203] ^ in2[203];
    assign G[29] = in[202] & in2[202];
    assign P[29] = in[202] ^ in2[202];
    assign G[30] = in[201] & in2[201];
    assign P[30] = in[201] ^ in2[201];
    assign G[31] = in[200] & in2[200];
    assign P[31] = in[200] ^ in2[200];
    assign G[32] = in[199] & in2[199];
    assign P[32] = in[199] ^ in2[199];
    assign G[33] = in[198] & in2[198];
    assign P[33] = in[198] ^ in2[198];
    assign G[34] = in[197] & in2[197];
    assign P[34] = in[197] ^ in2[197];
    assign G[35] = in[196] & in2[196];
    assign P[35] = in[196] ^ in2[196];
    assign G[36] = in[195] & in2[195];
    assign P[36] = in[195] ^ in2[195];
    assign G[37] = in[194] & in2[194];
    assign P[37] = in[194] ^ in2[194];
    assign G[38] = in[193] & in2[193];
    assign P[38] = in[193] ^ in2[193];
    assign G[39] = in[192] & in2[192];
    assign P[39] = in[192] ^ in2[192];
    assign G[40] = in[191] & in2[191];
    assign P[40] = in[191] ^ in2[191];
    assign G[41] = in[190] & in2[190];
    assign P[41] = in[190] ^ in2[190];
    assign G[42] = in[189] & in2[189];
    assign P[42] = in[189] ^ in2[189];
    assign G[43] = in[188] & in2[188];
    assign P[43] = in[188] ^ in2[188];
    assign G[44] = in[187] & in2[187];
    assign P[44] = in[187] ^ in2[187];
    assign G[45] = in[186] & in2[186];
    assign P[45] = in[186] ^ in2[186];
    assign G[46] = in[185] & in2[185];
    assign P[46] = in[185] ^ in2[185];
    assign G[47] = in[184] & in2[184];
    assign P[47] = in[184] ^ in2[184];
    assign G[48] = in[183] & in2[183];
    assign P[48] = in[183] ^ in2[183];
    assign G[49] = in[182] & in2[182];
    assign P[49] = in[182] ^ in2[182];
    assign G[50] = in[181] & in2[181];
    assign P[50] = in[181] ^ in2[181];
    assign G[51] = in[180] & in2[180];
    assign P[51] = in[180] ^ in2[180];
    assign G[52] = in[179] & in2[179];
    assign P[52] = in[179] ^ in2[179];
    assign G[53] = in[178] & in2[178];
    assign P[53] = in[178] ^ in2[178];
    assign G[54] = in[177] & in2[177];
    assign P[54] = in[177] ^ in2[177];
    assign G[55] = in[176] & in2[176];
    assign P[55] = in[176] ^ in2[176];
    assign G[56] = in[175] & in2[175];
    assign P[56] = in[175] ^ in2[175];
    assign G[57] = in[174] & in2[174];
    assign P[57] = in[174] ^ in2[174];
    assign G[58] = in[173] & in2[173];
    assign P[58] = in[173] ^ in2[173];
    assign G[59] = in[172] & in2[172];
    assign P[59] = in[172] ^ in2[172];
    assign G[60] = in[171] & in2[171];
    assign P[60] = in[171] ^ in2[171];
    assign G[61] = in[170] & in2[170];
    assign P[61] = in[170] ^ in2[170];
    assign G[62] = in[169] & in2[169];
    assign P[62] = in[169] ^ in2[169];
    assign G[63] = in[168] & in2[168];
    assign P[63] = in[168] ^ in2[168];
    assign G[64] = in[167] & in2[167];
    assign P[64] = in[167] ^ in2[167];
    assign G[65] = in[166] & in2[166];
    assign P[65] = in[166] ^ in2[166];
    assign G[66] = in[165] & in2[165];
    assign P[66] = in[165] ^ in2[165];
    assign G[67] = in[164] & in2[164];
    assign P[67] = in[164] ^ in2[164];
    assign G[68] = in[163] & in2[163];
    assign P[68] = in[163] ^ in2[163];
    assign G[69] = in[162] & in2[162];
    assign P[69] = in[162] ^ in2[162];
    assign G[70] = in[161] & in2[161];
    assign P[70] = in[161] ^ in2[161];
    assign G[71] = in[160] & in2[160];
    assign P[71] = in[160] ^ in2[160];
    assign G[72] = in[159] & in2[159];
    assign P[72] = in[159] ^ in2[159];
    assign G[73] = in[158] & in2[158];
    assign P[73] = in[158] ^ in2[158];
    assign G[74] = in[157] & in2[157];
    assign P[74] = in[157] ^ in2[157];
    assign G[75] = in[156] & in2[156];
    assign P[75] = in[156] ^ in2[156];
    assign G[76] = in[155] & in2[155];
    assign P[76] = in[155] ^ in2[155];
    assign G[77] = in[154] & in2[154];
    assign P[77] = in[154] ^ in2[154];
    assign G[78] = in[153] & in2[153];
    assign P[78] = in[153] ^ in2[153];
    assign G[79] = in[152] & in2[152];
    assign P[79] = in[152] ^ in2[152];
    assign G[80] = in[151] & in2[151];
    assign P[80] = in[151] ^ in2[151];
    assign G[81] = in[150] & in2[150];
    assign P[81] = in[150] ^ in2[150];
    assign G[82] = in[149] & in2[149];
    assign P[82] = in[149] ^ in2[149];
    assign G[83] = in[148] & in2[148];
    assign P[83] = in[148] ^ in2[148];
    assign G[84] = in[147] & in2[147];
    assign P[84] = in[147] ^ in2[147];
    assign G[85] = in[146] & in2[146];
    assign P[85] = in[146] ^ in2[146];
    assign G[86] = in[145] & in2[145];
    assign P[86] = in[145] ^ in2[145];
    assign G[87] = in[144] & in2[144];
    assign P[87] = in[144] ^ in2[144];
    assign G[88] = in[143] & in2[143];
    assign P[88] = in[143] ^ in2[143];
    assign G[89] = in[142] & in2[142];
    assign P[89] = in[142] ^ in2[142];
    assign G[90] = in[141] & in2[141];
    assign P[90] = in[141] ^ in2[141];
    assign G[91] = in[140] & in2[140];
    assign P[91] = in[140] ^ in2[140];
    assign G[92] = in[139] & in2[139];
    assign P[92] = in[139] ^ in2[139];
    assign G[93] = in[138] & in2[138];
    assign P[93] = in[138] ^ in2[138];
    assign G[94] = in[137] & in2[137];
    assign P[94] = in[137] ^ in2[137];
    assign G[95] = in[136] & in2[136];
    assign P[95] = in[136] ^ in2[136];
    assign G[96] = in[135] & in2[135];
    assign P[96] = in[135] ^ in2[135];
    assign G[97] = in[134] & in2[134];
    assign P[97] = in[134] ^ in2[134];
    assign G[98] = in[133] & in2[133];
    assign P[98] = in[133] ^ in2[133];
    assign G[99] = in[132] & in2[132];
    assign P[99] = in[132] ^ in2[132];
    assign G[100] = in[131] & in2[131];
    assign P[100] = in[131] ^ in2[131];
    assign G[101] = in[130] & in2[130];
    assign P[101] = in[130] ^ in2[130];
    assign G[102] = in[129] & in2[129];
    assign P[102] = in[129] ^ in2[129];
    assign G[103] = in[128] & in2[128];
    assign P[103] = in[128] ^ in2[128];
    assign G[104] = in[127] & in2[127];
    assign P[104] = in[127] ^ in2[127];
    assign G[105] = in[126] & in2[126];
    assign P[105] = in[126] ^ in2[126];
    assign G[106] = in[125] & in2[125];
    assign P[106] = in[125] ^ in2[125];
    assign G[107] = in[124] & in2[124];
    assign P[107] = in[124] ^ in2[124];
    assign G[108] = in[123] & in2[123];
    assign P[108] = in[123] ^ in2[123];
    assign G[109] = in[122] & in2[122];
    assign P[109] = in[122] ^ in2[122];
    assign G[110] = in[121] & in2[121];
    assign P[110] = in[121] ^ in2[121];
    assign G[111] = in[120] & in2[120];
    assign P[111] = in[120] ^ in2[120];
    assign G[112] = in[119] & in2[119];
    assign P[112] = in[119] ^ in2[119];
    assign G[113] = in[118] & in2[118];
    assign P[113] = in[118] ^ in2[118];
    assign G[114] = in[117] & in2[117];
    assign P[114] = in[117] ^ in2[117];
    assign G[115] = in[116] & in2[116];
    assign P[115] = in[116] ^ in2[116];
    assign G[116] = in[115] & in2[115];
    assign P[116] = in[115] ^ in2[115];
    assign G[117] = in[114] & in2[114];
    assign P[117] = in[114] ^ in2[114];
    assign G[118] = in[113] & in2[113];
    assign P[118] = in[113] ^ in2[113];
    assign G[119] = in[112] & in2[112];
    assign P[119] = in[112] ^ in2[112];
    assign G[120] = in[111] & in2[111];
    assign P[120] = in[111] ^ in2[111];
    assign G[121] = in[110] & in2[110];
    assign P[121] = in[110] ^ in2[110];
    assign G[122] = in[109] & in2[109];
    assign P[122] = in[109] ^ in2[109];
    assign G[123] = in[108] & in2[108];
    assign P[123] = in[108] ^ in2[108];
    assign G[124] = in[107] & in2[107];
    assign P[124] = in[107] ^ in2[107];
    assign G[125] = in[106] & in2[106];
    assign P[125] = in[106] ^ in2[106];
    assign G[126] = in[105] & in2[105];
    assign P[126] = in[105] ^ in2[105];
    assign G[127] = in[104] & in2[104];
    assign P[127] = in[104] ^ in2[104];
    assign G[128] = in[103] & in2[103];
    assign P[128] = in[103] ^ in2[103];
    assign G[129] = in[102] & in2[102];
    assign P[129] = in[102] ^ in2[102];
    assign G[130] = in[101] & in2[101];
    assign P[130] = in[101] ^ in2[101];
    assign G[131] = in[100] & in2[100];
    assign P[131] = in[100] ^ in2[100];
    assign G[132] = in[99] & in2[99];
    assign P[132] = in[99] ^ in2[99];
    assign G[133] = in[98] & in2[98];
    assign P[133] = in[98] ^ in2[98];
    assign G[134] = in[97] & in2[97];
    assign P[134] = in[97] ^ in2[97];
    assign G[135] = in[96] & in2[96];
    assign P[135] = in[96] ^ in2[96];
    assign G[136] = in[95] & in2[95];
    assign P[136] = in[95] ^ in2[95];
    assign G[137] = in[94] & in2[94];
    assign P[137] = in[94] ^ in2[94];
    assign G[138] = in[93] & in2[93];
    assign P[138] = in[93] ^ in2[93];
    assign G[139] = in[92] & in2[92];
    assign P[139] = in[92] ^ in2[92];
    assign G[140] = in[91] & in2[91];
    assign P[140] = in[91] ^ in2[91];
    assign G[141] = in[90] & in2[90];
    assign P[141] = in[90] ^ in2[90];
    assign G[142] = in[89] & in2[89];
    assign P[142] = in[89] ^ in2[89];
    assign G[143] = in[88] & in2[88];
    assign P[143] = in[88] ^ in2[88];
    assign G[144] = in[87] & in2[87];
    assign P[144] = in[87] ^ in2[87];
    assign G[145] = in[86] & in2[86];
    assign P[145] = in[86] ^ in2[86];
    assign G[146] = in[85] & in2[85];
    assign P[146] = in[85] ^ in2[85];
    assign G[147] = in[84] & in2[84];
    assign P[147] = in[84] ^ in2[84];
    assign G[148] = in[83] & in2[83];
    assign P[148] = in[83] ^ in2[83];
    assign G[149] = in[82] & in2[82];
    assign P[149] = in[82] ^ in2[82];
    assign G[150] = in[81] & in2[81];
    assign P[150] = in[81] ^ in2[81];
    assign G[151] = in[80] & in2[80];
    assign P[151] = in[80] ^ in2[80];
    assign G[152] = in[79] & in2[79];
    assign P[152] = in[79] ^ in2[79];
    assign G[153] = in[78] & in2[78];
    assign P[153] = in[78] ^ in2[78];
    assign G[154] = in[77] & in2[77];
    assign P[154] = in[77] ^ in2[77];
    assign G[155] = in[76] & in2[76];
    assign P[155] = in[76] ^ in2[76];
    assign G[156] = in[75] & in2[75];
    assign P[156] = in[75] ^ in2[75];
    assign G[157] = in[74] & in2[74];
    assign P[157] = in[74] ^ in2[74];
    assign G[158] = in[73] & in2[73];
    assign P[158] = in[73] ^ in2[73];
    assign G[159] = in[72] & in2[72];
    assign P[159] = in[72] ^ in2[72];
    assign G[160] = in[71] & in2[71];
    assign P[160] = in[71] ^ in2[71];
    assign G[161] = in[70] & in2[70];
    assign P[161] = in[70] ^ in2[70];
    assign G[162] = in[69] & in2[69];
    assign P[162] = in[69] ^ in2[69];
    assign G[163] = in[68] & in2[68];
    assign P[163] = in[68] ^ in2[68];
    assign G[164] = in[67] & in2[67];
    assign P[164] = in[67] ^ in2[67];
    assign G[165] = in[66] & in2[66];
    assign P[165] = in[66] ^ in2[66];
    assign G[166] = in[65] & in2[65];
    assign P[166] = in[65] ^ in2[65];
    assign G[167] = in[64] & in2[64];
    assign P[167] = in[64] ^ in2[64];
    assign G[168] = in[63] & in2[63];
    assign P[168] = in[63] ^ in2[63];
    assign G[169] = in[62] & in2[62];
    assign P[169] = in[62] ^ in2[62];
    assign G[170] = in[61] & in2[61];
    assign P[170] = in[61] ^ in2[61];
    assign G[171] = in[60] & in2[60];
    assign P[171] = in[60] ^ in2[60];
    assign G[172] = in[59] & in2[59];
    assign P[172] = in[59] ^ in2[59];
    assign G[173] = in[58] & in2[58];
    assign P[173] = in[58] ^ in2[58];
    assign G[174] = in[57] & in2[57];
    assign P[174] = in[57] ^ in2[57];
    assign G[175] = in[56] & in2[56];
    assign P[175] = in[56] ^ in2[56];
    assign G[176] = in[55] & in2[55];
    assign P[176] = in[55] ^ in2[55];
    assign G[177] = in[54] & in2[54];
    assign P[177] = in[54] ^ in2[54];
    assign G[178] = in[53] & in2[53];
    assign P[178] = in[53] ^ in2[53];
    assign G[179] = in[52] & in2[52];
    assign P[179] = in[52] ^ in2[52];
    assign G[180] = in[51] & in2[51];
    assign P[180] = in[51] ^ in2[51];
    assign G[181] = in[50] & in2[50];
    assign P[181] = in[50] ^ in2[50];
    assign G[182] = in[49] & in2[49];
    assign P[182] = in[49] ^ in2[49];
    assign G[183] = in[48] & in2[48];
    assign P[183] = in[48] ^ in2[48];
    assign G[184] = in[47] & in2[47];
    assign P[184] = in[47] ^ in2[47];
    assign G[185] = in[46] & in2[46];
    assign P[185] = in[46] ^ in2[46];
    assign G[186] = in[45] & in2[45];
    assign P[186] = in[45] ^ in2[45];
    assign G[187] = in[44] & in2[44];
    assign P[187] = in[44] ^ in2[44];
    assign G[188] = in[43] & in2[43];
    assign P[188] = in[43] ^ in2[43];
    assign G[189] = in[42] & in2[42];
    assign P[189] = in[42] ^ in2[42];
    assign G[190] = in[41] & in2[41];
    assign P[190] = in[41] ^ in2[41];
    assign G[191] = in[40] & in2[40];
    assign P[191] = in[40] ^ in2[40];
    assign G[192] = in[39] & in2[39];
    assign P[192] = in[39] ^ in2[39];
    assign G[193] = in[38] & in2[38];
    assign P[193] = in[38] ^ in2[38];
    assign G[194] = in[37] & in2[37];
    assign P[194] = in[37] ^ in2[37];
    assign G[195] = in[36] & in2[36];
    assign P[195] = in[36] ^ in2[36];
    assign G[196] = in[35] & in2[35];
    assign P[196] = in[35] ^ in2[35];
    assign G[197] = in[34] & in2[34];
    assign P[197] = in[34] ^ in2[34];
    assign G[198] = in[33] & in2[33];
    assign P[198] = in[33] ^ in2[33];
    assign G[199] = in[32] & in2[32];
    assign P[199] = in[32] ^ in2[32];
    assign G[200] = in[31] & in2[31];
    assign P[200] = in[31] ^ in2[31];
    assign G[201] = in[30] & in2[30];
    assign P[201] = in[30] ^ in2[30];
    assign G[202] = in[29] & in2[29];
    assign P[202] = in[29] ^ in2[29];
    assign G[203] = in[28] & in2[28];
    assign P[203] = in[28] ^ in2[28];
    assign G[204] = in[27] & in2[27];
    assign P[204] = in[27] ^ in2[27];
    assign G[205] = in[26] & in2[26];
    assign P[205] = in[26] ^ in2[26];
    assign G[206] = in[25] & in2[25];
    assign P[206] = in[25] ^ in2[25];
    assign G[207] = in[24] & in2[24];
    assign P[207] = in[24] ^ in2[24];
    assign G[208] = in[23] & in2[23];
    assign P[208] = in[23] ^ in2[23];
    assign G[209] = in[22] & in2[22];
    assign P[209] = in[22] ^ in2[22];
    assign G[210] = in[21] & in2[21];
    assign P[210] = in[21] ^ in2[21];
    assign G[211] = in[20] & in2[20];
    assign P[211] = in[20] ^ in2[20];
    assign G[212] = in[19] & in2[19];
    assign P[212] = in[19] ^ in2[19];
    assign G[213] = in[18] & in2[18];
    assign P[213] = in[18] ^ in2[18];
    assign G[214] = in[17] & in2[17];
    assign P[214] = in[17] ^ in2[17];
    assign G[215] = in[16] & in2[16];
    assign P[215] = in[16] ^ in2[16];
    assign G[216] = in[15] & in2[15];
    assign P[216] = in[15] ^ in2[15];
    assign G[217] = in[14] & in2[14];
    assign P[217] = in[14] ^ in2[14];
    assign G[218] = in[13] & in2[13];
    assign P[218] = in[13] ^ in2[13];
    assign G[219] = in[12] & in2[12];
    assign P[219] = in[12] ^ in2[12];
    assign G[220] = in[11] & in2[11];
    assign P[220] = in[11] ^ in2[11];
    assign G[221] = in[10] & in2[10];
    assign P[221] = in[10] ^ in2[10];
    assign G[222] = in[9] & in2[9];
    assign P[222] = in[9] ^ in2[9];
    assign G[223] = in[8] & in2[8];
    assign P[223] = in[8] ^ in2[8];
    assign G[224] = in[7] & in2[7];
    assign P[224] = in[7] ^ in2[7];
    assign G[225] = in[6] & in2[6];
    assign P[225] = in[6] ^ in2[6];
    assign G[226] = in[5] & in2[5];
    assign P[226] = in[5] ^ in2[5];
    assign G[227] = in[4] & in2[4];
    assign P[227] = in[4] ^ in2[4];
    assign G[228] = in[3] & in2[3];
    assign P[228] = in[3] ^ in2[3];
    assign G[229] = in[2] & in2[2];
    assign P[229] = in[2] ^ in2[2];
    assign G[230] = in[1] & in2[1];
    assign P[230] = in[1] ^ in2[1];
    assign G[231] = in[0] & in2[0];
    assign P[231] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign C[231] = G[230] | (P[230] & C[230]);
    assign cout = G[231] | (P[231] & C[231]);
    assign sum = P ^ C;
endmodule

module CLA231(output [230:0] sum, output cout, input [230:0] in1, input [230:0] in2;

    wire[230:0] G;
    wire[230:0] C;
    wire[230:0] P;

    assign G[0] = in[230] & in2[230];
    assign P[0] = in[230] ^ in2[230];
    assign G[1] = in[229] & in2[229];
    assign P[1] = in[229] ^ in2[229];
    assign G[2] = in[228] & in2[228];
    assign P[2] = in[228] ^ in2[228];
    assign G[3] = in[227] & in2[227];
    assign P[3] = in[227] ^ in2[227];
    assign G[4] = in[226] & in2[226];
    assign P[4] = in[226] ^ in2[226];
    assign G[5] = in[225] & in2[225];
    assign P[5] = in[225] ^ in2[225];
    assign G[6] = in[224] & in2[224];
    assign P[6] = in[224] ^ in2[224];
    assign G[7] = in[223] & in2[223];
    assign P[7] = in[223] ^ in2[223];
    assign G[8] = in[222] & in2[222];
    assign P[8] = in[222] ^ in2[222];
    assign G[9] = in[221] & in2[221];
    assign P[9] = in[221] ^ in2[221];
    assign G[10] = in[220] & in2[220];
    assign P[10] = in[220] ^ in2[220];
    assign G[11] = in[219] & in2[219];
    assign P[11] = in[219] ^ in2[219];
    assign G[12] = in[218] & in2[218];
    assign P[12] = in[218] ^ in2[218];
    assign G[13] = in[217] & in2[217];
    assign P[13] = in[217] ^ in2[217];
    assign G[14] = in[216] & in2[216];
    assign P[14] = in[216] ^ in2[216];
    assign G[15] = in[215] & in2[215];
    assign P[15] = in[215] ^ in2[215];
    assign G[16] = in[214] & in2[214];
    assign P[16] = in[214] ^ in2[214];
    assign G[17] = in[213] & in2[213];
    assign P[17] = in[213] ^ in2[213];
    assign G[18] = in[212] & in2[212];
    assign P[18] = in[212] ^ in2[212];
    assign G[19] = in[211] & in2[211];
    assign P[19] = in[211] ^ in2[211];
    assign G[20] = in[210] & in2[210];
    assign P[20] = in[210] ^ in2[210];
    assign G[21] = in[209] & in2[209];
    assign P[21] = in[209] ^ in2[209];
    assign G[22] = in[208] & in2[208];
    assign P[22] = in[208] ^ in2[208];
    assign G[23] = in[207] & in2[207];
    assign P[23] = in[207] ^ in2[207];
    assign G[24] = in[206] & in2[206];
    assign P[24] = in[206] ^ in2[206];
    assign G[25] = in[205] & in2[205];
    assign P[25] = in[205] ^ in2[205];
    assign G[26] = in[204] & in2[204];
    assign P[26] = in[204] ^ in2[204];
    assign G[27] = in[203] & in2[203];
    assign P[27] = in[203] ^ in2[203];
    assign G[28] = in[202] & in2[202];
    assign P[28] = in[202] ^ in2[202];
    assign G[29] = in[201] & in2[201];
    assign P[29] = in[201] ^ in2[201];
    assign G[30] = in[200] & in2[200];
    assign P[30] = in[200] ^ in2[200];
    assign G[31] = in[199] & in2[199];
    assign P[31] = in[199] ^ in2[199];
    assign G[32] = in[198] & in2[198];
    assign P[32] = in[198] ^ in2[198];
    assign G[33] = in[197] & in2[197];
    assign P[33] = in[197] ^ in2[197];
    assign G[34] = in[196] & in2[196];
    assign P[34] = in[196] ^ in2[196];
    assign G[35] = in[195] & in2[195];
    assign P[35] = in[195] ^ in2[195];
    assign G[36] = in[194] & in2[194];
    assign P[36] = in[194] ^ in2[194];
    assign G[37] = in[193] & in2[193];
    assign P[37] = in[193] ^ in2[193];
    assign G[38] = in[192] & in2[192];
    assign P[38] = in[192] ^ in2[192];
    assign G[39] = in[191] & in2[191];
    assign P[39] = in[191] ^ in2[191];
    assign G[40] = in[190] & in2[190];
    assign P[40] = in[190] ^ in2[190];
    assign G[41] = in[189] & in2[189];
    assign P[41] = in[189] ^ in2[189];
    assign G[42] = in[188] & in2[188];
    assign P[42] = in[188] ^ in2[188];
    assign G[43] = in[187] & in2[187];
    assign P[43] = in[187] ^ in2[187];
    assign G[44] = in[186] & in2[186];
    assign P[44] = in[186] ^ in2[186];
    assign G[45] = in[185] & in2[185];
    assign P[45] = in[185] ^ in2[185];
    assign G[46] = in[184] & in2[184];
    assign P[46] = in[184] ^ in2[184];
    assign G[47] = in[183] & in2[183];
    assign P[47] = in[183] ^ in2[183];
    assign G[48] = in[182] & in2[182];
    assign P[48] = in[182] ^ in2[182];
    assign G[49] = in[181] & in2[181];
    assign P[49] = in[181] ^ in2[181];
    assign G[50] = in[180] & in2[180];
    assign P[50] = in[180] ^ in2[180];
    assign G[51] = in[179] & in2[179];
    assign P[51] = in[179] ^ in2[179];
    assign G[52] = in[178] & in2[178];
    assign P[52] = in[178] ^ in2[178];
    assign G[53] = in[177] & in2[177];
    assign P[53] = in[177] ^ in2[177];
    assign G[54] = in[176] & in2[176];
    assign P[54] = in[176] ^ in2[176];
    assign G[55] = in[175] & in2[175];
    assign P[55] = in[175] ^ in2[175];
    assign G[56] = in[174] & in2[174];
    assign P[56] = in[174] ^ in2[174];
    assign G[57] = in[173] & in2[173];
    assign P[57] = in[173] ^ in2[173];
    assign G[58] = in[172] & in2[172];
    assign P[58] = in[172] ^ in2[172];
    assign G[59] = in[171] & in2[171];
    assign P[59] = in[171] ^ in2[171];
    assign G[60] = in[170] & in2[170];
    assign P[60] = in[170] ^ in2[170];
    assign G[61] = in[169] & in2[169];
    assign P[61] = in[169] ^ in2[169];
    assign G[62] = in[168] & in2[168];
    assign P[62] = in[168] ^ in2[168];
    assign G[63] = in[167] & in2[167];
    assign P[63] = in[167] ^ in2[167];
    assign G[64] = in[166] & in2[166];
    assign P[64] = in[166] ^ in2[166];
    assign G[65] = in[165] & in2[165];
    assign P[65] = in[165] ^ in2[165];
    assign G[66] = in[164] & in2[164];
    assign P[66] = in[164] ^ in2[164];
    assign G[67] = in[163] & in2[163];
    assign P[67] = in[163] ^ in2[163];
    assign G[68] = in[162] & in2[162];
    assign P[68] = in[162] ^ in2[162];
    assign G[69] = in[161] & in2[161];
    assign P[69] = in[161] ^ in2[161];
    assign G[70] = in[160] & in2[160];
    assign P[70] = in[160] ^ in2[160];
    assign G[71] = in[159] & in2[159];
    assign P[71] = in[159] ^ in2[159];
    assign G[72] = in[158] & in2[158];
    assign P[72] = in[158] ^ in2[158];
    assign G[73] = in[157] & in2[157];
    assign P[73] = in[157] ^ in2[157];
    assign G[74] = in[156] & in2[156];
    assign P[74] = in[156] ^ in2[156];
    assign G[75] = in[155] & in2[155];
    assign P[75] = in[155] ^ in2[155];
    assign G[76] = in[154] & in2[154];
    assign P[76] = in[154] ^ in2[154];
    assign G[77] = in[153] & in2[153];
    assign P[77] = in[153] ^ in2[153];
    assign G[78] = in[152] & in2[152];
    assign P[78] = in[152] ^ in2[152];
    assign G[79] = in[151] & in2[151];
    assign P[79] = in[151] ^ in2[151];
    assign G[80] = in[150] & in2[150];
    assign P[80] = in[150] ^ in2[150];
    assign G[81] = in[149] & in2[149];
    assign P[81] = in[149] ^ in2[149];
    assign G[82] = in[148] & in2[148];
    assign P[82] = in[148] ^ in2[148];
    assign G[83] = in[147] & in2[147];
    assign P[83] = in[147] ^ in2[147];
    assign G[84] = in[146] & in2[146];
    assign P[84] = in[146] ^ in2[146];
    assign G[85] = in[145] & in2[145];
    assign P[85] = in[145] ^ in2[145];
    assign G[86] = in[144] & in2[144];
    assign P[86] = in[144] ^ in2[144];
    assign G[87] = in[143] & in2[143];
    assign P[87] = in[143] ^ in2[143];
    assign G[88] = in[142] & in2[142];
    assign P[88] = in[142] ^ in2[142];
    assign G[89] = in[141] & in2[141];
    assign P[89] = in[141] ^ in2[141];
    assign G[90] = in[140] & in2[140];
    assign P[90] = in[140] ^ in2[140];
    assign G[91] = in[139] & in2[139];
    assign P[91] = in[139] ^ in2[139];
    assign G[92] = in[138] & in2[138];
    assign P[92] = in[138] ^ in2[138];
    assign G[93] = in[137] & in2[137];
    assign P[93] = in[137] ^ in2[137];
    assign G[94] = in[136] & in2[136];
    assign P[94] = in[136] ^ in2[136];
    assign G[95] = in[135] & in2[135];
    assign P[95] = in[135] ^ in2[135];
    assign G[96] = in[134] & in2[134];
    assign P[96] = in[134] ^ in2[134];
    assign G[97] = in[133] & in2[133];
    assign P[97] = in[133] ^ in2[133];
    assign G[98] = in[132] & in2[132];
    assign P[98] = in[132] ^ in2[132];
    assign G[99] = in[131] & in2[131];
    assign P[99] = in[131] ^ in2[131];
    assign G[100] = in[130] & in2[130];
    assign P[100] = in[130] ^ in2[130];
    assign G[101] = in[129] & in2[129];
    assign P[101] = in[129] ^ in2[129];
    assign G[102] = in[128] & in2[128];
    assign P[102] = in[128] ^ in2[128];
    assign G[103] = in[127] & in2[127];
    assign P[103] = in[127] ^ in2[127];
    assign G[104] = in[126] & in2[126];
    assign P[104] = in[126] ^ in2[126];
    assign G[105] = in[125] & in2[125];
    assign P[105] = in[125] ^ in2[125];
    assign G[106] = in[124] & in2[124];
    assign P[106] = in[124] ^ in2[124];
    assign G[107] = in[123] & in2[123];
    assign P[107] = in[123] ^ in2[123];
    assign G[108] = in[122] & in2[122];
    assign P[108] = in[122] ^ in2[122];
    assign G[109] = in[121] & in2[121];
    assign P[109] = in[121] ^ in2[121];
    assign G[110] = in[120] & in2[120];
    assign P[110] = in[120] ^ in2[120];
    assign G[111] = in[119] & in2[119];
    assign P[111] = in[119] ^ in2[119];
    assign G[112] = in[118] & in2[118];
    assign P[112] = in[118] ^ in2[118];
    assign G[113] = in[117] & in2[117];
    assign P[113] = in[117] ^ in2[117];
    assign G[114] = in[116] & in2[116];
    assign P[114] = in[116] ^ in2[116];
    assign G[115] = in[115] & in2[115];
    assign P[115] = in[115] ^ in2[115];
    assign G[116] = in[114] & in2[114];
    assign P[116] = in[114] ^ in2[114];
    assign G[117] = in[113] & in2[113];
    assign P[117] = in[113] ^ in2[113];
    assign G[118] = in[112] & in2[112];
    assign P[118] = in[112] ^ in2[112];
    assign G[119] = in[111] & in2[111];
    assign P[119] = in[111] ^ in2[111];
    assign G[120] = in[110] & in2[110];
    assign P[120] = in[110] ^ in2[110];
    assign G[121] = in[109] & in2[109];
    assign P[121] = in[109] ^ in2[109];
    assign G[122] = in[108] & in2[108];
    assign P[122] = in[108] ^ in2[108];
    assign G[123] = in[107] & in2[107];
    assign P[123] = in[107] ^ in2[107];
    assign G[124] = in[106] & in2[106];
    assign P[124] = in[106] ^ in2[106];
    assign G[125] = in[105] & in2[105];
    assign P[125] = in[105] ^ in2[105];
    assign G[126] = in[104] & in2[104];
    assign P[126] = in[104] ^ in2[104];
    assign G[127] = in[103] & in2[103];
    assign P[127] = in[103] ^ in2[103];
    assign G[128] = in[102] & in2[102];
    assign P[128] = in[102] ^ in2[102];
    assign G[129] = in[101] & in2[101];
    assign P[129] = in[101] ^ in2[101];
    assign G[130] = in[100] & in2[100];
    assign P[130] = in[100] ^ in2[100];
    assign G[131] = in[99] & in2[99];
    assign P[131] = in[99] ^ in2[99];
    assign G[132] = in[98] & in2[98];
    assign P[132] = in[98] ^ in2[98];
    assign G[133] = in[97] & in2[97];
    assign P[133] = in[97] ^ in2[97];
    assign G[134] = in[96] & in2[96];
    assign P[134] = in[96] ^ in2[96];
    assign G[135] = in[95] & in2[95];
    assign P[135] = in[95] ^ in2[95];
    assign G[136] = in[94] & in2[94];
    assign P[136] = in[94] ^ in2[94];
    assign G[137] = in[93] & in2[93];
    assign P[137] = in[93] ^ in2[93];
    assign G[138] = in[92] & in2[92];
    assign P[138] = in[92] ^ in2[92];
    assign G[139] = in[91] & in2[91];
    assign P[139] = in[91] ^ in2[91];
    assign G[140] = in[90] & in2[90];
    assign P[140] = in[90] ^ in2[90];
    assign G[141] = in[89] & in2[89];
    assign P[141] = in[89] ^ in2[89];
    assign G[142] = in[88] & in2[88];
    assign P[142] = in[88] ^ in2[88];
    assign G[143] = in[87] & in2[87];
    assign P[143] = in[87] ^ in2[87];
    assign G[144] = in[86] & in2[86];
    assign P[144] = in[86] ^ in2[86];
    assign G[145] = in[85] & in2[85];
    assign P[145] = in[85] ^ in2[85];
    assign G[146] = in[84] & in2[84];
    assign P[146] = in[84] ^ in2[84];
    assign G[147] = in[83] & in2[83];
    assign P[147] = in[83] ^ in2[83];
    assign G[148] = in[82] & in2[82];
    assign P[148] = in[82] ^ in2[82];
    assign G[149] = in[81] & in2[81];
    assign P[149] = in[81] ^ in2[81];
    assign G[150] = in[80] & in2[80];
    assign P[150] = in[80] ^ in2[80];
    assign G[151] = in[79] & in2[79];
    assign P[151] = in[79] ^ in2[79];
    assign G[152] = in[78] & in2[78];
    assign P[152] = in[78] ^ in2[78];
    assign G[153] = in[77] & in2[77];
    assign P[153] = in[77] ^ in2[77];
    assign G[154] = in[76] & in2[76];
    assign P[154] = in[76] ^ in2[76];
    assign G[155] = in[75] & in2[75];
    assign P[155] = in[75] ^ in2[75];
    assign G[156] = in[74] & in2[74];
    assign P[156] = in[74] ^ in2[74];
    assign G[157] = in[73] & in2[73];
    assign P[157] = in[73] ^ in2[73];
    assign G[158] = in[72] & in2[72];
    assign P[158] = in[72] ^ in2[72];
    assign G[159] = in[71] & in2[71];
    assign P[159] = in[71] ^ in2[71];
    assign G[160] = in[70] & in2[70];
    assign P[160] = in[70] ^ in2[70];
    assign G[161] = in[69] & in2[69];
    assign P[161] = in[69] ^ in2[69];
    assign G[162] = in[68] & in2[68];
    assign P[162] = in[68] ^ in2[68];
    assign G[163] = in[67] & in2[67];
    assign P[163] = in[67] ^ in2[67];
    assign G[164] = in[66] & in2[66];
    assign P[164] = in[66] ^ in2[66];
    assign G[165] = in[65] & in2[65];
    assign P[165] = in[65] ^ in2[65];
    assign G[166] = in[64] & in2[64];
    assign P[166] = in[64] ^ in2[64];
    assign G[167] = in[63] & in2[63];
    assign P[167] = in[63] ^ in2[63];
    assign G[168] = in[62] & in2[62];
    assign P[168] = in[62] ^ in2[62];
    assign G[169] = in[61] & in2[61];
    assign P[169] = in[61] ^ in2[61];
    assign G[170] = in[60] & in2[60];
    assign P[170] = in[60] ^ in2[60];
    assign G[171] = in[59] & in2[59];
    assign P[171] = in[59] ^ in2[59];
    assign G[172] = in[58] & in2[58];
    assign P[172] = in[58] ^ in2[58];
    assign G[173] = in[57] & in2[57];
    assign P[173] = in[57] ^ in2[57];
    assign G[174] = in[56] & in2[56];
    assign P[174] = in[56] ^ in2[56];
    assign G[175] = in[55] & in2[55];
    assign P[175] = in[55] ^ in2[55];
    assign G[176] = in[54] & in2[54];
    assign P[176] = in[54] ^ in2[54];
    assign G[177] = in[53] & in2[53];
    assign P[177] = in[53] ^ in2[53];
    assign G[178] = in[52] & in2[52];
    assign P[178] = in[52] ^ in2[52];
    assign G[179] = in[51] & in2[51];
    assign P[179] = in[51] ^ in2[51];
    assign G[180] = in[50] & in2[50];
    assign P[180] = in[50] ^ in2[50];
    assign G[181] = in[49] & in2[49];
    assign P[181] = in[49] ^ in2[49];
    assign G[182] = in[48] & in2[48];
    assign P[182] = in[48] ^ in2[48];
    assign G[183] = in[47] & in2[47];
    assign P[183] = in[47] ^ in2[47];
    assign G[184] = in[46] & in2[46];
    assign P[184] = in[46] ^ in2[46];
    assign G[185] = in[45] & in2[45];
    assign P[185] = in[45] ^ in2[45];
    assign G[186] = in[44] & in2[44];
    assign P[186] = in[44] ^ in2[44];
    assign G[187] = in[43] & in2[43];
    assign P[187] = in[43] ^ in2[43];
    assign G[188] = in[42] & in2[42];
    assign P[188] = in[42] ^ in2[42];
    assign G[189] = in[41] & in2[41];
    assign P[189] = in[41] ^ in2[41];
    assign G[190] = in[40] & in2[40];
    assign P[190] = in[40] ^ in2[40];
    assign G[191] = in[39] & in2[39];
    assign P[191] = in[39] ^ in2[39];
    assign G[192] = in[38] & in2[38];
    assign P[192] = in[38] ^ in2[38];
    assign G[193] = in[37] & in2[37];
    assign P[193] = in[37] ^ in2[37];
    assign G[194] = in[36] & in2[36];
    assign P[194] = in[36] ^ in2[36];
    assign G[195] = in[35] & in2[35];
    assign P[195] = in[35] ^ in2[35];
    assign G[196] = in[34] & in2[34];
    assign P[196] = in[34] ^ in2[34];
    assign G[197] = in[33] & in2[33];
    assign P[197] = in[33] ^ in2[33];
    assign G[198] = in[32] & in2[32];
    assign P[198] = in[32] ^ in2[32];
    assign G[199] = in[31] & in2[31];
    assign P[199] = in[31] ^ in2[31];
    assign G[200] = in[30] & in2[30];
    assign P[200] = in[30] ^ in2[30];
    assign G[201] = in[29] & in2[29];
    assign P[201] = in[29] ^ in2[29];
    assign G[202] = in[28] & in2[28];
    assign P[202] = in[28] ^ in2[28];
    assign G[203] = in[27] & in2[27];
    assign P[203] = in[27] ^ in2[27];
    assign G[204] = in[26] & in2[26];
    assign P[204] = in[26] ^ in2[26];
    assign G[205] = in[25] & in2[25];
    assign P[205] = in[25] ^ in2[25];
    assign G[206] = in[24] & in2[24];
    assign P[206] = in[24] ^ in2[24];
    assign G[207] = in[23] & in2[23];
    assign P[207] = in[23] ^ in2[23];
    assign G[208] = in[22] & in2[22];
    assign P[208] = in[22] ^ in2[22];
    assign G[209] = in[21] & in2[21];
    assign P[209] = in[21] ^ in2[21];
    assign G[210] = in[20] & in2[20];
    assign P[210] = in[20] ^ in2[20];
    assign G[211] = in[19] & in2[19];
    assign P[211] = in[19] ^ in2[19];
    assign G[212] = in[18] & in2[18];
    assign P[212] = in[18] ^ in2[18];
    assign G[213] = in[17] & in2[17];
    assign P[213] = in[17] ^ in2[17];
    assign G[214] = in[16] & in2[16];
    assign P[214] = in[16] ^ in2[16];
    assign G[215] = in[15] & in2[15];
    assign P[215] = in[15] ^ in2[15];
    assign G[216] = in[14] & in2[14];
    assign P[216] = in[14] ^ in2[14];
    assign G[217] = in[13] & in2[13];
    assign P[217] = in[13] ^ in2[13];
    assign G[218] = in[12] & in2[12];
    assign P[218] = in[12] ^ in2[12];
    assign G[219] = in[11] & in2[11];
    assign P[219] = in[11] ^ in2[11];
    assign G[220] = in[10] & in2[10];
    assign P[220] = in[10] ^ in2[10];
    assign G[221] = in[9] & in2[9];
    assign P[221] = in[9] ^ in2[9];
    assign G[222] = in[8] & in2[8];
    assign P[222] = in[8] ^ in2[8];
    assign G[223] = in[7] & in2[7];
    assign P[223] = in[7] ^ in2[7];
    assign G[224] = in[6] & in2[6];
    assign P[224] = in[6] ^ in2[6];
    assign G[225] = in[5] & in2[5];
    assign P[225] = in[5] ^ in2[5];
    assign G[226] = in[4] & in2[4];
    assign P[226] = in[4] ^ in2[4];
    assign G[227] = in[3] & in2[3];
    assign P[227] = in[3] ^ in2[3];
    assign G[228] = in[2] & in2[2];
    assign P[228] = in[2] ^ in2[2];
    assign G[229] = in[1] & in2[1];
    assign P[229] = in[1] ^ in2[1];
    assign G[230] = in[0] & in2[0];
    assign P[230] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign C[230] = G[229] | (P[229] & C[229]);
    assign cout = G[230] | (P[230] & C[230]);
    assign sum = P ^ C;
endmodule

module CLA230(output [229:0] sum, output cout, input [229:0] in1, input [229:0] in2;

    wire[229:0] G;
    wire[229:0] C;
    wire[229:0] P;

    assign G[0] = in[229] & in2[229];
    assign P[0] = in[229] ^ in2[229];
    assign G[1] = in[228] & in2[228];
    assign P[1] = in[228] ^ in2[228];
    assign G[2] = in[227] & in2[227];
    assign P[2] = in[227] ^ in2[227];
    assign G[3] = in[226] & in2[226];
    assign P[3] = in[226] ^ in2[226];
    assign G[4] = in[225] & in2[225];
    assign P[4] = in[225] ^ in2[225];
    assign G[5] = in[224] & in2[224];
    assign P[5] = in[224] ^ in2[224];
    assign G[6] = in[223] & in2[223];
    assign P[6] = in[223] ^ in2[223];
    assign G[7] = in[222] & in2[222];
    assign P[7] = in[222] ^ in2[222];
    assign G[8] = in[221] & in2[221];
    assign P[8] = in[221] ^ in2[221];
    assign G[9] = in[220] & in2[220];
    assign P[9] = in[220] ^ in2[220];
    assign G[10] = in[219] & in2[219];
    assign P[10] = in[219] ^ in2[219];
    assign G[11] = in[218] & in2[218];
    assign P[11] = in[218] ^ in2[218];
    assign G[12] = in[217] & in2[217];
    assign P[12] = in[217] ^ in2[217];
    assign G[13] = in[216] & in2[216];
    assign P[13] = in[216] ^ in2[216];
    assign G[14] = in[215] & in2[215];
    assign P[14] = in[215] ^ in2[215];
    assign G[15] = in[214] & in2[214];
    assign P[15] = in[214] ^ in2[214];
    assign G[16] = in[213] & in2[213];
    assign P[16] = in[213] ^ in2[213];
    assign G[17] = in[212] & in2[212];
    assign P[17] = in[212] ^ in2[212];
    assign G[18] = in[211] & in2[211];
    assign P[18] = in[211] ^ in2[211];
    assign G[19] = in[210] & in2[210];
    assign P[19] = in[210] ^ in2[210];
    assign G[20] = in[209] & in2[209];
    assign P[20] = in[209] ^ in2[209];
    assign G[21] = in[208] & in2[208];
    assign P[21] = in[208] ^ in2[208];
    assign G[22] = in[207] & in2[207];
    assign P[22] = in[207] ^ in2[207];
    assign G[23] = in[206] & in2[206];
    assign P[23] = in[206] ^ in2[206];
    assign G[24] = in[205] & in2[205];
    assign P[24] = in[205] ^ in2[205];
    assign G[25] = in[204] & in2[204];
    assign P[25] = in[204] ^ in2[204];
    assign G[26] = in[203] & in2[203];
    assign P[26] = in[203] ^ in2[203];
    assign G[27] = in[202] & in2[202];
    assign P[27] = in[202] ^ in2[202];
    assign G[28] = in[201] & in2[201];
    assign P[28] = in[201] ^ in2[201];
    assign G[29] = in[200] & in2[200];
    assign P[29] = in[200] ^ in2[200];
    assign G[30] = in[199] & in2[199];
    assign P[30] = in[199] ^ in2[199];
    assign G[31] = in[198] & in2[198];
    assign P[31] = in[198] ^ in2[198];
    assign G[32] = in[197] & in2[197];
    assign P[32] = in[197] ^ in2[197];
    assign G[33] = in[196] & in2[196];
    assign P[33] = in[196] ^ in2[196];
    assign G[34] = in[195] & in2[195];
    assign P[34] = in[195] ^ in2[195];
    assign G[35] = in[194] & in2[194];
    assign P[35] = in[194] ^ in2[194];
    assign G[36] = in[193] & in2[193];
    assign P[36] = in[193] ^ in2[193];
    assign G[37] = in[192] & in2[192];
    assign P[37] = in[192] ^ in2[192];
    assign G[38] = in[191] & in2[191];
    assign P[38] = in[191] ^ in2[191];
    assign G[39] = in[190] & in2[190];
    assign P[39] = in[190] ^ in2[190];
    assign G[40] = in[189] & in2[189];
    assign P[40] = in[189] ^ in2[189];
    assign G[41] = in[188] & in2[188];
    assign P[41] = in[188] ^ in2[188];
    assign G[42] = in[187] & in2[187];
    assign P[42] = in[187] ^ in2[187];
    assign G[43] = in[186] & in2[186];
    assign P[43] = in[186] ^ in2[186];
    assign G[44] = in[185] & in2[185];
    assign P[44] = in[185] ^ in2[185];
    assign G[45] = in[184] & in2[184];
    assign P[45] = in[184] ^ in2[184];
    assign G[46] = in[183] & in2[183];
    assign P[46] = in[183] ^ in2[183];
    assign G[47] = in[182] & in2[182];
    assign P[47] = in[182] ^ in2[182];
    assign G[48] = in[181] & in2[181];
    assign P[48] = in[181] ^ in2[181];
    assign G[49] = in[180] & in2[180];
    assign P[49] = in[180] ^ in2[180];
    assign G[50] = in[179] & in2[179];
    assign P[50] = in[179] ^ in2[179];
    assign G[51] = in[178] & in2[178];
    assign P[51] = in[178] ^ in2[178];
    assign G[52] = in[177] & in2[177];
    assign P[52] = in[177] ^ in2[177];
    assign G[53] = in[176] & in2[176];
    assign P[53] = in[176] ^ in2[176];
    assign G[54] = in[175] & in2[175];
    assign P[54] = in[175] ^ in2[175];
    assign G[55] = in[174] & in2[174];
    assign P[55] = in[174] ^ in2[174];
    assign G[56] = in[173] & in2[173];
    assign P[56] = in[173] ^ in2[173];
    assign G[57] = in[172] & in2[172];
    assign P[57] = in[172] ^ in2[172];
    assign G[58] = in[171] & in2[171];
    assign P[58] = in[171] ^ in2[171];
    assign G[59] = in[170] & in2[170];
    assign P[59] = in[170] ^ in2[170];
    assign G[60] = in[169] & in2[169];
    assign P[60] = in[169] ^ in2[169];
    assign G[61] = in[168] & in2[168];
    assign P[61] = in[168] ^ in2[168];
    assign G[62] = in[167] & in2[167];
    assign P[62] = in[167] ^ in2[167];
    assign G[63] = in[166] & in2[166];
    assign P[63] = in[166] ^ in2[166];
    assign G[64] = in[165] & in2[165];
    assign P[64] = in[165] ^ in2[165];
    assign G[65] = in[164] & in2[164];
    assign P[65] = in[164] ^ in2[164];
    assign G[66] = in[163] & in2[163];
    assign P[66] = in[163] ^ in2[163];
    assign G[67] = in[162] & in2[162];
    assign P[67] = in[162] ^ in2[162];
    assign G[68] = in[161] & in2[161];
    assign P[68] = in[161] ^ in2[161];
    assign G[69] = in[160] & in2[160];
    assign P[69] = in[160] ^ in2[160];
    assign G[70] = in[159] & in2[159];
    assign P[70] = in[159] ^ in2[159];
    assign G[71] = in[158] & in2[158];
    assign P[71] = in[158] ^ in2[158];
    assign G[72] = in[157] & in2[157];
    assign P[72] = in[157] ^ in2[157];
    assign G[73] = in[156] & in2[156];
    assign P[73] = in[156] ^ in2[156];
    assign G[74] = in[155] & in2[155];
    assign P[74] = in[155] ^ in2[155];
    assign G[75] = in[154] & in2[154];
    assign P[75] = in[154] ^ in2[154];
    assign G[76] = in[153] & in2[153];
    assign P[76] = in[153] ^ in2[153];
    assign G[77] = in[152] & in2[152];
    assign P[77] = in[152] ^ in2[152];
    assign G[78] = in[151] & in2[151];
    assign P[78] = in[151] ^ in2[151];
    assign G[79] = in[150] & in2[150];
    assign P[79] = in[150] ^ in2[150];
    assign G[80] = in[149] & in2[149];
    assign P[80] = in[149] ^ in2[149];
    assign G[81] = in[148] & in2[148];
    assign P[81] = in[148] ^ in2[148];
    assign G[82] = in[147] & in2[147];
    assign P[82] = in[147] ^ in2[147];
    assign G[83] = in[146] & in2[146];
    assign P[83] = in[146] ^ in2[146];
    assign G[84] = in[145] & in2[145];
    assign P[84] = in[145] ^ in2[145];
    assign G[85] = in[144] & in2[144];
    assign P[85] = in[144] ^ in2[144];
    assign G[86] = in[143] & in2[143];
    assign P[86] = in[143] ^ in2[143];
    assign G[87] = in[142] & in2[142];
    assign P[87] = in[142] ^ in2[142];
    assign G[88] = in[141] & in2[141];
    assign P[88] = in[141] ^ in2[141];
    assign G[89] = in[140] & in2[140];
    assign P[89] = in[140] ^ in2[140];
    assign G[90] = in[139] & in2[139];
    assign P[90] = in[139] ^ in2[139];
    assign G[91] = in[138] & in2[138];
    assign P[91] = in[138] ^ in2[138];
    assign G[92] = in[137] & in2[137];
    assign P[92] = in[137] ^ in2[137];
    assign G[93] = in[136] & in2[136];
    assign P[93] = in[136] ^ in2[136];
    assign G[94] = in[135] & in2[135];
    assign P[94] = in[135] ^ in2[135];
    assign G[95] = in[134] & in2[134];
    assign P[95] = in[134] ^ in2[134];
    assign G[96] = in[133] & in2[133];
    assign P[96] = in[133] ^ in2[133];
    assign G[97] = in[132] & in2[132];
    assign P[97] = in[132] ^ in2[132];
    assign G[98] = in[131] & in2[131];
    assign P[98] = in[131] ^ in2[131];
    assign G[99] = in[130] & in2[130];
    assign P[99] = in[130] ^ in2[130];
    assign G[100] = in[129] & in2[129];
    assign P[100] = in[129] ^ in2[129];
    assign G[101] = in[128] & in2[128];
    assign P[101] = in[128] ^ in2[128];
    assign G[102] = in[127] & in2[127];
    assign P[102] = in[127] ^ in2[127];
    assign G[103] = in[126] & in2[126];
    assign P[103] = in[126] ^ in2[126];
    assign G[104] = in[125] & in2[125];
    assign P[104] = in[125] ^ in2[125];
    assign G[105] = in[124] & in2[124];
    assign P[105] = in[124] ^ in2[124];
    assign G[106] = in[123] & in2[123];
    assign P[106] = in[123] ^ in2[123];
    assign G[107] = in[122] & in2[122];
    assign P[107] = in[122] ^ in2[122];
    assign G[108] = in[121] & in2[121];
    assign P[108] = in[121] ^ in2[121];
    assign G[109] = in[120] & in2[120];
    assign P[109] = in[120] ^ in2[120];
    assign G[110] = in[119] & in2[119];
    assign P[110] = in[119] ^ in2[119];
    assign G[111] = in[118] & in2[118];
    assign P[111] = in[118] ^ in2[118];
    assign G[112] = in[117] & in2[117];
    assign P[112] = in[117] ^ in2[117];
    assign G[113] = in[116] & in2[116];
    assign P[113] = in[116] ^ in2[116];
    assign G[114] = in[115] & in2[115];
    assign P[114] = in[115] ^ in2[115];
    assign G[115] = in[114] & in2[114];
    assign P[115] = in[114] ^ in2[114];
    assign G[116] = in[113] & in2[113];
    assign P[116] = in[113] ^ in2[113];
    assign G[117] = in[112] & in2[112];
    assign P[117] = in[112] ^ in2[112];
    assign G[118] = in[111] & in2[111];
    assign P[118] = in[111] ^ in2[111];
    assign G[119] = in[110] & in2[110];
    assign P[119] = in[110] ^ in2[110];
    assign G[120] = in[109] & in2[109];
    assign P[120] = in[109] ^ in2[109];
    assign G[121] = in[108] & in2[108];
    assign P[121] = in[108] ^ in2[108];
    assign G[122] = in[107] & in2[107];
    assign P[122] = in[107] ^ in2[107];
    assign G[123] = in[106] & in2[106];
    assign P[123] = in[106] ^ in2[106];
    assign G[124] = in[105] & in2[105];
    assign P[124] = in[105] ^ in2[105];
    assign G[125] = in[104] & in2[104];
    assign P[125] = in[104] ^ in2[104];
    assign G[126] = in[103] & in2[103];
    assign P[126] = in[103] ^ in2[103];
    assign G[127] = in[102] & in2[102];
    assign P[127] = in[102] ^ in2[102];
    assign G[128] = in[101] & in2[101];
    assign P[128] = in[101] ^ in2[101];
    assign G[129] = in[100] & in2[100];
    assign P[129] = in[100] ^ in2[100];
    assign G[130] = in[99] & in2[99];
    assign P[130] = in[99] ^ in2[99];
    assign G[131] = in[98] & in2[98];
    assign P[131] = in[98] ^ in2[98];
    assign G[132] = in[97] & in2[97];
    assign P[132] = in[97] ^ in2[97];
    assign G[133] = in[96] & in2[96];
    assign P[133] = in[96] ^ in2[96];
    assign G[134] = in[95] & in2[95];
    assign P[134] = in[95] ^ in2[95];
    assign G[135] = in[94] & in2[94];
    assign P[135] = in[94] ^ in2[94];
    assign G[136] = in[93] & in2[93];
    assign P[136] = in[93] ^ in2[93];
    assign G[137] = in[92] & in2[92];
    assign P[137] = in[92] ^ in2[92];
    assign G[138] = in[91] & in2[91];
    assign P[138] = in[91] ^ in2[91];
    assign G[139] = in[90] & in2[90];
    assign P[139] = in[90] ^ in2[90];
    assign G[140] = in[89] & in2[89];
    assign P[140] = in[89] ^ in2[89];
    assign G[141] = in[88] & in2[88];
    assign P[141] = in[88] ^ in2[88];
    assign G[142] = in[87] & in2[87];
    assign P[142] = in[87] ^ in2[87];
    assign G[143] = in[86] & in2[86];
    assign P[143] = in[86] ^ in2[86];
    assign G[144] = in[85] & in2[85];
    assign P[144] = in[85] ^ in2[85];
    assign G[145] = in[84] & in2[84];
    assign P[145] = in[84] ^ in2[84];
    assign G[146] = in[83] & in2[83];
    assign P[146] = in[83] ^ in2[83];
    assign G[147] = in[82] & in2[82];
    assign P[147] = in[82] ^ in2[82];
    assign G[148] = in[81] & in2[81];
    assign P[148] = in[81] ^ in2[81];
    assign G[149] = in[80] & in2[80];
    assign P[149] = in[80] ^ in2[80];
    assign G[150] = in[79] & in2[79];
    assign P[150] = in[79] ^ in2[79];
    assign G[151] = in[78] & in2[78];
    assign P[151] = in[78] ^ in2[78];
    assign G[152] = in[77] & in2[77];
    assign P[152] = in[77] ^ in2[77];
    assign G[153] = in[76] & in2[76];
    assign P[153] = in[76] ^ in2[76];
    assign G[154] = in[75] & in2[75];
    assign P[154] = in[75] ^ in2[75];
    assign G[155] = in[74] & in2[74];
    assign P[155] = in[74] ^ in2[74];
    assign G[156] = in[73] & in2[73];
    assign P[156] = in[73] ^ in2[73];
    assign G[157] = in[72] & in2[72];
    assign P[157] = in[72] ^ in2[72];
    assign G[158] = in[71] & in2[71];
    assign P[158] = in[71] ^ in2[71];
    assign G[159] = in[70] & in2[70];
    assign P[159] = in[70] ^ in2[70];
    assign G[160] = in[69] & in2[69];
    assign P[160] = in[69] ^ in2[69];
    assign G[161] = in[68] & in2[68];
    assign P[161] = in[68] ^ in2[68];
    assign G[162] = in[67] & in2[67];
    assign P[162] = in[67] ^ in2[67];
    assign G[163] = in[66] & in2[66];
    assign P[163] = in[66] ^ in2[66];
    assign G[164] = in[65] & in2[65];
    assign P[164] = in[65] ^ in2[65];
    assign G[165] = in[64] & in2[64];
    assign P[165] = in[64] ^ in2[64];
    assign G[166] = in[63] & in2[63];
    assign P[166] = in[63] ^ in2[63];
    assign G[167] = in[62] & in2[62];
    assign P[167] = in[62] ^ in2[62];
    assign G[168] = in[61] & in2[61];
    assign P[168] = in[61] ^ in2[61];
    assign G[169] = in[60] & in2[60];
    assign P[169] = in[60] ^ in2[60];
    assign G[170] = in[59] & in2[59];
    assign P[170] = in[59] ^ in2[59];
    assign G[171] = in[58] & in2[58];
    assign P[171] = in[58] ^ in2[58];
    assign G[172] = in[57] & in2[57];
    assign P[172] = in[57] ^ in2[57];
    assign G[173] = in[56] & in2[56];
    assign P[173] = in[56] ^ in2[56];
    assign G[174] = in[55] & in2[55];
    assign P[174] = in[55] ^ in2[55];
    assign G[175] = in[54] & in2[54];
    assign P[175] = in[54] ^ in2[54];
    assign G[176] = in[53] & in2[53];
    assign P[176] = in[53] ^ in2[53];
    assign G[177] = in[52] & in2[52];
    assign P[177] = in[52] ^ in2[52];
    assign G[178] = in[51] & in2[51];
    assign P[178] = in[51] ^ in2[51];
    assign G[179] = in[50] & in2[50];
    assign P[179] = in[50] ^ in2[50];
    assign G[180] = in[49] & in2[49];
    assign P[180] = in[49] ^ in2[49];
    assign G[181] = in[48] & in2[48];
    assign P[181] = in[48] ^ in2[48];
    assign G[182] = in[47] & in2[47];
    assign P[182] = in[47] ^ in2[47];
    assign G[183] = in[46] & in2[46];
    assign P[183] = in[46] ^ in2[46];
    assign G[184] = in[45] & in2[45];
    assign P[184] = in[45] ^ in2[45];
    assign G[185] = in[44] & in2[44];
    assign P[185] = in[44] ^ in2[44];
    assign G[186] = in[43] & in2[43];
    assign P[186] = in[43] ^ in2[43];
    assign G[187] = in[42] & in2[42];
    assign P[187] = in[42] ^ in2[42];
    assign G[188] = in[41] & in2[41];
    assign P[188] = in[41] ^ in2[41];
    assign G[189] = in[40] & in2[40];
    assign P[189] = in[40] ^ in2[40];
    assign G[190] = in[39] & in2[39];
    assign P[190] = in[39] ^ in2[39];
    assign G[191] = in[38] & in2[38];
    assign P[191] = in[38] ^ in2[38];
    assign G[192] = in[37] & in2[37];
    assign P[192] = in[37] ^ in2[37];
    assign G[193] = in[36] & in2[36];
    assign P[193] = in[36] ^ in2[36];
    assign G[194] = in[35] & in2[35];
    assign P[194] = in[35] ^ in2[35];
    assign G[195] = in[34] & in2[34];
    assign P[195] = in[34] ^ in2[34];
    assign G[196] = in[33] & in2[33];
    assign P[196] = in[33] ^ in2[33];
    assign G[197] = in[32] & in2[32];
    assign P[197] = in[32] ^ in2[32];
    assign G[198] = in[31] & in2[31];
    assign P[198] = in[31] ^ in2[31];
    assign G[199] = in[30] & in2[30];
    assign P[199] = in[30] ^ in2[30];
    assign G[200] = in[29] & in2[29];
    assign P[200] = in[29] ^ in2[29];
    assign G[201] = in[28] & in2[28];
    assign P[201] = in[28] ^ in2[28];
    assign G[202] = in[27] & in2[27];
    assign P[202] = in[27] ^ in2[27];
    assign G[203] = in[26] & in2[26];
    assign P[203] = in[26] ^ in2[26];
    assign G[204] = in[25] & in2[25];
    assign P[204] = in[25] ^ in2[25];
    assign G[205] = in[24] & in2[24];
    assign P[205] = in[24] ^ in2[24];
    assign G[206] = in[23] & in2[23];
    assign P[206] = in[23] ^ in2[23];
    assign G[207] = in[22] & in2[22];
    assign P[207] = in[22] ^ in2[22];
    assign G[208] = in[21] & in2[21];
    assign P[208] = in[21] ^ in2[21];
    assign G[209] = in[20] & in2[20];
    assign P[209] = in[20] ^ in2[20];
    assign G[210] = in[19] & in2[19];
    assign P[210] = in[19] ^ in2[19];
    assign G[211] = in[18] & in2[18];
    assign P[211] = in[18] ^ in2[18];
    assign G[212] = in[17] & in2[17];
    assign P[212] = in[17] ^ in2[17];
    assign G[213] = in[16] & in2[16];
    assign P[213] = in[16] ^ in2[16];
    assign G[214] = in[15] & in2[15];
    assign P[214] = in[15] ^ in2[15];
    assign G[215] = in[14] & in2[14];
    assign P[215] = in[14] ^ in2[14];
    assign G[216] = in[13] & in2[13];
    assign P[216] = in[13] ^ in2[13];
    assign G[217] = in[12] & in2[12];
    assign P[217] = in[12] ^ in2[12];
    assign G[218] = in[11] & in2[11];
    assign P[218] = in[11] ^ in2[11];
    assign G[219] = in[10] & in2[10];
    assign P[219] = in[10] ^ in2[10];
    assign G[220] = in[9] & in2[9];
    assign P[220] = in[9] ^ in2[9];
    assign G[221] = in[8] & in2[8];
    assign P[221] = in[8] ^ in2[8];
    assign G[222] = in[7] & in2[7];
    assign P[222] = in[7] ^ in2[7];
    assign G[223] = in[6] & in2[6];
    assign P[223] = in[6] ^ in2[6];
    assign G[224] = in[5] & in2[5];
    assign P[224] = in[5] ^ in2[5];
    assign G[225] = in[4] & in2[4];
    assign P[225] = in[4] ^ in2[4];
    assign G[226] = in[3] & in2[3];
    assign P[226] = in[3] ^ in2[3];
    assign G[227] = in[2] & in2[2];
    assign P[227] = in[2] ^ in2[2];
    assign G[228] = in[1] & in2[1];
    assign P[228] = in[1] ^ in2[1];
    assign G[229] = in[0] & in2[0];
    assign P[229] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign C[229] = G[228] | (P[228] & C[228]);
    assign cout = G[229] | (P[229] & C[229]);
    assign sum = P ^ C;
endmodule

module CLA229(output [228:0] sum, output cout, input [228:0] in1, input [228:0] in2;

    wire[228:0] G;
    wire[228:0] C;
    wire[228:0] P;

    assign G[0] = in[228] & in2[228];
    assign P[0] = in[228] ^ in2[228];
    assign G[1] = in[227] & in2[227];
    assign P[1] = in[227] ^ in2[227];
    assign G[2] = in[226] & in2[226];
    assign P[2] = in[226] ^ in2[226];
    assign G[3] = in[225] & in2[225];
    assign P[3] = in[225] ^ in2[225];
    assign G[4] = in[224] & in2[224];
    assign P[4] = in[224] ^ in2[224];
    assign G[5] = in[223] & in2[223];
    assign P[5] = in[223] ^ in2[223];
    assign G[6] = in[222] & in2[222];
    assign P[6] = in[222] ^ in2[222];
    assign G[7] = in[221] & in2[221];
    assign P[7] = in[221] ^ in2[221];
    assign G[8] = in[220] & in2[220];
    assign P[8] = in[220] ^ in2[220];
    assign G[9] = in[219] & in2[219];
    assign P[9] = in[219] ^ in2[219];
    assign G[10] = in[218] & in2[218];
    assign P[10] = in[218] ^ in2[218];
    assign G[11] = in[217] & in2[217];
    assign P[11] = in[217] ^ in2[217];
    assign G[12] = in[216] & in2[216];
    assign P[12] = in[216] ^ in2[216];
    assign G[13] = in[215] & in2[215];
    assign P[13] = in[215] ^ in2[215];
    assign G[14] = in[214] & in2[214];
    assign P[14] = in[214] ^ in2[214];
    assign G[15] = in[213] & in2[213];
    assign P[15] = in[213] ^ in2[213];
    assign G[16] = in[212] & in2[212];
    assign P[16] = in[212] ^ in2[212];
    assign G[17] = in[211] & in2[211];
    assign P[17] = in[211] ^ in2[211];
    assign G[18] = in[210] & in2[210];
    assign P[18] = in[210] ^ in2[210];
    assign G[19] = in[209] & in2[209];
    assign P[19] = in[209] ^ in2[209];
    assign G[20] = in[208] & in2[208];
    assign P[20] = in[208] ^ in2[208];
    assign G[21] = in[207] & in2[207];
    assign P[21] = in[207] ^ in2[207];
    assign G[22] = in[206] & in2[206];
    assign P[22] = in[206] ^ in2[206];
    assign G[23] = in[205] & in2[205];
    assign P[23] = in[205] ^ in2[205];
    assign G[24] = in[204] & in2[204];
    assign P[24] = in[204] ^ in2[204];
    assign G[25] = in[203] & in2[203];
    assign P[25] = in[203] ^ in2[203];
    assign G[26] = in[202] & in2[202];
    assign P[26] = in[202] ^ in2[202];
    assign G[27] = in[201] & in2[201];
    assign P[27] = in[201] ^ in2[201];
    assign G[28] = in[200] & in2[200];
    assign P[28] = in[200] ^ in2[200];
    assign G[29] = in[199] & in2[199];
    assign P[29] = in[199] ^ in2[199];
    assign G[30] = in[198] & in2[198];
    assign P[30] = in[198] ^ in2[198];
    assign G[31] = in[197] & in2[197];
    assign P[31] = in[197] ^ in2[197];
    assign G[32] = in[196] & in2[196];
    assign P[32] = in[196] ^ in2[196];
    assign G[33] = in[195] & in2[195];
    assign P[33] = in[195] ^ in2[195];
    assign G[34] = in[194] & in2[194];
    assign P[34] = in[194] ^ in2[194];
    assign G[35] = in[193] & in2[193];
    assign P[35] = in[193] ^ in2[193];
    assign G[36] = in[192] & in2[192];
    assign P[36] = in[192] ^ in2[192];
    assign G[37] = in[191] & in2[191];
    assign P[37] = in[191] ^ in2[191];
    assign G[38] = in[190] & in2[190];
    assign P[38] = in[190] ^ in2[190];
    assign G[39] = in[189] & in2[189];
    assign P[39] = in[189] ^ in2[189];
    assign G[40] = in[188] & in2[188];
    assign P[40] = in[188] ^ in2[188];
    assign G[41] = in[187] & in2[187];
    assign P[41] = in[187] ^ in2[187];
    assign G[42] = in[186] & in2[186];
    assign P[42] = in[186] ^ in2[186];
    assign G[43] = in[185] & in2[185];
    assign P[43] = in[185] ^ in2[185];
    assign G[44] = in[184] & in2[184];
    assign P[44] = in[184] ^ in2[184];
    assign G[45] = in[183] & in2[183];
    assign P[45] = in[183] ^ in2[183];
    assign G[46] = in[182] & in2[182];
    assign P[46] = in[182] ^ in2[182];
    assign G[47] = in[181] & in2[181];
    assign P[47] = in[181] ^ in2[181];
    assign G[48] = in[180] & in2[180];
    assign P[48] = in[180] ^ in2[180];
    assign G[49] = in[179] & in2[179];
    assign P[49] = in[179] ^ in2[179];
    assign G[50] = in[178] & in2[178];
    assign P[50] = in[178] ^ in2[178];
    assign G[51] = in[177] & in2[177];
    assign P[51] = in[177] ^ in2[177];
    assign G[52] = in[176] & in2[176];
    assign P[52] = in[176] ^ in2[176];
    assign G[53] = in[175] & in2[175];
    assign P[53] = in[175] ^ in2[175];
    assign G[54] = in[174] & in2[174];
    assign P[54] = in[174] ^ in2[174];
    assign G[55] = in[173] & in2[173];
    assign P[55] = in[173] ^ in2[173];
    assign G[56] = in[172] & in2[172];
    assign P[56] = in[172] ^ in2[172];
    assign G[57] = in[171] & in2[171];
    assign P[57] = in[171] ^ in2[171];
    assign G[58] = in[170] & in2[170];
    assign P[58] = in[170] ^ in2[170];
    assign G[59] = in[169] & in2[169];
    assign P[59] = in[169] ^ in2[169];
    assign G[60] = in[168] & in2[168];
    assign P[60] = in[168] ^ in2[168];
    assign G[61] = in[167] & in2[167];
    assign P[61] = in[167] ^ in2[167];
    assign G[62] = in[166] & in2[166];
    assign P[62] = in[166] ^ in2[166];
    assign G[63] = in[165] & in2[165];
    assign P[63] = in[165] ^ in2[165];
    assign G[64] = in[164] & in2[164];
    assign P[64] = in[164] ^ in2[164];
    assign G[65] = in[163] & in2[163];
    assign P[65] = in[163] ^ in2[163];
    assign G[66] = in[162] & in2[162];
    assign P[66] = in[162] ^ in2[162];
    assign G[67] = in[161] & in2[161];
    assign P[67] = in[161] ^ in2[161];
    assign G[68] = in[160] & in2[160];
    assign P[68] = in[160] ^ in2[160];
    assign G[69] = in[159] & in2[159];
    assign P[69] = in[159] ^ in2[159];
    assign G[70] = in[158] & in2[158];
    assign P[70] = in[158] ^ in2[158];
    assign G[71] = in[157] & in2[157];
    assign P[71] = in[157] ^ in2[157];
    assign G[72] = in[156] & in2[156];
    assign P[72] = in[156] ^ in2[156];
    assign G[73] = in[155] & in2[155];
    assign P[73] = in[155] ^ in2[155];
    assign G[74] = in[154] & in2[154];
    assign P[74] = in[154] ^ in2[154];
    assign G[75] = in[153] & in2[153];
    assign P[75] = in[153] ^ in2[153];
    assign G[76] = in[152] & in2[152];
    assign P[76] = in[152] ^ in2[152];
    assign G[77] = in[151] & in2[151];
    assign P[77] = in[151] ^ in2[151];
    assign G[78] = in[150] & in2[150];
    assign P[78] = in[150] ^ in2[150];
    assign G[79] = in[149] & in2[149];
    assign P[79] = in[149] ^ in2[149];
    assign G[80] = in[148] & in2[148];
    assign P[80] = in[148] ^ in2[148];
    assign G[81] = in[147] & in2[147];
    assign P[81] = in[147] ^ in2[147];
    assign G[82] = in[146] & in2[146];
    assign P[82] = in[146] ^ in2[146];
    assign G[83] = in[145] & in2[145];
    assign P[83] = in[145] ^ in2[145];
    assign G[84] = in[144] & in2[144];
    assign P[84] = in[144] ^ in2[144];
    assign G[85] = in[143] & in2[143];
    assign P[85] = in[143] ^ in2[143];
    assign G[86] = in[142] & in2[142];
    assign P[86] = in[142] ^ in2[142];
    assign G[87] = in[141] & in2[141];
    assign P[87] = in[141] ^ in2[141];
    assign G[88] = in[140] & in2[140];
    assign P[88] = in[140] ^ in2[140];
    assign G[89] = in[139] & in2[139];
    assign P[89] = in[139] ^ in2[139];
    assign G[90] = in[138] & in2[138];
    assign P[90] = in[138] ^ in2[138];
    assign G[91] = in[137] & in2[137];
    assign P[91] = in[137] ^ in2[137];
    assign G[92] = in[136] & in2[136];
    assign P[92] = in[136] ^ in2[136];
    assign G[93] = in[135] & in2[135];
    assign P[93] = in[135] ^ in2[135];
    assign G[94] = in[134] & in2[134];
    assign P[94] = in[134] ^ in2[134];
    assign G[95] = in[133] & in2[133];
    assign P[95] = in[133] ^ in2[133];
    assign G[96] = in[132] & in2[132];
    assign P[96] = in[132] ^ in2[132];
    assign G[97] = in[131] & in2[131];
    assign P[97] = in[131] ^ in2[131];
    assign G[98] = in[130] & in2[130];
    assign P[98] = in[130] ^ in2[130];
    assign G[99] = in[129] & in2[129];
    assign P[99] = in[129] ^ in2[129];
    assign G[100] = in[128] & in2[128];
    assign P[100] = in[128] ^ in2[128];
    assign G[101] = in[127] & in2[127];
    assign P[101] = in[127] ^ in2[127];
    assign G[102] = in[126] & in2[126];
    assign P[102] = in[126] ^ in2[126];
    assign G[103] = in[125] & in2[125];
    assign P[103] = in[125] ^ in2[125];
    assign G[104] = in[124] & in2[124];
    assign P[104] = in[124] ^ in2[124];
    assign G[105] = in[123] & in2[123];
    assign P[105] = in[123] ^ in2[123];
    assign G[106] = in[122] & in2[122];
    assign P[106] = in[122] ^ in2[122];
    assign G[107] = in[121] & in2[121];
    assign P[107] = in[121] ^ in2[121];
    assign G[108] = in[120] & in2[120];
    assign P[108] = in[120] ^ in2[120];
    assign G[109] = in[119] & in2[119];
    assign P[109] = in[119] ^ in2[119];
    assign G[110] = in[118] & in2[118];
    assign P[110] = in[118] ^ in2[118];
    assign G[111] = in[117] & in2[117];
    assign P[111] = in[117] ^ in2[117];
    assign G[112] = in[116] & in2[116];
    assign P[112] = in[116] ^ in2[116];
    assign G[113] = in[115] & in2[115];
    assign P[113] = in[115] ^ in2[115];
    assign G[114] = in[114] & in2[114];
    assign P[114] = in[114] ^ in2[114];
    assign G[115] = in[113] & in2[113];
    assign P[115] = in[113] ^ in2[113];
    assign G[116] = in[112] & in2[112];
    assign P[116] = in[112] ^ in2[112];
    assign G[117] = in[111] & in2[111];
    assign P[117] = in[111] ^ in2[111];
    assign G[118] = in[110] & in2[110];
    assign P[118] = in[110] ^ in2[110];
    assign G[119] = in[109] & in2[109];
    assign P[119] = in[109] ^ in2[109];
    assign G[120] = in[108] & in2[108];
    assign P[120] = in[108] ^ in2[108];
    assign G[121] = in[107] & in2[107];
    assign P[121] = in[107] ^ in2[107];
    assign G[122] = in[106] & in2[106];
    assign P[122] = in[106] ^ in2[106];
    assign G[123] = in[105] & in2[105];
    assign P[123] = in[105] ^ in2[105];
    assign G[124] = in[104] & in2[104];
    assign P[124] = in[104] ^ in2[104];
    assign G[125] = in[103] & in2[103];
    assign P[125] = in[103] ^ in2[103];
    assign G[126] = in[102] & in2[102];
    assign P[126] = in[102] ^ in2[102];
    assign G[127] = in[101] & in2[101];
    assign P[127] = in[101] ^ in2[101];
    assign G[128] = in[100] & in2[100];
    assign P[128] = in[100] ^ in2[100];
    assign G[129] = in[99] & in2[99];
    assign P[129] = in[99] ^ in2[99];
    assign G[130] = in[98] & in2[98];
    assign P[130] = in[98] ^ in2[98];
    assign G[131] = in[97] & in2[97];
    assign P[131] = in[97] ^ in2[97];
    assign G[132] = in[96] & in2[96];
    assign P[132] = in[96] ^ in2[96];
    assign G[133] = in[95] & in2[95];
    assign P[133] = in[95] ^ in2[95];
    assign G[134] = in[94] & in2[94];
    assign P[134] = in[94] ^ in2[94];
    assign G[135] = in[93] & in2[93];
    assign P[135] = in[93] ^ in2[93];
    assign G[136] = in[92] & in2[92];
    assign P[136] = in[92] ^ in2[92];
    assign G[137] = in[91] & in2[91];
    assign P[137] = in[91] ^ in2[91];
    assign G[138] = in[90] & in2[90];
    assign P[138] = in[90] ^ in2[90];
    assign G[139] = in[89] & in2[89];
    assign P[139] = in[89] ^ in2[89];
    assign G[140] = in[88] & in2[88];
    assign P[140] = in[88] ^ in2[88];
    assign G[141] = in[87] & in2[87];
    assign P[141] = in[87] ^ in2[87];
    assign G[142] = in[86] & in2[86];
    assign P[142] = in[86] ^ in2[86];
    assign G[143] = in[85] & in2[85];
    assign P[143] = in[85] ^ in2[85];
    assign G[144] = in[84] & in2[84];
    assign P[144] = in[84] ^ in2[84];
    assign G[145] = in[83] & in2[83];
    assign P[145] = in[83] ^ in2[83];
    assign G[146] = in[82] & in2[82];
    assign P[146] = in[82] ^ in2[82];
    assign G[147] = in[81] & in2[81];
    assign P[147] = in[81] ^ in2[81];
    assign G[148] = in[80] & in2[80];
    assign P[148] = in[80] ^ in2[80];
    assign G[149] = in[79] & in2[79];
    assign P[149] = in[79] ^ in2[79];
    assign G[150] = in[78] & in2[78];
    assign P[150] = in[78] ^ in2[78];
    assign G[151] = in[77] & in2[77];
    assign P[151] = in[77] ^ in2[77];
    assign G[152] = in[76] & in2[76];
    assign P[152] = in[76] ^ in2[76];
    assign G[153] = in[75] & in2[75];
    assign P[153] = in[75] ^ in2[75];
    assign G[154] = in[74] & in2[74];
    assign P[154] = in[74] ^ in2[74];
    assign G[155] = in[73] & in2[73];
    assign P[155] = in[73] ^ in2[73];
    assign G[156] = in[72] & in2[72];
    assign P[156] = in[72] ^ in2[72];
    assign G[157] = in[71] & in2[71];
    assign P[157] = in[71] ^ in2[71];
    assign G[158] = in[70] & in2[70];
    assign P[158] = in[70] ^ in2[70];
    assign G[159] = in[69] & in2[69];
    assign P[159] = in[69] ^ in2[69];
    assign G[160] = in[68] & in2[68];
    assign P[160] = in[68] ^ in2[68];
    assign G[161] = in[67] & in2[67];
    assign P[161] = in[67] ^ in2[67];
    assign G[162] = in[66] & in2[66];
    assign P[162] = in[66] ^ in2[66];
    assign G[163] = in[65] & in2[65];
    assign P[163] = in[65] ^ in2[65];
    assign G[164] = in[64] & in2[64];
    assign P[164] = in[64] ^ in2[64];
    assign G[165] = in[63] & in2[63];
    assign P[165] = in[63] ^ in2[63];
    assign G[166] = in[62] & in2[62];
    assign P[166] = in[62] ^ in2[62];
    assign G[167] = in[61] & in2[61];
    assign P[167] = in[61] ^ in2[61];
    assign G[168] = in[60] & in2[60];
    assign P[168] = in[60] ^ in2[60];
    assign G[169] = in[59] & in2[59];
    assign P[169] = in[59] ^ in2[59];
    assign G[170] = in[58] & in2[58];
    assign P[170] = in[58] ^ in2[58];
    assign G[171] = in[57] & in2[57];
    assign P[171] = in[57] ^ in2[57];
    assign G[172] = in[56] & in2[56];
    assign P[172] = in[56] ^ in2[56];
    assign G[173] = in[55] & in2[55];
    assign P[173] = in[55] ^ in2[55];
    assign G[174] = in[54] & in2[54];
    assign P[174] = in[54] ^ in2[54];
    assign G[175] = in[53] & in2[53];
    assign P[175] = in[53] ^ in2[53];
    assign G[176] = in[52] & in2[52];
    assign P[176] = in[52] ^ in2[52];
    assign G[177] = in[51] & in2[51];
    assign P[177] = in[51] ^ in2[51];
    assign G[178] = in[50] & in2[50];
    assign P[178] = in[50] ^ in2[50];
    assign G[179] = in[49] & in2[49];
    assign P[179] = in[49] ^ in2[49];
    assign G[180] = in[48] & in2[48];
    assign P[180] = in[48] ^ in2[48];
    assign G[181] = in[47] & in2[47];
    assign P[181] = in[47] ^ in2[47];
    assign G[182] = in[46] & in2[46];
    assign P[182] = in[46] ^ in2[46];
    assign G[183] = in[45] & in2[45];
    assign P[183] = in[45] ^ in2[45];
    assign G[184] = in[44] & in2[44];
    assign P[184] = in[44] ^ in2[44];
    assign G[185] = in[43] & in2[43];
    assign P[185] = in[43] ^ in2[43];
    assign G[186] = in[42] & in2[42];
    assign P[186] = in[42] ^ in2[42];
    assign G[187] = in[41] & in2[41];
    assign P[187] = in[41] ^ in2[41];
    assign G[188] = in[40] & in2[40];
    assign P[188] = in[40] ^ in2[40];
    assign G[189] = in[39] & in2[39];
    assign P[189] = in[39] ^ in2[39];
    assign G[190] = in[38] & in2[38];
    assign P[190] = in[38] ^ in2[38];
    assign G[191] = in[37] & in2[37];
    assign P[191] = in[37] ^ in2[37];
    assign G[192] = in[36] & in2[36];
    assign P[192] = in[36] ^ in2[36];
    assign G[193] = in[35] & in2[35];
    assign P[193] = in[35] ^ in2[35];
    assign G[194] = in[34] & in2[34];
    assign P[194] = in[34] ^ in2[34];
    assign G[195] = in[33] & in2[33];
    assign P[195] = in[33] ^ in2[33];
    assign G[196] = in[32] & in2[32];
    assign P[196] = in[32] ^ in2[32];
    assign G[197] = in[31] & in2[31];
    assign P[197] = in[31] ^ in2[31];
    assign G[198] = in[30] & in2[30];
    assign P[198] = in[30] ^ in2[30];
    assign G[199] = in[29] & in2[29];
    assign P[199] = in[29] ^ in2[29];
    assign G[200] = in[28] & in2[28];
    assign P[200] = in[28] ^ in2[28];
    assign G[201] = in[27] & in2[27];
    assign P[201] = in[27] ^ in2[27];
    assign G[202] = in[26] & in2[26];
    assign P[202] = in[26] ^ in2[26];
    assign G[203] = in[25] & in2[25];
    assign P[203] = in[25] ^ in2[25];
    assign G[204] = in[24] & in2[24];
    assign P[204] = in[24] ^ in2[24];
    assign G[205] = in[23] & in2[23];
    assign P[205] = in[23] ^ in2[23];
    assign G[206] = in[22] & in2[22];
    assign P[206] = in[22] ^ in2[22];
    assign G[207] = in[21] & in2[21];
    assign P[207] = in[21] ^ in2[21];
    assign G[208] = in[20] & in2[20];
    assign P[208] = in[20] ^ in2[20];
    assign G[209] = in[19] & in2[19];
    assign P[209] = in[19] ^ in2[19];
    assign G[210] = in[18] & in2[18];
    assign P[210] = in[18] ^ in2[18];
    assign G[211] = in[17] & in2[17];
    assign P[211] = in[17] ^ in2[17];
    assign G[212] = in[16] & in2[16];
    assign P[212] = in[16] ^ in2[16];
    assign G[213] = in[15] & in2[15];
    assign P[213] = in[15] ^ in2[15];
    assign G[214] = in[14] & in2[14];
    assign P[214] = in[14] ^ in2[14];
    assign G[215] = in[13] & in2[13];
    assign P[215] = in[13] ^ in2[13];
    assign G[216] = in[12] & in2[12];
    assign P[216] = in[12] ^ in2[12];
    assign G[217] = in[11] & in2[11];
    assign P[217] = in[11] ^ in2[11];
    assign G[218] = in[10] & in2[10];
    assign P[218] = in[10] ^ in2[10];
    assign G[219] = in[9] & in2[9];
    assign P[219] = in[9] ^ in2[9];
    assign G[220] = in[8] & in2[8];
    assign P[220] = in[8] ^ in2[8];
    assign G[221] = in[7] & in2[7];
    assign P[221] = in[7] ^ in2[7];
    assign G[222] = in[6] & in2[6];
    assign P[222] = in[6] ^ in2[6];
    assign G[223] = in[5] & in2[5];
    assign P[223] = in[5] ^ in2[5];
    assign G[224] = in[4] & in2[4];
    assign P[224] = in[4] ^ in2[4];
    assign G[225] = in[3] & in2[3];
    assign P[225] = in[3] ^ in2[3];
    assign G[226] = in[2] & in2[2];
    assign P[226] = in[2] ^ in2[2];
    assign G[227] = in[1] & in2[1];
    assign P[227] = in[1] ^ in2[1];
    assign G[228] = in[0] & in2[0];
    assign P[228] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign C[228] = G[227] | (P[227] & C[227]);
    assign cout = G[228] | (P[228] & C[228]);
    assign sum = P ^ C;
endmodule

module CLA228(output [227:0] sum, output cout, input [227:0] in1, input [227:0] in2;

    wire[227:0] G;
    wire[227:0] C;
    wire[227:0] P;

    assign G[0] = in[227] & in2[227];
    assign P[0] = in[227] ^ in2[227];
    assign G[1] = in[226] & in2[226];
    assign P[1] = in[226] ^ in2[226];
    assign G[2] = in[225] & in2[225];
    assign P[2] = in[225] ^ in2[225];
    assign G[3] = in[224] & in2[224];
    assign P[3] = in[224] ^ in2[224];
    assign G[4] = in[223] & in2[223];
    assign P[4] = in[223] ^ in2[223];
    assign G[5] = in[222] & in2[222];
    assign P[5] = in[222] ^ in2[222];
    assign G[6] = in[221] & in2[221];
    assign P[6] = in[221] ^ in2[221];
    assign G[7] = in[220] & in2[220];
    assign P[7] = in[220] ^ in2[220];
    assign G[8] = in[219] & in2[219];
    assign P[8] = in[219] ^ in2[219];
    assign G[9] = in[218] & in2[218];
    assign P[9] = in[218] ^ in2[218];
    assign G[10] = in[217] & in2[217];
    assign P[10] = in[217] ^ in2[217];
    assign G[11] = in[216] & in2[216];
    assign P[11] = in[216] ^ in2[216];
    assign G[12] = in[215] & in2[215];
    assign P[12] = in[215] ^ in2[215];
    assign G[13] = in[214] & in2[214];
    assign P[13] = in[214] ^ in2[214];
    assign G[14] = in[213] & in2[213];
    assign P[14] = in[213] ^ in2[213];
    assign G[15] = in[212] & in2[212];
    assign P[15] = in[212] ^ in2[212];
    assign G[16] = in[211] & in2[211];
    assign P[16] = in[211] ^ in2[211];
    assign G[17] = in[210] & in2[210];
    assign P[17] = in[210] ^ in2[210];
    assign G[18] = in[209] & in2[209];
    assign P[18] = in[209] ^ in2[209];
    assign G[19] = in[208] & in2[208];
    assign P[19] = in[208] ^ in2[208];
    assign G[20] = in[207] & in2[207];
    assign P[20] = in[207] ^ in2[207];
    assign G[21] = in[206] & in2[206];
    assign P[21] = in[206] ^ in2[206];
    assign G[22] = in[205] & in2[205];
    assign P[22] = in[205] ^ in2[205];
    assign G[23] = in[204] & in2[204];
    assign P[23] = in[204] ^ in2[204];
    assign G[24] = in[203] & in2[203];
    assign P[24] = in[203] ^ in2[203];
    assign G[25] = in[202] & in2[202];
    assign P[25] = in[202] ^ in2[202];
    assign G[26] = in[201] & in2[201];
    assign P[26] = in[201] ^ in2[201];
    assign G[27] = in[200] & in2[200];
    assign P[27] = in[200] ^ in2[200];
    assign G[28] = in[199] & in2[199];
    assign P[28] = in[199] ^ in2[199];
    assign G[29] = in[198] & in2[198];
    assign P[29] = in[198] ^ in2[198];
    assign G[30] = in[197] & in2[197];
    assign P[30] = in[197] ^ in2[197];
    assign G[31] = in[196] & in2[196];
    assign P[31] = in[196] ^ in2[196];
    assign G[32] = in[195] & in2[195];
    assign P[32] = in[195] ^ in2[195];
    assign G[33] = in[194] & in2[194];
    assign P[33] = in[194] ^ in2[194];
    assign G[34] = in[193] & in2[193];
    assign P[34] = in[193] ^ in2[193];
    assign G[35] = in[192] & in2[192];
    assign P[35] = in[192] ^ in2[192];
    assign G[36] = in[191] & in2[191];
    assign P[36] = in[191] ^ in2[191];
    assign G[37] = in[190] & in2[190];
    assign P[37] = in[190] ^ in2[190];
    assign G[38] = in[189] & in2[189];
    assign P[38] = in[189] ^ in2[189];
    assign G[39] = in[188] & in2[188];
    assign P[39] = in[188] ^ in2[188];
    assign G[40] = in[187] & in2[187];
    assign P[40] = in[187] ^ in2[187];
    assign G[41] = in[186] & in2[186];
    assign P[41] = in[186] ^ in2[186];
    assign G[42] = in[185] & in2[185];
    assign P[42] = in[185] ^ in2[185];
    assign G[43] = in[184] & in2[184];
    assign P[43] = in[184] ^ in2[184];
    assign G[44] = in[183] & in2[183];
    assign P[44] = in[183] ^ in2[183];
    assign G[45] = in[182] & in2[182];
    assign P[45] = in[182] ^ in2[182];
    assign G[46] = in[181] & in2[181];
    assign P[46] = in[181] ^ in2[181];
    assign G[47] = in[180] & in2[180];
    assign P[47] = in[180] ^ in2[180];
    assign G[48] = in[179] & in2[179];
    assign P[48] = in[179] ^ in2[179];
    assign G[49] = in[178] & in2[178];
    assign P[49] = in[178] ^ in2[178];
    assign G[50] = in[177] & in2[177];
    assign P[50] = in[177] ^ in2[177];
    assign G[51] = in[176] & in2[176];
    assign P[51] = in[176] ^ in2[176];
    assign G[52] = in[175] & in2[175];
    assign P[52] = in[175] ^ in2[175];
    assign G[53] = in[174] & in2[174];
    assign P[53] = in[174] ^ in2[174];
    assign G[54] = in[173] & in2[173];
    assign P[54] = in[173] ^ in2[173];
    assign G[55] = in[172] & in2[172];
    assign P[55] = in[172] ^ in2[172];
    assign G[56] = in[171] & in2[171];
    assign P[56] = in[171] ^ in2[171];
    assign G[57] = in[170] & in2[170];
    assign P[57] = in[170] ^ in2[170];
    assign G[58] = in[169] & in2[169];
    assign P[58] = in[169] ^ in2[169];
    assign G[59] = in[168] & in2[168];
    assign P[59] = in[168] ^ in2[168];
    assign G[60] = in[167] & in2[167];
    assign P[60] = in[167] ^ in2[167];
    assign G[61] = in[166] & in2[166];
    assign P[61] = in[166] ^ in2[166];
    assign G[62] = in[165] & in2[165];
    assign P[62] = in[165] ^ in2[165];
    assign G[63] = in[164] & in2[164];
    assign P[63] = in[164] ^ in2[164];
    assign G[64] = in[163] & in2[163];
    assign P[64] = in[163] ^ in2[163];
    assign G[65] = in[162] & in2[162];
    assign P[65] = in[162] ^ in2[162];
    assign G[66] = in[161] & in2[161];
    assign P[66] = in[161] ^ in2[161];
    assign G[67] = in[160] & in2[160];
    assign P[67] = in[160] ^ in2[160];
    assign G[68] = in[159] & in2[159];
    assign P[68] = in[159] ^ in2[159];
    assign G[69] = in[158] & in2[158];
    assign P[69] = in[158] ^ in2[158];
    assign G[70] = in[157] & in2[157];
    assign P[70] = in[157] ^ in2[157];
    assign G[71] = in[156] & in2[156];
    assign P[71] = in[156] ^ in2[156];
    assign G[72] = in[155] & in2[155];
    assign P[72] = in[155] ^ in2[155];
    assign G[73] = in[154] & in2[154];
    assign P[73] = in[154] ^ in2[154];
    assign G[74] = in[153] & in2[153];
    assign P[74] = in[153] ^ in2[153];
    assign G[75] = in[152] & in2[152];
    assign P[75] = in[152] ^ in2[152];
    assign G[76] = in[151] & in2[151];
    assign P[76] = in[151] ^ in2[151];
    assign G[77] = in[150] & in2[150];
    assign P[77] = in[150] ^ in2[150];
    assign G[78] = in[149] & in2[149];
    assign P[78] = in[149] ^ in2[149];
    assign G[79] = in[148] & in2[148];
    assign P[79] = in[148] ^ in2[148];
    assign G[80] = in[147] & in2[147];
    assign P[80] = in[147] ^ in2[147];
    assign G[81] = in[146] & in2[146];
    assign P[81] = in[146] ^ in2[146];
    assign G[82] = in[145] & in2[145];
    assign P[82] = in[145] ^ in2[145];
    assign G[83] = in[144] & in2[144];
    assign P[83] = in[144] ^ in2[144];
    assign G[84] = in[143] & in2[143];
    assign P[84] = in[143] ^ in2[143];
    assign G[85] = in[142] & in2[142];
    assign P[85] = in[142] ^ in2[142];
    assign G[86] = in[141] & in2[141];
    assign P[86] = in[141] ^ in2[141];
    assign G[87] = in[140] & in2[140];
    assign P[87] = in[140] ^ in2[140];
    assign G[88] = in[139] & in2[139];
    assign P[88] = in[139] ^ in2[139];
    assign G[89] = in[138] & in2[138];
    assign P[89] = in[138] ^ in2[138];
    assign G[90] = in[137] & in2[137];
    assign P[90] = in[137] ^ in2[137];
    assign G[91] = in[136] & in2[136];
    assign P[91] = in[136] ^ in2[136];
    assign G[92] = in[135] & in2[135];
    assign P[92] = in[135] ^ in2[135];
    assign G[93] = in[134] & in2[134];
    assign P[93] = in[134] ^ in2[134];
    assign G[94] = in[133] & in2[133];
    assign P[94] = in[133] ^ in2[133];
    assign G[95] = in[132] & in2[132];
    assign P[95] = in[132] ^ in2[132];
    assign G[96] = in[131] & in2[131];
    assign P[96] = in[131] ^ in2[131];
    assign G[97] = in[130] & in2[130];
    assign P[97] = in[130] ^ in2[130];
    assign G[98] = in[129] & in2[129];
    assign P[98] = in[129] ^ in2[129];
    assign G[99] = in[128] & in2[128];
    assign P[99] = in[128] ^ in2[128];
    assign G[100] = in[127] & in2[127];
    assign P[100] = in[127] ^ in2[127];
    assign G[101] = in[126] & in2[126];
    assign P[101] = in[126] ^ in2[126];
    assign G[102] = in[125] & in2[125];
    assign P[102] = in[125] ^ in2[125];
    assign G[103] = in[124] & in2[124];
    assign P[103] = in[124] ^ in2[124];
    assign G[104] = in[123] & in2[123];
    assign P[104] = in[123] ^ in2[123];
    assign G[105] = in[122] & in2[122];
    assign P[105] = in[122] ^ in2[122];
    assign G[106] = in[121] & in2[121];
    assign P[106] = in[121] ^ in2[121];
    assign G[107] = in[120] & in2[120];
    assign P[107] = in[120] ^ in2[120];
    assign G[108] = in[119] & in2[119];
    assign P[108] = in[119] ^ in2[119];
    assign G[109] = in[118] & in2[118];
    assign P[109] = in[118] ^ in2[118];
    assign G[110] = in[117] & in2[117];
    assign P[110] = in[117] ^ in2[117];
    assign G[111] = in[116] & in2[116];
    assign P[111] = in[116] ^ in2[116];
    assign G[112] = in[115] & in2[115];
    assign P[112] = in[115] ^ in2[115];
    assign G[113] = in[114] & in2[114];
    assign P[113] = in[114] ^ in2[114];
    assign G[114] = in[113] & in2[113];
    assign P[114] = in[113] ^ in2[113];
    assign G[115] = in[112] & in2[112];
    assign P[115] = in[112] ^ in2[112];
    assign G[116] = in[111] & in2[111];
    assign P[116] = in[111] ^ in2[111];
    assign G[117] = in[110] & in2[110];
    assign P[117] = in[110] ^ in2[110];
    assign G[118] = in[109] & in2[109];
    assign P[118] = in[109] ^ in2[109];
    assign G[119] = in[108] & in2[108];
    assign P[119] = in[108] ^ in2[108];
    assign G[120] = in[107] & in2[107];
    assign P[120] = in[107] ^ in2[107];
    assign G[121] = in[106] & in2[106];
    assign P[121] = in[106] ^ in2[106];
    assign G[122] = in[105] & in2[105];
    assign P[122] = in[105] ^ in2[105];
    assign G[123] = in[104] & in2[104];
    assign P[123] = in[104] ^ in2[104];
    assign G[124] = in[103] & in2[103];
    assign P[124] = in[103] ^ in2[103];
    assign G[125] = in[102] & in2[102];
    assign P[125] = in[102] ^ in2[102];
    assign G[126] = in[101] & in2[101];
    assign P[126] = in[101] ^ in2[101];
    assign G[127] = in[100] & in2[100];
    assign P[127] = in[100] ^ in2[100];
    assign G[128] = in[99] & in2[99];
    assign P[128] = in[99] ^ in2[99];
    assign G[129] = in[98] & in2[98];
    assign P[129] = in[98] ^ in2[98];
    assign G[130] = in[97] & in2[97];
    assign P[130] = in[97] ^ in2[97];
    assign G[131] = in[96] & in2[96];
    assign P[131] = in[96] ^ in2[96];
    assign G[132] = in[95] & in2[95];
    assign P[132] = in[95] ^ in2[95];
    assign G[133] = in[94] & in2[94];
    assign P[133] = in[94] ^ in2[94];
    assign G[134] = in[93] & in2[93];
    assign P[134] = in[93] ^ in2[93];
    assign G[135] = in[92] & in2[92];
    assign P[135] = in[92] ^ in2[92];
    assign G[136] = in[91] & in2[91];
    assign P[136] = in[91] ^ in2[91];
    assign G[137] = in[90] & in2[90];
    assign P[137] = in[90] ^ in2[90];
    assign G[138] = in[89] & in2[89];
    assign P[138] = in[89] ^ in2[89];
    assign G[139] = in[88] & in2[88];
    assign P[139] = in[88] ^ in2[88];
    assign G[140] = in[87] & in2[87];
    assign P[140] = in[87] ^ in2[87];
    assign G[141] = in[86] & in2[86];
    assign P[141] = in[86] ^ in2[86];
    assign G[142] = in[85] & in2[85];
    assign P[142] = in[85] ^ in2[85];
    assign G[143] = in[84] & in2[84];
    assign P[143] = in[84] ^ in2[84];
    assign G[144] = in[83] & in2[83];
    assign P[144] = in[83] ^ in2[83];
    assign G[145] = in[82] & in2[82];
    assign P[145] = in[82] ^ in2[82];
    assign G[146] = in[81] & in2[81];
    assign P[146] = in[81] ^ in2[81];
    assign G[147] = in[80] & in2[80];
    assign P[147] = in[80] ^ in2[80];
    assign G[148] = in[79] & in2[79];
    assign P[148] = in[79] ^ in2[79];
    assign G[149] = in[78] & in2[78];
    assign P[149] = in[78] ^ in2[78];
    assign G[150] = in[77] & in2[77];
    assign P[150] = in[77] ^ in2[77];
    assign G[151] = in[76] & in2[76];
    assign P[151] = in[76] ^ in2[76];
    assign G[152] = in[75] & in2[75];
    assign P[152] = in[75] ^ in2[75];
    assign G[153] = in[74] & in2[74];
    assign P[153] = in[74] ^ in2[74];
    assign G[154] = in[73] & in2[73];
    assign P[154] = in[73] ^ in2[73];
    assign G[155] = in[72] & in2[72];
    assign P[155] = in[72] ^ in2[72];
    assign G[156] = in[71] & in2[71];
    assign P[156] = in[71] ^ in2[71];
    assign G[157] = in[70] & in2[70];
    assign P[157] = in[70] ^ in2[70];
    assign G[158] = in[69] & in2[69];
    assign P[158] = in[69] ^ in2[69];
    assign G[159] = in[68] & in2[68];
    assign P[159] = in[68] ^ in2[68];
    assign G[160] = in[67] & in2[67];
    assign P[160] = in[67] ^ in2[67];
    assign G[161] = in[66] & in2[66];
    assign P[161] = in[66] ^ in2[66];
    assign G[162] = in[65] & in2[65];
    assign P[162] = in[65] ^ in2[65];
    assign G[163] = in[64] & in2[64];
    assign P[163] = in[64] ^ in2[64];
    assign G[164] = in[63] & in2[63];
    assign P[164] = in[63] ^ in2[63];
    assign G[165] = in[62] & in2[62];
    assign P[165] = in[62] ^ in2[62];
    assign G[166] = in[61] & in2[61];
    assign P[166] = in[61] ^ in2[61];
    assign G[167] = in[60] & in2[60];
    assign P[167] = in[60] ^ in2[60];
    assign G[168] = in[59] & in2[59];
    assign P[168] = in[59] ^ in2[59];
    assign G[169] = in[58] & in2[58];
    assign P[169] = in[58] ^ in2[58];
    assign G[170] = in[57] & in2[57];
    assign P[170] = in[57] ^ in2[57];
    assign G[171] = in[56] & in2[56];
    assign P[171] = in[56] ^ in2[56];
    assign G[172] = in[55] & in2[55];
    assign P[172] = in[55] ^ in2[55];
    assign G[173] = in[54] & in2[54];
    assign P[173] = in[54] ^ in2[54];
    assign G[174] = in[53] & in2[53];
    assign P[174] = in[53] ^ in2[53];
    assign G[175] = in[52] & in2[52];
    assign P[175] = in[52] ^ in2[52];
    assign G[176] = in[51] & in2[51];
    assign P[176] = in[51] ^ in2[51];
    assign G[177] = in[50] & in2[50];
    assign P[177] = in[50] ^ in2[50];
    assign G[178] = in[49] & in2[49];
    assign P[178] = in[49] ^ in2[49];
    assign G[179] = in[48] & in2[48];
    assign P[179] = in[48] ^ in2[48];
    assign G[180] = in[47] & in2[47];
    assign P[180] = in[47] ^ in2[47];
    assign G[181] = in[46] & in2[46];
    assign P[181] = in[46] ^ in2[46];
    assign G[182] = in[45] & in2[45];
    assign P[182] = in[45] ^ in2[45];
    assign G[183] = in[44] & in2[44];
    assign P[183] = in[44] ^ in2[44];
    assign G[184] = in[43] & in2[43];
    assign P[184] = in[43] ^ in2[43];
    assign G[185] = in[42] & in2[42];
    assign P[185] = in[42] ^ in2[42];
    assign G[186] = in[41] & in2[41];
    assign P[186] = in[41] ^ in2[41];
    assign G[187] = in[40] & in2[40];
    assign P[187] = in[40] ^ in2[40];
    assign G[188] = in[39] & in2[39];
    assign P[188] = in[39] ^ in2[39];
    assign G[189] = in[38] & in2[38];
    assign P[189] = in[38] ^ in2[38];
    assign G[190] = in[37] & in2[37];
    assign P[190] = in[37] ^ in2[37];
    assign G[191] = in[36] & in2[36];
    assign P[191] = in[36] ^ in2[36];
    assign G[192] = in[35] & in2[35];
    assign P[192] = in[35] ^ in2[35];
    assign G[193] = in[34] & in2[34];
    assign P[193] = in[34] ^ in2[34];
    assign G[194] = in[33] & in2[33];
    assign P[194] = in[33] ^ in2[33];
    assign G[195] = in[32] & in2[32];
    assign P[195] = in[32] ^ in2[32];
    assign G[196] = in[31] & in2[31];
    assign P[196] = in[31] ^ in2[31];
    assign G[197] = in[30] & in2[30];
    assign P[197] = in[30] ^ in2[30];
    assign G[198] = in[29] & in2[29];
    assign P[198] = in[29] ^ in2[29];
    assign G[199] = in[28] & in2[28];
    assign P[199] = in[28] ^ in2[28];
    assign G[200] = in[27] & in2[27];
    assign P[200] = in[27] ^ in2[27];
    assign G[201] = in[26] & in2[26];
    assign P[201] = in[26] ^ in2[26];
    assign G[202] = in[25] & in2[25];
    assign P[202] = in[25] ^ in2[25];
    assign G[203] = in[24] & in2[24];
    assign P[203] = in[24] ^ in2[24];
    assign G[204] = in[23] & in2[23];
    assign P[204] = in[23] ^ in2[23];
    assign G[205] = in[22] & in2[22];
    assign P[205] = in[22] ^ in2[22];
    assign G[206] = in[21] & in2[21];
    assign P[206] = in[21] ^ in2[21];
    assign G[207] = in[20] & in2[20];
    assign P[207] = in[20] ^ in2[20];
    assign G[208] = in[19] & in2[19];
    assign P[208] = in[19] ^ in2[19];
    assign G[209] = in[18] & in2[18];
    assign P[209] = in[18] ^ in2[18];
    assign G[210] = in[17] & in2[17];
    assign P[210] = in[17] ^ in2[17];
    assign G[211] = in[16] & in2[16];
    assign P[211] = in[16] ^ in2[16];
    assign G[212] = in[15] & in2[15];
    assign P[212] = in[15] ^ in2[15];
    assign G[213] = in[14] & in2[14];
    assign P[213] = in[14] ^ in2[14];
    assign G[214] = in[13] & in2[13];
    assign P[214] = in[13] ^ in2[13];
    assign G[215] = in[12] & in2[12];
    assign P[215] = in[12] ^ in2[12];
    assign G[216] = in[11] & in2[11];
    assign P[216] = in[11] ^ in2[11];
    assign G[217] = in[10] & in2[10];
    assign P[217] = in[10] ^ in2[10];
    assign G[218] = in[9] & in2[9];
    assign P[218] = in[9] ^ in2[9];
    assign G[219] = in[8] & in2[8];
    assign P[219] = in[8] ^ in2[8];
    assign G[220] = in[7] & in2[7];
    assign P[220] = in[7] ^ in2[7];
    assign G[221] = in[6] & in2[6];
    assign P[221] = in[6] ^ in2[6];
    assign G[222] = in[5] & in2[5];
    assign P[222] = in[5] ^ in2[5];
    assign G[223] = in[4] & in2[4];
    assign P[223] = in[4] ^ in2[4];
    assign G[224] = in[3] & in2[3];
    assign P[224] = in[3] ^ in2[3];
    assign G[225] = in[2] & in2[2];
    assign P[225] = in[2] ^ in2[2];
    assign G[226] = in[1] & in2[1];
    assign P[226] = in[1] ^ in2[1];
    assign G[227] = in[0] & in2[0];
    assign P[227] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign C[227] = G[226] | (P[226] & C[226]);
    assign cout = G[227] | (P[227] & C[227]);
    assign sum = P ^ C;
endmodule

module CLA227(output [226:0] sum, output cout, input [226:0] in1, input [226:0] in2;

    wire[226:0] G;
    wire[226:0] C;
    wire[226:0] P;

    assign G[0] = in[226] & in2[226];
    assign P[0] = in[226] ^ in2[226];
    assign G[1] = in[225] & in2[225];
    assign P[1] = in[225] ^ in2[225];
    assign G[2] = in[224] & in2[224];
    assign P[2] = in[224] ^ in2[224];
    assign G[3] = in[223] & in2[223];
    assign P[3] = in[223] ^ in2[223];
    assign G[4] = in[222] & in2[222];
    assign P[4] = in[222] ^ in2[222];
    assign G[5] = in[221] & in2[221];
    assign P[5] = in[221] ^ in2[221];
    assign G[6] = in[220] & in2[220];
    assign P[6] = in[220] ^ in2[220];
    assign G[7] = in[219] & in2[219];
    assign P[7] = in[219] ^ in2[219];
    assign G[8] = in[218] & in2[218];
    assign P[8] = in[218] ^ in2[218];
    assign G[9] = in[217] & in2[217];
    assign P[9] = in[217] ^ in2[217];
    assign G[10] = in[216] & in2[216];
    assign P[10] = in[216] ^ in2[216];
    assign G[11] = in[215] & in2[215];
    assign P[11] = in[215] ^ in2[215];
    assign G[12] = in[214] & in2[214];
    assign P[12] = in[214] ^ in2[214];
    assign G[13] = in[213] & in2[213];
    assign P[13] = in[213] ^ in2[213];
    assign G[14] = in[212] & in2[212];
    assign P[14] = in[212] ^ in2[212];
    assign G[15] = in[211] & in2[211];
    assign P[15] = in[211] ^ in2[211];
    assign G[16] = in[210] & in2[210];
    assign P[16] = in[210] ^ in2[210];
    assign G[17] = in[209] & in2[209];
    assign P[17] = in[209] ^ in2[209];
    assign G[18] = in[208] & in2[208];
    assign P[18] = in[208] ^ in2[208];
    assign G[19] = in[207] & in2[207];
    assign P[19] = in[207] ^ in2[207];
    assign G[20] = in[206] & in2[206];
    assign P[20] = in[206] ^ in2[206];
    assign G[21] = in[205] & in2[205];
    assign P[21] = in[205] ^ in2[205];
    assign G[22] = in[204] & in2[204];
    assign P[22] = in[204] ^ in2[204];
    assign G[23] = in[203] & in2[203];
    assign P[23] = in[203] ^ in2[203];
    assign G[24] = in[202] & in2[202];
    assign P[24] = in[202] ^ in2[202];
    assign G[25] = in[201] & in2[201];
    assign P[25] = in[201] ^ in2[201];
    assign G[26] = in[200] & in2[200];
    assign P[26] = in[200] ^ in2[200];
    assign G[27] = in[199] & in2[199];
    assign P[27] = in[199] ^ in2[199];
    assign G[28] = in[198] & in2[198];
    assign P[28] = in[198] ^ in2[198];
    assign G[29] = in[197] & in2[197];
    assign P[29] = in[197] ^ in2[197];
    assign G[30] = in[196] & in2[196];
    assign P[30] = in[196] ^ in2[196];
    assign G[31] = in[195] & in2[195];
    assign P[31] = in[195] ^ in2[195];
    assign G[32] = in[194] & in2[194];
    assign P[32] = in[194] ^ in2[194];
    assign G[33] = in[193] & in2[193];
    assign P[33] = in[193] ^ in2[193];
    assign G[34] = in[192] & in2[192];
    assign P[34] = in[192] ^ in2[192];
    assign G[35] = in[191] & in2[191];
    assign P[35] = in[191] ^ in2[191];
    assign G[36] = in[190] & in2[190];
    assign P[36] = in[190] ^ in2[190];
    assign G[37] = in[189] & in2[189];
    assign P[37] = in[189] ^ in2[189];
    assign G[38] = in[188] & in2[188];
    assign P[38] = in[188] ^ in2[188];
    assign G[39] = in[187] & in2[187];
    assign P[39] = in[187] ^ in2[187];
    assign G[40] = in[186] & in2[186];
    assign P[40] = in[186] ^ in2[186];
    assign G[41] = in[185] & in2[185];
    assign P[41] = in[185] ^ in2[185];
    assign G[42] = in[184] & in2[184];
    assign P[42] = in[184] ^ in2[184];
    assign G[43] = in[183] & in2[183];
    assign P[43] = in[183] ^ in2[183];
    assign G[44] = in[182] & in2[182];
    assign P[44] = in[182] ^ in2[182];
    assign G[45] = in[181] & in2[181];
    assign P[45] = in[181] ^ in2[181];
    assign G[46] = in[180] & in2[180];
    assign P[46] = in[180] ^ in2[180];
    assign G[47] = in[179] & in2[179];
    assign P[47] = in[179] ^ in2[179];
    assign G[48] = in[178] & in2[178];
    assign P[48] = in[178] ^ in2[178];
    assign G[49] = in[177] & in2[177];
    assign P[49] = in[177] ^ in2[177];
    assign G[50] = in[176] & in2[176];
    assign P[50] = in[176] ^ in2[176];
    assign G[51] = in[175] & in2[175];
    assign P[51] = in[175] ^ in2[175];
    assign G[52] = in[174] & in2[174];
    assign P[52] = in[174] ^ in2[174];
    assign G[53] = in[173] & in2[173];
    assign P[53] = in[173] ^ in2[173];
    assign G[54] = in[172] & in2[172];
    assign P[54] = in[172] ^ in2[172];
    assign G[55] = in[171] & in2[171];
    assign P[55] = in[171] ^ in2[171];
    assign G[56] = in[170] & in2[170];
    assign P[56] = in[170] ^ in2[170];
    assign G[57] = in[169] & in2[169];
    assign P[57] = in[169] ^ in2[169];
    assign G[58] = in[168] & in2[168];
    assign P[58] = in[168] ^ in2[168];
    assign G[59] = in[167] & in2[167];
    assign P[59] = in[167] ^ in2[167];
    assign G[60] = in[166] & in2[166];
    assign P[60] = in[166] ^ in2[166];
    assign G[61] = in[165] & in2[165];
    assign P[61] = in[165] ^ in2[165];
    assign G[62] = in[164] & in2[164];
    assign P[62] = in[164] ^ in2[164];
    assign G[63] = in[163] & in2[163];
    assign P[63] = in[163] ^ in2[163];
    assign G[64] = in[162] & in2[162];
    assign P[64] = in[162] ^ in2[162];
    assign G[65] = in[161] & in2[161];
    assign P[65] = in[161] ^ in2[161];
    assign G[66] = in[160] & in2[160];
    assign P[66] = in[160] ^ in2[160];
    assign G[67] = in[159] & in2[159];
    assign P[67] = in[159] ^ in2[159];
    assign G[68] = in[158] & in2[158];
    assign P[68] = in[158] ^ in2[158];
    assign G[69] = in[157] & in2[157];
    assign P[69] = in[157] ^ in2[157];
    assign G[70] = in[156] & in2[156];
    assign P[70] = in[156] ^ in2[156];
    assign G[71] = in[155] & in2[155];
    assign P[71] = in[155] ^ in2[155];
    assign G[72] = in[154] & in2[154];
    assign P[72] = in[154] ^ in2[154];
    assign G[73] = in[153] & in2[153];
    assign P[73] = in[153] ^ in2[153];
    assign G[74] = in[152] & in2[152];
    assign P[74] = in[152] ^ in2[152];
    assign G[75] = in[151] & in2[151];
    assign P[75] = in[151] ^ in2[151];
    assign G[76] = in[150] & in2[150];
    assign P[76] = in[150] ^ in2[150];
    assign G[77] = in[149] & in2[149];
    assign P[77] = in[149] ^ in2[149];
    assign G[78] = in[148] & in2[148];
    assign P[78] = in[148] ^ in2[148];
    assign G[79] = in[147] & in2[147];
    assign P[79] = in[147] ^ in2[147];
    assign G[80] = in[146] & in2[146];
    assign P[80] = in[146] ^ in2[146];
    assign G[81] = in[145] & in2[145];
    assign P[81] = in[145] ^ in2[145];
    assign G[82] = in[144] & in2[144];
    assign P[82] = in[144] ^ in2[144];
    assign G[83] = in[143] & in2[143];
    assign P[83] = in[143] ^ in2[143];
    assign G[84] = in[142] & in2[142];
    assign P[84] = in[142] ^ in2[142];
    assign G[85] = in[141] & in2[141];
    assign P[85] = in[141] ^ in2[141];
    assign G[86] = in[140] & in2[140];
    assign P[86] = in[140] ^ in2[140];
    assign G[87] = in[139] & in2[139];
    assign P[87] = in[139] ^ in2[139];
    assign G[88] = in[138] & in2[138];
    assign P[88] = in[138] ^ in2[138];
    assign G[89] = in[137] & in2[137];
    assign P[89] = in[137] ^ in2[137];
    assign G[90] = in[136] & in2[136];
    assign P[90] = in[136] ^ in2[136];
    assign G[91] = in[135] & in2[135];
    assign P[91] = in[135] ^ in2[135];
    assign G[92] = in[134] & in2[134];
    assign P[92] = in[134] ^ in2[134];
    assign G[93] = in[133] & in2[133];
    assign P[93] = in[133] ^ in2[133];
    assign G[94] = in[132] & in2[132];
    assign P[94] = in[132] ^ in2[132];
    assign G[95] = in[131] & in2[131];
    assign P[95] = in[131] ^ in2[131];
    assign G[96] = in[130] & in2[130];
    assign P[96] = in[130] ^ in2[130];
    assign G[97] = in[129] & in2[129];
    assign P[97] = in[129] ^ in2[129];
    assign G[98] = in[128] & in2[128];
    assign P[98] = in[128] ^ in2[128];
    assign G[99] = in[127] & in2[127];
    assign P[99] = in[127] ^ in2[127];
    assign G[100] = in[126] & in2[126];
    assign P[100] = in[126] ^ in2[126];
    assign G[101] = in[125] & in2[125];
    assign P[101] = in[125] ^ in2[125];
    assign G[102] = in[124] & in2[124];
    assign P[102] = in[124] ^ in2[124];
    assign G[103] = in[123] & in2[123];
    assign P[103] = in[123] ^ in2[123];
    assign G[104] = in[122] & in2[122];
    assign P[104] = in[122] ^ in2[122];
    assign G[105] = in[121] & in2[121];
    assign P[105] = in[121] ^ in2[121];
    assign G[106] = in[120] & in2[120];
    assign P[106] = in[120] ^ in2[120];
    assign G[107] = in[119] & in2[119];
    assign P[107] = in[119] ^ in2[119];
    assign G[108] = in[118] & in2[118];
    assign P[108] = in[118] ^ in2[118];
    assign G[109] = in[117] & in2[117];
    assign P[109] = in[117] ^ in2[117];
    assign G[110] = in[116] & in2[116];
    assign P[110] = in[116] ^ in2[116];
    assign G[111] = in[115] & in2[115];
    assign P[111] = in[115] ^ in2[115];
    assign G[112] = in[114] & in2[114];
    assign P[112] = in[114] ^ in2[114];
    assign G[113] = in[113] & in2[113];
    assign P[113] = in[113] ^ in2[113];
    assign G[114] = in[112] & in2[112];
    assign P[114] = in[112] ^ in2[112];
    assign G[115] = in[111] & in2[111];
    assign P[115] = in[111] ^ in2[111];
    assign G[116] = in[110] & in2[110];
    assign P[116] = in[110] ^ in2[110];
    assign G[117] = in[109] & in2[109];
    assign P[117] = in[109] ^ in2[109];
    assign G[118] = in[108] & in2[108];
    assign P[118] = in[108] ^ in2[108];
    assign G[119] = in[107] & in2[107];
    assign P[119] = in[107] ^ in2[107];
    assign G[120] = in[106] & in2[106];
    assign P[120] = in[106] ^ in2[106];
    assign G[121] = in[105] & in2[105];
    assign P[121] = in[105] ^ in2[105];
    assign G[122] = in[104] & in2[104];
    assign P[122] = in[104] ^ in2[104];
    assign G[123] = in[103] & in2[103];
    assign P[123] = in[103] ^ in2[103];
    assign G[124] = in[102] & in2[102];
    assign P[124] = in[102] ^ in2[102];
    assign G[125] = in[101] & in2[101];
    assign P[125] = in[101] ^ in2[101];
    assign G[126] = in[100] & in2[100];
    assign P[126] = in[100] ^ in2[100];
    assign G[127] = in[99] & in2[99];
    assign P[127] = in[99] ^ in2[99];
    assign G[128] = in[98] & in2[98];
    assign P[128] = in[98] ^ in2[98];
    assign G[129] = in[97] & in2[97];
    assign P[129] = in[97] ^ in2[97];
    assign G[130] = in[96] & in2[96];
    assign P[130] = in[96] ^ in2[96];
    assign G[131] = in[95] & in2[95];
    assign P[131] = in[95] ^ in2[95];
    assign G[132] = in[94] & in2[94];
    assign P[132] = in[94] ^ in2[94];
    assign G[133] = in[93] & in2[93];
    assign P[133] = in[93] ^ in2[93];
    assign G[134] = in[92] & in2[92];
    assign P[134] = in[92] ^ in2[92];
    assign G[135] = in[91] & in2[91];
    assign P[135] = in[91] ^ in2[91];
    assign G[136] = in[90] & in2[90];
    assign P[136] = in[90] ^ in2[90];
    assign G[137] = in[89] & in2[89];
    assign P[137] = in[89] ^ in2[89];
    assign G[138] = in[88] & in2[88];
    assign P[138] = in[88] ^ in2[88];
    assign G[139] = in[87] & in2[87];
    assign P[139] = in[87] ^ in2[87];
    assign G[140] = in[86] & in2[86];
    assign P[140] = in[86] ^ in2[86];
    assign G[141] = in[85] & in2[85];
    assign P[141] = in[85] ^ in2[85];
    assign G[142] = in[84] & in2[84];
    assign P[142] = in[84] ^ in2[84];
    assign G[143] = in[83] & in2[83];
    assign P[143] = in[83] ^ in2[83];
    assign G[144] = in[82] & in2[82];
    assign P[144] = in[82] ^ in2[82];
    assign G[145] = in[81] & in2[81];
    assign P[145] = in[81] ^ in2[81];
    assign G[146] = in[80] & in2[80];
    assign P[146] = in[80] ^ in2[80];
    assign G[147] = in[79] & in2[79];
    assign P[147] = in[79] ^ in2[79];
    assign G[148] = in[78] & in2[78];
    assign P[148] = in[78] ^ in2[78];
    assign G[149] = in[77] & in2[77];
    assign P[149] = in[77] ^ in2[77];
    assign G[150] = in[76] & in2[76];
    assign P[150] = in[76] ^ in2[76];
    assign G[151] = in[75] & in2[75];
    assign P[151] = in[75] ^ in2[75];
    assign G[152] = in[74] & in2[74];
    assign P[152] = in[74] ^ in2[74];
    assign G[153] = in[73] & in2[73];
    assign P[153] = in[73] ^ in2[73];
    assign G[154] = in[72] & in2[72];
    assign P[154] = in[72] ^ in2[72];
    assign G[155] = in[71] & in2[71];
    assign P[155] = in[71] ^ in2[71];
    assign G[156] = in[70] & in2[70];
    assign P[156] = in[70] ^ in2[70];
    assign G[157] = in[69] & in2[69];
    assign P[157] = in[69] ^ in2[69];
    assign G[158] = in[68] & in2[68];
    assign P[158] = in[68] ^ in2[68];
    assign G[159] = in[67] & in2[67];
    assign P[159] = in[67] ^ in2[67];
    assign G[160] = in[66] & in2[66];
    assign P[160] = in[66] ^ in2[66];
    assign G[161] = in[65] & in2[65];
    assign P[161] = in[65] ^ in2[65];
    assign G[162] = in[64] & in2[64];
    assign P[162] = in[64] ^ in2[64];
    assign G[163] = in[63] & in2[63];
    assign P[163] = in[63] ^ in2[63];
    assign G[164] = in[62] & in2[62];
    assign P[164] = in[62] ^ in2[62];
    assign G[165] = in[61] & in2[61];
    assign P[165] = in[61] ^ in2[61];
    assign G[166] = in[60] & in2[60];
    assign P[166] = in[60] ^ in2[60];
    assign G[167] = in[59] & in2[59];
    assign P[167] = in[59] ^ in2[59];
    assign G[168] = in[58] & in2[58];
    assign P[168] = in[58] ^ in2[58];
    assign G[169] = in[57] & in2[57];
    assign P[169] = in[57] ^ in2[57];
    assign G[170] = in[56] & in2[56];
    assign P[170] = in[56] ^ in2[56];
    assign G[171] = in[55] & in2[55];
    assign P[171] = in[55] ^ in2[55];
    assign G[172] = in[54] & in2[54];
    assign P[172] = in[54] ^ in2[54];
    assign G[173] = in[53] & in2[53];
    assign P[173] = in[53] ^ in2[53];
    assign G[174] = in[52] & in2[52];
    assign P[174] = in[52] ^ in2[52];
    assign G[175] = in[51] & in2[51];
    assign P[175] = in[51] ^ in2[51];
    assign G[176] = in[50] & in2[50];
    assign P[176] = in[50] ^ in2[50];
    assign G[177] = in[49] & in2[49];
    assign P[177] = in[49] ^ in2[49];
    assign G[178] = in[48] & in2[48];
    assign P[178] = in[48] ^ in2[48];
    assign G[179] = in[47] & in2[47];
    assign P[179] = in[47] ^ in2[47];
    assign G[180] = in[46] & in2[46];
    assign P[180] = in[46] ^ in2[46];
    assign G[181] = in[45] & in2[45];
    assign P[181] = in[45] ^ in2[45];
    assign G[182] = in[44] & in2[44];
    assign P[182] = in[44] ^ in2[44];
    assign G[183] = in[43] & in2[43];
    assign P[183] = in[43] ^ in2[43];
    assign G[184] = in[42] & in2[42];
    assign P[184] = in[42] ^ in2[42];
    assign G[185] = in[41] & in2[41];
    assign P[185] = in[41] ^ in2[41];
    assign G[186] = in[40] & in2[40];
    assign P[186] = in[40] ^ in2[40];
    assign G[187] = in[39] & in2[39];
    assign P[187] = in[39] ^ in2[39];
    assign G[188] = in[38] & in2[38];
    assign P[188] = in[38] ^ in2[38];
    assign G[189] = in[37] & in2[37];
    assign P[189] = in[37] ^ in2[37];
    assign G[190] = in[36] & in2[36];
    assign P[190] = in[36] ^ in2[36];
    assign G[191] = in[35] & in2[35];
    assign P[191] = in[35] ^ in2[35];
    assign G[192] = in[34] & in2[34];
    assign P[192] = in[34] ^ in2[34];
    assign G[193] = in[33] & in2[33];
    assign P[193] = in[33] ^ in2[33];
    assign G[194] = in[32] & in2[32];
    assign P[194] = in[32] ^ in2[32];
    assign G[195] = in[31] & in2[31];
    assign P[195] = in[31] ^ in2[31];
    assign G[196] = in[30] & in2[30];
    assign P[196] = in[30] ^ in2[30];
    assign G[197] = in[29] & in2[29];
    assign P[197] = in[29] ^ in2[29];
    assign G[198] = in[28] & in2[28];
    assign P[198] = in[28] ^ in2[28];
    assign G[199] = in[27] & in2[27];
    assign P[199] = in[27] ^ in2[27];
    assign G[200] = in[26] & in2[26];
    assign P[200] = in[26] ^ in2[26];
    assign G[201] = in[25] & in2[25];
    assign P[201] = in[25] ^ in2[25];
    assign G[202] = in[24] & in2[24];
    assign P[202] = in[24] ^ in2[24];
    assign G[203] = in[23] & in2[23];
    assign P[203] = in[23] ^ in2[23];
    assign G[204] = in[22] & in2[22];
    assign P[204] = in[22] ^ in2[22];
    assign G[205] = in[21] & in2[21];
    assign P[205] = in[21] ^ in2[21];
    assign G[206] = in[20] & in2[20];
    assign P[206] = in[20] ^ in2[20];
    assign G[207] = in[19] & in2[19];
    assign P[207] = in[19] ^ in2[19];
    assign G[208] = in[18] & in2[18];
    assign P[208] = in[18] ^ in2[18];
    assign G[209] = in[17] & in2[17];
    assign P[209] = in[17] ^ in2[17];
    assign G[210] = in[16] & in2[16];
    assign P[210] = in[16] ^ in2[16];
    assign G[211] = in[15] & in2[15];
    assign P[211] = in[15] ^ in2[15];
    assign G[212] = in[14] & in2[14];
    assign P[212] = in[14] ^ in2[14];
    assign G[213] = in[13] & in2[13];
    assign P[213] = in[13] ^ in2[13];
    assign G[214] = in[12] & in2[12];
    assign P[214] = in[12] ^ in2[12];
    assign G[215] = in[11] & in2[11];
    assign P[215] = in[11] ^ in2[11];
    assign G[216] = in[10] & in2[10];
    assign P[216] = in[10] ^ in2[10];
    assign G[217] = in[9] & in2[9];
    assign P[217] = in[9] ^ in2[9];
    assign G[218] = in[8] & in2[8];
    assign P[218] = in[8] ^ in2[8];
    assign G[219] = in[7] & in2[7];
    assign P[219] = in[7] ^ in2[7];
    assign G[220] = in[6] & in2[6];
    assign P[220] = in[6] ^ in2[6];
    assign G[221] = in[5] & in2[5];
    assign P[221] = in[5] ^ in2[5];
    assign G[222] = in[4] & in2[4];
    assign P[222] = in[4] ^ in2[4];
    assign G[223] = in[3] & in2[3];
    assign P[223] = in[3] ^ in2[3];
    assign G[224] = in[2] & in2[2];
    assign P[224] = in[2] ^ in2[2];
    assign G[225] = in[1] & in2[1];
    assign P[225] = in[1] ^ in2[1];
    assign G[226] = in[0] & in2[0];
    assign P[226] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign C[226] = G[225] | (P[225] & C[225]);
    assign cout = G[226] | (P[226] & C[226]);
    assign sum = P ^ C;
endmodule

module CLA226(output [225:0] sum, output cout, input [225:0] in1, input [225:0] in2;

    wire[225:0] G;
    wire[225:0] C;
    wire[225:0] P;

    assign G[0] = in[225] & in2[225];
    assign P[0] = in[225] ^ in2[225];
    assign G[1] = in[224] & in2[224];
    assign P[1] = in[224] ^ in2[224];
    assign G[2] = in[223] & in2[223];
    assign P[2] = in[223] ^ in2[223];
    assign G[3] = in[222] & in2[222];
    assign P[3] = in[222] ^ in2[222];
    assign G[4] = in[221] & in2[221];
    assign P[4] = in[221] ^ in2[221];
    assign G[5] = in[220] & in2[220];
    assign P[5] = in[220] ^ in2[220];
    assign G[6] = in[219] & in2[219];
    assign P[6] = in[219] ^ in2[219];
    assign G[7] = in[218] & in2[218];
    assign P[7] = in[218] ^ in2[218];
    assign G[8] = in[217] & in2[217];
    assign P[8] = in[217] ^ in2[217];
    assign G[9] = in[216] & in2[216];
    assign P[9] = in[216] ^ in2[216];
    assign G[10] = in[215] & in2[215];
    assign P[10] = in[215] ^ in2[215];
    assign G[11] = in[214] & in2[214];
    assign P[11] = in[214] ^ in2[214];
    assign G[12] = in[213] & in2[213];
    assign P[12] = in[213] ^ in2[213];
    assign G[13] = in[212] & in2[212];
    assign P[13] = in[212] ^ in2[212];
    assign G[14] = in[211] & in2[211];
    assign P[14] = in[211] ^ in2[211];
    assign G[15] = in[210] & in2[210];
    assign P[15] = in[210] ^ in2[210];
    assign G[16] = in[209] & in2[209];
    assign P[16] = in[209] ^ in2[209];
    assign G[17] = in[208] & in2[208];
    assign P[17] = in[208] ^ in2[208];
    assign G[18] = in[207] & in2[207];
    assign P[18] = in[207] ^ in2[207];
    assign G[19] = in[206] & in2[206];
    assign P[19] = in[206] ^ in2[206];
    assign G[20] = in[205] & in2[205];
    assign P[20] = in[205] ^ in2[205];
    assign G[21] = in[204] & in2[204];
    assign P[21] = in[204] ^ in2[204];
    assign G[22] = in[203] & in2[203];
    assign P[22] = in[203] ^ in2[203];
    assign G[23] = in[202] & in2[202];
    assign P[23] = in[202] ^ in2[202];
    assign G[24] = in[201] & in2[201];
    assign P[24] = in[201] ^ in2[201];
    assign G[25] = in[200] & in2[200];
    assign P[25] = in[200] ^ in2[200];
    assign G[26] = in[199] & in2[199];
    assign P[26] = in[199] ^ in2[199];
    assign G[27] = in[198] & in2[198];
    assign P[27] = in[198] ^ in2[198];
    assign G[28] = in[197] & in2[197];
    assign P[28] = in[197] ^ in2[197];
    assign G[29] = in[196] & in2[196];
    assign P[29] = in[196] ^ in2[196];
    assign G[30] = in[195] & in2[195];
    assign P[30] = in[195] ^ in2[195];
    assign G[31] = in[194] & in2[194];
    assign P[31] = in[194] ^ in2[194];
    assign G[32] = in[193] & in2[193];
    assign P[32] = in[193] ^ in2[193];
    assign G[33] = in[192] & in2[192];
    assign P[33] = in[192] ^ in2[192];
    assign G[34] = in[191] & in2[191];
    assign P[34] = in[191] ^ in2[191];
    assign G[35] = in[190] & in2[190];
    assign P[35] = in[190] ^ in2[190];
    assign G[36] = in[189] & in2[189];
    assign P[36] = in[189] ^ in2[189];
    assign G[37] = in[188] & in2[188];
    assign P[37] = in[188] ^ in2[188];
    assign G[38] = in[187] & in2[187];
    assign P[38] = in[187] ^ in2[187];
    assign G[39] = in[186] & in2[186];
    assign P[39] = in[186] ^ in2[186];
    assign G[40] = in[185] & in2[185];
    assign P[40] = in[185] ^ in2[185];
    assign G[41] = in[184] & in2[184];
    assign P[41] = in[184] ^ in2[184];
    assign G[42] = in[183] & in2[183];
    assign P[42] = in[183] ^ in2[183];
    assign G[43] = in[182] & in2[182];
    assign P[43] = in[182] ^ in2[182];
    assign G[44] = in[181] & in2[181];
    assign P[44] = in[181] ^ in2[181];
    assign G[45] = in[180] & in2[180];
    assign P[45] = in[180] ^ in2[180];
    assign G[46] = in[179] & in2[179];
    assign P[46] = in[179] ^ in2[179];
    assign G[47] = in[178] & in2[178];
    assign P[47] = in[178] ^ in2[178];
    assign G[48] = in[177] & in2[177];
    assign P[48] = in[177] ^ in2[177];
    assign G[49] = in[176] & in2[176];
    assign P[49] = in[176] ^ in2[176];
    assign G[50] = in[175] & in2[175];
    assign P[50] = in[175] ^ in2[175];
    assign G[51] = in[174] & in2[174];
    assign P[51] = in[174] ^ in2[174];
    assign G[52] = in[173] & in2[173];
    assign P[52] = in[173] ^ in2[173];
    assign G[53] = in[172] & in2[172];
    assign P[53] = in[172] ^ in2[172];
    assign G[54] = in[171] & in2[171];
    assign P[54] = in[171] ^ in2[171];
    assign G[55] = in[170] & in2[170];
    assign P[55] = in[170] ^ in2[170];
    assign G[56] = in[169] & in2[169];
    assign P[56] = in[169] ^ in2[169];
    assign G[57] = in[168] & in2[168];
    assign P[57] = in[168] ^ in2[168];
    assign G[58] = in[167] & in2[167];
    assign P[58] = in[167] ^ in2[167];
    assign G[59] = in[166] & in2[166];
    assign P[59] = in[166] ^ in2[166];
    assign G[60] = in[165] & in2[165];
    assign P[60] = in[165] ^ in2[165];
    assign G[61] = in[164] & in2[164];
    assign P[61] = in[164] ^ in2[164];
    assign G[62] = in[163] & in2[163];
    assign P[62] = in[163] ^ in2[163];
    assign G[63] = in[162] & in2[162];
    assign P[63] = in[162] ^ in2[162];
    assign G[64] = in[161] & in2[161];
    assign P[64] = in[161] ^ in2[161];
    assign G[65] = in[160] & in2[160];
    assign P[65] = in[160] ^ in2[160];
    assign G[66] = in[159] & in2[159];
    assign P[66] = in[159] ^ in2[159];
    assign G[67] = in[158] & in2[158];
    assign P[67] = in[158] ^ in2[158];
    assign G[68] = in[157] & in2[157];
    assign P[68] = in[157] ^ in2[157];
    assign G[69] = in[156] & in2[156];
    assign P[69] = in[156] ^ in2[156];
    assign G[70] = in[155] & in2[155];
    assign P[70] = in[155] ^ in2[155];
    assign G[71] = in[154] & in2[154];
    assign P[71] = in[154] ^ in2[154];
    assign G[72] = in[153] & in2[153];
    assign P[72] = in[153] ^ in2[153];
    assign G[73] = in[152] & in2[152];
    assign P[73] = in[152] ^ in2[152];
    assign G[74] = in[151] & in2[151];
    assign P[74] = in[151] ^ in2[151];
    assign G[75] = in[150] & in2[150];
    assign P[75] = in[150] ^ in2[150];
    assign G[76] = in[149] & in2[149];
    assign P[76] = in[149] ^ in2[149];
    assign G[77] = in[148] & in2[148];
    assign P[77] = in[148] ^ in2[148];
    assign G[78] = in[147] & in2[147];
    assign P[78] = in[147] ^ in2[147];
    assign G[79] = in[146] & in2[146];
    assign P[79] = in[146] ^ in2[146];
    assign G[80] = in[145] & in2[145];
    assign P[80] = in[145] ^ in2[145];
    assign G[81] = in[144] & in2[144];
    assign P[81] = in[144] ^ in2[144];
    assign G[82] = in[143] & in2[143];
    assign P[82] = in[143] ^ in2[143];
    assign G[83] = in[142] & in2[142];
    assign P[83] = in[142] ^ in2[142];
    assign G[84] = in[141] & in2[141];
    assign P[84] = in[141] ^ in2[141];
    assign G[85] = in[140] & in2[140];
    assign P[85] = in[140] ^ in2[140];
    assign G[86] = in[139] & in2[139];
    assign P[86] = in[139] ^ in2[139];
    assign G[87] = in[138] & in2[138];
    assign P[87] = in[138] ^ in2[138];
    assign G[88] = in[137] & in2[137];
    assign P[88] = in[137] ^ in2[137];
    assign G[89] = in[136] & in2[136];
    assign P[89] = in[136] ^ in2[136];
    assign G[90] = in[135] & in2[135];
    assign P[90] = in[135] ^ in2[135];
    assign G[91] = in[134] & in2[134];
    assign P[91] = in[134] ^ in2[134];
    assign G[92] = in[133] & in2[133];
    assign P[92] = in[133] ^ in2[133];
    assign G[93] = in[132] & in2[132];
    assign P[93] = in[132] ^ in2[132];
    assign G[94] = in[131] & in2[131];
    assign P[94] = in[131] ^ in2[131];
    assign G[95] = in[130] & in2[130];
    assign P[95] = in[130] ^ in2[130];
    assign G[96] = in[129] & in2[129];
    assign P[96] = in[129] ^ in2[129];
    assign G[97] = in[128] & in2[128];
    assign P[97] = in[128] ^ in2[128];
    assign G[98] = in[127] & in2[127];
    assign P[98] = in[127] ^ in2[127];
    assign G[99] = in[126] & in2[126];
    assign P[99] = in[126] ^ in2[126];
    assign G[100] = in[125] & in2[125];
    assign P[100] = in[125] ^ in2[125];
    assign G[101] = in[124] & in2[124];
    assign P[101] = in[124] ^ in2[124];
    assign G[102] = in[123] & in2[123];
    assign P[102] = in[123] ^ in2[123];
    assign G[103] = in[122] & in2[122];
    assign P[103] = in[122] ^ in2[122];
    assign G[104] = in[121] & in2[121];
    assign P[104] = in[121] ^ in2[121];
    assign G[105] = in[120] & in2[120];
    assign P[105] = in[120] ^ in2[120];
    assign G[106] = in[119] & in2[119];
    assign P[106] = in[119] ^ in2[119];
    assign G[107] = in[118] & in2[118];
    assign P[107] = in[118] ^ in2[118];
    assign G[108] = in[117] & in2[117];
    assign P[108] = in[117] ^ in2[117];
    assign G[109] = in[116] & in2[116];
    assign P[109] = in[116] ^ in2[116];
    assign G[110] = in[115] & in2[115];
    assign P[110] = in[115] ^ in2[115];
    assign G[111] = in[114] & in2[114];
    assign P[111] = in[114] ^ in2[114];
    assign G[112] = in[113] & in2[113];
    assign P[112] = in[113] ^ in2[113];
    assign G[113] = in[112] & in2[112];
    assign P[113] = in[112] ^ in2[112];
    assign G[114] = in[111] & in2[111];
    assign P[114] = in[111] ^ in2[111];
    assign G[115] = in[110] & in2[110];
    assign P[115] = in[110] ^ in2[110];
    assign G[116] = in[109] & in2[109];
    assign P[116] = in[109] ^ in2[109];
    assign G[117] = in[108] & in2[108];
    assign P[117] = in[108] ^ in2[108];
    assign G[118] = in[107] & in2[107];
    assign P[118] = in[107] ^ in2[107];
    assign G[119] = in[106] & in2[106];
    assign P[119] = in[106] ^ in2[106];
    assign G[120] = in[105] & in2[105];
    assign P[120] = in[105] ^ in2[105];
    assign G[121] = in[104] & in2[104];
    assign P[121] = in[104] ^ in2[104];
    assign G[122] = in[103] & in2[103];
    assign P[122] = in[103] ^ in2[103];
    assign G[123] = in[102] & in2[102];
    assign P[123] = in[102] ^ in2[102];
    assign G[124] = in[101] & in2[101];
    assign P[124] = in[101] ^ in2[101];
    assign G[125] = in[100] & in2[100];
    assign P[125] = in[100] ^ in2[100];
    assign G[126] = in[99] & in2[99];
    assign P[126] = in[99] ^ in2[99];
    assign G[127] = in[98] & in2[98];
    assign P[127] = in[98] ^ in2[98];
    assign G[128] = in[97] & in2[97];
    assign P[128] = in[97] ^ in2[97];
    assign G[129] = in[96] & in2[96];
    assign P[129] = in[96] ^ in2[96];
    assign G[130] = in[95] & in2[95];
    assign P[130] = in[95] ^ in2[95];
    assign G[131] = in[94] & in2[94];
    assign P[131] = in[94] ^ in2[94];
    assign G[132] = in[93] & in2[93];
    assign P[132] = in[93] ^ in2[93];
    assign G[133] = in[92] & in2[92];
    assign P[133] = in[92] ^ in2[92];
    assign G[134] = in[91] & in2[91];
    assign P[134] = in[91] ^ in2[91];
    assign G[135] = in[90] & in2[90];
    assign P[135] = in[90] ^ in2[90];
    assign G[136] = in[89] & in2[89];
    assign P[136] = in[89] ^ in2[89];
    assign G[137] = in[88] & in2[88];
    assign P[137] = in[88] ^ in2[88];
    assign G[138] = in[87] & in2[87];
    assign P[138] = in[87] ^ in2[87];
    assign G[139] = in[86] & in2[86];
    assign P[139] = in[86] ^ in2[86];
    assign G[140] = in[85] & in2[85];
    assign P[140] = in[85] ^ in2[85];
    assign G[141] = in[84] & in2[84];
    assign P[141] = in[84] ^ in2[84];
    assign G[142] = in[83] & in2[83];
    assign P[142] = in[83] ^ in2[83];
    assign G[143] = in[82] & in2[82];
    assign P[143] = in[82] ^ in2[82];
    assign G[144] = in[81] & in2[81];
    assign P[144] = in[81] ^ in2[81];
    assign G[145] = in[80] & in2[80];
    assign P[145] = in[80] ^ in2[80];
    assign G[146] = in[79] & in2[79];
    assign P[146] = in[79] ^ in2[79];
    assign G[147] = in[78] & in2[78];
    assign P[147] = in[78] ^ in2[78];
    assign G[148] = in[77] & in2[77];
    assign P[148] = in[77] ^ in2[77];
    assign G[149] = in[76] & in2[76];
    assign P[149] = in[76] ^ in2[76];
    assign G[150] = in[75] & in2[75];
    assign P[150] = in[75] ^ in2[75];
    assign G[151] = in[74] & in2[74];
    assign P[151] = in[74] ^ in2[74];
    assign G[152] = in[73] & in2[73];
    assign P[152] = in[73] ^ in2[73];
    assign G[153] = in[72] & in2[72];
    assign P[153] = in[72] ^ in2[72];
    assign G[154] = in[71] & in2[71];
    assign P[154] = in[71] ^ in2[71];
    assign G[155] = in[70] & in2[70];
    assign P[155] = in[70] ^ in2[70];
    assign G[156] = in[69] & in2[69];
    assign P[156] = in[69] ^ in2[69];
    assign G[157] = in[68] & in2[68];
    assign P[157] = in[68] ^ in2[68];
    assign G[158] = in[67] & in2[67];
    assign P[158] = in[67] ^ in2[67];
    assign G[159] = in[66] & in2[66];
    assign P[159] = in[66] ^ in2[66];
    assign G[160] = in[65] & in2[65];
    assign P[160] = in[65] ^ in2[65];
    assign G[161] = in[64] & in2[64];
    assign P[161] = in[64] ^ in2[64];
    assign G[162] = in[63] & in2[63];
    assign P[162] = in[63] ^ in2[63];
    assign G[163] = in[62] & in2[62];
    assign P[163] = in[62] ^ in2[62];
    assign G[164] = in[61] & in2[61];
    assign P[164] = in[61] ^ in2[61];
    assign G[165] = in[60] & in2[60];
    assign P[165] = in[60] ^ in2[60];
    assign G[166] = in[59] & in2[59];
    assign P[166] = in[59] ^ in2[59];
    assign G[167] = in[58] & in2[58];
    assign P[167] = in[58] ^ in2[58];
    assign G[168] = in[57] & in2[57];
    assign P[168] = in[57] ^ in2[57];
    assign G[169] = in[56] & in2[56];
    assign P[169] = in[56] ^ in2[56];
    assign G[170] = in[55] & in2[55];
    assign P[170] = in[55] ^ in2[55];
    assign G[171] = in[54] & in2[54];
    assign P[171] = in[54] ^ in2[54];
    assign G[172] = in[53] & in2[53];
    assign P[172] = in[53] ^ in2[53];
    assign G[173] = in[52] & in2[52];
    assign P[173] = in[52] ^ in2[52];
    assign G[174] = in[51] & in2[51];
    assign P[174] = in[51] ^ in2[51];
    assign G[175] = in[50] & in2[50];
    assign P[175] = in[50] ^ in2[50];
    assign G[176] = in[49] & in2[49];
    assign P[176] = in[49] ^ in2[49];
    assign G[177] = in[48] & in2[48];
    assign P[177] = in[48] ^ in2[48];
    assign G[178] = in[47] & in2[47];
    assign P[178] = in[47] ^ in2[47];
    assign G[179] = in[46] & in2[46];
    assign P[179] = in[46] ^ in2[46];
    assign G[180] = in[45] & in2[45];
    assign P[180] = in[45] ^ in2[45];
    assign G[181] = in[44] & in2[44];
    assign P[181] = in[44] ^ in2[44];
    assign G[182] = in[43] & in2[43];
    assign P[182] = in[43] ^ in2[43];
    assign G[183] = in[42] & in2[42];
    assign P[183] = in[42] ^ in2[42];
    assign G[184] = in[41] & in2[41];
    assign P[184] = in[41] ^ in2[41];
    assign G[185] = in[40] & in2[40];
    assign P[185] = in[40] ^ in2[40];
    assign G[186] = in[39] & in2[39];
    assign P[186] = in[39] ^ in2[39];
    assign G[187] = in[38] & in2[38];
    assign P[187] = in[38] ^ in2[38];
    assign G[188] = in[37] & in2[37];
    assign P[188] = in[37] ^ in2[37];
    assign G[189] = in[36] & in2[36];
    assign P[189] = in[36] ^ in2[36];
    assign G[190] = in[35] & in2[35];
    assign P[190] = in[35] ^ in2[35];
    assign G[191] = in[34] & in2[34];
    assign P[191] = in[34] ^ in2[34];
    assign G[192] = in[33] & in2[33];
    assign P[192] = in[33] ^ in2[33];
    assign G[193] = in[32] & in2[32];
    assign P[193] = in[32] ^ in2[32];
    assign G[194] = in[31] & in2[31];
    assign P[194] = in[31] ^ in2[31];
    assign G[195] = in[30] & in2[30];
    assign P[195] = in[30] ^ in2[30];
    assign G[196] = in[29] & in2[29];
    assign P[196] = in[29] ^ in2[29];
    assign G[197] = in[28] & in2[28];
    assign P[197] = in[28] ^ in2[28];
    assign G[198] = in[27] & in2[27];
    assign P[198] = in[27] ^ in2[27];
    assign G[199] = in[26] & in2[26];
    assign P[199] = in[26] ^ in2[26];
    assign G[200] = in[25] & in2[25];
    assign P[200] = in[25] ^ in2[25];
    assign G[201] = in[24] & in2[24];
    assign P[201] = in[24] ^ in2[24];
    assign G[202] = in[23] & in2[23];
    assign P[202] = in[23] ^ in2[23];
    assign G[203] = in[22] & in2[22];
    assign P[203] = in[22] ^ in2[22];
    assign G[204] = in[21] & in2[21];
    assign P[204] = in[21] ^ in2[21];
    assign G[205] = in[20] & in2[20];
    assign P[205] = in[20] ^ in2[20];
    assign G[206] = in[19] & in2[19];
    assign P[206] = in[19] ^ in2[19];
    assign G[207] = in[18] & in2[18];
    assign P[207] = in[18] ^ in2[18];
    assign G[208] = in[17] & in2[17];
    assign P[208] = in[17] ^ in2[17];
    assign G[209] = in[16] & in2[16];
    assign P[209] = in[16] ^ in2[16];
    assign G[210] = in[15] & in2[15];
    assign P[210] = in[15] ^ in2[15];
    assign G[211] = in[14] & in2[14];
    assign P[211] = in[14] ^ in2[14];
    assign G[212] = in[13] & in2[13];
    assign P[212] = in[13] ^ in2[13];
    assign G[213] = in[12] & in2[12];
    assign P[213] = in[12] ^ in2[12];
    assign G[214] = in[11] & in2[11];
    assign P[214] = in[11] ^ in2[11];
    assign G[215] = in[10] & in2[10];
    assign P[215] = in[10] ^ in2[10];
    assign G[216] = in[9] & in2[9];
    assign P[216] = in[9] ^ in2[9];
    assign G[217] = in[8] & in2[8];
    assign P[217] = in[8] ^ in2[8];
    assign G[218] = in[7] & in2[7];
    assign P[218] = in[7] ^ in2[7];
    assign G[219] = in[6] & in2[6];
    assign P[219] = in[6] ^ in2[6];
    assign G[220] = in[5] & in2[5];
    assign P[220] = in[5] ^ in2[5];
    assign G[221] = in[4] & in2[4];
    assign P[221] = in[4] ^ in2[4];
    assign G[222] = in[3] & in2[3];
    assign P[222] = in[3] ^ in2[3];
    assign G[223] = in[2] & in2[2];
    assign P[223] = in[2] ^ in2[2];
    assign G[224] = in[1] & in2[1];
    assign P[224] = in[1] ^ in2[1];
    assign G[225] = in[0] & in2[0];
    assign P[225] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign C[225] = G[224] | (P[224] & C[224]);
    assign cout = G[225] | (P[225] & C[225]);
    assign sum = P ^ C;
endmodule

module CLA225(output [224:0] sum, output cout, input [224:0] in1, input [224:0] in2;

    wire[224:0] G;
    wire[224:0] C;
    wire[224:0] P;

    assign G[0] = in[224] & in2[224];
    assign P[0] = in[224] ^ in2[224];
    assign G[1] = in[223] & in2[223];
    assign P[1] = in[223] ^ in2[223];
    assign G[2] = in[222] & in2[222];
    assign P[2] = in[222] ^ in2[222];
    assign G[3] = in[221] & in2[221];
    assign P[3] = in[221] ^ in2[221];
    assign G[4] = in[220] & in2[220];
    assign P[4] = in[220] ^ in2[220];
    assign G[5] = in[219] & in2[219];
    assign P[5] = in[219] ^ in2[219];
    assign G[6] = in[218] & in2[218];
    assign P[6] = in[218] ^ in2[218];
    assign G[7] = in[217] & in2[217];
    assign P[7] = in[217] ^ in2[217];
    assign G[8] = in[216] & in2[216];
    assign P[8] = in[216] ^ in2[216];
    assign G[9] = in[215] & in2[215];
    assign P[9] = in[215] ^ in2[215];
    assign G[10] = in[214] & in2[214];
    assign P[10] = in[214] ^ in2[214];
    assign G[11] = in[213] & in2[213];
    assign P[11] = in[213] ^ in2[213];
    assign G[12] = in[212] & in2[212];
    assign P[12] = in[212] ^ in2[212];
    assign G[13] = in[211] & in2[211];
    assign P[13] = in[211] ^ in2[211];
    assign G[14] = in[210] & in2[210];
    assign P[14] = in[210] ^ in2[210];
    assign G[15] = in[209] & in2[209];
    assign P[15] = in[209] ^ in2[209];
    assign G[16] = in[208] & in2[208];
    assign P[16] = in[208] ^ in2[208];
    assign G[17] = in[207] & in2[207];
    assign P[17] = in[207] ^ in2[207];
    assign G[18] = in[206] & in2[206];
    assign P[18] = in[206] ^ in2[206];
    assign G[19] = in[205] & in2[205];
    assign P[19] = in[205] ^ in2[205];
    assign G[20] = in[204] & in2[204];
    assign P[20] = in[204] ^ in2[204];
    assign G[21] = in[203] & in2[203];
    assign P[21] = in[203] ^ in2[203];
    assign G[22] = in[202] & in2[202];
    assign P[22] = in[202] ^ in2[202];
    assign G[23] = in[201] & in2[201];
    assign P[23] = in[201] ^ in2[201];
    assign G[24] = in[200] & in2[200];
    assign P[24] = in[200] ^ in2[200];
    assign G[25] = in[199] & in2[199];
    assign P[25] = in[199] ^ in2[199];
    assign G[26] = in[198] & in2[198];
    assign P[26] = in[198] ^ in2[198];
    assign G[27] = in[197] & in2[197];
    assign P[27] = in[197] ^ in2[197];
    assign G[28] = in[196] & in2[196];
    assign P[28] = in[196] ^ in2[196];
    assign G[29] = in[195] & in2[195];
    assign P[29] = in[195] ^ in2[195];
    assign G[30] = in[194] & in2[194];
    assign P[30] = in[194] ^ in2[194];
    assign G[31] = in[193] & in2[193];
    assign P[31] = in[193] ^ in2[193];
    assign G[32] = in[192] & in2[192];
    assign P[32] = in[192] ^ in2[192];
    assign G[33] = in[191] & in2[191];
    assign P[33] = in[191] ^ in2[191];
    assign G[34] = in[190] & in2[190];
    assign P[34] = in[190] ^ in2[190];
    assign G[35] = in[189] & in2[189];
    assign P[35] = in[189] ^ in2[189];
    assign G[36] = in[188] & in2[188];
    assign P[36] = in[188] ^ in2[188];
    assign G[37] = in[187] & in2[187];
    assign P[37] = in[187] ^ in2[187];
    assign G[38] = in[186] & in2[186];
    assign P[38] = in[186] ^ in2[186];
    assign G[39] = in[185] & in2[185];
    assign P[39] = in[185] ^ in2[185];
    assign G[40] = in[184] & in2[184];
    assign P[40] = in[184] ^ in2[184];
    assign G[41] = in[183] & in2[183];
    assign P[41] = in[183] ^ in2[183];
    assign G[42] = in[182] & in2[182];
    assign P[42] = in[182] ^ in2[182];
    assign G[43] = in[181] & in2[181];
    assign P[43] = in[181] ^ in2[181];
    assign G[44] = in[180] & in2[180];
    assign P[44] = in[180] ^ in2[180];
    assign G[45] = in[179] & in2[179];
    assign P[45] = in[179] ^ in2[179];
    assign G[46] = in[178] & in2[178];
    assign P[46] = in[178] ^ in2[178];
    assign G[47] = in[177] & in2[177];
    assign P[47] = in[177] ^ in2[177];
    assign G[48] = in[176] & in2[176];
    assign P[48] = in[176] ^ in2[176];
    assign G[49] = in[175] & in2[175];
    assign P[49] = in[175] ^ in2[175];
    assign G[50] = in[174] & in2[174];
    assign P[50] = in[174] ^ in2[174];
    assign G[51] = in[173] & in2[173];
    assign P[51] = in[173] ^ in2[173];
    assign G[52] = in[172] & in2[172];
    assign P[52] = in[172] ^ in2[172];
    assign G[53] = in[171] & in2[171];
    assign P[53] = in[171] ^ in2[171];
    assign G[54] = in[170] & in2[170];
    assign P[54] = in[170] ^ in2[170];
    assign G[55] = in[169] & in2[169];
    assign P[55] = in[169] ^ in2[169];
    assign G[56] = in[168] & in2[168];
    assign P[56] = in[168] ^ in2[168];
    assign G[57] = in[167] & in2[167];
    assign P[57] = in[167] ^ in2[167];
    assign G[58] = in[166] & in2[166];
    assign P[58] = in[166] ^ in2[166];
    assign G[59] = in[165] & in2[165];
    assign P[59] = in[165] ^ in2[165];
    assign G[60] = in[164] & in2[164];
    assign P[60] = in[164] ^ in2[164];
    assign G[61] = in[163] & in2[163];
    assign P[61] = in[163] ^ in2[163];
    assign G[62] = in[162] & in2[162];
    assign P[62] = in[162] ^ in2[162];
    assign G[63] = in[161] & in2[161];
    assign P[63] = in[161] ^ in2[161];
    assign G[64] = in[160] & in2[160];
    assign P[64] = in[160] ^ in2[160];
    assign G[65] = in[159] & in2[159];
    assign P[65] = in[159] ^ in2[159];
    assign G[66] = in[158] & in2[158];
    assign P[66] = in[158] ^ in2[158];
    assign G[67] = in[157] & in2[157];
    assign P[67] = in[157] ^ in2[157];
    assign G[68] = in[156] & in2[156];
    assign P[68] = in[156] ^ in2[156];
    assign G[69] = in[155] & in2[155];
    assign P[69] = in[155] ^ in2[155];
    assign G[70] = in[154] & in2[154];
    assign P[70] = in[154] ^ in2[154];
    assign G[71] = in[153] & in2[153];
    assign P[71] = in[153] ^ in2[153];
    assign G[72] = in[152] & in2[152];
    assign P[72] = in[152] ^ in2[152];
    assign G[73] = in[151] & in2[151];
    assign P[73] = in[151] ^ in2[151];
    assign G[74] = in[150] & in2[150];
    assign P[74] = in[150] ^ in2[150];
    assign G[75] = in[149] & in2[149];
    assign P[75] = in[149] ^ in2[149];
    assign G[76] = in[148] & in2[148];
    assign P[76] = in[148] ^ in2[148];
    assign G[77] = in[147] & in2[147];
    assign P[77] = in[147] ^ in2[147];
    assign G[78] = in[146] & in2[146];
    assign P[78] = in[146] ^ in2[146];
    assign G[79] = in[145] & in2[145];
    assign P[79] = in[145] ^ in2[145];
    assign G[80] = in[144] & in2[144];
    assign P[80] = in[144] ^ in2[144];
    assign G[81] = in[143] & in2[143];
    assign P[81] = in[143] ^ in2[143];
    assign G[82] = in[142] & in2[142];
    assign P[82] = in[142] ^ in2[142];
    assign G[83] = in[141] & in2[141];
    assign P[83] = in[141] ^ in2[141];
    assign G[84] = in[140] & in2[140];
    assign P[84] = in[140] ^ in2[140];
    assign G[85] = in[139] & in2[139];
    assign P[85] = in[139] ^ in2[139];
    assign G[86] = in[138] & in2[138];
    assign P[86] = in[138] ^ in2[138];
    assign G[87] = in[137] & in2[137];
    assign P[87] = in[137] ^ in2[137];
    assign G[88] = in[136] & in2[136];
    assign P[88] = in[136] ^ in2[136];
    assign G[89] = in[135] & in2[135];
    assign P[89] = in[135] ^ in2[135];
    assign G[90] = in[134] & in2[134];
    assign P[90] = in[134] ^ in2[134];
    assign G[91] = in[133] & in2[133];
    assign P[91] = in[133] ^ in2[133];
    assign G[92] = in[132] & in2[132];
    assign P[92] = in[132] ^ in2[132];
    assign G[93] = in[131] & in2[131];
    assign P[93] = in[131] ^ in2[131];
    assign G[94] = in[130] & in2[130];
    assign P[94] = in[130] ^ in2[130];
    assign G[95] = in[129] & in2[129];
    assign P[95] = in[129] ^ in2[129];
    assign G[96] = in[128] & in2[128];
    assign P[96] = in[128] ^ in2[128];
    assign G[97] = in[127] & in2[127];
    assign P[97] = in[127] ^ in2[127];
    assign G[98] = in[126] & in2[126];
    assign P[98] = in[126] ^ in2[126];
    assign G[99] = in[125] & in2[125];
    assign P[99] = in[125] ^ in2[125];
    assign G[100] = in[124] & in2[124];
    assign P[100] = in[124] ^ in2[124];
    assign G[101] = in[123] & in2[123];
    assign P[101] = in[123] ^ in2[123];
    assign G[102] = in[122] & in2[122];
    assign P[102] = in[122] ^ in2[122];
    assign G[103] = in[121] & in2[121];
    assign P[103] = in[121] ^ in2[121];
    assign G[104] = in[120] & in2[120];
    assign P[104] = in[120] ^ in2[120];
    assign G[105] = in[119] & in2[119];
    assign P[105] = in[119] ^ in2[119];
    assign G[106] = in[118] & in2[118];
    assign P[106] = in[118] ^ in2[118];
    assign G[107] = in[117] & in2[117];
    assign P[107] = in[117] ^ in2[117];
    assign G[108] = in[116] & in2[116];
    assign P[108] = in[116] ^ in2[116];
    assign G[109] = in[115] & in2[115];
    assign P[109] = in[115] ^ in2[115];
    assign G[110] = in[114] & in2[114];
    assign P[110] = in[114] ^ in2[114];
    assign G[111] = in[113] & in2[113];
    assign P[111] = in[113] ^ in2[113];
    assign G[112] = in[112] & in2[112];
    assign P[112] = in[112] ^ in2[112];
    assign G[113] = in[111] & in2[111];
    assign P[113] = in[111] ^ in2[111];
    assign G[114] = in[110] & in2[110];
    assign P[114] = in[110] ^ in2[110];
    assign G[115] = in[109] & in2[109];
    assign P[115] = in[109] ^ in2[109];
    assign G[116] = in[108] & in2[108];
    assign P[116] = in[108] ^ in2[108];
    assign G[117] = in[107] & in2[107];
    assign P[117] = in[107] ^ in2[107];
    assign G[118] = in[106] & in2[106];
    assign P[118] = in[106] ^ in2[106];
    assign G[119] = in[105] & in2[105];
    assign P[119] = in[105] ^ in2[105];
    assign G[120] = in[104] & in2[104];
    assign P[120] = in[104] ^ in2[104];
    assign G[121] = in[103] & in2[103];
    assign P[121] = in[103] ^ in2[103];
    assign G[122] = in[102] & in2[102];
    assign P[122] = in[102] ^ in2[102];
    assign G[123] = in[101] & in2[101];
    assign P[123] = in[101] ^ in2[101];
    assign G[124] = in[100] & in2[100];
    assign P[124] = in[100] ^ in2[100];
    assign G[125] = in[99] & in2[99];
    assign P[125] = in[99] ^ in2[99];
    assign G[126] = in[98] & in2[98];
    assign P[126] = in[98] ^ in2[98];
    assign G[127] = in[97] & in2[97];
    assign P[127] = in[97] ^ in2[97];
    assign G[128] = in[96] & in2[96];
    assign P[128] = in[96] ^ in2[96];
    assign G[129] = in[95] & in2[95];
    assign P[129] = in[95] ^ in2[95];
    assign G[130] = in[94] & in2[94];
    assign P[130] = in[94] ^ in2[94];
    assign G[131] = in[93] & in2[93];
    assign P[131] = in[93] ^ in2[93];
    assign G[132] = in[92] & in2[92];
    assign P[132] = in[92] ^ in2[92];
    assign G[133] = in[91] & in2[91];
    assign P[133] = in[91] ^ in2[91];
    assign G[134] = in[90] & in2[90];
    assign P[134] = in[90] ^ in2[90];
    assign G[135] = in[89] & in2[89];
    assign P[135] = in[89] ^ in2[89];
    assign G[136] = in[88] & in2[88];
    assign P[136] = in[88] ^ in2[88];
    assign G[137] = in[87] & in2[87];
    assign P[137] = in[87] ^ in2[87];
    assign G[138] = in[86] & in2[86];
    assign P[138] = in[86] ^ in2[86];
    assign G[139] = in[85] & in2[85];
    assign P[139] = in[85] ^ in2[85];
    assign G[140] = in[84] & in2[84];
    assign P[140] = in[84] ^ in2[84];
    assign G[141] = in[83] & in2[83];
    assign P[141] = in[83] ^ in2[83];
    assign G[142] = in[82] & in2[82];
    assign P[142] = in[82] ^ in2[82];
    assign G[143] = in[81] & in2[81];
    assign P[143] = in[81] ^ in2[81];
    assign G[144] = in[80] & in2[80];
    assign P[144] = in[80] ^ in2[80];
    assign G[145] = in[79] & in2[79];
    assign P[145] = in[79] ^ in2[79];
    assign G[146] = in[78] & in2[78];
    assign P[146] = in[78] ^ in2[78];
    assign G[147] = in[77] & in2[77];
    assign P[147] = in[77] ^ in2[77];
    assign G[148] = in[76] & in2[76];
    assign P[148] = in[76] ^ in2[76];
    assign G[149] = in[75] & in2[75];
    assign P[149] = in[75] ^ in2[75];
    assign G[150] = in[74] & in2[74];
    assign P[150] = in[74] ^ in2[74];
    assign G[151] = in[73] & in2[73];
    assign P[151] = in[73] ^ in2[73];
    assign G[152] = in[72] & in2[72];
    assign P[152] = in[72] ^ in2[72];
    assign G[153] = in[71] & in2[71];
    assign P[153] = in[71] ^ in2[71];
    assign G[154] = in[70] & in2[70];
    assign P[154] = in[70] ^ in2[70];
    assign G[155] = in[69] & in2[69];
    assign P[155] = in[69] ^ in2[69];
    assign G[156] = in[68] & in2[68];
    assign P[156] = in[68] ^ in2[68];
    assign G[157] = in[67] & in2[67];
    assign P[157] = in[67] ^ in2[67];
    assign G[158] = in[66] & in2[66];
    assign P[158] = in[66] ^ in2[66];
    assign G[159] = in[65] & in2[65];
    assign P[159] = in[65] ^ in2[65];
    assign G[160] = in[64] & in2[64];
    assign P[160] = in[64] ^ in2[64];
    assign G[161] = in[63] & in2[63];
    assign P[161] = in[63] ^ in2[63];
    assign G[162] = in[62] & in2[62];
    assign P[162] = in[62] ^ in2[62];
    assign G[163] = in[61] & in2[61];
    assign P[163] = in[61] ^ in2[61];
    assign G[164] = in[60] & in2[60];
    assign P[164] = in[60] ^ in2[60];
    assign G[165] = in[59] & in2[59];
    assign P[165] = in[59] ^ in2[59];
    assign G[166] = in[58] & in2[58];
    assign P[166] = in[58] ^ in2[58];
    assign G[167] = in[57] & in2[57];
    assign P[167] = in[57] ^ in2[57];
    assign G[168] = in[56] & in2[56];
    assign P[168] = in[56] ^ in2[56];
    assign G[169] = in[55] & in2[55];
    assign P[169] = in[55] ^ in2[55];
    assign G[170] = in[54] & in2[54];
    assign P[170] = in[54] ^ in2[54];
    assign G[171] = in[53] & in2[53];
    assign P[171] = in[53] ^ in2[53];
    assign G[172] = in[52] & in2[52];
    assign P[172] = in[52] ^ in2[52];
    assign G[173] = in[51] & in2[51];
    assign P[173] = in[51] ^ in2[51];
    assign G[174] = in[50] & in2[50];
    assign P[174] = in[50] ^ in2[50];
    assign G[175] = in[49] & in2[49];
    assign P[175] = in[49] ^ in2[49];
    assign G[176] = in[48] & in2[48];
    assign P[176] = in[48] ^ in2[48];
    assign G[177] = in[47] & in2[47];
    assign P[177] = in[47] ^ in2[47];
    assign G[178] = in[46] & in2[46];
    assign P[178] = in[46] ^ in2[46];
    assign G[179] = in[45] & in2[45];
    assign P[179] = in[45] ^ in2[45];
    assign G[180] = in[44] & in2[44];
    assign P[180] = in[44] ^ in2[44];
    assign G[181] = in[43] & in2[43];
    assign P[181] = in[43] ^ in2[43];
    assign G[182] = in[42] & in2[42];
    assign P[182] = in[42] ^ in2[42];
    assign G[183] = in[41] & in2[41];
    assign P[183] = in[41] ^ in2[41];
    assign G[184] = in[40] & in2[40];
    assign P[184] = in[40] ^ in2[40];
    assign G[185] = in[39] & in2[39];
    assign P[185] = in[39] ^ in2[39];
    assign G[186] = in[38] & in2[38];
    assign P[186] = in[38] ^ in2[38];
    assign G[187] = in[37] & in2[37];
    assign P[187] = in[37] ^ in2[37];
    assign G[188] = in[36] & in2[36];
    assign P[188] = in[36] ^ in2[36];
    assign G[189] = in[35] & in2[35];
    assign P[189] = in[35] ^ in2[35];
    assign G[190] = in[34] & in2[34];
    assign P[190] = in[34] ^ in2[34];
    assign G[191] = in[33] & in2[33];
    assign P[191] = in[33] ^ in2[33];
    assign G[192] = in[32] & in2[32];
    assign P[192] = in[32] ^ in2[32];
    assign G[193] = in[31] & in2[31];
    assign P[193] = in[31] ^ in2[31];
    assign G[194] = in[30] & in2[30];
    assign P[194] = in[30] ^ in2[30];
    assign G[195] = in[29] & in2[29];
    assign P[195] = in[29] ^ in2[29];
    assign G[196] = in[28] & in2[28];
    assign P[196] = in[28] ^ in2[28];
    assign G[197] = in[27] & in2[27];
    assign P[197] = in[27] ^ in2[27];
    assign G[198] = in[26] & in2[26];
    assign P[198] = in[26] ^ in2[26];
    assign G[199] = in[25] & in2[25];
    assign P[199] = in[25] ^ in2[25];
    assign G[200] = in[24] & in2[24];
    assign P[200] = in[24] ^ in2[24];
    assign G[201] = in[23] & in2[23];
    assign P[201] = in[23] ^ in2[23];
    assign G[202] = in[22] & in2[22];
    assign P[202] = in[22] ^ in2[22];
    assign G[203] = in[21] & in2[21];
    assign P[203] = in[21] ^ in2[21];
    assign G[204] = in[20] & in2[20];
    assign P[204] = in[20] ^ in2[20];
    assign G[205] = in[19] & in2[19];
    assign P[205] = in[19] ^ in2[19];
    assign G[206] = in[18] & in2[18];
    assign P[206] = in[18] ^ in2[18];
    assign G[207] = in[17] & in2[17];
    assign P[207] = in[17] ^ in2[17];
    assign G[208] = in[16] & in2[16];
    assign P[208] = in[16] ^ in2[16];
    assign G[209] = in[15] & in2[15];
    assign P[209] = in[15] ^ in2[15];
    assign G[210] = in[14] & in2[14];
    assign P[210] = in[14] ^ in2[14];
    assign G[211] = in[13] & in2[13];
    assign P[211] = in[13] ^ in2[13];
    assign G[212] = in[12] & in2[12];
    assign P[212] = in[12] ^ in2[12];
    assign G[213] = in[11] & in2[11];
    assign P[213] = in[11] ^ in2[11];
    assign G[214] = in[10] & in2[10];
    assign P[214] = in[10] ^ in2[10];
    assign G[215] = in[9] & in2[9];
    assign P[215] = in[9] ^ in2[9];
    assign G[216] = in[8] & in2[8];
    assign P[216] = in[8] ^ in2[8];
    assign G[217] = in[7] & in2[7];
    assign P[217] = in[7] ^ in2[7];
    assign G[218] = in[6] & in2[6];
    assign P[218] = in[6] ^ in2[6];
    assign G[219] = in[5] & in2[5];
    assign P[219] = in[5] ^ in2[5];
    assign G[220] = in[4] & in2[4];
    assign P[220] = in[4] ^ in2[4];
    assign G[221] = in[3] & in2[3];
    assign P[221] = in[3] ^ in2[3];
    assign G[222] = in[2] & in2[2];
    assign P[222] = in[2] ^ in2[2];
    assign G[223] = in[1] & in2[1];
    assign P[223] = in[1] ^ in2[1];
    assign G[224] = in[0] & in2[0];
    assign P[224] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign C[224] = G[223] | (P[223] & C[223]);
    assign cout = G[224] | (P[224] & C[224]);
    assign sum = P ^ C;
endmodule

module CLA224(output [223:0] sum, output cout, input [223:0] in1, input [223:0] in2;

    wire[223:0] G;
    wire[223:0] C;
    wire[223:0] P;

    assign G[0] = in[223] & in2[223];
    assign P[0] = in[223] ^ in2[223];
    assign G[1] = in[222] & in2[222];
    assign P[1] = in[222] ^ in2[222];
    assign G[2] = in[221] & in2[221];
    assign P[2] = in[221] ^ in2[221];
    assign G[3] = in[220] & in2[220];
    assign P[3] = in[220] ^ in2[220];
    assign G[4] = in[219] & in2[219];
    assign P[4] = in[219] ^ in2[219];
    assign G[5] = in[218] & in2[218];
    assign P[5] = in[218] ^ in2[218];
    assign G[6] = in[217] & in2[217];
    assign P[6] = in[217] ^ in2[217];
    assign G[7] = in[216] & in2[216];
    assign P[7] = in[216] ^ in2[216];
    assign G[8] = in[215] & in2[215];
    assign P[8] = in[215] ^ in2[215];
    assign G[9] = in[214] & in2[214];
    assign P[9] = in[214] ^ in2[214];
    assign G[10] = in[213] & in2[213];
    assign P[10] = in[213] ^ in2[213];
    assign G[11] = in[212] & in2[212];
    assign P[11] = in[212] ^ in2[212];
    assign G[12] = in[211] & in2[211];
    assign P[12] = in[211] ^ in2[211];
    assign G[13] = in[210] & in2[210];
    assign P[13] = in[210] ^ in2[210];
    assign G[14] = in[209] & in2[209];
    assign P[14] = in[209] ^ in2[209];
    assign G[15] = in[208] & in2[208];
    assign P[15] = in[208] ^ in2[208];
    assign G[16] = in[207] & in2[207];
    assign P[16] = in[207] ^ in2[207];
    assign G[17] = in[206] & in2[206];
    assign P[17] = in[206] ^ in2[206];
    assign G[18] = in[205] & in2[205];
    assign P[18] = in[205] ^ in2[205];
    assign G[19] = in[204] & in2[204];
    assign P[19] = in[204] ^ in2[204];
    assign G[20] = in[203] & in2[203];
    assign P[20] = in[203] ^ in2[203];
    assign G[21] = in[202] & in2[202];
    assign P[21] = in[202] ^ in2[202];
    assign G[22] = in[201] & in2[201];
    assign P[22] = in[201] ^ in2[201];
    assign G[23] = in[200] & in2[200];
    assign P[23] = in[200] ^ in2[200];
    assign G[24] = in[199] & in2[199];
    assign P[24] = in[199] ^ in2[199];
    assign G[25] = in[198] & in2[198];
    assign P[25] = in[198] ^ in2[198];
    assign G[26] = in[197] & in2[197];
    assign P[26] = in[197] ^ in2[197];
    assign G[27] = in[196] & in2[196];
    assign P[27] = in[196] ^ in2[196];
    assign G[28] = in[195] & in2[195];
    assign P[28] = in[195] ^ in2[195];
    assign G[29] = in[194] & in2[194];
    assign P[29] = in[194] ^ in2[194];
    assign G[30] = in[193] & in2[193];
    assign P[30] = in[193] ^ in2[193];
    assign G[31] = in[192] & in2[192];
    assign P[31] = in[192] ^ in2[192];
    assign G[32] = in[191] & in2[191];
    assign P[32] = in[191] ^ in2[191];
    assign G[33] = in[190] & in2[190];
    assign P[33] = in[190] ^ in2[190];
    assign G[34] = in[189] & in2[189];
    assign P[34] = in[189] ^ in2[189];
    assign G[35] = in[188] & in2[188];
    assign P[35] = in[188] ^ in2[188];
    assign G[36] = in[187] & in2[187];
    assign P[36] = in[187] ^ in2[187];
    assign G[37] = in[186] & in2[186];
    assign P[37] = in[186] ^ in2[186];
    assign G[38] = in[185] & in2[185];
    assign P[38] = in[185] ^ in2[185];
    assign G[39] = in[184] & in2[184];
    assign P[39] = in[184] ^ in2[184];
    assign G[40] = in[183] & in2[183];
    assign P[40] = in[183] ^ in2[183];
    assign G[41] = in[182] & in2[182];
    assign P[41] = in[182] ^ in2[182];
    assign G[42] = in[181] & in2[181];
    assign P[42] = in[181] ^ in2[181];
    assign G[43] = in[180] & in2[180];
    assign P[43] = in[180] ^ in2[180];
    assign G[44] = in[179] & in2[179];
    assign P[44] = in[179] ^ in2[179];
    assign G[45] = in[178] & in2[178];
    assign P[45] = in[178] ^ in2[178];
    assign G[46] = in[177] & in2[177];
    assign P[46] = in[177] ^ in2[177];
    assign G[47] = in[176] & in2[176];
    assign P[47] = in[176] ^ in2[176];
    assign G[48] = in[175] & in2[175];
    assign P[48] = in[175] ^ in2[175];
    assign G[49] = in[174] & in2[174];
    assign P[49] = in[174] ^ in2[174];
    assign G[50] = in[173] & in2[173];
    assign P[50] = in[173] ^ in2[173];
    assign G[51] = in[172] & in2[172];
    assign P[51] = in[172] ^ in2[172];
    assign G[52] = in[171] & in2[171];
    assign P[52] = in[171] ^ in2[171];
    assign G[53] = in[170] & in2[170];
    assign P[53] = in[170] ^ in2[170];
    assign G[54] = in[169] & in2[169];
    assign P[54] = in[169] ^ in2[169];
    assign G[55] = in[168] & in2[168];
    assign P[55] = in[168] ^ in2[168];
    assign G[56] = in[167] & in2[167];
    assign P[56] = in[167] ^ in2[167];
    assign G[57] = in[166] & in2[166];
    assign P[57] = in[166] ^ in2[166];
    assign G[58] = in[165] & in2[165];
    assign P[58] = in[165] ^ in2[165];
    assign G[59] = in[164] & in2[164];
    assign P[59] = in[164] ^ in2[164];
    assign G[60] = in[163] & in2[163];
    assign P[60] = in[163] ^ in2[163];
    assign G[61] = in[162] & in2[162];
    assign P[61] = in[162] ^ in2[162];
    assign G[62] = in[161] & in2[161];
    assign P[62] = in[161] ^ in2[161];
    assign G[63] = in[160] & in2[160];
    assign P[63] = in[160] ^ in2[160];
    assign G[64] = in[159] & in2[159];
    assign P[64] = in[159] ^ in2[159];
    assign G[65] = in[158] & in2[158];
    assign P[65] = in[158] ^ in2[158];
    assign G[66] = in[157] & in2[157];
    assign P[66] = in[157] ^ in2[157];
    assign G[67] = in[156] & in2[156];
    assign P[67] = in[156] ^ in2[156];
    assign G[68] = in[155] & in2[155];
    assign P[68] = in[155] ^ in2[155];
    assign G[69] = in[154] & in2[154];
    assign P[69] = in[154] ^ in2[154];
    assign G[70] = in[153] & in2[153];
    assign P[70] = in[153] ^ in2[153];
    assign G[71] = in[152] & in2[152];
    assign P[71] = in[152] ^ in2[152];
    assign G[72] = in[151] & in2[151];
    assign P[72] = in[151] ^ in2[151];
    assign G[73] = in[150] & in2[150];
    assign P[73] = in[150] ^ in2[150];
    assign G[74] = in[149] & in2[149];
    assign P[74] = in[149] ^ in2[149];
    assign G[75] = in[148] & in2[148];
    assign P[75] = in[148] ^ in2[148];
    assign G[76] = in[147] & in2[147];
    assign P[76] = in[147] ^ in2[147];
    assign G[77] = in[146] & in2[146];
    assign P[77] = in[146] ^ in2[146];
    assign G[78] = in[145] & in2[145];
    assign P[78] = in[145] ^ in2[145];
    assign G[79] = in[144] & in2[144];
    assign P[79] = in[144] ^ in2[144];
    assign G[80] = in[143] & in2[143];
    assign P[80] = in[143] ^ in2[143];
    assign G[81] = in[142] & in2[142];
    assign P[81] = in[142] ^ in2[142];
    assign G[82] = in[141] & in2[141];
    assign P[82] = in[141] ^ in2[141];
    assign G[83] = in[140] & in2[140];
    assign P[83] = in[140] ^ in2[140];
    assign G[84] = in[139] & in2[139];
    assign P[84] = in[139] ^ in2[139];
    assign G[85] = in[138] & in2[138];
    assign P[85] = in[138] ^ in2[138];
    assign G[86] = in[137] & in2[137];
    assign P[86] = in[137] ^ in2[137];
    assign G[87] = in[136] & in2[136];
    assign P[87] = in[136] ^ in2[136];
    assign G[88] = in[135] & in2[135];
    assign P[88] = in[135] ^ in2[135];
    assign G[89] = in[134] & in2[134];
    assign P[89] = in[134] ^ in2[134];
    assign G[90] = in[133] & in2[133];
    assign P[90] = in[133] ^ in2[133];
    assign G[91] = in[132] & in2[132];
    assign P[91] = in[132] ^ in2[132];
    assign G[92] = in[131] & in2[131];
    assign P[92] = in[131] ^ in2[131];
    assign G[93] = in[130] & in2[130];
    assign P[93] = in[130] ^ in2[130];
    assign G[94] = in[129] & in2[129];
    assign P[94] = in[129] ^ in2[129];
    assign G[95] = in[128] & in2[128];
    assign P[95] = in[128] ^ in2[128];
    assign G[96] = in[127] & in2[127];
    assign P[96] = in[127] ^ in2[127];
    assign G[97] = in[126] & in2[126];
    assign P[97] = in[126] ^ in2[126];
    assign G[98] = in[125] & in2[125];
    assign P[98] = in[125] ^ in2[125];
    assign G[99] = in[124] & in2[124];
    assign P[99] = in[124] ^ in2[124];
    assign G[100] = in[123] & in2[123];
    assign P[100] = in[123] ^ in2[123];
    assign G[101] = in[122] & in2[122];
    assign P[101] = in[122] ^ in2[122];
    assign G[102] = in[121] & in2[121];
    assign P[102] = in[121] ^ in2[121];
    assign G[103] = in[120] & in2[120];
    assign P[103] = in[120] ^ in2[120];
    assign G[104] = in[119] & in2[119];
    assign P[104] = in[119] ^ in2[119];
    assign G[105] = in[118] & in2[118];
    assign P[105] = in[118] ^ in2[118];
    assign G[106] = in[117] & in2[117];
    assign P[106] = in[117] ^ in2[117];
    assign G[107] = in[116] & in2[116];
    assign P[107] = in[116] ^ in2[116];
    assign G[108] = in[115] & in2[115];
    assign P[108] = in[115] ^ in2[115];
    assign G[109] = in[114] & in2[114];
    assign P[109] = in[114] ^ in2[114];
    assign G[110] = in[113] & in2[113];
    assign P[110] = in[113] ^ in2[113];
    assign G[111] = in[112] & in2[112];
    assign P[111] = in[112] ^ in2[112];
    assign G[112] = in[111] & in2[111];
    assign P[112] = in[111] ^ in2[111];
    assign G[113] = in[110] & in2[110];
    assign P[113] = in[110] ^ in2[110];
    assign G[114] = in[109] & in2[109];
    assign P[114] = in[109] ^ in2[109];
    assign G[115] = in[108] & in2[108];
    assign P[115] = in[108] ^ in2[108];
    assign G[116] = in[107] & in2[107];
    assign P[116] = in[107] ^ in2[107];
    assign G[117] = in[106] & in2[106];
    assign P[117] = in[106] ^ in2[106];
    assign G[118] = in[105] & in2[105];
    assign P[118] = in[105] ^ in2[105];
    assign G[119] = in[104] & in2[104];
    assign P[119] = in[104] ^ in2[104];
    assign G[120] = in[103] & in2[103];
    assign P[120] = in[103] ^ in2[103];
    assign G[121] = in[102] & in2[102];
    assign P[121] = in[102] ^ in2[102];
    assign G[122] = in[101] & in2[101];
    assign P[122] = in[101] ^ in2[101];
    assign G[123] = in[100] & in2[100];
    assign P[123] = in[100] ^ in2[100];
    assign G[124] = in[99] & in2[99];
    assign P[124] = in[99] ^ in2[99];
    assign G[125] = in[98] & in2[98];
    assign P[125] = in[98] ^ in2[98];
    assign G[126] = in[97] & in2[97];
    assign P[126] = in[97] ^ in2[97];
    assign G[127] = in[96] & in2[96];
    assign P[127] = in[96] ^ in2[96];
    assign G[128] = in[95] & in2[95];
    assign P[128] = in[95] ^ in2[95];
    assign G[129] = in[94] & in2[94];
    assign P[129] = in[94] ^ in2[94];
    assign G[130] = in[93] & in2[93];
    assign P[130] = in[93] ^ in2[93];
    assign G[131] = in[92] & in2[92];
    assign P[131] = in[92] ^ in2[92];
    assign G[132] = in[91] & in2[91];
    assign P[132] = in[91] ^ in2[91];
    assign G[133] = in[90] & in2[90];
    assign P[133] = in[90] ^ in2[90];
    assign G[134] = in[89] & in2[89];
    assign P[134] = in[89] ^ in2[89];
    assign G[135] = in[88] & in2[88];
    assign P[135] = in[88] ^ in2[88];
    assign G[136] = in[87] & in2[87];
    assign P[136] = in[87] ^ in2[87];
    assign G[137] = in[86] & in2[86];
    assign P[137] = in[86] ^ in2[86];
    assign G[138] = in[85] & in2[85];
    assign P[138] = in[85] ^ in2[85];
    assign G[139] = in[84] & in2[84];
    assign P[139] = in[84] ^ in2[84];
    assign G[140] = in[83] & in2[83];
    assign P[140] = in[83] ^ in2[83];
    assign G[141] = in[82] & in2[82];
    assign P[141] = in[82] ^ in2[82];
    assign G[142] = in[81] & in2[81];
    assign P[142] = in[81] ^ in2[81];
    assign G[143] = in[80] & in2[80];
    assign P[143] = in[80] ^ in2[80];
    assign G[144] = in[79] & in2[79];
    assign P[144] = in[79] ^ in2[79];
    assign G[145] = in[78] & in2[78];
    assign P[145] = in[78] ^ in2[78];
    assign G[146] = in[77] & in2[77];
    assign P[146] = in[77] ^ in2[77];
    assign G[147] = in[76] & in2[76];
    assign P[147] = in[76] ^ in2[76];
    assign G[148] = in[75] & in2[75];
    assign P[148] = in[75] ^ in2[75];
    assign G[149] = in[74] & in2[74];
    assign P[149] = in[74] ^ in2[74];
    assign G[150] = in[73] & in2[73];
    assign P[150] = in[73] ^ in2[73];
    assign G[151] = in[72] & in2[72];
    assign P[151] = in[72] ^ in2[72];
    assign G[152] = in[71] & in2[71];
    assign P[152] = in[71] ^ in2[71];
    assign G[153] = in[70] & in2[70];
    assign P[153] = in[70] ^ in2[70];
    assign G[154] = in[69] & in2[69];
    assign P[154] = in[69] ^ in2[69];
    assign G[155] = in[68] & in2[68];
    assign P[155] = in[68] ^ in2[68];
    assign G[156] = in[67] & in2[67];
    assign P[156] = in[67] ^ in2[67];
    assign G[157] = in[66] & in2[66];
    assign P[157] = in[66] ^ in2[66];
    assign G[158] = in[65] & in2[65];
    assign P[158] = in[65] ^ in2[65];
    assign G[159] = in[64] & in2[64];
    assign P[159] = in[64] ^ in2[64];
    assign G[160] = in[63] & in2[63];
    assign P[160] = in[63] ^ in2[63];
    assign G[161] = in[62] & in2[62];
    assign P[161] = in[62] ^ in2[62];
    assign G[162] = in[61] & in2[61];
    assign P[162] = in[61] ^ in2[61];
    assign G[163] = in[60] & in2[60];
    assign P[163] = in[60] ^ in2[60];
    assign G[164] = in[59] & in2[59];
    assign P[164] = in[59] ^ in2[59];
    assign G[165] = in[58] & in2[58];
    assign P[165] = in[58] ^ in2[58];
    assign G[166] = in[57] & in2[57];
    assign P[166] = in[57] ^ in2[57];
    assign G[167] = in[56] & in2[56];
    assign P[167] = in[56] ^ in2[56];
    assign G[168] = in[55] & in2[55];
    assign P[168] = in[55] ^ in2[55];
    assign G[169] = in[54] & in2[54];
    assign P[169] = in[54] ^ in2[54];
    assign G[170] = in[53] & in2[53];
    assign P[170] = in[53] ^ in2[53];
    assign G[171] = in[52] & in2[52];
    assign P[171] = in[52] ^ in2[52];
    assign G[172] = in[51] & in2[51];
    assign P[172] = in[51] ^ in2[51];
    assign G[173] = in[50] & in2[50];
    assign P[173] = in[50] ^ in2[50];
    assign G[174] = in[49] & in2[49];
    assign P[174] = in[49] ^ in2[49];
    assign G[175] = in[48] & in2[48];
    assign P[175] = in[48] ^ in2[48];
    assign G[176] = in[47] & in2[47];
    assign P[176] = in[47] ^ in2[47];
    assign G[177] = in[46] & in2[46];
    assign P[177] = in[46] ^ in2[46];
    assign G[178] = in[45] & in2[45];
    assign P[178] = in[45] ^ in2[45];
    assign G[179] = in[44] & in2[44];
    assign P[179] = in[44] ^ in2[44];
    assign G[180] = in[43] & in2[43];
    assign P[180] = in[43] ^ in2[43];
    assign G[181] = in[42] & in2[42];
    assign P[181] = in[42] ^ in2[42];
    assign G[182] = in[41] & in2[41];
    assign P[182] = in[41] ^ in2[41];
    assign G[183] = in[40] & in2[40];
    assign P[183] = in[40] ^ in2[40];
    assign G[184] = in[39] & in2[39];
    assign P[184] = in[39] ^ in2[39];
    assign G[185] = in[38] & in2[38];
    assign P[185] = in[38] ^ in2[38];
    assign G[186] = in[37] & in2[37];
    assign P[186] = in[37] ^ in2[37];
    assign G[187] = in[36] & in2[36];
    assign P[187] = in[36] ^ in2[36];
    assign G[188] = in[35] & in2[35];
    assign P[188] = in[35] ^ in2[35];
    assign G[189] = in[34] & in2[34];
    assign P[189] = in[34] ^ in2[34];
    assign G[190] = in[33] & in2[33];
    assign P[190] = in[33] ^ in2[33];
    assign G[191] = in[32] & in2[32];
    assign P[191] = in[32] ^ in2[32];
    assign G[192] = in[31] & in2[31];
    assign P[192] = in[31] ^ in2[31];
    assign G[193] = in[30] & in2[30];
    assign P[193] = in[30] ^ in2[30];
    assign G[194] = in[29] & in2[29];
    assign P[194] = in[29] ^ in2[29];
    assign G[195] = in[28] & in2[28];
    assign P[195] = in[28] ^ in2[28];
    assign G[196] = in[27] & in2[27];
    assign P[196] = in[27] ^ in2[27];
    assign G[197] = in[26] & in2[26];
    assign P[197] = in[26] ^ in2[26];
    assign G[198] = in[25] & in2[25];
    assign P[198] = in[25] ^ in2[25];
    assign G[199] = in[24] & in2[24];
    assign P[199] = in[24] ^ in2[24];
    assign G[200] = in[23] & in2[23];
    assign P[200] = in[23] ^ in2[23];
    assign G[201] = in[22] & in2[22];
    assign P[201] = in[22] ^ in2[22];
    assign G[202] = in[21] & in2[21];
    assign P[202] = in[21] ^ in2[21];
    assign G[203] = in[20] & in2[20];
    assign P[203] = in[20] ^ in2[20];
    assign G[204] = in[19] & in2[19];
    assign P[204] = in[19] ^ in2[19];
    assign G[205] = in[18] & in2[18];
    assign P[205] = in[18] ^ in2[18];
    assign G[206] = in[17] & in2[17];
    assign P[206] = in[17] ^ in2[17];
    assign G[207] = in[16] & in2[16];
    assign P[207] = in[16] ^ in2[16];
    assign G[208] = in[15] & in2[15];
    assign P[208] = in[15] ^ in2[15];
    assign G[209] = in[14] & in2[14];
    assign P[209] = in[14] ^ in2[14];
    assign G[210] = in[13] & in2[13];
    assign P[210] = in[13] ^ in2[13];
    assign G[211] = in[12] & in2[12];
    assign P[211] = in[12] ^ in2[12];
    assign G[212] = in[11] & in2[11];
    assign P[212] = in[11] ^ in2[11];
    assign G[213] = in[10] & in2[10];
    assign P[213] = in[10] ^ in2[10];
    assign G[214] = in[9] & in2[9];
    assign P[214] = in[9] ^ in2[9];
    assign G[215] = in[8] & in2[8];
    assign P[215] = in[8] ^ in2[8];
    assign G[216] = in[7] & in2[7];
    assign P[216] = in[7] ^ in2[7];
    assign G[217] = in[6] & in2[6];
    assign P[217] = in[6] ^ in2[6];
    assign G[218] = in[5] & in2[5];
    assign P[218] = in[5] ^ in2[5];
    assign G[219] = in[4] & in2[4];
    assign P[219] = in[4] ^ in2[4];
    assign G[220] = in[3] & in2[3];
    assign P[220] = in[3] ^ in2[3];
    assign G[221] = in[2] & in2[2];
    assign P[221] = in[2] ^ in2[2];
    assign G[222] = in[1] & in2[1];
    assign P[222] = in[1] ^ in2[1];
    assign G[223] = in[0] & in2[0];
    assign P[223] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign C[223] = G[222] | (P[222] & C[222]);
    assign cout = G[223] | (P[223] & C[223]);
    assign sum = P ^ C;
endmodule

module CLA223(output [222:0] sum, output cout, input [222:0] in1, input [222:0] in2;

    wire[222:0] G;
    wire[222:0] C;
    wire[222:0] P;

    assign G[0] = in[222] & in2[222];
    assign P[0] = in[222] ^ in2[222];
    assign G[1] = in[221] & in2[221];
    assign P[1] = in[221] ^ in2[221];
    assign G[2] = in[220] & in2[220];
    assign P[2] = in[220] ^ in2[220];
    assign G[3] = in[219] & in2[219];
    assign P[3] = in[219] ^ in2[219];
    assign G[4] = in[218] & in2[218];
    assign P[4] = in[218] ^ in2[218];
    assign G[5] = in[217] & in2[217];
    assign P[5] = in[217] ^ in2[217];
    assign G[6] = in[216] & in2[216];
    assign P[6] = in[216] ^ in2[216];
    assign G[7] = in[215] & in2[215];
    assign P[7] = in[215] ^ in2[215];
    assign G[8] = in[214] & in2[214];
    assign P[8] = in[214] ^ in2[214];
    assign G[9] = in[213] & in2[213];
    assign P[9] = in[213] ^ in2[213];
    assign G[10] = in[212] & in2[212];
    assign P[10] = in[212] ^ in2[212];
    assign G[11] = in[211] & in2[211];
    assign P[11] = in[211] ^ in2[211];
    assign G[12] = in[210] & in2[210];
    assign P[12] = in[210] ^ in2[210];
    assign G[13] = in[209] & in2[209];
    assign P[13] = in[209] ^ in2[209];
    assign G[14] = in[208] & in2[208];
    assign P[14] = in[208] ^ in2[208];
    assign G[15] = in[207] & in2[207];
    assign P[15] = in[207] ^ in2[207];
    assign G[16] = in[206] & in2[206];
    assign P[16] = in[206] ^ in2[206];
    assign G[17] = in[205] & in2[205];
    assign P[17] = in[205] ^ in2[205];
    assign G[18] = in[204] & in2[204];
    assign P[18] = in[204] ^ in2[204];
    assign G[19] = in[203] & in2[203];
    assign P[19] = in[203] ^ in2[203];
    assign G[20] = in[202] & in2[202];
    assign P[20] = in[202] ^ in2[202];
    assign G[21] = in[201] & in2[201];
    assign P[21] = in[201] ^ in2[201];
    assign G[22] = in[200] & in2[200];
    assign P[22] = in[200] ^ in2[200];
    assign G[23] = in[199] & in2[199];
    assign P[23] = in[199] ^ in2[199];
    assign G[24] = in[198] & in2[198];
    assign P[24] = in[198] ^ in2[198];
    assign G[25] = in[197] & in2[197];
    assign P[25] = in[197] ^ in2[197];
    assign G[26] = in[196] & in2[196];
    assign P[26] = in[196] ^ in2[196];
    assign G[27] = in[195] & in2[195];
    assign P[27] = in[195] ^ in2[195];
    assign G[28] = in[194] & in2[194];
    assign P[28] = in[194] ^ in2[194];
    assign G[29] = in[193] & in2[193];
    assign P[29] = in[193] ^ in2[193];
    assign G[30] = in[192] & in2[192];
    assign P[30] = in[192] ^ in2[192];
    assign G[31] = in[191] & in2[191];
    assign P[31] = in[191] ^ in2[191];
    assign G[32] = in[190] & in2[190];
    assign P[32] = in[190] ^ in2[190];
    assign G[33] = in[189] & in2[189];
    assign P[33] = in[189] ^ in2[189];
    assign G[34] = in[188] & in2[188];
    assign P[34] = in[188] ^ in2[188];
    assign G[35] = in[187] & in2[187];
    assign P[35] = in[187] ^ in2[187];
    assign G[36] = in[186] & in2[186];
    assign P[36] = in[186] ^ in2[186];
    assign G[37] = in[185] & in2[185];
    assign P[37] = in[185] ^ in2[185];
    assign G[38] = in[184] & in2[184];
    assign P[38] = in[184] ^ in2[184];
    assign G[39] = in[183] & in2[183];
    assign P[39] = in[183] ^ in2[183];
    assign G[40] = in[182] & in2[182];
    assign P[40] = in[182] ^ in2[182];
    assign G[41] = in[181] & in2[181];
    assign P[41] = in[181] ^ in2[181];
    assign G[42] = in[180] & in2[180];
    assign P[42] = in[180] ^ in2[180];
    assign G[43] = in[179] & in2[179];
    assign P[43] = in[179] ^ in2[179];
    assign G[44] = in[178] & in2[178];
    assign P[44] = in[178] ^ in2[178];
    assign G[45] = in[177] & in2[177];
    assign P[45] = in[177] ^ in2[177];
    assign G[46] = in[176] & in2[176];
    assign P[46] = in[176] ^ in2[176];
    assign G[47] = in[175] & in2[175];
    assign P[47] = in[175] ^ in2[175];
    assign G[48] = in[174] & in2[174];
    assign P[48] = in[174] ^ in2[174];
    assign G[49] = in[173] & in2[173];
    assign P[49] = in[173] ^ in2[173];
    assign G[50] = in[172] & in2[172];
    assign P[50] = in[172] ^ in2[172];
    assign G[51] = in[171] & in2[171];
    assign P[51] = in[171] ^ in2[171];
    assign G[52] = in[170] & in2[170];
    assign P[52] = in[170] ^ in2[170];
    assign G[53] = in[169] & in2[169];
    assign P[53] = in[169] ^ in2[169];
    assign G[54] = in[168] & in2[168];
    assign P[54] = in[168] ^ in2[168];
    assign G[55] = in[167] & in2[167];
    assign P[55] = in[167] ^ in2[167];
    assign G[56] = in[166] & in2[166];
    assign P[56] = in[166] ^ in2[166];
    assign G[57] = in[165] & in2[165];
    assign P[57] = in[165] ^ in2[165];
    assign G[58] = in[164] & in2[164];
    assign P[58] = in[164] ^ in2[164];
    assign G[59] = in[163] & in2[163];
    assign P[59] = in[163] ^ in2[163];
    assign G[60] = in[162] & in2[162];
    assign P[60] = in[162] ^ in2[162];
    assign G[61] = in[161] & in2[161];
    assign P[61] = in[161] ^ in2[161];
    assign G[62] = in[160] & in2[160];
    assign P[62] = in[160] ^ in2[160];
    assign G[63] = in[159] & in2[159];
    assign P[63] = in[159] ^ in2[159];
    assign G[64] = in[158] & in2[158];
    assign P[64] = in[158] ^ in2[158];
    assign G[65] = in[157] & in2[157];
    assign P[65] = in[157] ^ in2[157];
    assign G[66] = in[156] & in2[156];
    assign P[66] = in[156] ^ in2[156];
    assign G[67] = in[155] & in2[155];
    assign P[67] = in[155] ^ in2[155];
    assign G[68] = in[154] & in2[154];
    assign P[68] = in[154] ^ in2[154];
    assign G[69] = in[153] & in2[153];
    assign P[69] = in[153] ^ in2[153];
    assign G[70] = in[152] & in2[152];
    assign P[70] = in[152] ^ in2[152];
    assign G[71] = in[151] & in2[151];
    assign P[71] = in[151] ^ in2[151];
    assign G[72] = in[150] & in2[150];
    assign P[72] = in[150] ^ in2[150];
    assign G[73] = in[149] & in2[149];
    assign P[73] = in[149] ^ in2[149];
    assign G[74] = in[148] & in2[148];
    assign P[74] = in[148] ^ in2[148];
    assign G[75] = in[147] & in2[147];
    assign P[75] = in[147] ^ in2[147];
    assign G[76] = in[146] & in2[146];
    assign P[76] = in[146] ^ in2[146];
    assign G[77] = in[145] & in2[145];
    assign P[77] = in[145] ^ in2[145];
    assign G[78] = in[144] & in2[144];
    assign P[78] = in[144] ^ in2[144];
    assign G[79] = in[143] & in2[143];
    assign P[79] = in[143] ^ in2[143];
    assign G[80] = in[142] & in2[142];
    assign P[80] = in[142] ^ in2[142];
    assign G[81] = in[141] & in2[141];
    assign P[81] = in[141] ^ in2[141];
    assign G[82] = in[140] & in2[140];
    assign P[82] = in[140] ^ in2[140];
    assign G[83] = in[139] & in2[139];
    assign P[83] = in[139] ^ in2[139];
    assign G[84] = in[138] & in2[138];
    assign P[84] = in[138] ^ in2[138];
    assign G[85] = in[137] & in2[137];
    assign P[85] = in[137] ^ in2[137];
    assign G[86] = in[136] & in2[136];
    assign P[86] = in[136] ^ in2[136];
    assign G[87] = in[135] & in2[135];
    assign P[87] = in[135] ^ in2[135];
    assign G[88] = in[134] & in2[134];
    assign P[88] = in[134] ^ in2[134];
    assign G[89] = in[133] & in2[133];
    assign P[89] = in[133] ^ in2[133];
    assign G[90] = in[132] & in2[132];
    assign P[90] = in[132] ^ in2[132];
    assign G[91] = in[131] & in2[131];
    assign P[91] = in[131] ^ in2[131];
    assign G[92] = in[130] & in2[130];
    assign P[92] = in[130] ^ in2[130];
    assign G[93] = in[129] & in2[129];
    assign P[93] = in[129] ^ in2[129];
    assign G[94] = in[128] & in2[128];
    assign P[94] = in[128] ^ in2[128];
    assign G[95] = in[127] & in2[127];
    assign P[95] = in[127] ^ in2[127];
    assign G[96] = in[126] & in2[126];
    assign P[96] = in[126] ^ in2[126];
    assign G[97] = in[125] & in2[125];
    assign P[97] = in[125] ^ in2[125];
    assign G[98] = in[124] & in2[124];
    assign P[98] = in[124] ^ in2[124];
    assign G[99] = in[123] & in2[123];
    assign P[99] = in[123] ^ in2[123];
    assign G[100] = in[122] & in2[122];
    assign P[100] = in[122] ^ in2[122];
    assign G[101] = in[121] & in2[121];
    assign P[101] = in[121] ^ in2[121];
    assign G[102] = in[120] & in2[120];
    assign P[102] = in[120] ^ in2[120];
    assign G[103] = in[119] & in2[119];
    assign P[103] = in[119] ^ in2[119];
    assign G[104] = in[118] & in2[118];
    assign P[104] = in[118] ^ in2[118];
    assign G[105] = in[117] & in2[117];
    assign P[105] = in[117] ^ in2[117];
    assign G[106] = in[116] & in2[116];
    assign P[106] = in[116] ^ in2[116];
    assign G[107] = in[115] & in2[115];
    assign P[107] = in[115] ^ in2[115];
    assign G[108] = in[114] & in2[114];
    assign P[108] = in[114] ^ in2[114];
    assign G[109] = in[113] & in2[113];
    assign P[109] = in[113] ^ in2[113];
    assign G[110] = in[112] & in2[112];
    assign P[110] = in[112] ^ in2[112];
    assign G[111] = in[111] & in2[111];
    assign P[111] = in[111] ^ in2[111];
    assign G[112] = in[110] & in2[110];
    assign P[112] = in[110] ^ in2[110];
    assign G[113] = in[109] & in2[109];
    assign P[113] = in[109] ^ in2[109];
    assign G[114] = in[108] & in2[108];
    assign P[114] = in[108] ^ in2[108];
    assign G[115] = in[107] & in2[107];
    assign P[115] = in[107] ^ in2[107];
    assign G[116] = in[106] & in2[106];
    assign P[116] = in[106] ^ in2[106];
    assign G[117] = in[105] & in2[105];
    assign P[117] = in[105] ^ in2[105];
    assign G[118] = in[104] & in2[104];
    assign P[118] = in[104] ^ in2[104];
    assign G[119] = in[103] & in2[103];
    assign P[119] = in[103] ^ in2[103];
    assign G[120] = in[102] & in2[102];
    assign P[120] = in[102] ^ in2[102];
    assign G[121] = in[101] & in2[101];
    assign P[121] = in[101] ^ in2[101];
    assign G[122] = in[100] & in2[100];
    assign P[122] = in[100] ^ in2[100];
    assign G[123] = in[99] & in2[99];
    assign P[123] = in[99] ^ in2[99];
    assign G[124] = in[98] & in2[98];
    assign P[124] = in[98] ^ in2[98];
    assign G[125] = in[97] & in2[97];
    assign P[125] = in[97] ^ in2[97];
    assign G[126] = in[96] & in2[96];
    assign P[126] = in[96] ^ in2[96];
    assign G[127] = in[95] & in2[95];
    assign P[127] = in[95] ^ in2[95];
    assign G[128] = in[94] & in2[94];
    assign P[128] = in[94] ^ in2[94];
    assign G[129] = in[93] & in2[93];
    assign P[129] = in[93] ^ in2[93];
    assign G[130] = in[92] & in2[92];
    assign P[130] = in[92] ^ in2[92];
    assign G[131] = in[91] & in2[91];
    assign P[131] = in[91] ^ in2[91];
    assign G[132] = in[90] & in2[90];
    assign P[132] = in[90] ^ in2[90];
    assign G[133] = in[89] & in2[89];
    assign P[133] = in[89] ^ in2[89];
    assign G[134] = in[88] & in2[88];
    assign P[134] = in[88] ^ in2[88];
    assign G[135] = in[87] & in2[87];
    assign P[135] = in[87] ^ in2[87];
    assign G[136] = in[86] & in2[86];
    assign P[136] = in[86] ^ in2[86];
    assign G[137] = in[85] & in2[85];
    assign P[137] = in[85] ^ in2[85];
    assign G[138] = in[84] & in2[84];
    assign P[138] = in[84] ^ in2[84];
    assign G[139] = in[83] & in2[83];
    assign P[139] = in[83] ^ in2[83];
    assign G[140] = in[82] & in2[82];
    assign P[140] = in[82] ^ in2[82];
    assign G[141] = in[81] & in2[81];
    assign P[141] = in[81] ^ in2[81];
    assign G[142] = in[80] & in2[80];
    assign P[142] = in[80] ^ in2[80];
    assign G[143] = in[79] & in2[79];
    assign P[143] = in[79] ^ in2[79];
    assign G[144] = in[78] & in2[78];
    assign P[144] = in[78] ^ in2[78];
    assign G[145] = in[77] & in2[77];
    assign P[145] = in[77] ^ in2[77];
    assign G[146] = in[76] & in2[76];
    assign P[146] = in[76] ^ in2[76];
    assign G[147] = in[75] & in2[75];
    assign P[147] = in[75] ^ in2[75];
    assign G[148] = in[74] & in2[74];
    assign P[148] = in[74] ^ in2[74];
    assign G[149] = in[73] & in2[73];
    assign P[149] = in[73] ^ in2[73];
    assign G[150] = in[72] & in2[72];
    assign P[150] = in[72] ^ in2[72];
    assign G[151] = in[71] & in2[71];
    assign P[151] = in[71] ^ in2[71];
    assign G[152] = in[70] & in2[70];
    assign P[152] = in[70] ^ in2[70];
    assign G[153] = in[69] & in2[69];
    assign P[153] = in[69] ^ in2[69];
    assign G[154] = in[68] & in2[68];
    assign P[154] = in[68] ^ in2[68];
    assign G[155] = in[67] & in2[67];
    assign P[155] = in[67] ^ in2[67];
    assign G[156] = in[66] & in2[66];
    assign P[156] = in[66] ^ in2[66];
    assign G[157] = in[65] & in2[65];
    assign P[157] = in[65] ^ in2[65];
    assign G[158] = in[64] & in2[64];
    assign P[158] = in[64] ^ in2[64];
    assign G[159] = in[63] & in2[63];
    assign P[159] = in[63] ^ in2[63];
    assign G[160] = in[62] & in2[62];
    assign P[160] = in[62] ^ in2[62];
    assign G[161] = in[61] & in2[61];
    assign P[161] = in[61] ^ in2[61];
    assign G[162] = in[60] & in2[60];
    assign P[162] = in[60] ^ in2[60];
    assign G[163] = in[59] & in2[59];
    assign P[163] = in[59] ^ in2[59];
    assign G[164] = in[58] & in2[58];
    assign P[164] = in[58] ^ in2[58];
    assign G[165] = in[57] & in2[57];
    assign P[165] = in[57] ^ in2[57];
    assign G[166] = in[56] & in2[56];
    assign P[166] = in[56] ^ in2[56];
    assign G[167] = in[55] & in2[55];
    assign P[167] = in[55] ^ in2[55];
    assign G[168] = in[54] & in2[54];
    assign P[168] = in[54] ^ in2[54];
    assign G[169] = in[53] & in2[53];
    assign P[169] = in[53] ^ in2[53];
    assign G[170] = in[52] & in2[52];
    assign P[170] = in[52] ^ in2[52];
    assign G[171] = in[51] & in2[51];
    assign P[171] = in[51] ^ in2[51];
    assign G[172] = in[50] & in2[50];
    assign P[172] = in[50] ^ in2[50];
    assign G[173] = in[49] & in2[49];
    assign P[173] = in[49] ^ in2[49];
    assign G[174] = in[48] & in2[48];
    assign P[174] = in[48] ^ in2[48];
    assign G[175] = in[47] & in2[47];
    assign P[175] = in[47] ^ in2[47];
    assign G[176] = in[46] & in2[46];
    assign P[176] = in[46] ^ in2[46];
    assign G[177] = in[45] & in2[45];
    assign P[177] = in[45] ^ in2[45];
    assign G[178] = in[44] & in2[44];
    assign P[178] = in[44] ^ in2[44];
    assign G[179] = in[43] & in2[43];
    assign P[179] = in[43] ^ in2[43];
    assign G[180] = in[42] & in2[42];
    assign P[180] = in[42] ^ in2[42];
    assign G[181] = in[41] & in2[41];
    assign P[181] = in[41] ^ in2[41];
    assign G[182] = in[40] & in2[40];
    assign P[182] = in[40] ^ in2[40];
    assign G[183] = in[39] & in2[39];
    assign P[183] = in[39] ^ in2[39];
    assign G[184] = in[38] & in2[38];
    assign P[184] = in[38] ^ in2[38];
    assign G[185] = in[37] & in2[37];
    assign P[185] = in[37] ^ in2[37];
    assign G[186] = in[36] & in2[36];
    assign P[186] = in[36] ^ in2[36];
    assign G[187] = in[35] & in2[35];
    assign P[187] = in[35] ^ in2[35];
    assign G[188] = in[34] & in2[34];
    assign P[188] = in[34] ^ in2[34];
    assign G[189] = in[33] & in2[33];
    assign P[189] = in[33] ^ in2[33];
    assign G[190] = in[32] & in2[32];
    assign P[190] = in[32] ^ in2[32];
    assign G[191] = in[31] & in2[31];
    assign P[191] = in[31] ^ in2[31];
    assign G[192] = in[30] & in2[30];
    assign P[192] = in[30] ^ in2[30];
    assign G[193] = in[29] & in2[29];
    assign P[193] = in[29] ^ in2[29];
    assign G[194] = in[28] & in2[28];
    assign P[194] = in[28] ^ in2[28];
    assign G[195] = in[27] & in2[27];
    assign P[195] = in[27] ^ in2[27];
    assign G[196] = in[26] & in2[26];
    assign P[196] = in[26] ^ in2[26];
    assign G[197] = in[25] & in2[25];
    assign P[197] = in[25] ^ in2[25];
    assign G[198] = in[24] & in2[24];
    assign P[198] = in[24] ^ in2[24];
    assign G[199] = in[23] & in2[23];
    assign P[199] = in[23] ^ in2[23];
    assign G[200] = in[22] & in2[22];
    assign P[200] = in[22] ^ in2[22];
    assign G[201] = in[21] & in2[21];
    assign P[201] = in[21] ^ in2[21];
    assign G[202] = in[20] & in2[20];
    assign P[202] = in[20] ^ in2[20];
    assign G[203] = in[19] & in2[19];
    assign P[203] = in[19] ^ in2[19];
    assign G[204] = in[18] & in2[18];
    assign P[204] = in[18] ^ in2[18];
    assign G[205] = in[17] & in2[17];
    assign P[205] = in[17] ^ in2[17];
    assign G[206] = in[16] & in2[16];
    assign P[206] = in[16] ^ in2[16];
    assign G[207] = in[15] & in2[15];
    assign P[207] = in[15] ^ in2[15];
    assign G[208] = in[14] & in2[14];
    assign P[208] = in[14] ^ in2[14];
    assign G[209] = in[13] & in2[13];
    assign P[209] = in[13] ^ in2[13];
    assign G[210] = in[12] & in2[12];
    assign P[210] = in[12] ^ in2[12];
    assign G[211] = in[11] & in2[11];
    assign P[211] = in[11] ^ in2[11];
    assign G[212] = in[10] & in2[10];
    assign P[212] = in[10] ^ in2[10];
    assign G[213] = in[9] & in2[9];
    assign P[213] = in[9] ^ in2[9];
    assign G[214] = in[8] & in2[8];
    assign P[214] = in[8] ^ in2[8];
    assign G[215] = in[7] & in2[7];
    assign P[215] = in[7] ^ in2[7];
    assign G[216] = in[6] & in2[6];
    assign P[216] = in[6] ^ in2[6];
    assign G[217] = in[5] & in2[5];
    assign P[217] = in[5] ^ in2[5];
    assign G[218] = in[4] & in2[4];
    assign P[218] = in[4] ^ in2[4];
    assign G[219] = in[3] & in2[3];
    assign P[219] = in[3] ^ in2[3];
    assign G[220] = in[2] & in2[2];
    assign P[220] = in[2] ^ in2[2];
    assign G[221] = in[1] & in2[1];
    assign P[221] = in[1] ^ in2[1];
    assign G[222] = in[0] & in2[0];
    assign P[222] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign C[222] = G[221] | (P[221] & C[221]);
    assign cout = G[222] | (P[222] & C[222]);
    assign sum = P ^ C;
endmodule

module CLA222(output [221:0] sum, output cout, input [221:0] in1, input [221:0] in2;

    wire[221:0] G;
    wire[221:0] C;
    wire[221:0] P;

    assign G[0] = in[221] & in2[221];
    assign P[0] = in[221] ^ in2[221];
    assign G[1] = in[220] & in2[220];
    assign P[1] = in[220] ^ in2[220];
    assign G[2] = in[219] & in2[219];
    assign P[2] = in[219] ^ in2[219];
    assign G[3] = in[218] & in2[218];
    assign P[3] = in[218] ^ in2[218];
    assign G[4] = in[217] & in2[217];
    assign P[4] = in[217] ^ in2[217];
    assign G[5] = in[216] & in2[216];
    assign P[5] = in[216] ^ in2[216];
    assign G[6] = in[215] & in2[215];
    assign P[6] = in[215] ^ in2[215];
    assign G[7] = in[214] & in2[214];
    assign P[7] = in[214] ^ in2[214];
    assign G[8] = in[213] & in2[213];
    assign P[8] = in[213] ^ in2[213];
    assign G[9] = in[212] & in2[212];
    assign P[9] = in[212] ^ in2[212];
    assign G[10] = in[211] & in2[211];
    assign P[10] = in[211] ^ in2[211];
    assign G[11] = in[210] & in2[210];
    assign P[11] = in[210] ^ in2[210];
    assign G[12] = in[209] & in2[209];
    assign P[12] = in[209] ^ in2[209];
    assign G[13] = in[208] & in2[208];
    assign P[13] = in[208] ^ in2[208];
    assign G[14] = in[207] & in2[207];
    assign P[14] = in[207] ^ in2[207];
    assign G[15] = in[206] & in2[206];
    assign P[15] = in[206] ^ in2[206];
    assign G[16] = in[205] & in2[205];
    assign P[16] = in[205] ^ in2[205];
    assign G[17] = in[204] & in2[204];
    assign P[17] = in[204] ^ in2[204];
    assign G[18] = in[203] & in2[203];
    assign P[18] = in[203] ^ in2[203];
    assign G[19] = in[202] & in2[202];
    assign P[19] = in[202] ^ in2[202];
    assign G[20] = in[201] & in2[201];
    assign P[20] = in[201] ^ in2[201];
    assign G[21] = in[200] & in2[200];
    assign P[21] = in[200] ^ in2[200];
    assign G[22] = in[199] & in2[199];
    assign P[22] = in[199] ^ in2[199];
    assign G[23] = in[198] & in2[198];
    assign P[23] = in[198] ^ in2[198];
    assign G[24] = in[197] & in2[197];
    assign P[24] = in[197] ^ in2[197];
    assign G[25] = in[196] & in2[196];
    assign P[25] = in[196] ^ in2[196];
    assign G[26] = in[195] & in2[195];
    assign P[26] = in[195] ^ in2[195];
    assign G[27] = in[194] & in2[194];
    assign P[27] = in[194] ^ in2[194];
    assign G[28] = in[193] & in2[193];
    assign P[28] = in[193] ^ in2[193];
    assign G[29] = in[192] & in2[192];
    assign P[29] = in[192] ^ in2[192];
    assign G[30] = in[191] & in2[191];
    assign P[30] = in[191] ^ in2[191];
    assign G[31] = in[190] & in2[190];
    assign P[31] = in[190] ^ in2[190];
    assign G[32] = in[189] & in2[189];
    assign P[32] = in[189] ^ in2[189];
    assign G[33] = in[188] & in2[188];
    assign P[33] = in[188] ^ in2[188];
    assign G[34] = in[187] & in2[187];
    assign P[34] = in[187] ^ in2[187];
    assign G[35] = in[186] & in2[186];
    assign P[35] = in[186] ^ in2[186];
    assign G[36] = in[185] & in2[185];
    assign P[36] = in[185] ^ in2[185];
    assign G[37] = in[184] & in2[184];
    assign P[37] = in[184] ^ in2[184];
    assign G[38] = in[183] & in2[183];
    assign P[38] = in[183] ^ in2[183];
    assign G[39] = in[182] & in2[182];
    assign P[39] = in[182] ^ in2[182];
    assign G[40] = in[181] & in2[181];
    assign P[40] = in[181] ^ in2[181];
    assign G[41] = in[180] & in2[180];
    assign P[41] = in[180] ^ in2[180];
    assign G[42] = in[179] & in2[179];
    assign P[42] = in[179] ^ in2[179];
    assign G[43] = in[178] & in2[178];
    assign P[43] = in[178] ^ in2[178];
    assign G[44] = in[177] & in2[177];
    assign P[44] = in[177] ^ in2[177];
    assign G[45] = in[176] & in2[176];
    assign P[45] = in[176] ^ in2[176];
    assign G[46] = in[175] & in2[175];
    assign P[46] = in[175] ^ in2[175];
    assign G[47] = in[174] & in2[174];
    assign P[47] = in[174] ^ in2[174];
    assign G[48] = in[173] & in2[173];
    assign P[48] = in[173] ^ in2[173];
    assign G[49] = in[172] & in2[172];
    assign P[49] = in[172] ^ in2[172];
    assign G[50] = in[171] & in2[171];
    assign P[50] = in[171] ^ in2[171];
    assign G[51] = in[170] & in2[170];
    assign P[51] = in[170] ^ in2[170];
    assign G[52] = in[169] & in2[169];
    assign P[52] = in[169] ^ in2[169];
    assign G[53] = in[168] & in2[168];
    assign P[53] = in[168] ^ in2[168];
    assign G[54] = in[167] & in2[167];
    assign P[54] = in[167] ^ in2[167];
    assign G[55] = in[166] & in2[166];
    assign P[55] = in[166] ^ in2[166];
    assign G[56] = in[165] & in2[165];
    assign P[56] = in[165] ^ in2[165];
    assign G[57] = in[164] & in2[164];
    assign P[57] = in[164] ^ in2[164];
    assign G[58] = in[163] & in2[163];
    assign P[58] = in[163] ^ in2[163];
    assign G[59] = in[162] & in2[162];
    assign P[59] = in[162] ^ in2[162];
    assign G[60] = in[161] & in2[161];
    assign P[60] = in[161] ^ in2[161];
    assign G[61] = in[160] & in2[160];
    assign P[61] = in[160] ^ in2[160];
    assign G[62] = in[159] & in2[159];
    assign P[62] = in[159] ^ in2[159];
    assign G[63] = in[158] & in2[158];
    assign P[63] = in[158] ^ in2[158];
    assign G[64] = in[157] & in2[157];
    assign P[64] = in[157] ^ in2[157];
    assign G[65] = in[156] & in2[156];
    assign P[65] = in[156] ^ in2[156];
    assign G[66] = in[155] & in2[155];
    assign P[66] = in[155] ^ in2[155];
    assign G[67] = in[154] & in2[154];
    assign P[67] = in[154] ^ in2[154];
    assign G[68] = in[153] & in2[153];
    assign P[68] = in[153] ^ in2[153];
    assign G[69] = in[152] & in2[152];
    assign P[69] = in[152] ^ in2[152];
    assign G[70] = in[151] & in2[151];
    assign P[70] = in[151] ^ in2[151];
    assign G[71] = in[150] & in2[150];
    assign P[71] = in[150] ^ in2[150];
    assign G[72] = in[149] & in2[149];
    assign P[72] = in[149] ^ in2[149];
    assign G[73] = in[148] & in2[148];
    assign P[73] = in[148] ^ in2[148];
    assign G[74] = in[147] & in2[147];
    assign P[74] = in[147] ^ in2[147];
    assign G[75] = in[146] & in2[146];
    assign P[75] = in[146] ^ in2[146];
    assign G[76] = in[145] & in2[145];
    assign P[76] = in[145] ^ in2[145];
    assign G[77] = in[144] & in2[144];
    assign P[77] = in[144] ^ in2[144];
    assign G[78] = in[143] & in2[143];
    assign P[78] = in[143] ^ in2[143];
    assign G[79] = in[142] & in2[142];
    assign P[79] = in[142] ^ in2[142];
    assign G[80] = in[141] & in2[141];
    assign P[80] = in[141] ^ in2[141];
    assign G[81] = in[140] & in2[140];
    assign P[81] = in[140] ^ in2[140];
    assign G[82] = in[139] & in2[139];
    assign P[82] = in[139] ^ in2[139];
    assign G[83] = in[138] & in2[138];
    assign P[83] = in[138] ^ in2[138];
    assign G[84] = in[137] & in2[137];
    assign P[84] = in[137] ^ in2[137];
    assign G[85] = in[136] & in2[136];
    assign P[85] = in[136] ^ in2[136];
    assign G[86] = in[135] & in2[135];
    assign P[86] = in[135] ^ in2[135];
    assign G[87] = in[134] & in2[134];
    assign P[87] = in[134] ^ in2[134];
    assign G[88] = in[133] & in2[133];
    assign P[88] = in[133] ^ in2[133];
    assign G[89] = in[132] & in2[132];
    assign P[89] = in[132] ^ in2[132];
    assign G[90] = in[131] & in2[131];
    assign P[90] = in[131] ^ in2[131];
    assign G[91] = in[130] & in2[130];
    assign P[91] = in[130] ^ in2[130];
    assign G[92] = in[129] & in2[129];
    assign P[92] = in[129] ^ in2[129];
    assign G[93] = in[128] & in2[128];
    assign P[93] = in[128] ^ in2[128];
    assign G[94] = in[127] & in2[127];
    assign P[94] = in[127] ^ in2[127];
    assign G[95] = in[126] & in2[126];
    assign P[95] = in[126] ^ in2[126];
    assign G[96] = in[125] & in2[125];
    assign P[96] = in[125] ^ in2[125];
    assign G[97] = in[124] & in2[124];
    assign P[97] = in[124] ^ in2[124];
    assign G[98] = in[123] & in2[123];
    assign P[98] = in[123] ^ in2[123];
    assign G[99] = in[122] & in2[122];
    assign P[99] = in[122] ^ in2[122];
    assign G[100] = in[121] & in2[121];
    assign P[100] = in[121] ^ in2[121];
    assign G[101] = in[120] & in2[120];
    assign P[101] = in[120] ^ in2[120];
    assign G[102] = in[119] & in2[119];
    assign P[102] = in[119] ^ in2[119];
    assign G[103] = in[118] & in2[118];
    assign P[103] = in[118] ^ in2[118];
    assign G[104] = in[117] & in2[117];
    assign P[104] = in[117] ^ in2[117];
    assign G[105] = in[116] & in2[116];
    assign P[105] = in[116] ^ in2[116];
    assign G[106] = in[115] & in2[115];
    assign P[106] = in[115] ^ in2[115];
    assign G[107] = in[114] & in2[114];
    assign P[107] = in[114] ^ in2[114];
    assign G[108] = in[113] & in2[113];
    assign P[108] = in[113] ^ in2[113];
    assign G[109] = in[112] & in2[112];
    assign P[109] = in[112] ^ in2[112];
    assign G[110] = in[111] & in2[111];
    assign P[110] = in[111] ^ in2[111];
    assign G[111] = in[110] & in2[110];
    assign P[111] = in[110] ^ in2[110];
    assign G[112] = in[109] & in2[109];
    assign P[112] = in[109] ^ in2[109];
    assign G[113] = in[108] & in2[108];
    assign P[113] = in[108] ^ in2[108];
    assign G[114] = in[107] & in2[107];
    assign P[114] = in[107] ^ in2[107];
    assign G[115] = in[106] & in2[106];
    assign P[115] = in[106] ^ in2[106];
    assign G[116] = in[105] & in2[105];
    assign P[116] = in[105] ^ in2[105];
    assign G[117] = in[104] & in2[104];
    assign P[117] = in[104] ^ in2[104];
    assign G[118] = in[103] & in2[103];
    assign P[118] = in[103] ^ in2[103];
    assign G[119] = in[102] & in2[102];
    assign P[119] = in[102] ^ in2[102];
    assign G[120] = in[101] & in2[101];
    assign P[120] = in[101] ^ in2[101];
    assign G[121] = in[100] & in2[100];
    assign P[121] = in[100] ^ in2[100];
    assign G[122] = in[99] & in2[99];
    assign P[122] = in[99] ^ in2[99];
    assign G[123] = in[98] & in2[98];
    assign P[123] = in[98] ^ in2[98];
    assign G[124] = in[97] & in2[97];
    assign P[124] = in[97] ^ in2[97];
    assign G[125] = in[96] & in2[96];
    assign P[125] = in[96] ^ in2[96];
    assign G[126] = in[95] & in2[95];
    assign P[126] = in[95] ^ in2[95];
    assign G[127] = in[94] & in2[94];
    assign P[127] = in[94] ^ in2[94];
    assign G[128] = in[93] & in2[93];
    assign P[128] = in[93] ^ in2[93];
    assign G[129] = in[92] & in2[92];
    assign P[129] = in[92] ^ in2[92];
    assign G[130] = in[91] & in2[91];
    assign P[130] = in[91] ^ in2[91];
    assign G[131] = in[90] & in2[90];
    assign P[131] = in[90] ^ in2[90];
    assign G[132] = in[89] & in2[89];
    assign P[132] = in[89] ^ in2[89];
    assign G[133] = in[88] & in2[88];
    assign P[133] = in[88] ^ in2[88];
    assign G[134] = in[87] & in2[87];
    assign P[134] = in[87] ^ in2[87];
    assign G[135] = in[86] & in2[86];
    assign P[135] = in[86] ^ in2[86];
    assign G[136] = in[85] & in2[85];
    assign P[136] = in[85] ^ in2[85];
    assign G[137] = in[84] & in2[84];
    assign P[137] = in[84] ^ in2[84];
    assign G[138] = in[83] & in2[83];
    assign P[138] = in[83] ^ in2[83];
    assign G[139] = in[82] & in2[82];
    assign P[139] = in[82] ^ in2[82];
    assign G[140] = in[81] & in2[81];
    assign P[140] = in[81] ^ in2[81];
    assign G[141] = in[80] & in2[80];
    assign P[141] = in[80] ^ in2[80];
    assign G[142] = in[79] & in2[79];
    assign P[142] = in[79] ^ in2[79];
    assign G[143] = in[78] & in2[78];
    assign P[143] = in[78] ^ in2[78];
    assign G[144] = in[77] & in2[77];
    assign P[144] = in[77] ^ in2[77];
    assign G[145] = in[76] & in2[76];
    assign P[145] = in[76] ^ in2[76];
    assign G[146] = in[75] & in2[75];
    assign P[146] = in[75] ^ in2[75];
    assign G[147] = in[74] & in2[74];
    assign P[147] = in[74] ^ in2[74];
    assign G[148] = in[73] & in2[73];
    assign P[148] = in[73] ^ in2[73];
    assign G[149] = in[72] & in2[72];
    assign P[149] = in[72] ^ in2[72];
    assign G[150] = in[71] & in2[71];
    assign P[150] = in[71] ^ in2[71];
    assign G[151] = in[70] & in2[70];
    assign P[151] = in[70] ^ in2[70];
    assign G[152] = in[69] & in2[69];
    assign P[152] = in[69] ^ in2[69];
    assign G[153] = in[68] & in2[68];
    assign P[153] = in[68] ^ in2[68];
    assign G[154] = in[67] & in2[67];
    assign P[154] = in[67] ^ in2[67];
    assign G[155] = in[66] & in2[66];
    assign P[155] = in[66] ^ in2[66];
    assign G[156] = in[65] & in2[65];
    assign P[156] = in[65] ^ in2[65];
    assign G[157] = in[64] & in2[64];
    assign P[157] = in[64] ^ in2[64];
    assign G[158] = in[63] & in2[63];
    assign P[158] = in[63] ^ in2[63];
    assign G[159] = in[62] & in2[62];
    assign P[159] = in[62] ^ in2[62];
    assign G[160] = in[61] & in2[61];
    assign P[160] = in[61] ^ in2[61];
    assign G[161] = in[60] & in2[60];
    assign P[161] = in[60] ^ in2[60];
    assign G[162] = in[59] & in2[59];
    assign P[162] = in[59] ^ in2[59];
    assign G[163] = in[58] & in2[58];
    assign P[163] = in[58] ^ in2[58];
    assign G[164] = in[57] & in2[57];
    assign P[164] = in[57] ^ in2[57];
    assign G[165] = in[56] & in2[56];
    assign P[165] = in[56] ^ in2[56];
    assign G[166] = in[55] & in2[55];
    assign P[166] = in[55] ^ in2[55];
    assign G[167] = in[54] & in2[54];
    assign P[167] = in[54] ^ in2[54];
    assign G[168] = in[53] & in2[53];
    assign P[168] = in[53] ^ in2[53];
    assign G[169] = in[52] & in2[52];
    assign P[169] = in[52] ^ in2[52];
    assign G[170] = in[51] & in2[51];
    assign P[170] = in[51] ^ in2[51];
    assign G[171] = in[50] & in2[50];
    assign P[171] = in[50] ^ in2[50];
    assign G[172] = in[49] & in2[49];
    assign P[172] = in[49] ^ in2[49];
    assign G[173] = in[48] & in2[48];
    assign P[173] = in[48] ^ in2[48];
    assign G[174] = in[47] & in2[47];
    assign P[174] = in[47] ^ in2[47];
    assign G[175] = in[46] & in2[46];
    assign P[175] = in[46] ^ in2[46];
    assign G[176] = in[45] & in2[45];
    assign P[176] = in[45] ^ in2[45];
    assign G[177] = in[44] & in2[44];
    assign P[177] = in[44] ^ in2[44];
    assign G[178] = in[43] & in2[43];
    assign P[178] = in[43] ^ in2[43];
    assign G[179] = in[42] & in2[42];
    assign P[179] = in[42] ^ in2[42];
    assign G[180] = in[41] & in2[41];
    assign P[180] = in[41] ^ in2[41];
    assign G[181] = in[40] & in2[40];
    assign P[181] = in[40] ^ in2[40];
    assign G[182] = in[39] & in2[39];
    assign P[182] = in[39] ^ in2[39];
    assign G[183] = in[38] & in2[38];
    assign P[183] = in[38] ^ in2[38];
    assign G[184] = in[37] & in2[37];
    assign P[184] = in[37] ^ in2[37];
    assign G[185] = in[36] & in2[36];
    assign P[185] = in[36] ^ in2[36];
    assign G[186] = in[35] & in2[35];
    assign P[186] = in[35] ^ in2[35];
    assign G[187] = in[34] & in2[34];
    assign P[187] = in[34] ^ in2[34];
    assign G[188] = in[33] & in2[33];
    assign P[188] = in[33] ^ in2[33];
    assign G[189] = in[32] & in2[32];
    assign P[189] = in[32] ^ in2[32];
    assign G[190] = in[31] & in2[31];
    assign P[190] = in[31] ^ in2[31];
    assign G[191] = in[30] & in2[30];
    assign P[191] = in[30] ^ in2[30];
    assign G[192] = in[29] & in2[29];
    assign P[192] = in[29] ^ in2[29];
    assign G[193] = in[28] & in2[28];
    assign P[193] = in[28] ^ in2[28];
    assign G[194] = in[27] & in2[27];
    assign P[194] = in[27] ^ in2[27];
    assign G[195] = in[26] & in2[26];
    assign P[195] = in[26] ^ in2[26];
    assign G[196] = in[25] & in2[25];
    assign P[196] = in[25] ^ in2[25];
    assign G[197] = in[24] & in2[24];
    assign P[197] = in[24] ^ in2[24];
    assign G[198] = in[23] & in2[23];
    assign P[198] = in[23] ^ in2[23];
    assign G[199] = in[22] & in2[22];
    assign P[199] = in[22] ^ in2[22];
    assign G[200] = in[21] & in2[21];
    assign P[200] = in[21] ^ in2[21];
    assign G[201] = in[20] & in2[20];
    assign P[201] = in[20] ^ in2[20];
    assign G[202] = in[19] & in2[19];
    assign P[202] = in[19] ^ in2[19];
    assign G[203] = in[18] & in2[18];
    assign P[203] = in[18] ^ in2[18];
    assign G[204] = in[17] & in2[17];
    assign P[204] = in[17] ^ in2[17];
    assign G[205] = in[16] & in2[16];
    assign P[205] = in[16] ^ in2[16];
    assign G[206] = in[15] & in2[15];
    assign P[206] = in[15] ^ in2[15];
    assign G[207] = in[14] & in2[14];
    assign P[207] = in[14] ^ in2[14];
    assign G[208] = in[13] & in2[13];
    assign P[208] = in[13] ^ in2[13];
    assign G[209] = in[12] & in2[12];
    assign P[209] = in[12] ^ in2[12];
    assign G[210] = in[11] & in2[11];
    assign P[210] = in[11] ^ in2[11];
    assign G[211] = in[10] & in2[10];
    assign P[211] = in[10] ^ in2[10];
    assign G[212] = in[9] & in2[9];
    assign P[212] = in[9] ^ in2[9];
    assign G[213] = in[8] & in2[8];
    assign P[213] = in[8] ^ in2[8];
    assign G[214] = in[7] & in2[7];
    assign P[214] = in[7] ^ in2[7];
    assign G[215] = in[6] & in2[6];
    assign P[215] = in[6] ^ in2[6];
    assign G[216] = in[5] & in2[5];
    assign P[216] = in[5] ^ in2[5];
    assign G[217] = in[4] & in2[4];
    assign P[217] = in[4] ^ in2[4];
    assign G[218] = in[3] & in2[3];
    assign P[218] = in[3] ^ in2[3];
    assign G[219] = in[2] & in2[2];
    assign P[219] = in[2] ^ in2[2];
    assign G[220] = in[1] & in2[1];
    assign P[220] = in[1] ^ in2[1];
    assign G[221] = in[0] & in2[0];
    assign P[221] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign C[221] = G[220] | (P[220] & C[220]);
    assign cout = G[221] | (P[221] & C[221]);
    assign sum = P ^ C;
endmodule

module CLA221(output [220:0] sum, output cout, input [220:0] in1, input [220:0] in2;

    wire[220:0] G;
    wire[220:0] C;
    wire[220:0] P;

    assign G[0] = in[220] & in2[220];
    assign P[0] = in[220] ^ in2[220];
    assign G[1] = in[219] & in2[219];
    assign P[1] = in[219] ^ in2[219];
    assign G[2] = in[218] & in2[218];
    assign P[2] = in[218] ^ in2[218];
    assign G[3] = in[217] & in2[217];
    assign P[3] = in[217] ^ in2[217];
    assign G[4] = in[216] & in2[216];
    assign P[4] = in[216] ^ in2[216];
    assign G[5] = in[215] & in2[215];
    assign P[5] = in[215] ^ in2[215];
    assign G[6] = in[214] & in2[214];
    assign P[6] = in[214] ^ in2[214];
    assign G[7] = in[213] & in2[213];
    assign P[7] = in[213] ^ in2[213];
    assign G[8] = in[212] & in2[212];
    assign P[8] = in[212] ^ in2[212];
    assign G[9] = in[211] & in2[211];
    assign P[9] = in[211] ^ in2[211];
    assign G[10] = in[210] & in2[210];
    assign P[10] = in[210] ^ in2[210];
    assign G[11] = in[209] & in2[209];
    assign P[11] = in[209] ^ in2[209];
    assign G[12] = in[208] & in2[208];
    assign P[12] = in[208] ^ in2[208];
    assign G[13] = in[207] & in2[207];
    assign P[13] = in[207] ^ in2[207];
    assign G[14] = in[206] & in2[206];
    assign P[14] = in[206] ^ in2[206];
    assign G[15] = in[205] & in2[205];
    assign P[15] = in[205] ^ in2[205];
    assign G[16] = in[204] & in2[204];
    assign P[16] = in[204] ^ in2[204];
    assign G[17] = in[203] & in2[203];
    assign P[17] = in[203] ^ in2[203];
    assign G[18] = in[202] & in2[202];
    assign P[18] = in[202] ^ in2[202];
    assign G[19] = in[201] & in2[201];
    assign P[19] = in[201] ^ in2[201];
    assign G[20] = in[200] & in2[200];
    assign P[20] = in[200] ^ in2[200];
    assign G[21] = in[199] & in2[199];
    assign P[21] = in[199] ^ in2[199];
    assign G[22] = in[198] & in2[198];
    assign P[22] = in[198] ^ in2[198];
    assign G[23] = in[197] & in2[197];
    assign P[23] = in[197] ^ in2[197];
    assign G[24] = in[196] & in2[196];
    assign P[24] = in[196] ^ in2[196];
    assign G[25] = in[195] & in2[195];
    assign P[25] = in[195] ^ in2[195];
    assign G[26] = in[194] & in2[194];
    assign P[26] = in[194] ^ in2[194];
    assign G[27] = in[193] & in2[193];
    assign P[27] = in[193] ^ in2[193];
    assign G[28] = in[192] & in2[192];
    assign P[28] = in[192] ^ in2[192];
    assign G[29] = in[191] & in2[191];
    assign P[29] = in[191] ^ in2[191];
    assign G[30] = in[190] & in2[190];
    assign P[30] = in[190] ^ in2[190];
    assign G[31] = in[189] & in2[189];
    assign P[31] = in[189] ^ in2[189];
    assign G[32] = in[188] & in2[188];
    assign P[32] = in[188] ^ in2[188];
    assign G[33] = in[187] & in2[187];
    assign P[33] = in[187] ^ in2[187];
    assign G[34] = in[186] & in2[186];
    assign P[34] = in[186] ^ in2[186];
    assign G[35] = in[185] & in2[185];
    assign P[35] = in[185] ^ in2[185];
    assign G[36] = in[184] & in2[184];
    assign P[36] = in[184] ^ in2[184];
    assign G[37] = in[183] & in2[183];
    assign P[37] = in[183] ^ in2[183];
    assign G[38] = in[182] & in2[182];
    assign P[38] = in[182] ^ in2[182];
    assign G[39] = in[181] & in2[181];
    assign P[39] = in[181] ^ in2[181];
    assign G[40] = in[180] & in2[180];
    assign P[40] = in[180] ^ in2[180];
    assign G[41] = in[179] & in2[179];
    assign P[41] = in[179] ^ in2[179];
    assign G[42] = in[178] & in2[178];
    assign P[42] = in[178] ^ in2[178];
    assign G[43] = in[177] & in2[177];
    assign P[43] = in[177] ^ in2[177];
    assign G[44] = in[176] & in2[176];
    assign P[44] = in[176] ^ in2[176];
    assign G[45] = in[175] & in2[175];
    assign P[45] = in[175] ^ in2[175];
    assign G[46] = in[174] & in2[174];
    assign P[46] = in[174] ^ in2[174];
    assign G[47] = in[173] & in2[173];
    assign P[47] = in[173] ^ in2[173];
    assign G[48] = in[172] & in2[172];
    assign P[48] = in[172] ^ in2[172];
    assign G[49] = in[171] & in2[171];
    assign P[49] = in[171] ^ in2[171];
    assign G[50] = in[170] & in2[170];
    assign P[50] = in[170] ^ in2[170];
    assign G[51] = in[169] & in2[169];
    assign P[51] = in[169] ^ in2[169];
    assign G[52] = in[168] & in2[168];
    assign P[52] = in[168] ^ in2[168];
    assign G[53] = in[167] & in2[167];
    assign P[53] = in[167] ^ in2[167];
    assign G[54] = in[166] & in2[166];
    assign P[54] = in[166] ^ in2[166];
    assign G[55] = in[165] & in2[165];
    assign P[55] = in[165] ^ in2[165];
    assign G[56] = in[164] & in2[164];
    assign P[56] = in[164] ^ in2[164];
    assign G[57] = in[163] & in2[163];
    assign P[57] = in[163] ^ in2[163];
    assign G[58] = in[162] & in2[162];
    assign P[58] = in[162] ^ in2[162];
    assign G[59] = in[161] & in2[161];
    assign P[59] = in[161] ^ in2[161];
    assign G[60] = in[160] & in2[160];
    assign P[60] = in[160] ^ in2[160];
    assign G[61] = in[159] & in2[159];
    assign P[61] = in[159] ^ in2[159];
    assign G[62] = in[158] & in2[158];
    assign P[62] = in[158] ^ in2[158];
    assign G[63] = in[157] & in2[157];
    assign P[63] = in[157] ^ in2[157];
    assign G[64] = in[156] & in2[156];
    assign P[64] = in[156] ^ in2[156];
    assign G[65] = in[155] & in2[155];
    assign P[65] = in[155] ^ in2[155];
    assign G[66] = in[154] & in2[154];
    assign P[66] = in[154] ^ in2[154];
    assign G[67] = in[153] & in2[153];
    assign P[67] = in[153] ^ in2[153];
    assign G[68] = in[152] & in2[152];
    assign P[68] = in[152] ^ in2[152];
    assign G[69] = in[151] & in2[151];
    assign P[69] = in[151] ^ in2[151];
    assign G[70] = in[150] & in2[150];
    assign P[70] = in[150] ^ in2[150];
    assign G[71] = in[149] & in2[149];
    assign P[71] = in[149] ^ in2[149];
    assign G[72] = in[148] & in2[148];
    assign P[72] = in[148] ^ in2[148];
    assign G[73] = in[147] & in2[147];
    assign P[73] = in[147] ^ in2[147];
    assign G[74] = in[146] & in2[146];
    assign P[74] = in[146] ^ in2[146];
    assign G[75] = in[145] & in2[145];
    assign P[75] = in[145] ^ in2[145];
    assign G[76] = in[144] & in2[144];
    assign P[76] = in[144] ^ in2[144];
    assign G[77] = in[143] & in2[143];
    assign P[77] = in[143] ^ in2[143];
    assign G[78] = in[142] & in2[142];
    assign P[78] = in[142] ^ in2[142];
    assign G[79] = in[141] & in2[141];
    assign P[79] = in[141] ^ in2[141];
    assign G[80] = in[140] & in2[140];
    assign P[80] = in[140] ^ in2[140];
    assign G[81] = in[139] & in2[139];
    assign P[81] = in[139] ^ in2[139];
    assign G[82] = in[138] & in2[138];
    assign P[82] = in[138] ^ in2[138];
    assign G[83] = in[137] & in2[137];
    assign P[83] = in[137] ^ in2[137];
    assign G[84] = in[136] & in2[136];
    assign P[84] = in[136] ^ in2[136];
    assign G[85] = in[135] & in2[135];
    assign P[85] = in[135] ^ in2[135];
    assign G[86] = in[134] & in2[134];
    assign P[86] = in[134] ^ in2[134];
    assign G[87] = in[133] & in2[133];
    assign P[87] = in[133] ^ in2[133];
    assign G[88] = in[132] & in2[132];
    assign P[88] = in[132] ^ in2[132];
    assign G[89] = in[131] & in2[131];
    assign P[89] = in[131] ^ in2[131];
    assign G[90] = in[130] & in2[130];
    assign P[90] = in[130] ^ in2[130];
    assign G[91] = in[129] & in2[129];
    assign P[91] = in[129] ^ in2[129];
    assign G[92] = in[128] & in2[128];
    assign P[92] = in[128] ^ in2[128];
    assign G[93] = in[127] & in2[127];
    assign P[93] = in[127] ^ in2[127];
    assign G[94] = in[126] & in2[126];
    assign P[94] = in[126] ^ in2[126];
    assign G[95] = in[125] & in2[125];
    assign P[95] = in[125] ^ in2[125];
    assign G[96] = in[124] & in2[124];
    assign P[96] = in[124] ^ in2[124];
    assign G[97] = in[123] & in2[123];
    assign P[97] = in[123] ^ in2[123];
    assign G[98] = in[122] & in2[122];
    assign P[98] = in[122] ^ in2[122];
    assign G[99] = in[121] & in2[121];
    assign P[99] = in[121] ^ in2[121];
    assign G[100] = in[120] & in2[120];
    assign P[100] = in[120] ^ in2[120];
    assign G[101] = in[119] & in2[119];
    assign P[101] = in[119] ^ in2[119];
    assign G[102] = in[118] & in2[118];
    assign P[102] = in[118] ^ in2[118];
    assign G[103] = in[117] & in2[117];
    assign P[103] = in[117] ^ in2[117];
    assign G[104] = in[116] & in2[116];
    assign P[104] = in[116] ^ in2[116];
    assign G[105] = in[115] & in2[115];
    assign P[105] = in[115] ^ in2[115];
    assign G[106] = in[114] & in2[114];
    assign P[106] = in[114] ^ in2[114];
    assign G[107] = in[113] & in2[113];
    assign P[107] = in[113] ^ in2[113];
    assign G[108] = in[112] & in2[112];
    assign P[108] = in[112] ^ in2[112];
    assign G[109] = in[111] & in2[111];
    assign P[109] = in[111] ^ in2[111];
    assign G[110] = in[110] & in2[110];
    assign P[110] = in[110] ^ in2[110];
    assign G[111] = in[109] & in2[109];
    assign P[111] = in[109] ^ in2[109];
    assign G[112] = in[108] & in2[108];
    assign P[112] = in[108] ^ in2[108];
    assign G[113] = in[107] & in2[107];
    assign P[113] = in[107] ^ in2[107];
    assign G[114] = in[106] & in2[106];
    assign P[114] = in[106] ^ in2[106];
    assign G[115] = in[105] & in2[105];
    assign P[115] = in[105] ^ in2[105];
    assign G[116] = in[104] & in2[104];
    assign P[116] = in[104] ^ in2[104];
    assign G[117] = in[103] & in2[103];
    assign P[117] = in[103] ^ in2[103];
    assign G[118] = in[102] & in2[102];
    assign P[118] = in[102] ^ in2[102];
    assign G[119] = in[101] & in2[101];
    assign P[119] = in[101] ^ in2[101];
    assign G[120] = in[100] & in2[100];
    assign P[120] = in[100] ^ in2[100];
    assign G[121] = in[99] & in2[99];
    assign P[121] = in[99] ^ in2[99];
    assign G[122] = in[98] & in2[98];
    assign P[122] = in[98] ^ in2[98];
    assign G[123] = in[97] & in2[97];
    assign P[123] = in[97] ^ in2[97];
    assign G[124] = in[96] & in2[96];
    assign P[124] = in[96] ^ in2[96];
    assign G[125] = in[95] & in2[95];
    assign P[125] = in[95] ^ in2[95];
    assign G[126] = in[94] & in2[94];
    assign P[126] = in[94] ^ in2[94];
    assign G[127] = in[93] & in2[93];
    assign P[127] = in[93] ^ in2[93];
    assign G[128] = in[92] & in2[92];
    assign P[128] = in[92] ^ in2[92];
    assign G[129] = in[91] & in2[91];
    assign P[129] = in[91] ^ in2[91];
    assign G[130] = in[90] & in2[90];
    assign P[130] = in[90] ^ in2[90];
    assign G[131] = in[89] & in2[89];
    assign P[131] = in[89] ^ in2[89];
    assign G[132] = in[88] & in2[88];
    assign P[132] = in[88] ^ in2[88];
    assign G[133] = in[87] & in2[87];
    assign P[133] = in[87] ^ in2[87];
    assign G[134] = in[86] & in2[86];
    assign P[134] = in[86] ^ in2[86];
    assign G[135] = in[85] & in2[85];
    assign P[135] = in[85] ^ in2[85];
    assign G[136] = in[84] & in2[84];
    assign P[136] = in[84] ^ in2[84];
    assign G[137] = in[83] & in2[83];
    assign P[137] = in[83] ^ in2[83];
    assign G[138] = in[82] & in2[82];
    assign P[138] = in[82] ^ in2[82];
    assign G[139] = in[81] & in2[81];
    assign P[139] = in[81] ^ in2[81];
    assign G[140] = in[80] & in2[80];
    assign P[140] = in[80] ^ in2[80];
    assign G[141] = in[79] & in2[79];
    assign P[141] = in[79] ^ in2[79];
    assign G[142] = in[78] & in2[78];
    assign P[142] = in[78] ^ in2[78];
    assign G[143] = in[77] & in2[77];
    assign P[143] = in[77] ^ in2[77];
    assign G[144] = in[76] & in2[76];
    assign P[144] = in[76] ^ in2[76];
    assign G[145] = in[75] & in2[75];
    assign P[145] = in[75] ^ in2[75];
    assign G[146] = in[74] & in2[74];
    assign P[146] = in[74] ^ in2[74];
    assign G[147] = in[73] & in2[73];
    assign P[147] = in[73] ^ in2[73];
    assign G[148] = in[72] & in2[72];
    assign P[148] = in[72] ^ in2[72];
    assign G[149] = in[71] & in2[71];
    assign P[149] = in[71] ^ in2[71];
    assign G[150] = in[70] & in2[70];
    assign P[150] = in[70] ^ in2[70];
    assign G[151] = in[69] & in2[69];
    assign P[151] = in[69] ^ in2[69];
    assign G[152] = in[68] & in2[68];
    assign P[152] = in[68] ^ in2[68];
    assign G[153] = in[67] & in2[67];
    assign P[153] = in[67] ^ in2[67];
    assign G[154] = in[66] & in2[66];
    assign P[154] = in[66] ^ in2[66];
    assign G[155] = in[65] & in2[65];
    assign P[155] = in[65] ^ in2[65];
    assign G[156] = in[64] & in2[64];
    assign P[156] = in[64] ^ in2[64];
    assign G[157] = in[63] & in2[63];
    assign P[157] = in[63] ^ in2[63];
    assign G[158] = in[62] & in2[62];
    assign P[158] = in[62] ^ in2[62];
    assign G[159] = in[61] & in2[61];
    assign P[159] = in[61] ^ in2[61];
    assign G[160] = in[60] & in2[60];
    assign P[160] = in[60] ^ in2[60];
    assign G[161] = in[59] & in2[59];
    assign P[161] = in[59] ^ in2[59];
    assign G[162] = in[58] & in2[58];
    assign P[162] = in[58] ^ in2[58];
    assign G[163] = in[57] & in2[57];
    assign P[163] = in[57] ^ in2[57];
    assign G[164] = in[56] & in2[56];
    assign P[164] = in[56] ^ in2[56];
    assign G[165] = in[55] & in2[55];
    assign P[165] = in[55] ^ in2[55];
    assign G[166] = in[54] & in2[54];
    assign P[166] = in[54] ^ in2[54];
    assign G[167] = in[53] & in2[53];
    assign P[167] = in[53] ^ in2[53];
    assign G[168] = in[52] & in2[52];
    assign P[168] = in[52] ^ in2[52];
    assign G[169] = in[51] & in2[51];
    assign P[169] = in[51] ^ in2[51];
    assign G[170] = in[50] & in2[50];
    assign P[170] = in[50] ^ in2[50];
    assign G[171] = in[49] & in2[49];
    assign P[171] = in[49] ^ in2[49];
    assign G[172] = in[48] & in2[48];
    assign P[172] = in[48] ^ in2[48];
    assign G[173] = in[47] & in2[47];
    assign P[173] = in[47] ^ in2[47];
    assign G[174] = in[46] & in2[46];
    assign P[174] = in[46] ^ in2[46];
    assign G[175] = in[45] & in2[45];
    assign P[175] = in[45] ^ in2[45];
    assign G[176] = in[44] & in2[44];
    assign P[176] = in[44] ^ in2[44];
    assign G[177] = in[43] & in2[43];
    assign P[177] = in[43] ^ in2[43];
    assign G[178] = in[42] & in2[42];
    assign P[178] = in[42] ^ in2[42];
    assign G[179] = in[41] & in2[41];
    assign P[179] = in[41] ^ in2[41];
    assign G[180] = in[40] & in2[40];
    assign P[180] = in[40] ^ in2[40];
    assign G[181] = in[39] & in2[39];
    assign P[181] = in[39] ^ in2[39];
    assign G[182] = in[38] & in2[38];
    assign P[182] = in[38] ^ in2[38];
    assign G[183] = in[37] & in2[37];
    assign P[183] = in[37] ^ in2[37];
    assign G[184] = in[36] & in2[36];
    assign P[184] = in[36] ^ in2[36];
    assign G[185] = in[35] & in2[35];
    assign P[185] = in[35] ^ in2[35];
    assign G[186] = in[34] & in2[34];
    assign P[186] = in[34] ^ in2[34];
    assign G[187] = in[33] & in2[33];
    assign P[187] = in[33] ^ in2[33];
    assign G[188] = in[32] & in2[32];
    assign P[188] = in[32] ^ in2[32];
    assign G[189] = in[31] & in2[31];
    assign P[189] = in[31] ^ in2[31];
    assign G[190] = in[30] & in2[30];
    assign P[190] = in[30] ^ in2[30];
    assign G[191] = in[29] & in2[29];
    assign P[191] = in[29] ^ in2[29];
    assign G[192] = in[28] & in2[28];
    assign P[192] = in[28] ^ in2[28];
    assign G[193] = in[27] & in2[27];
    assign P[193] = in[27] ^ in2[27];
    assign G[194] = in[26] & in2[26];
    assign P[194] = in[26] ^ in2[26];
    assign G[195] = in[25] & in2[25];
    assign P[195] = in[25] ^ in2[25];
    assign G[196] = in[24] & in2[24];
    assign P[196] = in[24] ^ in2[24];
    assign G[197] = in[23] & in2[23];
    assign P[197] = in[23] ^ in2[23];
    assign G[198] = in[22] & in2[22];
    assign P[198] = in[22] ^ in2[22];
    assign G[199] = in[21] & in2[21];
    assign P[199] = in[21] ^ in2[21];
    assign G[200] = in[20] & in2[20];
    assign P[200] = in[20] ^ in2[20];
    assign G[201] = in[19] & in2[19];
    assign P[201] = in[19] ^ in2[19];
    assign G[202] = in[18] & in2[18];
    assign P[202] = in[18] ^ in2[18];
    assign G[203] = in[17] & in2[17];
    assign P[203] = in[17] ^ in2[17];
    assign G[204] = in[16] & in2[16];
    assign P[204] = in[16] ^ in2[16];
    assign G[205] = in[15] & in2[15];
    assign P[205] = in[15] ^ in2[15];
    assign G[206] = in[14] & in2[14];
    assign P[206] = in[14] ^ in2[14];
    assign G[207] = in[13] & in2[13];
    assign P[207] = in[13] ^ in2[13];
    assign G[208] = in[12] & in2[12];
    assign P[208] = in[12] ^ in2[12];
    assign G[209] = in[11] & in2[11];
    assign P[209] = in[11] ^ in2[11];
    assign G[210] = in[10] & in2[10];
    assign P[210] = in[10] ^ in2[10];
    assign G[211] = in[9] & in2[9];
    assign P[211] = in[9] ^ in2[9];
    assign G[212] = in[8] & in2[8];
    assign P[212] = in[8] ^ in2[8];
    assign G[213] = in[7] & in2[7];
    assign P[213] = in[7] ^ in2[7];
    assign G[214] = in[6] & in2[6];
    assign P[214] = in[6] ^ in2[6];
    assign G[215] = in[5] & in2[5];
    assign P[215] = in[5] ^ in2[5];
    assign G[216] = in[4] & in2[4];
    assign P[216] = in[4] ^ in2[4];
    assign G[217] = in[3] & in2[3];
    assign P[217] = in[3] ^ in2[3];
    assign G[218] = in[2] & in2[2];
    assign P[218] = in[2] ^ in2[2];
    assign G[219] = in[1] & in2[1];
    assign P[219] = in[1] ^ in2[1];
    assign G[220] = in[0] & in2[0];
    assign P[220] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign C[220] = G[219] | (P[219] & C[219]);
    assign cout = G[220] | (P[220] & C[220]);
    assign sum = P ^ C;
endmodule

module CLA220(output [219:0] sum, output cout, input [219:0] in1, input [219:0] in2;

    wire[219:0] G;
    wire[219:0] C;
    wire[219:0] P;

    assign G[0] = in[219] & in2[219];
    assign P[0] = in[219] ^ in2[219];
    assign G[1] = in[218] & in2[218];
    assign P[1] = in[218] ^ in2[218];
    assign G[2] = in[217] & in2[217];
    assign P[2] = in[217] ^ in2[217];
    assign G[3] = in[216] & in2[216];
    assign P[3] = in[216] ^ in2[216];
    assign G[4] = in[215] & in2[215];
    assign P[4] = in[215] ^ in2[215];
    assign G[5] = in[214] & in2[214];
    assign P[5] = in[214] ^ in2[214];
    assign G[6] = in[213] & in2[213];
    assign P[6] = in[213] ^ in2[213];
    assign G[7] = in[212] & in2[212];
    assign P[7] = in[212] ^ in2[212];
    assign G[8] = in[211] & in2[211];
    assign P[8] = in[211] ^ in2[211];
    assign G[9] = in[210] & in2[210];
    assign P[9] = in[210] ^ in2[210];
    assign G[10] = in[209] & in2[209];
    assign P[10] = in[209] ^ in2[209];
    assign G[11] = in[208] & in2[208];
    assign P[11] = in[208] ^ in2[208];
    assign G[12] = in[207] & in2[207];
    assign P[12] = in[207] ^ in2[207];
    assign G[13] = in[206] & in2[206];
    assign P[13] = in[206] ^ in2[206];
    assign G[14] = in[205] & in2[205];
    assign P[14] = in[205] ^ in2[205];
    assign G[15] = in[204] & in2[204];
    assign P[15] = in[204] ^ in2[204];
    assign G[16] = in[203] & in2[203];
    assign P[16] = in[203] ^ in2[203];
    assign G[17] = in[202] & in2[202];
    assign P[17] = in[202] ^ in2[202];
    assign G[18] = in[201] & in2[201];
    assign P[18] = in[201] ^ in2[201];
    assign G[19] = in[200] & in2[200];
    assign P[19] = in[200] ^ in2[200];
    assign G[20] = in[199] & in2[199];
    assign P[20] = in[199] ^ in2[199];
    assign G[21] = in[198] & in2[198];
    assign P[21] = in[198] ^ in2[198];
    assign G[22] = in[197] & in2[197];
    assign P[22] = in[197] ^ in2[197];
    assign G[23] = in[196] & in2[196];
    assign P[23] = in[196] ^ in2[196];
    assign G[24] = in[195] & in2[195];
    assign P[24] = in[195] ^ in2[195];
    assign G[25] = in[194] & in2[194];
    assign P[25] = in[194] ^ in2[194];
    assign G[26] = in[193] & in2[193];
    assign P[26] = in[193] ^ in2[193];
    assign G[27] = in[192] & in2[192];
    assign P[27] = in[192] ^ in2[192];
    assign G[28] = in[191] & in2[191];
    assign P[28] = in[191] ^ in2[191];
    assign G[29] = in[190] & in2[190];
    assign P[29] = in[190] ^ in2[190];
    assign G[30] = in[189] & in2[189];
    assign P[30] = in[189] ^ in2[189];
    assign G[31] = in[188] & in2[188];
    assign P[31] = in[188] ^ in2[188];
    assign G[32] = in[187] & in2[187];
    assign P[32] = in[187] ^ in2[187];
    assign G[33] = in[186] & in2[186];
    assign P[33] = in[186] ^ in2[186];
    assign G[34] = in[185] & in2[185];
    assign P[34] = in[185] ^ in2[185];
    assign G[35] = in[184] & in2[184];
    assign P[35] = in[184] ^ in2[184];
    assign G[36] = in[183] & in2[183];
    assign P[36] = in[183] ^ in2[183];
    assign G[37] = in[182] & in2[182];
    assign P[37] = in[182] ^ in2[182];
    assign G[38] = in[181] & in2[181];
    assign P[38] = in[181] ^ in2[181];
    assign G[39] = in[180] & in2[180];
    assign P[39] = in[180] ^ in2[180];
    assign G[40] = in[179] & in2[179];
    assign P[40] = in[179] ^ in2[179];
    assign G[41] = in[178] & in2[178];
    assign P[41] = in[178] ^ in2[178];
    assign G[42] = in[177] & in2[177];
    assign P[42] = in[177] ^ in2[177];
    assign G[43] = in[176] & in2[176];
    assign P[43] = in[176] ^ in2[176];
    assign G[44] = in[175] & in2[175];
    assign P[44] = in[175] ^ in2[175];
    assign G[45] = in[174] & in2[174];
    assign P[45] = in[174] ^ in2[174];
    assign G[46] = in[173] & in2[173];
    assign P[46] = in[173] ^ in2[173];
    assign G[47] = in[172] & in2[172];
    assign P[47] = in[172] ^ in2[172];
    assign G[48] = in[171] & in2[171];
    assign P[48] = in[171] ^ in2[171];
    assign G[49] = in[170] & in2[170];
    assign P[49] = in[170] ^ in2[170];
    assign G[50] = in[169] & in2[169];
    assign P[50] = in[169] ^ in2[169];
    assign G[51] = in[168] & in2[168];
    assign P[51] = in[168] ^ in2[168];
    assign G[52] = in[167] & in2[167];
    assign P[52] = in[167] ^ in2[167];
    assign G[53] = in[166] & in2[166];
    assign P[53] = in[166] ^ in2[166];
    assign G[54] = in[165] & in2[165];
    assign P[54] = in[165] ^ in2[165];
    assign G[55] = in[164] & in2[164];
    assign P[55] = in[164] ^ in2[164];
    assign G[56] = in[163] & in2[163];
    assign P[56] = in[163] ^ in2[163];
    assign G[57] = in[162] & in2[162];
    assign P[57] = in[162] ^ in2[162];
    assign G[58] = in[161] & in2[161];
    assign P[58] = in[161] ^ in2[161];
    assign G[59] = in[160] & in2[160];
    assign P[59] = in[160] ^ in2[160];
    assign G[60] = in[159] & in2[159];
    assign P[60] = in[159] ^ in2[159];
    assign G[61] = in[158] & in2[158];
    assign P[61] = in[158] ^ in2[158];
    assign G[62] = in[157] & in2[157];
    assign P[62] = in[157] ^ in2[157];
    assign G[63] = in[156] & in2[156];
    assign P[63] = in[156] ^ in2[156];
    assign G[64] = in[155] & in2[155];
    assign P[64] = in[155] ^ in2[155];
    assign G[65] = in[154] & in2[154];
    assign P[65] = in[154] ^ in2[154];
    assign G[66] = in[153] & in2[153];
    assign P[66] = in[153] ^ in2[153];
    assign G[67] = in[152] & in2[152];
    assign P[67] = in[152] ^ in2[152];
    assign G[68] = in[151] & in2[151];
    assign P[68] = in[151] ^ in2[151];
    assign G[69] = in[150] & in2[150];
    assign P[69] = in[150] ^ in2[150];
    assign G[70] = in[149] & in2[149];
    assign P[70] = in[149] ^ in2[149];
    assign G[71] = in[148] & in2[148];
    assign P[71] = in[148] ^ in2[148];
    assign G[72] = in[147] & in2[147];
    assign P[72] = in[147] ^ in2[147];
    assign G[73] = in[146] & in2[146];
    assign P[73] = in[146] ^ in2[146];
    assign G[74] = in[145] & in2[145];
    assign P[74] = in[145] ^ in2[145];
    assign G[75] = in[144] & in2[144];
    assign P[75] = in[144] ^ in2[144];
    assign G[76] = in[143] & in2[143];
    assign P[76] = in[143] ^ in2[143];
    assign G[77] = in[142] & in2[142];
    assign P[77] = in[142] ^ in2[142];
    assign G[78] = in[141] & in2[141];
    assign P[78] = in[141] ^ in2[141];
    assign G[79] = in[140] & in2[140];
    assign P[79] = in[140] ^ in2[140];
    assign G[80] = in[139] & in2[139];
    assign P[80] = in[139] ^ in2[139];
    assign G[81] = in[138] & in2[138];
    assign P[81] = in[138] ^ in2[138];
    assign G[82] = in[137] & in2[137];
    assign P[82] = in[137] ^ in2[137];
    assign G[83] = in[136] & in2[136];
    assign P[83] = in[136] ^ in2[136];
    assign G[84] = in[135] & in2[135];
    assign P[84] = in[135] ^ in2[135];
    assign G[85] = in[134] & in2[134];
    assign P[85] = in[134] ^ in2[134];
    assign G[86] = in[133] & in2[133];
    assign P[86] = in[133] ^ in2[133];
    assign G[87] = in[132] & in2[132];
    assign P[87] = in[132] ^ in2[132];
    assign G[88] = in[131] & in2[131];
    assign P[88] = in[131] ^ in2[131];
    assign G[89] = in[130] & in2[130];
    assign P[89] = in[130] ^ in2[130];
    assign G[90] = in[129] & in2[129];
    assign P[90] = in[129] ^ in2[129];
    assign G[91] = in[128] & in2[128];
    assign P[91] = in[128] ^ in2[128];
    assign G[92] = in[127] & in2[127];
    assign P[92] = in[127] ^ in2[127];
    assign G[93] = in[126] & in2[126];
    assign P[93] = in[126] ^ in2[126];
    assign G[94] = in[125] & in2[125];
    assign P[94] = in[125] ^ in2[125];
    assign G[95] = in[124] & in2[124];
    assign P[95] = in[124] ^ in2[124];
    assign G[96] = in[123] & in2[123];
    assign P[96] = in[123] ^ in2[123];
    assign G[97] = in[122] & in2[122];
    assign P[97] = in[122] ^ in2[122];
    assign G[98] = in[121] & in2[121];
    assign P[98] = in[121] ^ in2[121];
    assign G[99] = in[120] & in2[120];
    assign P[99] = in[120] ^ in2[120];
    assign G[100] = in[119] & in2[119];
    assign P[100] = in[119] ^ in2[119];
    assign G[101] = in[118] & in2[118];
    assign P[101] = in[118] ^ in2[118];
    assign G[102] = in[117] & in2[117];
    assign P[102] = in[117] ^ in2[117];
    assign G[103] = in[116] & in2[116];
    assign P[103] = in[116] ^ in2[116];
    assign G[104] = in[115] & in2[115];
    assign P[104] = in[115] ^ in2[115];
    assign G[105] = in[114] & in2[114];
    assign P[105] = in[114] ^ in2[114];
    assign G[106] = in[113] & in2[113];
    assign P[106] = in[113] ^ in2[113];
    assign G[107] = in[112] & in2[112];
    assign P[107] = in[112] ^ in2[112];
    assign G[108] = in[111] & in2[111];
    assign P[108] = in[111] ^ in2[111];
    assign G[109] = in[110] & in2[110];
    assign P[109] = in[110] ^ in2[110];
    assign G[110] = in[109] & in2[109];
    assign P[110] = in[109] ^ in2[109];
    assign G[111] = in[108] & in2[108];
    assign P[111] = in[108] ^ in2[108];
    assign G[112] = in[107] & in2[107];
    assign P[112] = in[107] ^ in2[107];
    assign G[113] = in[106] & in2[106];
    assign P[113] = in[106] ^ in2[106];
    assign G[114] = in[105] & in2[105];
    assign P[114] = in[105] ^ in2[105];
    assign G[115] = in[104] & in2[104];
    assign P[115] = in[104] ^ in2[104];
    assign G[116] = in[103] & in2[103];
    assign P[116] = in[103] ^ in2[103];
    assign G[117] = in[102] & in2[102];
    assign P[117] = in[102] ^ in2[102];
    assign G[118] = in[101] & in2[101];
    assign P[118] = in[101] ^ in2[101];
    assign G[119] = in[100] & in2[100];
    assign P[119] = in[100] ^ in2[100];
    assign G[120] = in[99] & in2[99];
    assign P[120] = in[99] ^ in2[99];
    assign G[121] = in[98] & in2[98];
    assign P[121] = in[98] ^ in2[98];
    assign G[122] = in[97] & in2[97];
    assign P[122] = in[97] ^ in2[97];
    assign G[123] = in[96] & in2[96];
    assign P[123] = in[96] ^ in2[96];
    assign G[124] = in[95] & in2[95];
    assign P[124] = in[95] ^ in2[95];
    assign G[125] = in[94] & in2[94];
    assign P[125] = in[94] ^ in2[94];
    assign G[126] = in[93] & in2[93];
    assign P[126] = in[93] ^ in2[93];
    assign G[127] = in[92] & in2[92];
    assign P[127] = in[92] ^ in2[92];
    assign G[128] = in[91] & in2[91];
    assign P[128] = in[91] ^ in2[91];
    assign G[129] = in[90] & in2[90];
    assign P[129] = in[90] ^ in2[90];
    assign G[130] = in[89] & in2[89];
    assign P[130] = in[89] ^ in2[89];
    assign G[131] = in[88] & in2[88];
    assign P[131] = in[88] ^ in2[88];
    assign G[132] = in[87] & in2[87];
    assign P[132] = in[87] ^ in2[87];
    assign G[133] = in[86] & in2[86];
    assign P[133] = in[86] ^ in2[86];
    assign G[134] = in[85] & in2[85];
    assign P[134] = in[85] ^ in2[85];
    assign G[135] = in[84] & in2[84];
    assign P[135] = in[84] ^ in2[84];
    assign G[136] = in[83] & in2[83];
    assign P[136] = in[83] ^ in2[83];
    assign G[137] = in[82] & in2[82];
    assign P[137] = in[82] ^ in2[82];
    assign G[138] = in[81] & in2[81];
    assign P[138] = in[81] ^ in2[81];
    assign G[139] = in[80] & in2[80];
    assign P[139] = in[80] ^ in2[80];
    assign G[140] = in[79] & in2[79];
    assign P[140] = in[79] ^ in2[79];
    assign G[141] = in[78] & in2[78];
    assign P[141] = in[78] ^ in2[78];
    assign G[142] = in[77] & in2[77];
    assign P[142] = in[77] ^ in2[77];
    assign G[143] = in[76] & in2[76];
    assign P[143] = in[76] ^ in2[76];
    assign G[144] = in[75] & in2[75];
    assign P[144] = in[75] ^ in2[75];
    assign G[145] = in[74] & in2[74];
    assign P[145] = in[74] ^ in2[74];
    assign G[146] = in[73] & in2[73];
    assign P[146] = in[73] ^ in2[73];
    assign G[147] = in[72] & in2[72];
    assign P[147] = in[72] ^ in2[72];
    assign G[148] = in[71] & in2[71];
    assign P[148] = in[71] ^ in2[71];
    assign G[149] = in[70] & in2[70];
    assign P[149] = in[70] ^ in2[70];
    assign G[150] = in[69] & in2[69];
    assign P[150] = in[69] ^ in2[69];
    assign G[151] = in[68] & in2[68];
    assign P[151] = in[68] ^ in2[68];
    assign G[152] = in[67] & in2[67];
    assign P[152] = in[67] ^ in2[67];
    assign G[153] = in[66] & in2[66];
    assign P[153] = in[66] ^ in2[66];
    assign G[154] = in[65] & in2[65];
    assign P[154] = in[65] ^ in2[65];
    assign G[155] = in[64] & in2[64];
    assign P[155] = in[64] ^ in2[64];
    assign G[156] = in[63] & in2[63];
    assign P[156] = in[63] ^ in2[63];
    assign G[157] = in[62] & in2[62];
    assign P[157] = in[62] ^ in2[62];
    assign G[158] = in[61] & in2[61];
    assign P[158] = in[61] ^ in2[61];
    assign G[159] = in[60] & in2[60];
    assign P[159] = in[60] ^ in2[60];
    assign G[160] = in[59] & in2[59];
    assign P[160] = in[59] ^ in2[59];
    assign G[161] = in[58] & in2[58];
    assign P[161] = in[58] ^ in2[58];
    assign G[162] = in[57] & in2[57];
    assign P[162] = in[57] ^ in2[57];
    assign G[163] = in[56] & in2[56];
    assign P[163] = in[56] ^ in2[56];
    assign G[164] = in[55] & in2[55];
    assign P[164] = in[55] ^ in2[55];
    assign G[165] = in[54] & in2[54];
    assign P[165] = in[54] ^ in2[54];
    assign G[166] = in[53] & in2[53];
    assign P[166] = in[53] ^ in2[53];
    assign G[167] = in[52] & in2[52];
    assign P[167] = in[52] ^ in2[52];
    assign G[168] = in[51] & in2[51];
    assign P[168] = in[51] ^ in2[51];
    assign G[169] = in[50] & in2[50];
    assign P[169] = in[50] ^ in2[50];
    assign G[170] = in[49] & in2[49];
    assign P[170] = in[49] ^ in2[49];
    assign G[171] = in[48] & in2[48];
    assign P[171] = in[48] ^ in2[48];
    assign G[172] = in[47] & in2[47];
    assign P[172] = in[47] ^ in2[47];
    assign G[173] = in[46] & in2[46];
    assign P[173] = in[46] ^ in2[46];
    assign G[174] = in[45] & in2[45];
    assign P[174] = in[45] ^ in2[45];
    assign G[175] = in[44] & in2[44];
    assign P[175] = in[44] ^ in2[44];
    assign G[176] = in[43] & in2[43];
    assign P[176] = in[43] ^ in2[43];
    assign G[177] = in[42] & in2[42];
    assign P[177] = in[42] ^ in2[42];
    assign G[178] = in[41] & in2[41];
    assign P[178] = in[41] ^ in2[41];
    assign G[179] = in[40] & in2[40];
    assign P[179] = in[40] ^ in2[40];
    assign G[180] = in[39] & in2[39];
    assign P[180] = in[39] ^ in2[39];
    assign G[181] = in[38] & in2[38];
    assign P[181] = in[38] ^ in2[38];
    assign G[182] = in[37] & in2[37];
    assign P[182] = in[37] ^ in2[37];
    assign G[183] = in[36] & in2[36];
    assign P[183] = in[36] ^ in2[36];
    assign G[184] = in[35] & in2[35];
    assign P[184] = in[35] ^ in2[35];
    assign G[185] = in[34] & in2[34];
    assign P[185] = in[34] ^ in2[34];
    assign G[186] = in[33] & in2[33];
    assign P[186] = in[33] ^ in2[33];
    assign G[187] = in[32] & in2[32];
    assign P[187] = in[32] ^ in2[32];
    assign G[188] = in[31] & in2[31];
    assign P[188] = in[31] ^ in2[31];
    assign G[189] = in[30] & in2[30];
    assign P[189] = in[30] ^ in2[30];
    assign G[190] = in[29] & in2[29];
    assign P[190] = in[29] ^ in2[29];
    assign G[191] = in[28] & in2[28];
    assign P[191] = in[28] ^ in2[28];
    assign G[192] = in[27] & in2[27];
    assign P[192] = in[27] ^ in2[27];
    assign G[193] = in[26] & in2[26];
    assign P[193] = in[26] ^ in2[26];
    assign G[194] = in[25] & in2[25];
    assign P[194] = in[25] ^ in2[25];
    assign G[195] = in[24] & in2[24];
    assign P[195] = in[24] ^ in2[24];
    assign G[196] = in[23] & in2[23];
    assign P[196] = in[23] ^ in2[23];
    assign G[197] = in[22] & in2[22];
    assign P[197] = in[22] ^ in2[22];
    assign G[198] = in[21] & in2[21];
    assign P[198] = in[21] ^ in2[21];
    assign G[199] = in[20] & in2[20];
    assign P[199] = in[20] ^ in2[20];
    assign G[200] = in[19] & in2[19];
    assign P[200] = in[19] ^ in2[19];
    assign G[201] = in[18] & in2[18];
    assign P[201] = in[18] ^ in2[18];
    assign G[202] = in[17] & in2[17];
    assign P[202] = in[17] ^ in2[17];
    assign G[203] = in[16] & in2[16];
    assign P[203] = in[16] ^ in2[16];
    assign G[204] = in[15] & in2[15];
    assign P[204] = in[15] ^ in2[15];
    assign G[205] = in[14] & in2[14];
    assign P[205] = in[14] ^ in2[14];
    assign G[206] = in[13] & in2[13];
    assign P[206] = in[13] ^ in2[13];
    assign G[207] = in[12] & in2[12];
    assign P[207] = in[12] ^ in2[12];
    assign G[208] = in[11] & in2[11];
    assign P[208] = in[11] ^ in2[11];
    assign G[209] = in[10] & in2[10];
    assign P[209] = in[10] ^ in2[10];
    assign G[210] = in[9] & in2[9];
    assign P[210] = in[9] ^ in2[9];
    assign G[211] = in[8] & in2[8];
    assign P[211] = in[8] ^ in2[8];
    assign G[212] = in[7] & in2[7];
    assign P[212] = in[7] ^ in2[7];
    assign G[213] = in[6] & in2[6];
    assign P[213] = in[6] ^ in2[6];
    assign G[214] = in[5] & in2[5];
    assign P[214] = in[5] ^ in2[5];
    assign G[215] = in[4] & in2[4];
    assign P[215] = in[4] ^ in2[4];
    assign G[216] = in[3] & in2[3];
    assign P[216] = in[3] ^ in2[3];
    assign G[217] = in[2] & in2[2];
    assign P[217] = in[2] ^ in2[2];
    assign G[218] = in[1] & in2[1];
    assign P[218] = in[1] ^ in2[1];
    assign G[219] = in[0] & in2[0];
    assign P[219] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign C[219] = G[218] | (P[218] & C[218]);
    assign cout = G[219] | (P[219] & C[219]);
    assign sum = P ^ C;
endmodule

module CLA219(output [218:0] sum, output cout, input [218:0] in1, input [218:0] in2;

    wire[218:0] G;
    wire[218:0] C;
    wire[218:0] P;

    assign G[0] = in[218] & in2[218];
    assign P[0] = in[218] ^ in2[218];
    assign G[1] = in[217] & in2[217];
    assign P[1] = in[217] ^ in2[217];
    assign G[2] = in[216] & in2[216];
    assign P[2] = in[216] ^ in2[216];
    assign G[3] = in[215] & in2[215];
    assign P[3] = in[215] ^ in2[215];
    assign G[4] = in[214] & in2[214];
    assign P[4] = in[214] ^ in2[214];
    assign G[5] = in[213] & in2[213];
    assign P[5] = in[213] ^ in2[213];
    assign G[6] = in[212] & in2[212];
    assign P[6] = in[212] ^ in2[212];
    assign G[7] = in[211] & in2[211];
    assign P[7] = in[211] ^ in2[211];
    assign G[8] = in[210] & in2[210];
    assign P[8] = in[210] ^ in2[210];
    assign G[9] = in[209] & in2[209];
    assign P[9] = in[209] ^ in2[209];
    assign G[10] = in[208] & in2[208];
    assign P[10] = in[208] ^ in2[208];
    assign G[11] = in[207] & in2[207];
    assign P[11] = in[207] ^ in2[207];
    assign G[12] = in[206] & in2[206];
    assign P[12] = in[206] ^ in2[206];
    assign G[13] = in[205] & in2[205];
    assign P[13] = in[205] ^ in2[205];
    assign G[14] = in[204] & in2[204];
    assign P[14] = in[204] ^ in2[204];
    assign G[15] = in[203] & in2[203];
    assign P[15] = in[203] ^ in2[203];
    assign G[16] = in[202] & in2[202];
    assign P[16] = in[202] ^ in2[202];
    assign G[17] = in[201] & in2[201];
    assign P[17] = in[201] ^ in2[201];
    assign G[18] = in[200] & in2[200];
    assign P[18] = in[200] ^ in2[200];
    assign G[19] = in[199] & in2[199];
    assign P[19] = in[199] ^ in2[199];
    assign G[20] = in[198] & in2[198];
    assign P[20] = in[198] ^ in2[198];
    assign G[21] = in[197] & in2[197];
    assign P[21] = in[197] ^ in2[197];
    assign G[22] = in[196] & in2[196];
    assign P[22] = in[196] ^ in2[196];
    assign G[23] = in[195] & in2[195];
    assign P[23] = in[195] ^ in2[195];
    assign G[24] = in[194] & in2[194];
    assign P[24] = in[194] ^ in2[194];
    assign G[25] = in[193] & in2[193];
    assign P[25] = in[193] ^ in2[193];
    assign G[26] = in[192] & in2[192];
    assign P[26] = in[192] ^ in2[192];
    assign G[27] = in[191] & in2[191];
    assign P[27] = in[191] ^ in2[191];
    assign G[28] = in[190] & in2[190];
    assign P[28] = in[190] ^ in2[190];
    assign G[29] = in[189] & in2[189];
    assign P[29] = in[189] ^ in2[189];
    assign G[30] = in[188] & in2[188];
    assign P[30] = in[188] ^ in2[188];
    assign G[31] = in[187] & in2[187];
    assign P[31] = in[187] ^ in2[187];
    assign G[32] = in[186] & in2[186];
    assign P[32] = in[186] ^ in2[186];
    assign G[33] = in[185] & in2[185];
    assign P[33] = in[185] ^ in2[185];
    assign G[34] = in[184] & in2[184];
    assign P[34] = in[184] ^ in2[184];
    assign G[35] = in[183] & in2[183];
    assign P[35] = in[183] ^ in2[183];
    assign G[36] = in[182] & in2[182];
    assign P[36] = in[182] ^ in2[182];
    assign G[37] = in[181] & in2[181];
    assign P[37] = in[181] ^ in2[181];
    assign G[38] = in[180] & in2[180];
    assign P[38] = in[180] ^ in2[180];
    assign G[39] = in[179] & in2[179];
    assign P[39] = in[179] ^ in2[179];
    assign G[40] = in[178] & in2[178];
    assign P[40] = in[178] ^ in2[178];
    assign G[41] = in[177] & in2[177];
    assign P[41] = in[177] ^ in2[177];
    assign G[42] = in[176] & in2[176];
    assign P[42] = in[176] ^ in2[176];
    assign G[43] = in[175] & in2[175];
    assign P[43] = in[175] ^ in2[175];
    assign G[44] = in[174] & in2[174];
    assign P[44] = in[174] ^ in2[174];
    assign G[45] = in[173] & in2[173];
    assign P[45] = in[173] ^ in2[173];
    assign G[46] = in[172] & in2[172];
    assign P[46] = in[172] ^ in2[172];
    assign G[47] = in[171] & in2[171];
    assign P[47] = in[171] ^ in2[171];
    assign G[48] = in[170] & in2[170];
    assign P[48] = in[170] ^ in2[170];
    assign G[49] = in[169] & in2[169];
    assign P[49] = in[169] ^ in2[169];
    assign G[50] = in[168] & in2[168];
    assign P[50] = in[168] ^ in2[168];
    assign G[51] = in[167] & in2[167];
    assign P[51] = in[167] ^ in2[167];
    assign G[52] = in[166] & in2[166];
    assign P[52] = in[166] ^ in2[166];
    assign G[53] = in[165] & in2[165];
    assign P[53] = in[165] ^ in2[165];
    assign G[54] = in[164] & in2[164];
    assign P[54] = in[164] ^ in2[164];
    assign G[55] = in[163] & in2[163];
    assign P[55] = in[163] ^ in2[163];
    assign G[56] = in[162] & in2[162];
    assign P[56] = in[162] ^ in2[162];
    assign G[57] = in[161] & in2[161];
    assign P[57] = in[161] ^ in2[161];
    assign G[58] = in[160] & in2[160];
    assign P[58] = in[160] ^ in2[160];
    assign G[59] = in[159] & in2[159];
    assign P[59] = in[159] ^ in2[159];
    assign G[60] = in[158] & in2[158];
    assign P[60] = in[158] ^ in2[158];
    assign G[61] = in[157] & in2[157];
    assign P[61] = in[157] ^ in2[157];
    assign G[62] = in[156] & in2[156];
    assign P[62] = in[156] ^ in2[156];
    assign G[63] = in[155] & in2[155];
    assign P[63] = in[155] ^ in2[155];
    assign G[64] = in[154] & in2[154];
    assign P[64] = in[154] ^ in2[154];
    assign G[65] = in[153] & in2[153];
    assign P[65] = in[153] ^ in2[153];
    assign G[66] = in[152] & in2[152];
    assign P[66] = in[152] ^ in2[152];
    assign G[67] = in[151] & in2[151];
    assign P[67] = in[151] ^ in2[151];
    assign G[68] = in[150] & in2[150];
    assign P[68] = in[150] ^ in2[150];
    assign G[69] = in[149] & in2[149];
    assign P[69] = in[149] ^ in2[149];
    assign G[70] = in[148] & in2[148];
    assign P[70] = in[148] ^ in2[148];
    assign G[71] = in[147] & in2[147];
    assign P[71] = in[147] ^ in2[147];
    assign G[72] = in[146] & in2[146];
    assign P[72] = in[146] ^ in2[146];
    assign G[73] = in[145] & in2[145];
    assign P[73] = in[145] ^ in2[145];
    assign G[74] = in[144] & in2[144];
    assign P[74] = in[144] ^ in2[144];
    assign G[75] = in[143] & in2[143];
    assign P[75] = in[143] ^ in2[143];
    assign G[76] = in[142] & in2[142];
    assign P[76] = in[142] ^ in2[142];
    assign G[77] = in[141] & in2[141];
    assign P[77] = in[141] ^ in2[141];
    assign G[78] = in[140] & in2[140];
    assign P[78] = in[140] ^ in2[140];
    assign G[79] = in[139] & in2[139];
    assign P[79] = in[139] ^ in2[139];
    assign G[80] = in[138] & in2[138];
    assign P[80] = in[138] ^ in2[138];
    assign G[81] = in[137] & in2[137];
    assign P[81] = in[137] ^ in2[137];
    assign G[82] = in[136] & in2[136];
    assign P[82] = in[136] ^ in2[136];
    assign G[83] = in[135] & in2[135];
    assign P[83] = in[135] ^ in2[135];
    assign G[84] = in[134] & in2[134];
    assign P[84] = in[134] ^ in2[134];
    assign G[85] = in[133] & in2[133];
    assign P[85] = in[133] ^ in2[133];
    assign G[86] = in[132] & in2[132];
    assign P[86] = in[132] ^ in2[132];
    assign G[87] = in[131] & in2[131];
    assign P[87] = in[131] ^ in2[131];
    assign G[88] = in[130] & in2[130];
    assign P[88] = in[130] ^ in2[130];
    assign G[89] = in[129] & in2[129];
    assign P[89] = in[129] ^ in2[129];
    assign G[90] = in[128] & in2[128];
    assign P[90] = in[128] ^ in2[128];
    assign G[91] = in[127] & in2[127];
    assign P[91] = in[127] ^ in2[127];
    assign G[92] = in[126] & in2[126];
    assign P[92] = in[126] ^ in2[126];
    assign G[93] = in[125] & in2[125];
    assign P[93] = in[125] ^ in2[125];
    assign G[94] = in[124] & in2[124];
    assign P[94] = in[124] ^ in2[124];
    assign G[95] = in[123] & in2[123];
    assign P[95] = in[123] ^ in2[123];
    assign G[96] = in[122] & in2[122];
    assign P[96] = in[122] ^ in2[122];
    assign G[97] = in[121] & in2[121];
    assign P[97] = in[121] ^ in2[121];
    assign G[98] = in[120] & in2[120];
    assign P[98] = in[120] ^ in2[120];
    assign G[99] = in[119] & in2[119];
    assign P[99] = in[119] ^ in2[119];
    assign G[100] = in[118] & in2[118];
    assign P[100] = in[118] ^ in2[118];
    assign G[101] = in[117] & in2[117];
    assign P[101] = in[117] ^ in2[117];
    assign G[102] = in[116] & in2[116];
    assign P[102] = in[116] ^ in2[116];
    assign G[103] = in[115] & in2[115];
    assign P[103] = in[115] ^ in2[115];
    assign G[104] = in[114] & in2[114];
    assign P[104] = in[114] ^ in2[114];
    assign G[105] = in[113] & in2[113];
    assign P[105] = in[113] ^ in2[113];
    assign G[106] = in[112] & in2[112];
    assign P[106] = in[112] ^ in2[112];
    assign G[107] = in[111] & in2[111];
    assign P[107] = in[111] ^ in2[111];
    assign G[108] = in[110] & in2[110];
    assign P[108] = in[110] ^ in2[110];
    assign G[109] = in[109] & in2[109];
    assign P[109] = in[109] ^ in2[109];
    assign G[110] = in[108] & in2[108];
    assign P[110] = in[108] ^ in2[108];
    assign G[111] = in[107] & in2[107];
    assign P[111] = in[107] ^ in2[107];
    assign G[112] = in[106] & in2[106];
    assign P[112] = in[106] ^ in2[106];
    assign G[113] = in[105] & in2[105];
    assign P[113] = in[105] ^ in2[105];
    assign G[114] = in[104] & in2[104];
    assign P[114] = in[104] ^ in2[104];
    assign G[115] = in[103] & in2[103];
    assign P[115] = in[103] ^ in2[103];
    assign G[116] = in[102] & in2[102];
    assign P[116] = in[102] ^ in2[102];
    assign G[117] = in[101] & in2[101];
    assign P[117] = in[101] ^ in2[101];
    assign G[118] = in[100] & in2[100];
    assign P[118] = in[100] ^ in2[100];
    assign G[119] = in[99] & in2[99];
    assign P[119] = in[99] ^ in2[99];
    assign G[120] = in[98] & in2[98];
    assign P[120] = in[98] ^ in2[98];
    assign G[121] = in[97] & in2[97];
    assign P[121] = in[97] ^ in2[97];
    assign G[122] = in[96] & in2[96];
    assign P[122] = in[96] ^ in2[96];
    assign G[123] = in[95] & in2[95];
    assign P[123] = in[95] ^ in2[95];
    assign G[124] = in[94] & in2[94];
    assign P[124] = in[94] ^ in2[94];
    assign G[125] = in[93] & in2[93];
    assign P[125] = in[93] ^ in2[93];
    assign G[126] = in[92] & in2[92];
    assign P[126] = in[92] ^ in2[92];
    assign G[127] = in[91] & in2[91];
    assign P[127] = in[91] ^ in2[91];
    assign G[128] = in[90] & in2[90];
    assign P[128] = in[90] ^ in2[90];
    assign G[129] = in[89] & in2[89];
    assign P[129] = in[89] ^ in2[89];
    assign G[130] = in[88] & in2[88];
    assign P[130] = in[88] ^ in2[88];
    assign G[131] = in[87] & in2[87];
    assign P[131] = in[87] ^ in2[87];
    assign G[132] = in[86] & in2[86];
    assign P[132] = in[86] ^ in2[86];
    assign G[133] = in[85] & in2[85];
    assign P[133] = in[85] ^ in2[85];
    assign G[134] = in[84] & in2[84];
    assign P[134] = in[84] ^ in2[84];
    assign G[135] = in[83] & in2[83];
    assign P[135] = in[83] ^ in2[83];
    assign G[136] = in[82] & in2[82];
    assign P[136] = in[82] ^ in2[82];
    assign G[137] = in[81] & in2[81];
    assign P[137] = in[81] ^ in2[81];
    assign G[138] = in[80] & in2[80];
    assign P[138] = in[80] ^ in2[80];
    assign G[139] = in[79] & in2[79];
    assign P[139] = in[79] ^ in2[79];
    assign G[140] = in[78] & in2[78];
    assign P[140] = in[78] ^ in2[78];
    assign G[141] = in[77] & in2[77];
    assign P[141] = in[77] ^ in2[77];
    assign G[142] = in[76] & in2[76];
    assign P[142] = in[76] ^ in2[76];
    assign G[143] = in[75] & in2[75];
    assign P[143] = in[75] ^ in2[75];
    assign G[144] = in[74] & in2[74];
    assign P[144] = in[74] ^ in2[74];
    assign G[145] = in[73] & in2[73];
    assign P[145] = in[73] ^ in2[73];
    assign G[146] = in[72] & in2[72];
    assign P[146] = in[72] ^ in2[72];
    assign G[147] = in[71] & in2[71];
    assign P[147] = in[71] ^ in2[71];
    assign G[148] = in[70] & in2[70];
    assign P[148] = in[70] ^ in2[70];
    assign G[149] = in[69] & in2[69];
    assign P[149] = in[69] ^ in2[69];
    assign G[150] = in[68] & in2[68];
    assign P[150] = in[68] ^ in2[68];
    assign G[151] = in[67] & in2[67];
    assign P[151] = in[67] ^ in2[67];
    assign G[152] = in[66] & in2[66];
    assign P[152] = in[66] ^ in2[66];
    assign G[153] = in[65] & in2[65];
    assign P[153] = in[65] ^ in2[65];
    assign G[154] = in[64] & in2[64];
    assign P[154] = in[64] ^ in2[64];
    assign G[155] = in[63] & in2[63];
    assign P[155] = in[63] ^ in2[63];
    assign G[156] = in[62] & in2[62];
    assign P[156] = in[62] ^ in2[62];
    assign G[157] = in[61] & in2[61];
    assign P[157] = in[61] ^ in2[61];
    assign G[158] = in[60] & in2[60];
    assign P[158] = in[60] ^ in2[60];
    assign G[159] = in[59] & in2[59];
    assign P[159] = in[59] ^ in2[59];
    assign G[160] = in[58] & in2[58];
    assign P[160] = in[58] ^ in2[58];
    assign G[161] = in[57] & in2[57];
    assign P[161] = in[57] ^ in2[57];
    assign G[162] = in[56] & in2[56];
    assign P[162] = in[56] ^ in2[56];
    assign G[163] = in[55] & in2[55];
    assign P[163] = in[55] ^ in2[55];
    assign G[164] = in[54] & in2[54];
    assign P[164] = in[54] ^ in2[54];
    assign G[165] = in[53] & in2[53];
    assign P[165] = in[53] ^ in2[53];
    assign G[166] = in[52] & in2[52];
    assign P[166] = in[52] ^ in2[52];
    assign G[167] = in[51] & in2[51];
    assign P[167] = in[51] ^ in2[51];
    assign G[168] = in[50] & in2[50];
    assign P[168] = in[50] ^ in2[50];
    assign G[169] = in[49] & in2[49];
    assign P[169] = in[49] ^ in2[49];
    assign G[170] = in[48] & in2[48];
    assign P[170] = in[48] ^ in2[48];
    assign G[171] = in[47] & in2[47];
    assign P[171] = in[47] ^ in2[47];
    assign G[172] = in[46] & in2[46];
    assign P[172] = in[46] ^ in2[46];
    assign G[173] = in[45] & in2[45];
    assign P[173] = in[45] ^ in2[45];
    assign G[174] = in[44] & in2[44];
    assign P[174] = in[44] ^ in2[44];
    assign G[175] = in[43] & in2[43];
    assign P[175] = in[43] ^ in2[43];
    assign G[176] = in[42] & in2[42];
    assign P[176] = in[42] ^ in2[42];
    assign G[177] = in[41] & in2[41];
    assign P[177] = in[41] ^ in2[41];
    assign G[178] = in[40] & in2[40];
    assign P[178] = in[40] ^ in2[40];
    assign G[179] = in[39] & in2[39];
    assign P[179] = in[39] ^ in2[39];
    assign G[180] = in[38] & in2[38];
    assign P[180] = in[38] ^ in2[38];
    assign G[181] = in[37] & in2[37];
    assign P[181] = in[37] ^ in2[37];
    assign G[182] = in[36] & in2[36];
    assign P[182] = in[36] ^ in2[36];
    assign G[183] = in[35] & in2[35];
    assign P[183] = in[35] ^ in2[35];
    assign G[184] = in[34] & in2[34];
    assign P[184] = in[34] ^ in2[34];
    assign G[185] = in[33] & in2[33];
    assign P[185] = in[33] ^ in2[33];
    assign G[186] = in[32] & in2[32];
    assign P[186] = in[32] ^ in2[32];
    assign G[187] = in[31] & in2[31];
    assign P[187] = in[31] ^ in2[31];
    assign G[188] = in[30] & in2[30];
    assign P[188] = in[30] ^ in2[30];
    assign G[189] = in[29] & in2[29];
    assign P[189] = in[29] ^ in2[29];
    assign G[190] = in[28] & in2[28];
    assign P[190] = in[28] ^ in2[28];
    assign G[191] = in[27] & in2[27];
    assign P[191] = in[27] ^ in2[27];
    assign G[192] = in[26] & in2[26];
    assign P[192] = in[26] ^ in2[26];
    assign G[193] = in[25] & in2[25];
    assign P[193] = in[25] ^ in2[25];
    assign G[194] = in[24] & in2[24];
    assign P[194] = in[24] ^ in2[24];
    assign G[195] = in[23] & in2[23];
    assign P[195] = in[23] ^ in2[23];
    assign G[196] = in[22] & in2[22];
    assign P[196] = in[22] ^ in2[22];
    assign G[197] = in[21] & in2[21];
    assign P[197] = in[21] ^ in2[21];
    assign G[198] = in[20] & in2[20];
    assign P[198] = in[20] ^ in2[20];
    assign G[199] = in[19] & in2[19];
    assign P[199] = in[19] ^ in2[19];
    assign G[200] = in[18] & in2[18];
    assign P[200] = in[18] ^ in2[18];
    assign G[201] = in[17] & in2[17];
    assign P[201] = in[17] ^ in2[17];
    assign G[202] = in[16] & in2[16];
    assign P[202] = in[16] ^ in2[16];
    assign G[203] = in[15] & in2[15];
    assign P[203] = in[15] ^ in2[15];
    assign G[204] = in[14] & in2[14];
    assign P[204] = in[14] ^ in2[14];
    assign G[205] = in[13] & in2[13];
    assign P[205] = in[13] ^ in2[13];
    assign G[206] = in[12] & in2[12];
    assign P[206] = in[12] ^ in2[12];
    assign G[207] = in[11] & in2[11];
    assign P[207] = in[11] ^ in2[11];
    assign G[208] = in[10] & in2[10];
    assign P[208] = in[10] ^ in2[10];
    assign G[209] = in[9] & in2[9];
    assign P[209] = in[9] ^ in2[9];
    assign G[210] = in[8] & in2[8];
    assign P[210] = in[8] ^ in2[8];
    assign G[211] = in[7] & in2[7];
    assign P[211] = in[7] ^ in2[7];
    assign G[212] = in[6] & in2[6];
    assign P[212] = in[6] ^ in2[6];
    assign G[213] = in[5] & in2[5];
    assign P[213] = in[5] ^ in2[5];
    assign G[214] = in[4] & in2[4];
    assign P[214] = in[4] ^ in2[4];
    assign G[215] = in[3] & in2[3];
    assign P[215] = in[3] ^ in2[3];
    assign G[216] = in[2] & in2[2];
    assign P[216] = in[2] ^ in2[2];
    assign G[217] = in[1] & in2[1];
    assign P[217] = in[1] ^ in2[1];
    assign G[218] = in[0] & in2[0];
    assign P[218] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign C[218] = G[217] | (P[217] & C[217]);
    assign cout = G[218] | (P[218] & C[218]);
    assign sum = P ^ C;
endmodule

module CLA218(output [217:0] sum, output cout, input [217:0] in1, input [217:0] in2;

    wire[217:0] G;
    wire[217:0] C;
    wire[217:0] P;

    assign G[0] = in[217] & in2[217];
    assign P[0] = in[217] ^ in2[217];
    assign G[1] = in[216] & in2[216];
    assign P[1] = in[216] ^ in2[216];
    assign G[2] = in[215] & in2[215];
    assign P[2] = in[215] ^ in2[215];
    assign G[3] = in[214] & in2[214];
    assign P[3] = in[214] ^ in2[214];
    assign G[4] = in[213] & in2[213];
    assign P[4] = in[213] ^ in2[213];
    assign G[5] = in[212] & in2[212];
    assign P[5] = in[212] ^ in2[212];
    assign G[6] = in[211] & in2[211];
    assign P[6] = in[211] ^ in2[211];
    assign G[7] = in[210] & in2[210];
    assign P[7] = in[210] ^ in2[210];
    assign G[8] = in[209] & in2[209];
    assign P[8] = in[209] ^ in2[209];
    assign G[9] = in[208] & in2[208];
    assign P[9] = in[208] ^ in2[208];
    assign G[10] = in[207] & in2[207];
    assign P[10] = in[207] ^ in2[207];
    assign G[11] = in[206] & in2[206];
    assign P[11] = in[206] ^ in2[206];
    assign G[12] = in[205] & in2[205];
    assign P[12] = in[205] ^ in2[205];
    assign G[13] = in[204] & in2[204];
    assign P[13] = in[204] ^ in2[204];
    assign G[14] = in[203] & in2[203];
    assign P[14] = in[203] ^ in2[203];
    assign G[15] = in[202] & in2[202];
    assign P[15] = in[202] ^ in2[202];
    assign G[16] = in[201] & in2[201];
    assign P[16] = in[201] ^ in2[201];
    assign G[17] = in[200] & in2[200];
    assign P[17] = in[200] ^ in2[200];
    assign G[18] = in[199] & in2[199];
    assign P[18] = in[199] ^ in2[199];
    assign G[19] = in[198] & in2[198];
    assign P[19] = in[198] ^ in2[198];
    assign G[20] = in[197] & in2[197];
    assign P[20] = in[197] ^ in2[197];
    assign G[21] = in[196] & in2[196];
    assign P[21] = in[196] ^ in2[196];
    assign G[22] = in[195] & in2[195];
    assign P[22] = in[195] ^ in2[195];
    assign G[23] = in[194] & in2[194];
    assign P[23] = in[194] ^ in2[194];
    assign G[24] = in[193] & in2[193];
    assign P[24] = in[193] ^ in2[193];
    assign G[25] = in[192] & in2[192];
    assign P[25] = in[192] ^ in2[192];
    assign G[26] = in[191] & in2[191];
    assign P[26] = in[191] ^ in2[191];
    assign G[27] = in[190] & in2[190];
    assign P[27] = in[190] ^ in2[190];
    assign G[28] = in[189] & in2[189];
    assign P[28] = in[189] ^ in2[189];
    assign G[29] = in[188] & in2[188];
    assign P[29] = in[188] ^ in2[188];
    assign G[30] = in[187] & in2[187];
    assign P[30] = in[187] ^ in2[187];
    assign G[31] = in[186] & in2[186];
    assign P[31] = in[186] ^ in2[186];
    assign G[32] = in[185] & in2[185];
    assign P[32] = in[185] ^ in2[185];
    assign G[33] = in[184] & in2[184];
    assign P[33] = in[184] ^ in2[184];
    assign G[34] = in[183] & in2[183];
    assign P[34] = in[183] ^ in2[183];
    assign G[35] = in[182] & in2[182];
    assign P[35] = in[182] ^ in2[182];
    assign G[36] = in[181] & in2[181];
    assign P[36] = in[181] ^ in2[181];
    assign G[37] = in[180] & in2[180];
    assign P[37] = in[180] ^ in2[180];
    assign G[38] = in[179] & in2[179];
    assign P[38] = in[179] ^ in2[179];
    assign G[39] = in[178] & in2[178];
    assign P[39] = in[178] ^ in2[178];
    assign G[40] = in[177] & in2[177];
    assign P[40] = in[177] ^ in2[177];
    assign G[41] = in[176] & in2[176];
    assign P[41] = in[176] ^ in2[176];
    assign G[42] = in[175] & in2[175];
    assign P[42] = in[175] ^ in2[175];
    assign G[43] = in[174] & in2[174];
    assign P[43] = in[174] ^ in2[174];
    assign G[44] = in[173] & in2[173];
    assign P[44] = in[173] ^ in2[173];
    assign G[45] = in[172] & in2[172];
    assign P[45] = in[172] ^ in2[172];
    assign G[46] = in[171] & in2[171];
    assign P[46] = in[171] ^ in2[171];
    assign G[47] = in[170] & in2[170];
    assign P[47] = in[170] ^ in2[170];
    assign G[48] = in[169] & in2[169];
    assign P[48] = in[169] ^ in2[169];
    assign G[49] = in[168] & in2[168];
    assign P[49] = in[168] ^ in2[168];
    assign G[50] = in[167] & in2[167];
    assign P[50] = in[167] ^ in2[167];
    assign G[51] = in[166] & in2[166];
    assign P[51] = in[166] ^ in2[166];
    assign G[52] = in[165] & in2[165];
    assign P[52] = in[165] ^ in2[165];
    assign G[53] = in[164] & in2[164];
    assign P[53] = in[164] ^ in2[164];
    assign G[54] = in[163] & in2[163];
    assign P[54] = in[163] ^ in2[163];
    assign G[55] = in[162] & in2[162];
    assign P[55] = in[162] ^ in2[162];
    assign G[56] = in[161] & in2[161];
    assign P[56] = in[161] ^ in2[161];
    assign G[57] = in[160] & in2[160];
    assign P[57] = in[160] ^ in2[160];
    assign G[58] = in[159] & in2[159];
    assign P[58] = in[159] ^ in2[159];
    assign G[59] = in[158] & in2[158];
    assign P[59] = in[158] ^ in2[158];
    assign G[60] = in[157] & in2[157];
    assign P[60] = in[157] ^ in2[157];
    assign G[61] = in[156] & in2[156];
    assign P[61] = in[156] ^ in2[156];
    assign G[62] = in[155] & in2[155];
    assign P[62] = in[155] ^ in2[155];
    assign G[63] = in[154] & in2[154];
    assign P[63] = in[154] ^ in2[154];
    assign G[64] = in[153] & in2[153];
    assign P[64] = in[153] ^ in2[153];
    assign G[65] = in[152] & in2[152];
    assign P[65] = in[152] ^ in2[152];
    assign G[66] = in[151] & in2[151];
    assign P[66] = in[151] ^ in2[151];
    assign G[67] = in[150] & in2[150];
    assign P[67] = in[150] ^ in2[150];
    assign G[68] = in[149] & in2[149];
    assign P[68] = in[149] ^ in2[149];
    assign G[69] = in[148] & in2[148];
    assign P[69] = in[148] ^ in2[148];
    assign G[70] = in[147] & in2[147];
    assign P[70] = in[147] ^ in2[147];
    assign G[71] = in[146] & in2[146];
    assign P[71] = in[146] ^ in2[146];
    assign G[72] = in[145] & in2[145];
    assign P[72] = in[145] ^ in2[145];
    assign G[73] = in[144] & in2[144];
    assign P[73] = in[144] ^ in2[144];
    assign G[74] = in[143] & in2[143];
    assign P[74] = in[143] ^ in2[143];
    assign G[75] = in[142] & in2[142];
    assign P[75] = in[142] ^ in2[142];
    assign G[76] = in[141] & in2[141];
    assign P[76] = in[141] ^ in2[141];
    assign G[77] = in[140] & in2[140];
    assign P[77] = in[140] ^ in2[140];
    assign G[78] = in[139] & in2[139];
    assign P[78] = in[139] ^ in2[139];
    assign G[79] = in[138] & in2[138];
    assign P[79] = in[138] ^ in2[138];
    assign G[80] = in[137] & in2[137];
    assign P[80] = in[137] ^ in2[137];
    assign G[81] = in[136] & in2[136];
    assign P[81] = in[136] ^ in2[136];
    assign G[82] = in[135] & in2[135];
    assign P[82] = in[135] ^ in2[135];
    assign G[83] = in[134] & in2[134];
    assign P[83] = in[134] ^ in2[134];
    assign G[84] = in[133] & in2[133];
    assign P[84] = in[133] ^ in2[133];
    assign G[85] = in[132] & in2[132];
    assign P[85] = in[132] ^ in2[132];
    assign G[86] = in[131] & in2[131];
    assign P[86] = in[131] ^ in2[131];
    assign G[87] = in[130] & in2[130];
    assign P[87] = in[130] ^ in2[130];
    assign G[88] = in[129] & in2[129];
    assign P[88] = in[129] ^ in2[129];
    assign G[89] = in[128] & in2[128];
    assign P[89] = in[128] ^ in2[128];
    assign G[90] = in[127] & in2[127];
    assign P[90] = in[127] ^ in2[127];
    assign G[91] = in[126] & in2[126];
    assign P[91] = in[126] ^ in2[126];
    assign G[92] = in[125] & in2[125];
    assign P[92] = in[125] ^ in2[125];
    assign G[93] = in[124] & in2[124];
    assign P[93] = in[124] ^ in2[124];
    assign G[94] = in[123] & in2[123];
    assign P[94] = in[123] ^ in2[123];
    assign G[95] = in[122] & in2[122];
    assign P[95] = in[122] ^ in2[122];
    assign G[96] = in[121] & in2[121];
    assign P[96] = in[121] ^ in2[121];
    assign G[97] = in[120] & in2[120];
    assign P[97] = in[120] ^ in2[120];
    assign G[98] = in[119] & in2[119];
    assign P[98] = in[119] ^ in2[119];
    assign G[99] = in[118] & in2[118];
    assign P[99] = in[118] ^ in2[118];
    assign G[100] = in[117] & in2[117];
    assign P[100] = in[117] ^ in2[117];
    assign G[101] = in[116] & in2[116];
    assign P[101] = in[116] ^ in2[116];
    assign G[102] = in[115] & in2[115];
    assign P[102] = in[115] ^ in2[115];
    assign G[103] = in[114] & in2[114];
    assign P[103] = in[114] ^ in2[114];
    assign G[104] = in[113] & in2[113];
    assign P[104] = in[113] ^ in2[113];
    assign G[105] = in[112] & in2[112];
    assign P[105] = in[112] ^ in2[112];
    assign G[106] = in[111] & in2[111];
    assign P[106] = in[111] ^ in2[111];
    assign G[107] = in[110] & in2[110];
    assign P[107] = in[110] ^ in2[110];
    assign G[108] = in[109] & in2[109];
    assign P[108] = in[109] ^ in2[109];
    assign G[109] = in[108] & in2[108];
    assign P[109] = in[108] ^ in2[108];
    assign G[110] = in[107] & in2[107];
    assign P[110] = in[107] ^ in2[107];
    assign G[111] = in[106] & in2[106];
    assign P[111] = in[106] ^ in2[106];
    assign G[112] = in[105] & in2[105];
    assign P[112] = in[105] ^ in2[105];
    assign G[113] = in[104] & in2[104];
    assign P[113] = in[104] ^ in2[104];
    assign G[114] = in[103] & in2[103];
    assign P[114] = in[103] ^ in2[103];
    assign G[115] = in[102] & in2[102];
    assign P[115] = in[102] ^ in2[102];
    assign G[116] = in[101] & in2[101];
    assign P[116] = in[101] ^ in2[101];
    assign G[117] = in[100] & in2[100];
    assign P[117] = in[100] ^ in2[100];
    assign G[118] = in[99] & in2[99];
    assign P[118] = in[99] ^ in2[99];
    assign G[119] = in[98] & in2[98];
    assign P[119] = in[98] ^ in2[98];
    assign G[120] = in[97] & in2[97];
    assign P[120] = in[97] ^ in2[97];
    assign G[121] = in[96] & in2[96];
    assign P[121] = in[96] ^ in2[96];
    assign G[122] = in[95] & in2[95];
    assign P[122] = in[95] ^ in2[95];
    assign G[123] = in[94] & in2[94];
    assign P[123] = in[94] ^ in2[94];
    assign G[124] = in[93] & in2[93];
    assign P[124] = in[93] ^ in2[93];
    assign G[125] = in[92] & in2[92];
    assign P[125] = in[92] ^ in2[92];
    assign G[126] = in[91] & in2[91];
    assign P[126] = in[91] ^ in2[91];
    assign G[127] = in[90] & in2[90];
    assign P[127] = in[90] ^ in2[90];
    assign G[128] = in[89] & in2[89];
    assign P[128] = in[89] ^ in2[89];
    assign G[129] = in[88] & in2[88];
    assign P[129] = in[88] ^ in2[88];
    assign G[130] = in[87] & in2[87];
    assign P[130] = in[87] ^ in2[87];
    assign G[131] = in[86] & in2[86];
    assign P[131] = in[86] ^ in2[86];
    assign G[132] = in[85] & in2[85];
    assign P[132] = in[85] ^ in2[85];
    assign G[133] = in[84] & in2[84];
    assign P[133] = in[84] ^ in2[84];
    assign G[134] = in[83] & in2[83];
    assign P[134] = in[83] ^ in2[83];
    assign G[135] = in[82] & in2[82];
    assign P[135] = in[82] ^ in2[82];
    assign G[136] = in[81] & in2[81];
    assign P[136] = in[81] ^ in2[81];
    assign G[137] = in[80] & in2[80];
    assign P[137] = in[80] ^ in2[80];
    assign G[138] = in[79] & in2[79];
    assign P[138] = in[79] ^ in2[79];
    assign G[139] = in[78] & in2[78];
    assign P[139] = in[78] ^ in2[78];
    assign G[140] = in[77] & in2[77];
    assign P[140] = in[77] ^ in2[77];
    assign G[141] = in[76] & in2[76];
    assign P[141] = in[76] ^ in2[76];
    assign G[142] = in[75] & in2[75];
    assign P[142] = in[75] ^ in2[75];
    assign G[143] = in[74] & in2[74];
    assign P[143] = in[74] ^ in2[74];
    assign G[144] = in[73] & in2[73];
    assign P[144] = in[73] ^ in2[73];
    assign G[145] = in[72] & in2[72];
    assign P[145] = in[72] ^ in2[72];
    assign G[146] = in[71] & in2[71];
    assign P[146] = in[71] ^ in2[71];
    assign G[147] = in[70] & in2[70];
    assign P[147] = in[70] ^ in2[70];
    assign G[148] = in[69] & in2[69];
    assign P[148] = in[69] ^ in2[69];
    assign G[149] = in[68] & in2[68];
    assign P[149] = in[68] ^ in2[68];
    assign G[150] = in[67] & in2[67];
    assign P[150] = in[67] ^ in2[67];
    assign G[151] = in[66] & in2[66];
    assign P[151] = in[66] ^ in2[66];
    assign G[152] = in[65] & in2[65];
    assign P[152] = in[65] ^ in2[65];
    assign G[153] = in[64] & in2[64];
    assign P[153] = in[64] ^ in2[64];
    assign G[154] = in[63] & in2[63];
    assign P[154] = in[63] ^ in2[63];
    assign G[155] = in[62] & in2[62];
    assign P[155] = in[62] ^ in2[62];
    assign G[156] = in[61] & in2[61];
    assign P[156] = in[61] ^ in2[61];
    assign G[157] = in[60] & in2[60];
    assign P[157] = in[60] ^ in2[60];
    assign G[158] = in[59] & in2[59];
    assign P[158] = in[59] ^ in2[59];
    assign G[159] = in[58] & in2[58];
    assign P[159] = in[58] ^ in2[58];
    assign G[160] = in[57] & in2[57];
    assign P[160] = in[57] ^ in2[57];
    assign G[161] = in[56] & in2[56];
    assign P[161] = in[56] ^ in2[56];
    assign G[162] = in[55] & in2[55];
    assign P[162] = in[55] ^ in2[55];
    assign G[163] = in[54] & in2[54];
    assign P[163] = in[54] ^ in2[54];
    assign G[164] = in[53] & in2[53];
    assign P[164] = in[53] ^ in2[53];
    assign G[165] = in[52] & in2[52];
    assign P[165] = in[52] ^ in2[52];
    assign G[166] = in[51] & in2[51];
    assign P[166] = in[51] ^ in2[51];
    assign G[167] = in[50] & in2[50];
    assign P[167] = in[50] ^ in2[50];
    assign G[168] = in[49] & in2[49];
    assign P[168] = in[49] ^ in2[49];
    assign G[169] = in[48] & in2[48];
    assign P[169] = in[48] ^ in2[48];
    assign G[170] = in[47] & in2[47];
    assign P[170] = in[47] ^ in2[47];
    assign G[171] = in[46] & in2[46];
    assign P[171] = in[46] ^ in2[46];
    assign G[172] = in[45] & in2[45];
    assign P[172] = in[45] ^ in2[45];
    assign G[173] = in[44] & in2[44];
    assign P[173] = in[44] ^ in2[44];
    assign G[174] = in[43] & in2[43];
    assign P[174] = in[43] ^ in2[43];
    assign G[175] = in[42] & in2[42];
    assign P[175] = in[42] ^ in2[42];
    assign G[176] = in[41] & in2[41];
    assign P[176] = in[41] ^ in2[41];
    assign G[177] = in[40] & in2[40];
    assign P[177] = in[40] ^ in2[40];
    assign G[178] = in[39] & in2[39];
    assign P[178] = in[39] ^ in2[39];
    assign G[179] = in[38] & in2[38];
    assign P[179] = in[38] ^ in2[38];
    assign G[180] = in[37] & in2[37];
    assign P[180] = in[37] ^ in2[37];
    assign G[181] = in[36] & in2[36];
    assign P[181] = in[36] ^ in2[36];
    assign G[182] = in[35] & in2[35];
    assign P[182] = in[35] ^ in2[35];
    assign G[183] = in[34] & in2[34];
    assign P[183] = in[34] ^ in2[34];
    assign G[184] = in[33] & in2[33];
    assign P[184] = in[33] ^ in2[33];
    assign G[185] = in[32] & in2[32];
    assign P[185] = in[32] ^ in2[32];
    assign G[186] = in[31] & in2[31];
    assign P[186] = in[31] ^ in2[31];
    assign G[187] = in[30] & in2[30];
    assign P[187] = in[30] ^ in2[30];
    assign G[188] = in[29] & in2[29];
    assign P[188] = in[29] ^ in2[29];
    assign G[189] = in[28] & in2[28];
    assign P[189] = in[28] ^ in2[28];
    assign G[190] = in[27] & in2[27];
    assign P[190] = in[27] ^ in2[27];
    assign G[191] = in[26] & in2[26];
    assign P[191] = in[26] ^ in2[26];
    assign G[192] = in[25] & in2[25];
    assign P[192] = in[25] ^ in2[25];
    assign G[193] = in[24] & in2[24];
    assign P[193] = in[24] ^ in2[24];
    assign G[194] = in[23] & in2[23];
    assign P[194] = in[23] ^ in2[23];
    assign G[195] = in[22] & in2[22];
    assign P[195] = in[22] ^ in2[22];
    assign G[196] = in[21] & in2[21];
    assign P[196] = in[21] ^ in2[21];
    assign G[197] = in[20] & in2[20];
    assign P[197] = in[20] ^ in2[20];
    assign G[198] = in[19] & in2[19];
    assign P[198] = in[19] ^ in2[19];
    assign G[199] = in[18] & in2[18];
    assign P[199] = in[18] ^ in2[18];
    assign G[200] = in[17] & in2[17];
    assign P[200] = in[17] ^ in2[17];
    assign G[201] = in[16] & in2[16];
    assign P[201] = in[16] ^ in2[16];
    assign G[202] = in[15] & in2[15];
    assign P[202] = in[15] ^ in2[15];
    assign G[203] = in[14] & in2[14];
    assign P[203] = in[14] ^ in2[14];
    assign G[204] = in[13] & in2[13];
    assign P[204] = in[13] ^ in2[13];
    assign G[205] = in[12] & in2[12];
    assign P[205] = in[12] ^ in2[12];
    assign G[206] = in[11] & in2[11];
    assign P[206] = in[11] ^ in2[11];
    assign G[207] = in[10] & in2[10];
    assign P[207] = in[10] ^ in2[10];
    assign G[208] = in[9] & in2[9];
    assign P[208] = in[9] ^ in2[9];
    assign G[209] = in[8] & in2[8];
    assign P[209] = in[8] ^ in2[8];
    assign G[210] = in[7] & in2[7];
    assign P[210] = in[7] ^ in2[7];
    assign G[211] = in[6] & in2[6];
    assign P[211] = in[6] ^ in2[6];
    assign G[212] = in[5] & in2[5];
    assign P[212] = in[5] ^ in2[5];
    assign G[213] = in[4] & in2[4];
    assign P[213] = in[4] ^ in2[4];
    assign G[214] = in[3] & in2[3];
    assign P[214] = in[3] ^ in2[3];
    assign G[215] = in[2] & in2[2];
    assign P[215] = in[2] ^ in2[2];
    assign G[216] = in[1] & in2[1];
    assign P[216] = in[1] ^ in2[1];
    assign G[217] = in[0] & in2[0];
    assign P[217] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign C[217] = G[216] | (P[216] & C[216]);
    assign cout = G[217] | (P[217] & C[217]);
    assign sum = P ^ C;
endmodule

module CLA217(output [216:0] sum, output cout, input [216:0] in1, input [216:0] in2;

    wire[216:0] G;
    wire[216:0] C;
    wire[216:0] P;

    assign G[0] = in[216] & in2[216];
    assign P[0] = in[216] ^ in2[216];
    assign G[1] = in[215] & in2[215];
    assign P[1] = in[215] ^ in2[215];
    assign G[2] = in[214] & in2[214];
    assign P[2] = in[214] ^ in2[214];
    assign G[3] = in[213] & in2[213];
    assign P[3] = in[213] ^ in2[213];
    assign G[4] = in[212] & in2[212];
    assign P[4] = in[212] ^ in2[212];
    assign G[5] = in[211] & in2[211];
    assign P[5] = in[211] ^ in2[211];
    assign G[6] = in[210] & in2[210];
    assign P[6] = in[210] ^ in2[210];
    assign G[7] = in[209] & in2[209];
    assign P[7] = in[209] ^ in2[209];
    assign G[8] = in[208] & in2[208];
    assign P[8] = in[208] ^ in2[208];
    assign G[9] = in[207] & in2[207];
    assign P[9] = in[207] ^ in2[207];
    assign G[10] = in[206] & in2[206];
    assign P[10] = in[206] ^ in2[206];
    assign G[11] = in[205] & in2[205];
    assign P[11] = in[205] ^ in2[205];
    assign G[12] = in[204] & in2[204];
    assign P[12] = in[204] ^ in2[204];
    assign G[13] = in[203] & in2[203];
    assign P[13] = in[203] ^ in2[203];
    assign G[14] = in[202] & in2[202];
    assign P[14] = in[202] ^ in2[202];
    assign G[15] = in[201] & in2[201];
    assign P[15] = in[201] ^ in2[201];
    assign G[16] = in[200] & in2[200];
    assign P[16] = in[200] ^ in2[200];
    assign G[17] = in[199] & in2[199];
    assign P[17] = in[199] ^ in2[199];
    assign G[18] = in[198] & in2[198];
    assign P[18] = in[198] ^ in2[198];
    assign G[19] = in[197] & in2[197];
    assign P[19] = in[197] ^ in2[197];
    assign G[20] = in[196] & in2[196];
    assign P[20] = in[196] ^ in2[196];
    assign G[21] = in[195] & in2[195];
    assign P[21] = in[195] ^ in2[195];
    assign G[22] = in[194] & in2[194];
    assign P[22] = in[194] ^ in2[194];
    assign G[23] = in[193] & in2[193];
    assign P[23] = in[193] ^ in2[193];
    assign G[24] = in[192] & in2[192];
    assign P[24] = in[192] ^ in2[192];
    assign G[25] = in[191] & in2[191];
    assign P[25] = in[191] ^ in2[191];
    assign G[26] = in[190] & in2[190];
    assign P[26] = in[190] ^ in2[190];
    assign G[27] = in[189] & in2[189];
    assign P[27] = in[189] ^ in2[189];
    assign G[28] = in[188] & in2[188];
    assign P[28] = in[188] ^ in2[188];
    assign G[29] = in[187] & in2[187];
    assign P[29] = in[187] ^ in2[187];
    assign G[30] = in[186] & in2[186];
    assign P[30] = in[186] ^ in2[186];
    assign G[31] = in[185] & in2[185];
    assign P[31] = in[185] ^ in2[185];
    assign G[32] = in[184] & in2[184];
    assign P[32] = in[184] ^ in2[184];
    assign G[33] = in[183] & in2[183];
    assign P[33] = in[183] ^ in2[183];
    assign G[34] = in[182] & in2[182];
    assign P[34] = in[182] ^ in2[182];
    assign G[35] = in[181] & in2[181];
    assign P[35] = in[181] ^ in2[181];
    assign G[36] = in[180] & in2[180];
    assign P[36] = in[180] ^ in2[180];
    assign G[37] = in[179] & in2[179];
    assign P[37] = in[179] ^ in2[179];
    assign G[38] = in[178] & in2[178];
    assign P[38] = in[178] ^ in2[178];
    assign G[39] = in[177] & in2[177];
    assign P[39] = in[177] ^ in2[177];
    assign G[40] = in[176] & in2[176];
    assign P[40] = in[176] ^ in2[176];
    assign G[41] = in[175] & in2[175];
    assign P[41] = in[175] ^ in2[175];
    assign G[42] = in[174] & in2[174];
    assign P[42] = in[174] ^ in2[174];
    assign G[43] = in[173] & in2[173];
    assign P[43] = in[173] ^ in2[173];
    assign G[44] = in[172] & in2[172];
    assign P[44] = in[172] ^ in2[172];
    assign G[45] = in[171] & in2[171];
    assign P[45] = in[171] ^ in2[171];
    assign G[46] = in[170] & in2[170];
    assign P[46] = in[170] ^ in2[170];
    assign G[47] = in[169] & in2[169];
    assign P[47] = in[169] ^ in2[169];
    assign G[48] = in[168] & in2[168];
    assign P[48] = in[168] ^ in2[168];
    assign G[49] = in[167] & in2[167];
    assign P[49] = in[167] ^ in2[167];
    assign G[50] = in[166] & in2[166];
    assign P[50] = in[166] ^ in2[166];
    assign G[51] = in[165] & in2[165];
    assign P[51] = in[165] ^ in2[165];
    assign G[52] = in[164] & in2[164];
    assign P[52] = in[164] ^ in2[164];
    assign G[53] = in[163] & in2[163];
    assign P[53] = in[163] ^ in2[163];
    assign G[54] = in[162] & in2[162];
    assign P[54] = in[162] ^ in2[162];
    assign G[55] = in[161] & in2[161];
    assign P[55] = in[161] ^ in2[161];
    assign G[56] = in[160] & in2[160];
    assign P[56] = in[160] ^ in2[160];
    assign G[57] = in[159] & in2[159];
    assign P[57] = in[159] ^ in2[159];
    assign G[58] = in[158] & in2[158];
    assign P[58] = in[158] ^ in2[158];
    assign G[59] = in[157] & in2[157];
    assign P[59] = in[157] ^ in2[157];
    assign G[60] = in[156] & in2[156];
    assign P[60] = in[156] ^ in2[156];
    assign G[61] = in[155] & in2[155];
    assign P[61] = in[155] ^ in2[155];
    assign G[62] = in[154] & in2[154];
    assign P[62] = in[154] ^ in2[154];
    assign G[63] = in[153] & in2[153];
    assign P[63] = in[153] ^ in2[153];
    assign G[64] = in[152] & in2[152];
    assign P[64] = in[152] ^ in2[152];
    assign G[65] = in[151] & in2[151];
    assign P[65] = in[151] ^ in2[151];
    assign G[66] = in[150] & in2[150];
    assign P[66] = in[150] ^ in2[150];
    assign G[67] = in[149] & in2[149];
    assign P[67] = in[149] ^ in2[149];
    assign G[68] = in[148] & in2[148];
    assign P[68] = in[148] ^ in2[148];
    assign G[69] = in[147] & in2[147];
    assign P[69] = in[147] ^ in2[147];
    assign G[70] = in[146] & in2[146];
    assign P[70] = in[146] ^ in2[146];
    assign G[71] = in[145] & in2[145];
    assign P[71] = in[145] ^ in2[145];
    assign G[72] = in[144] & in2[144];
    assign P[72] = in[144] ^ in2[144];
    assign G[73] = in[143] & in2[143];
    assign P[73] = in[143] ^ in2[143];
    assign G[74] = in[142] & in2[142];
    assign P[74] = in[142] ^ in2[142];
    assign G[75] = in[141] & in2[141];
    assign P[75] = in[141] ^ in2[141];
    assign G[76] = in[140] & in2[140];
    assign P[76] = in[140] ^ in2[140];
    assign G[77] = in[139] & in2[139];
    assign P[77] = in[139] ^ in2[139];
    assign G[78] = in[138] & in2[138];
    assign P[78] = in[138] ^ in2[138];
    assign G[79] = in[137] & in2[137];
    assign P[79] = in[137] ^ in2[137];
    assign G[80] = in[136] & in2[136];
    assign P[80] = in[136] ^ in2[136];
    assign G[81] = in[135] & in2[135];
    assign P[81] = in[135] ^ in2[135];
    assign G[82] = in[134] & in2[134];
    assign P[82] = in[134] ^ in2[134];
    assign G[83] = in[133] & in2[133];
    assign P[83] = in[133] ^ in2[133];
    assign G[84] = in[132] & in2[132];
    assign P[84] = in[132] ^ in2[132];
    assign G[85] = in[131] & in2[131];
    assign P[85] = in[131] ^ in2[131];
    assign G[86] = in[130] & in2[130];
    assign P[86] = in[130] ^ in2[130];
    assign G[87] = in[129] & in2[129];
    assign P[87] = in[129] ^ in2[129];
    assign G[88] = in[128] & in2[128];
    assign P[88] = in[128] ^ in2[128];
    assign G[89] = in[127] & in2[127];
    assign P[89] = in[127] ^ in2[127];
    assign G[90] = in[126] & in2[126];
    assign P[90] = in[126] ^ in2[126];
    assign G[91] = in[125] & in2[125];
    assign P[91] = in[125] ^ in2[125];
    assign G[92] = in[124] & in2[124];
    assign P[92] = in[124] ^ in2[124];
    assign G[93] = in[123] & in2[123];
    assign P[93] = in[123] ^ in2[123];
    assign G[94] = in[122] & in2[122];
    assign P[94] = in[122] ^ in2[122];
    assign G[95] = in[121] & in2[121];
    assign P[95] = in[121] ^ in2[121];
    assign G[96] = in[120] & in2[120];
    assign P[96] = in[120] ^ in2[120];
    assign G[97] = in[119] & in2[119];
    assign P[97] = in[119] ^ in2[119];
    assign G[98] = in[118] & in2[118];
    assign P[98] = in[118] ^ in2[118];
    assign G[99] = in[117] & in2[117];
    assign P[99] = in[117] ^ in2[117];
    assign G[100] = in[116] & in2[116];
    assign P[100] = in[116] ^ in2[116];
    assign G[101] = in[115] & in2[115];
    assign P[101] = in[115] ^ in2[115];
    assign G[102] = in[114] & in2[114];
    assign P[102] = in[114] ^ in2[114];
    assign G[103] = in[113] & in2[113];
    assign P[103] = in[113] ^ in2[113];
    assign G[104] = in[112] & in2[112];
    assign P[104] = in[112] ^ in2[112];
    assign G[105] = in[111] & in2[111];
    assign P[105] = in[111] ^ in2[111];
    assign G[106] = in[110] & in2[110];
    assign P[106] = in[110] ^ in2[110];
    assign G[107] = in[109] & in2[109];
    assign P[107] = in[109] ^ in2[109];
    assign G[108] = in[108] & in2[108];
    assign P[108] = in[108] ^ in2[108];
    assign G[109] = in[107] & in2[107];
    assign P[109] = in[107] ^ in2[107];
    assign G[110] = in[106] & in2[106];
    assign P[110] = in[106] ^ in2[106];
    assign G[111] = in[105] & in2[105];
    assign P[111] = in[105] ^ in2[105];
    assign G[112] = in[104] & in2[104];
    assign P[112] = in[104] ^ in2[104];
    assign G[113] = in[103] & in2[103];
    assign P[113] = in[103] ^ in2[103];
    assign G[114] = in[102] & in2[102];
    assign P[114] = in[102] ^ in2[102];
    assign G[115] = in[101] & in2[101];
    assign P[115] = in[101] ^ in2[101];
    assign G[116] = in[100] & in2[100];
    assign P[116] = in[100] ^ in2[100];
    assign G[117] = in[99] & in2[99];
    assign P[117] = in[99] ^ in2[99];
    assign G[118] = in[98] & in2[98];
    assign P[118] = in[98] ^ in2[98];
    assign G[119] = in[97] & in2[97];
    assign P[119] = in[97] ^ in2[97];
    assign G[120] = in[96] & in2[96];
    assign P[120] = in[96] ^ in2[96];
    assign G[121] = in[95] & in2[95];
    assign P[121] = in[95] ^ in2[95];
    assign G[122] = in[94] & in2[94];
    assign P[122] = in[94] ^ in2[94];
    assign G[123] = in[93] & in2[93];
    assign P[123] = in[93] ^ in2[93];
    assign G[124] = in[92] & in2[92];
    assign P[124] = in[92] ^ in2[92];
    assign G[125] = in[91] & in2[91];
    assign P[125] = in[91] ^ in2[91];
    assign G[126] = in[90] & in2[90];
    assign P[126] = in[90] ^ in2[90];
    assign G[127] = in[89] & in2[89];
    assign P[127] = in[89] ^ in2[89];
    assign G[128] = in[88] & in2[88];
    assign P[128] = in[88] ^ in2[88];
    assign G[129] = in[87] & in2[87];
    assign P[129] = in[87] ^ in2[87];
    assign G[130] = in[86] & in2[86];
    assign P[130] = in[86] ^ in2[86];
    assign G[131] = in[85] & in2[85];
    assign P[131] = in[85] ^ in2[85];
    assign G[132] = in[84] & in2[84];
    assign P[132] = in[84] ^ in2[84];
    assign G[133] = in[83] & in2[83];
    assign P[133] = in[83] ^ in2[83];
    assign G[134] = in[82] & in2[82];
    assign P[134] = in[82] ^ in2[82];
    assign G[135] = in[81] & in2[81];
    assign P[135] = in[81] ^ in2[81];
    assign G[136] = in[80] & in2[80];
    assign P[136] = in[80] ^ in2[80];
    assign G[137] = in[79] & in2[79];
    assign P[137] = in[79] ^ in2[79];
    assign G[138] = in[78] & in2[78];
    assign P[138] = in[78] ^ in2[78];
    assign G[139] = in[77] & in2[77];
    assign P[139] = in[77] ^ in2[77];
    assign G[140] = in[76] & in2[76];
    assign P[140] = in[76] ^ in2[76];
    assign G[141] = in[75] & in2[75];
    assign P[141] = in[75] ^ in2[75];
    assign G[142] = in[74] & in2[74];
    assign P[142] = in[74] ^ in2[74];
    assign G[143] = in[73] & in2[73];
    assign P[143] = in[73] ^ in2[73];
    assign G[144] = in[72] & in2[72];
    assign P[144] = in[72] ^ in2[72];
    assign G[145] = in[71] & in2[71];
    assign P[145] = in[71] ^ in2[71];
    assign G[146] = in[70] & in2[70];
    assign P[146] = in[70] ^ in2[70];
    assign G[147] = in[69] & in2[69];
    assign P[147] = in[69] ^ in2[69];
    assign G[148] = in[68] & in2[68];
    assign P[148] = in[68] ^ in2[68];
    assign G[149] = in[67] & in2[67];
    assign P[149] = in[67] ^ in2[67];
    assign G[150] = in[66] & in2[66];
    assign P[150] = in[66] ^ in2[66];
    assign G[151] = in[65] & in2[65];
    assign P[151] = in[65] ^ in2[65];
    assign G[152] = in[64] & in2[64];
    assign P[152] = in[64] ^ in2[64];
    assign G[153] = in[63] & in2[63];
    assign P[153] = in[63] ^ in2[63];
    assign G[154] = in[62] & in2[62];
    assign P[154] = in[62] ^ in2[62];
    assign G[155] = in[61] & in2[61];
    assign P[155] = in[61] ^ in2[61];
    assign G[156] = in[60] & in2[60];
    assign P[156] = in[60] ^ in2[60];
    assign G[157] = in[59] & in2[59];
    assign P[157] = in[59] ^ in2[59];
    assign G[158] = in[58] & in2[58];
    assign P[158] = in[58] ^ in2[58];
    assign G[159] = in[57] & in2[57];
    assign P[159] = in[57] ^ in2[57];
    assign G[160] = in[56] & in2[56];
    assign P[160] = in[56] ^ in2[56];
    assign G[161] = in[55] & in2[55];
    assign P[161] = in[55] ^ in2[55];
    assign G[162] = in[54] & in2[54];
    assign P[162] = in[54] ^ in2[54];
    assign G[163] = in[53] & in2[53];
    assign P[163] = in[53] ^ in2[53];
    assign G[164] = in[52] & in2[52];
    assign P[164] = in[52] ^ in2[52];
    assign G[165] = in[51] & in2[51];
    assign P[165] = in[51] ^ in2[51];
    assign G[166] = in[50] & in2[50];
    assign P[166] = in[50] ^ in2[50];
    assign G[167] = in[49] & in2[49];
    assign P[167] = in[49] ^ in2[49];
    assign G[168] = in[48] & in2[48];
    assign P[168] = in[48] ^ in2[48];
    assign G[169] = in[47] & in2[47];
    assign P[169] = in[47] ^ in2[47];
    assign G[170] = in[46] & in2[46];
    assign P[170] = in[46] ^ in2[46];
    assign G[171] = in[45] & in2[45];
    assign P[171] = in[45] ^ in2[45];
    assign G[172] = in[44] & in2[44];
    assign P[172] = in[44] ^ in2[44];
    assign G[173] = in[43] & in2[43];
    assign P[173] = in[43] ^ in2[43];
    assign G[174] = in[42] & in2[42];
    assign P[174] = in[42] ^ in2[42];
    assign G[175] = in[41] & in2[41];
    assign P[175] = in[41] ^ in2[41];
    assign G[176] = in[40] & in2[40];
    assign P[176] = in[40] ^ in2[40];
    assign G[177] = in[39] & in2[39];
    assign P[177] = in[39] ^ in2[39];
    assign G[178] = in[38] & in2[38];
    assign P[178] = in[38] ^ in2[38];
    assign G[179] = in[37] & in2[37];
    assign P[179] = in[37] ^ in2[37];
    assign G[180] = in[36] & in2[36];
    assign P[180] = in[36] ^ in2[36];
    assign G[181] = in[35] & in2[35];
    assign P[181] = in[35] ^ in2[35];
    assign G[182] = in[34] & in2[34];
    assign P[182] = in[34] ^ in2[34];
    assign G[183] = in[33] & in2[33];
    assign P[183] = in[33] ^ in2[33];
    assign G[184] = in[32] & in2[32];
    assign P[184] = in[32] ^ in2[32];
    assign G[185] = in[31] & in2[31];
    assign P[185] = in[31] ^ in2[31];
    assign G[186] = in[30] & in2[30];
    assign P[186] = in[30] ^ in2[30];
    assign G[187] = in[29] & in2[29];
    assign P[187] = in[29] ^ in2[29];
    assign G[188] = in[28] & in2[28];
    assign P[188] = in[28] ^ in2[28];
    assign G[189] = in[27] & in2[27];
    assign P[189] = in[27] ^ in2[27];
    assign G[190] = in[26] & in2[26];
    assign P[190] = in[26] ^ in2[26];
    assign G[191] = in[25] & in2[25];
    assign P[191] = in[25] ^ in2[25];
    assign G[192] = in[24] & in2[24];
    assign P[192] = in[24] ^ in2[24];
    assign G[193] = in[23] & in2[23];
    assign P[193] = in[23] ^ in2[23];
    assign G[194] = in[22] & in2[22];
    assign P[194] = in[22] ^ in2[22];
    assign G[195] = in[21] & in2[21];
    assign P[195] = in[21] ^ in2[21];
    assign G[196] = in[20] & in2[20];
    assign P[196] = in[20] ^ in2[20];
    assign G[197] = in[19] & in2[19];
    assign P[197] = in[19] ^ in2[19];
    assign G[198] = in[18] & in2[18];
    assign P[198] = in[18] ^ in2[18];
    assign G[199] = in[17] & in2[17];
    assign P[199] = in[17] ^ in2[17];
    assign G[200] = in[16] & in2[16];
    assign P[200] = in[16] ^ in2[16];
    assign G[201] = in[15] & in2[15];
    assign P[201] = in[15] ^ in2[15];
    assign G[202] = in[14] & in2[14];
    assign P[202] = in[14] ^ in2[14];
    assign G[203] = in[13] & in2[13];
    assign P[203] = in[13] ^ in2[13];
    assign G[204] = in[12] & in2[12];
    assign P[204] = in[12] ^ in2[12];
    assign G[205] = in[11] & in2[11];
    assign P[205] = in[11] ^ in2[11];
    assign G[206] = in[10] & in2[10];
    assign P[206] = in[10] ^ in2[10];
    assign G[207] = in[9] & in2[9];
    assign P[207] = in[9] ^ in2[9];
    assign G[208] = in[8] & in2[8];
    assign P[208] = in[8] ^ in2[8];
    assign G[209] = in[7] & in2[7];
    assign P[209] = in[7] ^ in2[7];
    assign G[210] = in[6] & in2[6];
    assign P[210] = in[6] ^ in2[6];
    assign G[211] = in[5] & in2[5];
    assign P[211] = in[5] ^ in2[5];
    assign G[212] = in[4] & in2[4];
    assign P[212] = in[4] ^ in2[4];
    assign G[213] = in[3] & in2[3];
    assign P[213] = in[3] ^ in2[3];
    assign G[214] = in[2] & in2[2];
    assign P[214] = in[2] ^ in2[2];
    assign G[215] = in[1] & in2[1];
    assign P[215] = in[1] ^ in2[1];
    assign G[216] = in[0] & in2[0];
    assign P[216] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign C[216] = G[215] | (P[215] & C[215]);
    assign cout = G[216] | (P[216] & C[216]);
    assign sum = P ^ C;
endmodule

module CLA216(output [215:0] sum, output cout, input [215:0] in1, input [215:0] in2;

    wire[215:0] G;
    wire[215:0] C;
    wire[215:0] P;

    assign G[0] = in[215] & in2[215];
    assign P[0] = in[215] ^ in2[215];
    assign G[1] = in[214] & in2[214];
    assign P[1] = in[214] ^ in2[214];
    assign G[2] = in[213] & in2[213];
    assign P[2] = in[213] ^ in2[213];
    assign G[3] = in[212] & in2[212];
    assign P[3] = in[212] ^ in2[212];
    assign G[4] = in[211] & in2[211];
    assign P[4] = in[211] ^ in2[211];
    assign G[5] = in[210] & in2[210];
    assign P[5] = in[210] ^ in2[210];
    assign G[6] = in[209] & in2[209];
    assign P[6] = in[209] ^ in2[209];
    assign G[7] = in[208] & in2[208];
    assign P[7] = in[208] ^ in2[208];
    assign G[8] = in[207] & in2[207];
    assign P[8] = in[207] ^ in2[207];
    assign G[9] = in[206] & in2[206];
    assign P[9] = in[206] ^ in2[206];
    assign G[10] = in[205] & in2[205];
    assign P[10] = in[205] ^ in2[205];
    assign G[11] = in[204] & in2[204];
    assign P[11] = in[204] ^ in2[204];
    assign G[12] = in[203] & in2[203];
    assign P[12] = in[203] ^ in2[203];
    assign G[13] = in[202] & in2[202];
    assign P[13] = in[202] ^ in2[202];
    assign G[14] = in[201] & in2[201];
    assign P[14] = in[201] ^ in2[201];
    assign G[15] = in[200] & in2[200];
    assign P[15] = in[200] ^ in2[200];
    assign G[16] = in[199] & in2[199];
    assign P[16] = in[199] ^ in2[199];
    assign G[17] = in[198] & in2[198];
    assign P[17] = in[198] ^ in2[198];
    assign G[18] = in[197] & in2[197];
    assign P[18] = in[197] ^ in2[197];
    assign G[19] = in[196] & in2[196];
    assign P[19] = in[196] ^ in2[196];
    assign G[20] = in[195] & in2[195];
    assign P[20] = in[195] ^ in2[195];
    assign G[21] = in[194] & in2[194];
    assign P[21] = in[194] ^ in2[194];
    assign G[22] = in[193] & in2[193];
    assign P[22] = in[193] ^ in2[193];
    assign G[23] = in[192] & in2[192];
    assign P[23] = in[192] ^ in2[192];
    assign G[24] = in[191] & in2[191];
    assign P[24] = in[191] ^ in2[191];
    assign G[25] = in[190] & in2[190];
    assign P[25] = in[190] ^ in2[190];
    assign G[26] = in[189] & in2[189];
    assign P[26] = in[189] ^ in2[189];
    assign G[27] = in[188] & in2[188];
    assign P[27] = in[188] ^ in2[188];
    assign G[28] = in[187] & in2[187];
    assign P[28] = in[187] ^ in2[187];
    assign G[29] = in[186] & in2[186];
    assign P[29] = in[186] ^ in2[186];
    assign G[30] = in[185] & in2[185];
    assign P[30] = in[185] ^ in2[185];
    assign G[31] = in[184] & in2[184];
    assign P[31] = in[184] ^ in2[184];
    assign G[32] = in[183] & in2[183];
    assign P[32] = in[183] ^ in2[183];
    assign G[33] = in[182] & in2[182];
    assign P[33] = in[182] ^ in2[182];
    assign G[34] = in[181] & in2[181];
    assign P[34] = in[181] ^ in2[181];
    assign G[35] = in[180] & in2[180];
    assign P[35] = in[180] ^ in2[180];
    assign G[36] = in[179] & in2[179];
    assign P[36] = in[179] ^ in2[179];
    assign G[37] = in[178] & in2[178];
    assign P[37] = in[178] ^ in2[178];
    assign G[38] = in[177] & in2[177];
    assign P[38] = in[177] ^ in2[177];
    assign G[39] = in[176] & in2[176];
    assign P[39] = in[176] ^ in2[176];
    assign G[40] = in[175] & in2[175];
    assign P[40] = in[175] ^ in2[175];
    assign G[41] = in[174] & in2[174];
    assign P[41] = in[174] ^ in2[174];
    assign G[42] = in[173] & in2[173];
    assign P[42] = in[173] ^ in2[173];
    assign G[43] = in[172] & in2[172];
    assign P[43] = in[172] ^ in2[172];
    assign G[44] = in[171] & in2[171];
    assign P[44] = in[171] ^ in2[171];
    assign G[45] = in[170] & in2[170];
    assign P[45] = in[170] ^ in2[170];
    assign G[46] = in[169] & in2[169];
    assign P[46] = in[169] ^ in2[169];
    assign G[47] = in[168] & in2[168];
    assign P[47] = in[168] ^ in2[168];
    assign G[48] = in[167] & in2[167];
    assign P[48] = in[167] ^ in2[167];
    assign G[49] = in[166] & in2[166];
    assign P[49] = in[166] ^ in2[166];
    assign G[50] = in[165] & in2[165];
    assign P[50] = in[165] ^ in2[165];
    assign G[51] = in[164] & in2[164];
    assign P[51] = in[164] ^ in2[164];
    assign G[52] = in[163] & in2[163];
    assign P[52] = in[163] ^ in2[163];
    assign G[53] = in[162] & in2[162];
    assign P[53] = in[162] ^ in2[162];
    assign G[54] = in[161] & in2[161];
    assign P[54] = in[161] ^ in2[161];
    assign G[55] = in[160] & in2[160];
    assign P[55] = in[160] ^ in2[160];
    assign G[56] = in[159] & in2[159];
    assign P[56] = in[159] ^ in2[159];
    assign G[57] = in[158] & in2[158];
    assign P[57] = in[158] ^ in2[158];
    assign G[58] = in[157] & in2[157];
    assign P[58] = in[157] ^ in2[157];
    assign G[59] = in[156] & in2[156];
    assign P[59] = in[156] ^ in2[156];
    assign G[60] = in[155] & in2[155];
    assign P[60] = in[155] ^ in2[155];
    assign G[61] = in[154] & in2[154];
    assign P[61] = in[154] ^ in2[154];
    assign G[62] = in[153] & in2[153];
    assign P[62] = in[153] ^ in2[153];
    assign G[63] = in[152] & in2[152];
    assign P[63] = in[152] ^ in2[152];
    assign G[64] = in[151] & in2[151];
    assign P[64] = in[151] ^ in2[151];
    assign G[65] = in[150] & in2[150];
    assign P[65] = in[150] ^ in2[150];
    assign G[66] = in[149] & in2[149];
    assign P[66] = in[149] ^ in2[149];
    assign G[67] = in[148] & in2[148];
    assign P[67] = in[148] ^ in2[148];
    assign G[68] = in[147] & in2[147];
    assign P[68] = in[147] ^ in2[147];
    assign G[69] = in[146] & in2[146];
    assign P[69] = in[146] ^ in2[146];
    assign G[70] = in[145] & in2[145];
    assign P[70] = in[145] ^ in2[145];
    assign G[71] = in[144] & in2[144];
    assign P[71] = in[144] ^ in2[144];
    assign G[72] = in[143] & in2[143];
    assign P[72] = in[143] ^ in2[143];
    assign G[73] = in[142] & in2[142];
    assign P[73] = in[142] ^ in2[142];
    assign G[74] = in[141] & in2[141];
    assign P[74] = in[141] ^ in2[141];
    assign G[75] = in[140] & in2[140];
    assign P[75] = in[140] ^ in2[140];
    assign G[76] = in[139] & in2[139];
    assign P[76] = in[139] ^ in2[139];
    assign G[77] = in[138] & in2[138];
    assign P[77] = in[138] ^ in2[138];
    assign G[78] = in[137] & in2[137];
    assign P[78] = in[137] ^ in2[137];
    assign G[79] = in[136] & in2[136];
    assign P[79] = in[136] ^ in2[136];
    assign G[80] = in[135] & in2[135];
    assign P[80] = in[135] ^ in2[135];
    assign G[81] = in[134] & in2[134];
    assign P[81] = in[134] ^ in2[134];
    assign G[82] = in[133] & in2[133];
    assign P[82] = in[133] ^ in2[133];
    assign G[83] = in[132] & in2[132];
    assign P[83] = in[132] ^ in2[132];
    assign G[84] = in[131] & in2[131];
    assign P[84] = in[131] ^ in2[131];
    assign G[85] = in[130] & in2[130];
    assign P[85] = in[130] ^ in2[130];
    assign G[86] = in[129] & in2[129];
    assign P[86] = in[129] ^ in2[129];
    assign G[87] = in[128] & in2[128];
    assign P[87] = in[128] ^ in2[128];
    assign G[88] = in[127] & in2[127];
    assign P[88] = in[127] ^ in2[127];
    assign G[89] = in[126] & in2[126];
    assign P[89] = in[126] ^ in2[126];
    assign G[90] = in[125] & in2[125];
    assign P[90] = in[125] ^ in2[125];
    assign G[91] = in[124] & in2[124];
    assign P[91] = in[124] ^ in2[124];
    assign G[92] = in[123] & in2[123];
    assign P[92] = in[123] ^ in2[123];
    assign G[93] = in[122] & in2[122];
    assign P[93] = in[122] ^ in2[122];
    assign G[94] = in[121] & in2[121];
    assign P[94] = in[121] ^ in2[121];
    assign G[95] = in[120] & in2[120];
    assign P[95] = in[120] ^ in2[120];
    assign G[96] = in[119] & in2[119];
    assign P[96] = in[119] ^ in2[119];
    assign G[97] = in[118] & in2[118];
    assign P[97] = in[118] ^ in2[118];
    assign G[98] = in[117] & in2[117];
    assign P[98] = in[117] ^ in2[117];
    assign G[99] = in[116] & in2[116];
    assign P[99] = in[116] ^ in2[116];
    assign G[100] = in[115] & in2[115];
    assign P[100] = in[115] ^ in2[115];
    assign G[101] = in[114] & in2[114];
    assign P[101] = in[114] ^ in2[114];
    assign G[102] = in[113] & in2[113];
    assign P[102] = in[113] ^ in2[113];
    assign G[103] = in[112] & in2[112];
    assign P[103] = in[112] ^ in2[112];
    assign G[104] = in[111] & in2[111];
    assign P[104] = in[111] ^ in2[111];
    assign G[105] = in[110] & in2[110];
    assign P[105] = in[110] ^ in2[110];
    assign G[106] = in[109] & in2[109];
    assign P[106] = in[109] ^ in2[109];
    assign G[107] = in[108] & in2[108];
    assign P[107] = in[108] ^ in2[108];
    assign G[108] = in[107] & in2[107];
    assign P[108] = in[107] ^ in2[107];
    assign G[109] = in[106] & in2[106];
    assign P[109] = in[106] ^ in2[106];
    assign G[110] = in[105] & in2[105];
    assign P[110] = in[105] ^ in2[105];
    assign G[111] = in[104] & in2[104];
    assign P[111] = in[104] ^ in2[104];
    assign G[112] = in[103] & in2[103];
    assign P[112] = in[103] ^ in2[103];
    assign G[113] = in[102] & in2[102];
    assign P[113] = in[102] ^ in2[102];
    assign G[114] = in[101] & in2[101];
    assign P[114] = in[101] ^ in2[101];
    assign G[115] = in[100] & in2[100];
    assign P[115] = in[100] ^ in2[100];
    assign G[116] = in[99] & in2[99];
    assign P[116] = in[99] ^ in2[99];
    assign G[117] = in[98] & in2[98];
    assign P[117] = in[98] ^ in2[98];
    assign G[118] = in[97] & in2[97];
    assign P[118] = in[97] ^ in2[97];
    assign G[119] = in[96] & in2[96];
    assign P[119] = in[96] ^ in2[96];
    assign G[120] = in[95] & in2[95];
    assign P[120] = in[95] ^ in2[95];
    assign G[121] = in[94] & in2[94];
    assign P[121] = in[94] ^ in2[94];
    assign G[122] = in[93] & in2[93];
    assign P[122] = in[93] ^ in2[93];
    assign G[123] = in[92] & in2[92];
    assign P[123] = in[92] ^ in2[92];
    assign G[124] = in[91] & in2[91];
    assign P[124] = in[91] ^ in2[91];
    assign G[125] = in[90] & in2[90];
    assign P[125] = in[90] ^ in2[90];
    assign G[126] = in[89] & in2[89];
    assign P[126] = in[89] ^ in2[89];
    assign G[127] = in[88] & in2[88];
    assign P[127] = in[88] ^ in2[88];
    assign G[128] = in[87] & in2[87];
    assign P[128] = in[87] ^ in2[87];
    assign G[129] = in[86] & in2[86];
    assign P[129] = in[86] ^ in2[86];
    assign G[130] = in[85] & in2[85];
    assign P[130] = in[85] ^ in2[85];
    assign G[131] = in[84] & in2[84];
    assign P[131] = in[84] ^ in2[84];
    assign G[132] = in[83] & in2[83];
    assign P[132] = in[83] ^ in2[83];
    assign G[133] = in[82] & in2[82];
    assign P[133] = in[82] ^ in2[82];
    assign G[134] = in[81] & in2[81];
    assign P[134] = in[81] ^ in2[81];
    assign G[135] = in[80] & in2[80];
    assign P[135] = in[80] ^ in2[80];
    assign G[136] = in[79] & in2[79];
    assign P[136] = in[79] ^ in2[79];
    assign G[137] = in[78] & in2[78];
    assign P[137] = in[78] ^ in2[78];
    assign G[138] = in[77] & in2[77];
    assign P[138] = in[77] ^ in2[77];
    assign G[139] = in[76] & in2[76];
    assign P[139] = in[76] ^ in2[76];
    assign G[140] = in[75] & in2[75];
    assign P[140] = in[75] ^ in2[75];
    assign G[141] = in[74] & in2[74];
    assign P[141] = in[74] ^ in2[74];
    assign G[142] = in[73] & in2[73];
    assign P[142] = in[73] ^ in2[73];
    assign G[143] = in[72] & in2[72];
    assign P[143] = in[72] ^ in2[72];
    assign G[144] = in[71] & in2[71];
    assign P[144] = in[71] ^ in2[71];
    assign G[145] = in[70] & in2[70];
    assign P[145] = in[70] ^ in2[70];
    assign G[146] = in[69] & in2[69];
    assign P[146] = in[69] ^ in2[69];
    assign G[147] = in[68] & in2[68];
    assign P[147] = in[68] ^ in2[68];
    assign G[148] = in[67] & in2[67];
    assign P[148] = in[67] ^ in2[67];
    assign G[149] = in[66] & in2[66];
    assign P[149] = in[66] ^ in2[66];
    assign G[150] = in[65] & in2[65];
    assign P[150] = in[65] ^ in2[65];
    assign G[151] = in[64] & in2[64];
    assign P[151] = in[64] ^ in2[64];
    assign G[152] = in[63] & in2[63];
    assign P[152] = in[63] ^ in2[63];
    assign G[153] = in[62] & in2[62];
    assign P[153] = in[62] ^ in2[62];
    assign G[154] = in[61] & in2[61];
    assign P[154] = in[61] ^ in2[61];
    assign G[155] = in[60] & in2[60];
    assign P[155] = in[60] ^ in2[60];
    assign G[156] = in[59] & in2[59];
    assign P[156] = in[59] ^ in2[59];
    assign G[157] = in[58] & in2[58];
    assign P[157] = in[58] ^ in2[58];
    assign G[158] = in[57] & in2[57];
    assign P[158] = in[57] ^ in2[57];
    assign G[159] = in[56] & in2[56];
    assign P[159] = in[56] ^ in2[56];
    assign G[160] = in[55] & in2[55];
    assign P[160] = in[55] ^ in2[55];
    assign G[161] = in[54] & in2[54];
    assign P[161] = in[54] ^ in2[54];
    assign G[162] = in[53] & in2[53];
    assign P[162] = in[53] ^ in2[53];
    assign G[163] = in[52] & in2[52];
    assign P[163] = in[52] ^ in2[52];
    assign G[164] = in[51] & in2[51];
    assign P[164] = in[51] ^ in2[51];
    assign G[165] = in[50] & in2[50];
    assign P[165] = in[50] ^ in2[50];
    assign G[166] = in[49] & in2[49];
    assign P[166] = in[49] ^ in2[49];
    assign G[167] = in[48] & in2[48];
    assign P[167] = in[48] ^ in2[48];
    assign G[168] = in[47] & in2[47];
    assign P[168] = in[47] ^ in2[47];
    assign G[169] = in[46] & in2[46];
    assign P[169] = in[46] ^ in2[46];
    assign G[170] = in[45] & in2[45];
    assign P[170] = in[45] ^ in2[45];
    assign G[171] = in[44] & in2[44];
    assign P[171] = in[44] ^ in2[44];
    assign G[172] = in[43] & in2[43];
    assign P[172] = in[43] ^ in2[43];
    assign G[173] = in[42] & in2[42];
    assign P[173] = in[42] ^ in2[42];
    assign G[174] = in[41] & in2[41];
    assign P[174] = in[41] ^ in2[41];
    assign G[175] = in[40] & in2[40];
    assign P[175] = in[40] ^ in2[40];
    assign G[176] = in[39] & in2[39];
    assign P[176] = in[39] ^ in2[39];
    assign G[177] = in[38] & in2[38];
    assign P[177] = in[38] ^ in2[38];
    assign G[178] = in[37] & in2[37];
    assign P[178] = in[37] ^ in2[37];
    assign G[179] = in[36] & in2[36];
    assign P[179] = in[36] ^ in2[36];
    assign G[180] = in[35] & in2[35];
    assign P[180] = in[35] ^ in2[35];
    assign G[181] = in[34] & in2[34];
    assign P[181] = in[34] ^ in2[34];
    assign G[182] = in[33] & in2[33];
    assign P[182] = in[33] ^ in2[33];
    assign G[183] = in[32] & in2[32];
    assign P[183] = in[32] ^ in2[32];
    assign G[184] = in[31] & in2[31];
    assign P[184] = in[31] ^ in2[31];
    assign G[185] = in[30] & in2[30];
    assign P[185] = in[30] ^ in2[30];
    assign G[186] = in[29] & in2[29];
    assign P[186] = in[29] ^ in2[29];
    assign G[187] = in[28] & in2[28];
    assign P[187] = in[28] ^ in2[28];
    assign G[188] = in[27] & in2[27];
    assign P[188] = in[27] ^ in2[27];
    assign G[189] = in[26] & in2[26];
    assign P[189] = in[26] ^ in2[26];
    assign G[190] = in[25] & in2[25];
    assign P[190] = in[25] ^ in2[25];
    assign G[191] = in[24] & in2[24];
    assign P[191] = in[24] ^ in2[24];
    assign G[192] = in[23] & in2[23];
    assign P[192] = in[23] ^ in2[23];
    assign G[193] = in[22] & in2[22];
    assign P[193] = in[22] ^ in2[22];
    assign G[194] = in[21] & in2[21];
    assign P[194] = in[21] ^ in2[21];
    assign G[195] = in[20] & in2[20];
    assign P[195] = in[20] ^ in2[20];
    assign G[196] = in[19] & in2[19];
    assign P[196] = in[19] ^ in2[19];
    assign G[197] = in[18] & in2[18];
    assign P[197] = in[18] ^ in2[18];
    assign G[198] = in[17] & in2[17];
    assign P[198] = in[17] ^ in2[17];
    assign G[199] = in[16] & in2[16];
    assign P[199] = in[16] ^ in2[16];
    assign G[200] = in[15] & in2[15];
    assign P[200] = in[15] ^ in2[15];
    assign G[201] = in[14] & in2[14];
    assign P[201] = in[14] ^ in2[14];
    assign G[202] = in[13] & in2[13];
    assign P[202] = in[13] ^ in2[13];
    assign G[203] = in[12] & in2[12];
    assign P[203] = in[12] ^ in2[12];
    assign G[204] = in[11] & in2[11];
    assign P[204] = in[11] ^ in2[11];
    assign G[205] = in[10] & in2[10];
    assign P[205] = in[10] ^ in2[10];
    assign G[206] = in[9] & in2[9];
    assign P[206] = in[9] ^ in2[9];
    assign G[207] = in[8] & in2[8];
    assign P[207] = in[8] ^ in2[8];
    assign G[208] = in[7] & in2[7];
    assign P[208] = in[7] ^ in2[7];
    assign G[209] = in[6] & in2[6];
    assign P[209] = in[6] ^ in2[6];
    assign G[210] = in[5] & in2[5];
    assign P[210] = in[5] ^ in2[5];
    assign G[211] = in[4] & in2[4];
    assign P[211] = in[4] ^ in2[4];
    assign G[212] = in[3] & in2[3];
    assign P[212] = in[3] ^ in2[3];
    assign G[213] = in[2] & in2[2];
    assign P[213] = in[2] ^ in2[2];
    assign G[214] = in[1] & in2[1];
    assign P[214] = in[1] ^ in2[1];
    assign G[215] = in[0] & in2[0];
    assign P[215] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign C[215] = G[214] | (P[214] & C[214]);
    assign cout = G[215] | (P[215] & C[215]);
    assign sum = P ^ C;
endmodule

module CLA215(output [214:0] sum, output cout, input [214:0] in1, input [214:0] in2;

    wire[214:0] G;
    wire[214:0] C;
    wire[214:0] P;

    assign G[0] = in[214] & in2[214];
    assign P[0] = in[214] ^ in2[214];
    assign G[1] = in[213] & in2[213];
    assign P[1] = in[213] ^ in2[213];
    assign G[2] = in[212] & in2[212];
    assign P[2] = in[212] ^ in2[212];
    assign G[3] = in[211] & in2[211];
    assign P[3] = in[211] ^ in2[211];
    assign G[4] = in[210] & in2[210];
    assign P[4] = in[210] ^ in2[210];
    assign G[5] = in[209] & in2[209];
    assign P[5] = in[209] ^ in2[209];
    assign G[6] = in[208] & in2[208];
    assign P[6] = in[208] ^ in2[208];
    assign G[7] = in[207] & in2[207];
    assign P[7] = in[207] ^ in2[207];
    assign G[8] = in[206] & in2[206];
    assign P[8] = in[206] ^ in2[206];
    assign G[9] = in[205] & in2[205];
    assign P[9] = in[205] ^ in2[205];
    assign G[10] = in[204] & in2[204];
    assign P[10] = in[204] ^ in2[204];
    assign G[11] = in[203] & in2[203];
    assign P[11] = in[203] ^ in2[203];
    assign G[12] = in[202] & in2[202];
    assign P[12] = in[202] ^ in2[202];
    assign G[13] = in[201] & in2[201];
    assign P[13] = in[201] ^ in2[201];
    assign G[14] = in[200] & in2[200];
    assign P[14] = in[200] ^ in2[200];
    assign G[15] = in[199] & in2[199];
    assign P[15] = in[199] ^ in2[199];
    assign G[16] = in[198] & in2[198];
    assign P[16] = in[198] ^ in2[198];
    assign G[17] = in[197] & in2[197];
    assign P[17] = in[197] ^ in2[197];
    assign G[18] = in[196] & in2[196];
    assign P[18] = in[196] ^ in2[196];
    assign G[19] = in[195] & in2[195];
    assign P[19] = in[195] ^ in2[195];
    assign G[20] = in[194] & in2[194];
    assign P[20] = in[194] ^ in2[194];
    assign G[21] = in[193] & in2[193];
    assign P[21] = in[193] ^ in2[193];
    assign G[22] = in[192] & in2[192];
    assign P[22] = in[192] ^ in2[192];
    assign G[23] = in[191] & in2[191];
    assign P[23] = in[191] ^ in2[191];
    assign G[24] = in[190] & in2[190];
    assign P[24] = in[190] ^ in2[190];
    assign G[25] = in[189] & in2[189];
    assign P[25] = in[189] ^ in2[189];
    assign G[26] = in[188] & in2[188];
    assign P[26] = in[188] ^ in2[188];
    assign G[27] = in[187] & in2[187];
    assign P[27] = in[187] ^ in2[187];
    assign G[28] = in[186] & in2[186];
    assign P[28] = in[186] ^ in2[186];
    assign G[29] = in[185] & in2[185];
    assign P[29] = in[185] ^ in2[185];
    assign G[30] = in[184] & in2[184];
    assign P[30] = in[184] ^ in2[184];
    assign G[31] = in[183] & in2[183];
    assign P[31] = in[183] ^ in2[183];
    assign G[32] = in[182] & in2[182];
    assign P[32] = in[182] ^ in2[182];
    assign G[33] = in[181] & in2[181];
    assign P[33] = in[181] ^ in2[181];
    assign G[34] = in[180] & in2[180];
    assign P[34] = in[180] ^ in2[180];
    assign G[35] = in[179] & in2[179];
    assign P[35] = in[179] ^ in2[179];
    assign G[36] = in[178] & in2[178];
    assign P[36] = in[178] ^ in2[178];
    assign G[37] = in[177] & in2[177];
    assign P[37] = in[177] ^ in2[177];
    assign G[38] = in[176] & in2[176];
    assign P[38] = in[176] ^ in2[176];
    assign G[39] = in[175] & in2[175];
    assign P[39] = in[175] ^ in2[175];
    assign G[40] = in[174] & in2[174];
    assign P[40] = in[174] ^ in2[174];
    assign G[41] = in[173] & in2[173];
    assign P[41] = in[173] ^ in2[173];
    assign G[42] = in[172] & in2[172];
    assign P[42] = in[172] ^ in2[172];
    assign G[43] = in[171] & in2[171];
    assign P[43] = in[171] ^ in2[171];
    assign G[44] = in[170] & in2[170];
    assign P[44] = in[170] ^ in2[170];
    assign G[45] = in[169] & in2[169];
    assign P[45] = in[169] ^ in2[169];
    assign G[46] = in[168] & in2[168];
    assign P[46] = in[168] ^ in2[168];
    assign G[47] = in[167] & in2[167];
    assign P[47] = in[167] ^ in2[167];
    assign G[48] = in[166] & in2[166];
    assign P[48] = in[166] ^ in2[166];
    assign G[49] = in[165] & in2[165];
    assign P[49] = in[165] ^ in2[165];
    assign G[50] = in[164] & in2[164];
    assign P[50] = in[164] ^ in2[164];
    assign G[51] = in[163] & in2[163];
    assign P[51] = in[163] ^ in2[163];
    assign G[52] = in[162] & in2[162];
    assign P[52] = in[162] ^ in2[162];
    assign G[53] = in[161] & in2[161];
    assign P[53] = in[161] ^ in2[161];
    assign G[54] = in[160] & in2[160];
    assign P[54] = in[160] ^ in2[160];
    assign G[55] = in[159] & in2[159];
    assign P[55] = in[159] ^ in2[159];
    assign G[56] = in[158] & in2[158];
    assign P[56] = in[158] ^ in2[158];
    assign G[57] = in[157] & in2[157];
    assign P[57] = in[157] ^ in2[157];
    assign G[58] = in[156] & in2[156];
    assign P[58] = in[156] ^ in2[156];
    assign G[59] = in[155] & in2[155];
    assign P[59] = in[155] ^ in2[155];
    assign G[60] = in[154] & in2[154];
    assign P[60] = in[154] ^ in2[154];
    assign G[61] = in[153] & in2[153];
    assign P[61] = in[153] ^ in2[153];
    assign G[62] = in[152] & in2[152];
    assign P[62] = in[152] ^ in2[152];
    assign G[63] = in[151] & in2[151];
    assign P[63] = in[151] ^ in2[151];
    assign G[64] = in[150] & in2[150];
    assign P[64] = in[150] ^ in2[150];
    assign G[65] = in[149] & in2[149];
    assign P[65] = in[149] ^ in2[149];
    assign G[66] = in[148] & in2[148];
    assign P[66] = in[148] ^ in2[148];
    assign G[67] = in[147] & in2[147];
    assign P[67] = in[147] ^ in2[147];
    assign G[68] = in[146] & in2[146];
    assign P[68] = in[146] ^ in2[146];
    assign G[69] = in[145] & in2[145];
    assign P[69] = in[145] ^ in2[145];
    assign G[70] = in[144] & in2[144];
    assign P[70] = in[144] ^ in2[144];
    assign G[71] = in[143] & in2[143];
    assign P[71] = in[143] ^ in2[143];
    assign G[72] = in[142] & in2[142];
    assign P[72] = in[142] ^ in2[142];
    assign G[73] = in[141] & in2[141];
    assign P[73] = in[141] ^ in2[141];
    assign G[74] = in[140] & in2[140];
    assign P[74] = in[140] ^ in2[140];
    assign G[75] = in[139] & in2[139];
    assign P[75] = in[139] ^ in2[139];
    assign G[76] = in[138] & in2[138];
    assign P[76] = in[138] ^ in2[138];
    assign G[77] = in[137] & in2[137];
    assign P[77] = in[137] ^ in2[137];
    assign G[78] = in[136] & in2[136];
    assign P[78] = in[136] ^ in2[136];
    assign G[79] = in[135] & in2[135];
    assign P[79] = in[135] ^ in2[135];
    assign G[80] = in[134] & in2[134];
    assign P[80] = in[134] ^ in2[134];
    assign G[81] = in[133] & in2[133];
    assign P[81] = in[133] ^ in2[133];
    assign G[82] = in[132] & in2[132];
    assign P[82] = in[132] ^ in2[132];
    assign G[83] = in[131] & in2[131];
    assign P[83] = in[131] ^ in2[131];
    assign G[84] = in[130] & in2[130];
    assign P[84] = in[130] ^ in2[130];
    assign G[85] = in[129] & in2[129];
    assign P[85] = in[129] ^ in2[129];
    assign G[86] = in[128] & in2[128];
    assign P[86] = in[128] ^ in2[128];
    assign G[87] = in[127] & in2[127];
    assign P[87] = in[127] ^ in2[127];
    assign G[88] = in[126] & in2[126];
    assign P[88] = in[126] ^ in2[126];
    assign G[89] = in[125] & in2[125];
    assign P[89] = in[125] ^ in2[125];
    assign G[90] = in[124] & in2[124];
    assign P[90] = in[124] ^ in2[124];
    assign G[91] = in[123] & in2[123];
    assign P[91] = in[123] ^ in2[123];
    assign G[92] = in[122] & in2[122];
    assign P[92] = in[122] ^ in2[122];
    assign G[93] = in[121] & in2[121];
    assign P[93] = in[121] ^ in2[121];
    assign G[94] = in[120] & in2[120];
    assign P[94] = in[120] ^ in2[120];
    assign G[95] = in[119] & in2[119];
    assign P[95] = in[119] ^ in2[119];
    assign G[96] = in[118] & in2[118];
    assign P[96] = in[118] ^ in2[118];
    assign G[97] = in[117] & in2[117];
    assign P[97] = in[117] ^ in2[117];
    assign G[98] = in[116] & in2[116];
    assign P[98] = in[116] ^ in2[116];
    assign G[99] = in[115] & in2[115];
    assign P[99] = in[115] ^ in2[115];
    assign G[100] = in[114] & in2[114];
    assign P[100] = in[114] ^ in2[114];
    assign G[101] = in[113] & in2[113];
    assign P[101] = in[113] ^ in2[113];
    assign G[102] = in[112] & in2[112];
    assign P[102] = in[112] ^ in2[112];
    assign G[103] = in[111] & in2[111];
    assign P[103] = in[111] ^ in2[111];
    assign G[104] = in[110] & in2[110];
    assign P[104] = in[110] ^ in2[110];
    assign G[105] = in[109] & in2[109];
    assign P[105] = in[109] ^ in2[109];
    assign G[106] = in[108] & in2[108];
    assign P[106] = in[108] ^ in2[108];
    assign G[107] = in[107] & in2[107];
    assign P[107] = in[107] ^ in2[107];
    assign G[108] = in[106] & in2[106];
    assign P[108] = in[106] ^ in2[106];
    assign G[109] = in[105] & in2[105];
    assign P[109] = in[105] ^ in2[105];
    assign G[110] = in[104] & in2[104];
    assign P[110] = in[104] ^ in2[104];
    assign G[111] = in[103] & in2[103];
    assign P[111] = in[103] ^ in2[103];
    assign G[112] = in[102] & in2[102];
    assign P[112] = in[102] ^ in2[102];
    assign G[113] = in[101] & in2[101];
    assign P[113] = in[101] ^ in2[101];
    assign G[114] = in[100] & in2[100];
    assign P[114] = in[100] ^ in2[100];
    assign G[115] = in[99] & in2[99];
    assign P[115] = in[99] ^ in2[99];
    assign G[116] = in[98] & in2[98];
    assign P[116] = in[98] ^ in2[98];
    assign G[117] = in[97] & in2[97];
    assign P[117] = in[97] ^ in2[97];
    assign G[118] = in[96] & in2[96];
    assign P[118] = in[96] ^ in2[96];
    assign G[119] = in[95] & in2[95];
    assign P[119] = in[95] ^ in2[95];
    assign G[120] = in[94] & in2[94];
    assign P[120] = in[94] ^ in2[94];
    assign G[121] = in[93] & in2[93];
    assign P[121] = in[93] ^ in2[93];
    assign G[122] = in[92] & in2[92];
    assign P[122] = in[92] ^ in2[92];
    assign G[123] = in[91] & in2[91];
    assign P[123] = in[91] ^ in2[91];
    assign G[124] = in[90] & in2[90];
    assign P[124] = in[90] ^ in2[90];
    assign G[125] = in[89] & in2[89];
    assign P[125] = in[89] ^ in2[89];
    assign G[126] = in[88] & in2[88];
    assign P[126] = in[88] ^ in2[88];
    assign G[127] = in[87] & in2[87];
    assign P[127] = in[87] ^ in2[87];
    assign G[128] = in[86] & in2[86];
    assign P[128] = in[86] ^ in2[86];
    assign G[129] = in[85] & in2[85];
    assign P[129] = in[85] ^ in2[85];
    assign G[130] = in[84] & in2[84];
    assign P[130] = in[84] ^ in2[84];
    assign G[131] = in[83] & in2[83];
    assign P[131] = in[83] ^ in2[83];
    assign G[132] = in[82] & in2[82];
    assign P[132] = in[82] ^ in2[82];
    assign G[133] = in[81] & in2[81];
    assign P[133] = in[81] ^ in2[81];
    assign G[134] = in[80] & in2[80];
    assign P[134] = in[80] ^ in2[80];
    assign G[135] = in[79] & in2[79];
    assign P[135] = in[79] ^ in2[79];
    assign G[136] = in[78] & in2[78];
    assign P[136] = in[78] ^ in2[78];
    assign G[137] = in[77] & in2[77];
    assign P[137] = in[77] ^ in2[77];
    assign G[138] = in[76] & in2[76];
    assign P[138] = in[76] ^ in2[76];
    assign G[139] = in[75] & in2[75];
    assign P[139] = in[75] ^ in2[75];
    assign G[140] = in[74] & in2[74];
    assign P[140] = in[74] ^ in2[74];
    assign G[141] = in[73] & in2[73];
    assign P[141] = in[73] ^ in2[73];
    assign G[142] = in[72] & in2[72];
    assign P[142] = in[72] ^ in2[72];
    assign G[143] = in[71] & in2[71];
    assign P[143] = in[71] ^ in2[71];
    assign G[144] = in[70] & in2[70];
    assign P[144] = in[70] ^ in2[70];
    assign G[145] = in[69] & in2[69];
    assign P[145] = in[69] ^ in2[69];
    assign G[146] = in[68] & in2[68];
    assign P[146] = in[68] ^ in2[68];
    assign G[147] = in[67] & in2[67];
    assign P[147] = in[67] ^ in2[67];
    assign G[148] = in[66] & in2[66];
    assign P[148] = in[66] ^ in2[66];
    assign G[149] = in[65] & in2[65];
    assign P[149] = in[65] ^ in2[65];
    assign G[150] = in[64] & in2[64];
    assign P[150] = in[64] ^ in2[64];
    assign G[151] = in[63] & in2[63];
    assign P[151] = in[63] ^ in2[63];
    assign G[152] = in[62] & in2[62];
    assign P[152] = in[62] ^ in2[62];
    assign G[153] = in[61] & in2[61];
    assign P[153] = in[61] ^ in2[61];
    assign G[154] = in[60] & in2[60];
    assign P[154] = in[60] ^ in2[60];
    assign G[155] = in[59] & in2[59];
    assign P[155] = in[59] ^ in2[59];
    assign G[156] = in[58] & in2[58];
    assign P[156] = in[58] ^ in2[58];
    assign G[157] = in[57] & in2[57];
    assign P[157] = in[57] ^ in2[57];
    assign G[158] = in[56] & in2[56];
    assign P[158] = in[56] ^ in2[56];
    assign G[159] = in[55] & in2[55];
    assign P[159] = in[55] ^ in2[55];
    assign G[160] = in[54] & in2[54];
    assign P[160] = in[54] ^ in2[54];
    assign G[161] = in[53] & in2[53];
    assign P[161] = in[53] ^ in2[53];
    assign G[162] = in[52] & in2[52];
    assign P[162] = in[52] ^ in2[52];
    assign G[163] = in[51] & in2[51];
    assign P[163] = in[51] ^ in2[51];
    assign G[164] = in[50] & in2[50];
    assign P[164] = in[50] ^ in2[50];
    assign G[165] = in[49] & in2[49];
    assign P[165] = in[49] ^ in2[49];
    assign G[166] = in[48] & in2[48];
    assign P[166] = in[48] ^ in2[48];
    assign G[167] = in[47] & in2[47];
    assign P[167] = in[47] ^ in2[47];
    assign G[168] = in[46] & in2[46];
    assign P[168] = in[46] ^ in2[46];
    assign G[169] = in[45] & in2[45];
    assign P[169] = in[45] ^ in2[45];
    assign G[170] = in[44] & in2[44];
    assign P[170] = in[44] ^ in2[44];
    assign G[171] = in[43] & in2[43];
    assign P[171] = in[43] ^ in2[43];
    assign G[172] = in[42] & in2[42];
    assign P[172] = in[42] ^ in2[42];
    assign G[173] = in[41] & in2[41];
    assign P[173] = in[41] ^ in2[41];
    assign G[174] = in[40] & in2[40];
    assign P[174] = in[40] ^ in2[40];
    assign G[175] = in[39] & in2[39];
    assign P[175] = in[39] ^ in2[39];
    assign G[176] = in[38] & in2[38];
    assign P[176] = in[38] ^ in2[38];
    assign G[177] = in[37] & in2[37];
    assign P[177] = in[37] ^ in2[37];
    assign G[178] = in[36] & in2[36];
    assign P[178] = in[36] ^ in2[36];
    assign G[179] = in[35] & in2[35];
    assign P[179] = in[35] ^ in2[35];
    assign G[180] = in[34] & in2[34];
    assign P[180] = in[34] ^ in2[34];
    assign G[181] = in[33] & in2[33];
    assign P[181] = in[33] ^ in2[33];
    assign G[182] = in[32] & in2[32];
    assign P[182] = in[32] ^ in2[32];
    assign G[183] = in[31] & in2[31];
    assign P[183] = in[31] ^ in2[31];
    assign G[184] = in[30] & in2[30];
    assign P[184] = in[30] ^ in2[30];
    assign G[185] = in[29] & in2[29];
    assign P[185] = in[29] ^ in2[29];
    assign G[186] = in[28] & in2[28];
    assign P[186] = in[28] ^ in2[28];
    assign G[187] = in[27] & in2[27];
    assign P[187] = in[27] ^ in2[27];
    assign G[188] = in[26] & in2[26];
    assign P[188] = in[26] ^ in2[26];
    assign G[189] = in[25] & in2[25];
    assign P[189] = in[25] ^ in2[25];
    assign G[190] = in[24] & in2[24];
    assign P[190] = in[24] ^ in2[24];
    assign G[191] = in[23] & in2[23];
    assign P[191] = in[23] ^ in2[23];
    assign G[192] = in[22] & in2[22];
    assign P[192] = in[22] ^ in2[22];
    assign G[193] = in[21] & in2[21];
    assign P[193] = in[21] ^ in2[21];
    assign G[194] = in[20] & in2[20];
    assign P[194] = in[20] ^ in2[20];
    assign G[195] = in[19] & in2[19];
    assign P[195] = in[19] ^ in2[19];
    assign G[196] = in[18] & in2[18];
    assign P[196] = in[18] ^ in2[18];
    assign G[197] = in[17] & in2[17];
    assign P[197] = in[17] ^ in2[17];
    assign G[198] = in[16] & in2[16];
    assign P[198] = in[16] ^ in2[16];
    assign G[199] = in[15] & in2[15];
    assign P[199] = in[15] ^ in2[15];
    assign G[200] = in[14] & in2[14];
    assign P[200] = in[14] ^ in2[14];
    assign G[201] = in[13] & in2[13];
    assign P[201] = in[13] ^ in2[13];
    assign G[202] = in[12] & in2[12];
    assign P[202] = in[12] ^ in2[12];
    assign G[203] = in[11] & in2[11];
    assign P[203] = in[11] ^ in2[11];
    assign G[204] = in[10] & in2[10];
    assign P[204] = in[10] ^ in2[10];
    assign G[205] = in[9] & in2[9];
    assign P[205] = in[9] ^ in2[9];
    assign G[206] = in[8] & in2[8];
    assign P[206] = in[8] ^ in2[8];
    assign G[207] = in[7] & in2[7];
    assign P[207] = in[7] ^ in2[7];
    assign G[208] = in[6] & in2[6];
    assign P[208] = in[6] ^ in2[6];
    assign G[209] = in[5] & in2[5];
    assign P[209] = in[5] ^ in2[5];
    assign G[210] = in[4] & in2[4];
    assign P[210] = in[4] ^ in2[4];
    assign G[211] = in[3] & in2[3];
    assign P[211] = in[3] ^ in2[3];
    assign G[212] = in[2] & in2[2];
    assign P[212] = in[2] ^ in2[2];
    assign G[213] = in[1] & in2[1];
    assign P[213] = in[1] ^ in2[1];
    assign G[214] = in[0] & in2[0];
    assign P[214] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign C[214] = G[213] | (P[213] & C[213]);
    assign cout = G[214] | (P[214] & C[214]);
    assign sum = P ^ C;
endmodule

module CLA214(output [213:0] sum, output cout, input [213:0] in1, input [213:0] in2;

    wire[213:0] G;
    wire[213:0] C;
    wire[213:0] P;

    assign G[0] = in[213] & in2[213];
    assign P[0] = in[213] ^ in2[213];
    assign G[1] = in[212] & in2[212];
    assign P[1] = in[212] ^ in2[212];
    assign G[2] = in[211] & in2[211];
    assign P[2] = in[211] ^ in2[211];
    assign G[3] = in[210] & in2[210];
    assign P[3] = in[210] ^ in2[210];
    assign G[4] = in[209] & in2[209];
    assign P[4] = in[209] ^ in2[209];
    assign G[5] = in[208] & in2[208];
    assign P[5] = in[208] ^ in2[208];
    assign G[6] = in[207] & in2[207];
    assign P[6] = in[207] ^ in2[207];
    assign G[7] = in[206] & in2[206];
    assign P[7] = in[206] ^ in2[206];
    assign G[8] = in[205] & in2[205];
    assign P[8] = in[205] ^ in2[205];
    assign G[9] = in[204] & in2[204];
    assign P[9] = in[204] ^ in2[204];
    assign G[10] = in[203] & in2[203];
    assign P[10] = in[203] ^ in2[203];
    assign G[11] = in[202] & in2[202];
    assign P[11] = in[202] ^ in2[202];
    assign G[12] = in[201] & in2[201];
    assign P[12] = in[201] ^ in2[201];
    assign G[13] = in[200] & in2[200];
    assign P[13] = in[200] ^ in2[200];
    assign G[14] = in[199] & in2[199];
    assign P[14] = in[199] ^ in2[199];
    assign G[15] = in[198] & in2[198];
    assign P[15] = in[198] ^ in2[198];
    assign G[16] = in[197] & in2[197];
    assign P[16] = in[197] ^ in2[197];
    assign G[17] = in[196] & in2[196];
    assign P[17] = in[196] ^ in2[196];
    assign G[18] = in[195] & in2[195];
    assign P[18] = in[195] ^ in2[195];
    assign G[19] = in[194] & in2[194];
    assign P[19] = in[194] ^ in2[194];
    assign G[20] = in[193] & in2[193];
    assign P[20] = in[193] ^ in2[193];
    assign G[21] = in[192] & in2[192];
    assign P[21] = in[192] ^ in2[192];
    assign G[22] = in[191] & in2[191];
    assign P[22] = in[191] ^ in2[191];
    assign G[23] = in[190] & in2[190];
    assign P[23] = in[190] ^ in2[190];
    assign G[24] = in[189] & in2[189];
    assign P[24] = in[189] ^ in2[189];
    assign G[25] = in[188] & in2[188];
    assign P[25] = in[188] ^ in2[188];
    assign G[26] = in[187] & in2[187];
    assign P[26] = in[187] ^ in2[187];
    assign G[27] = in[186] & in2[186];
    assign P[27] = in[186] ^ in2[186];
    assign G[28] = in[185] & in2[185];
    assign P[28] = in[185] ^ in2[185];
    assign G[29] = in[184] & in2[184];
    assign P[29] = in[184] ^ in2[184];
    assign G[30] = in[183] & in2[183];
    assign P[30] = in[183] ^ in2[183];
    assign G[31] = in[182] & in2[182];
    assign P[31] = in[182] ^ in2[182];
    assign G[32] = in[181] & in2[181];
    assign P[32] = in[181] ^ in2[181];
    assign G[33] = in[180] & in2[180];
    assign P[33] = in[180] ^ in2[180];
    assign G[34] = in[179] & in2[179];
    assign P[34] = in[179] ^ in2[179];
    assign G[35] = in[178] & in2[178];
    assign P[35] = in[178] ^ in2[178];
    assign G[36] = in[177] & in2[177];
    assign P[36] = in[177] ^ in2[177];
    assign G[37] = in[176] & in2[176];
    assign P[37] = in[176] ^ in2[176];
    assign G[38] = in[175] & in2[175];
    assign P[38] = in[175] ^ in2[175];
    assign G[39] = in[174] & in2[174];
    assign P[39] = in[174] ^ in2[174];
    assign G[40] = in[173] & in2[173];
    assign P[40] = in[173] ^ in2[173];
    assign G[41] = in[172] & in2[172];
    assign P[41] = in[172] ^ in2[172];
    assign G[42] = in[171] & in2[171];
    assign P[42] = in[171] ^ in2[171];
    assign G[43] = in[170] & in2[170];
    assign P[43] = in[170] ^ in2[170];
    assign G[44] = in[169] & in2[169];
    assign P[44] = in[169] ^ in2[169];
    assign G[45] = in[168] & in2[168];
    assign P[45] = in[168] ^ in2[168];
    assign G[46] = in[167] & in2[167];
    assign P[46] = in[167] ^ in2[167];
    assign G[47] = in[166] & in2[166];
    assign P[47] = in[166] ^ in2[166];
    assign G[48] = in[165] & in2[165];
    assign P[48] = in[165] ^ in2[165];
    assign G[49] = in[164] & in2[164];
    assign P[49] = in[164] ^ in2[164];
    assign G[50] = in[163] & in2[163];
    assign P[50] = in[163] ^ in2[163];
    assign G[51] = in[162] & in2[162];
    assign P[51] = in[162] ^ in2[162];
    assign G[52] = in[161] & in2[161];
    assign P[52] = in[161] ^ in2[161];
    assign G[53] = in[160] & in2[160];
    assign P[53] = in[160] ^ in2[160];
    assign G[54] = in[159] & in2[159];
    assign P[54] = in[159] ^ in2[159];
    assign G[55] = in[158] & in2[158];
    assign P[55] = in[158] ^ in2[158];
    assign G[56] = in[157] & in2[157];
    assign P[56] = in[157] ^ in2[157];
    assign G[57] = in[156] & in2[156];
    assign P[57] = in[156] ^ in2[156];
    assign G[58] = in[155] & in2[155];
    assign P[58] = in[155] ^ in2[155];
    assign G[59] = in[154] & in2[154];
    assign P[59] = in[154] ^ in2[154];
    assign G[60] = in[153] & in2[153];
    assign P[60] = in[153] ^ in2[153];
    assign G[61] = in[152] & in2[152];
    assign P[61] = in[152] ^ in2[152];
    assign G[62] = in[151] & in2[151];
    assign P[62] = in[151] ^ in2[151];
    assign G[63] = in[150] & in2[150];
    assign P[63] = in[150] ^ in2[150];
    assign G[64] = in[149] & in2[149];
    assign P[64] = in[149] ^ in2[149];
    assign G[65] = in[148] & in2[148];
    assign P[65] = in[148] ^ in2[148];
    assign G[66] = in[147] & in2[147];
    assign P[66] = in[147] ^ in2[147];
    assign G[67] = in[146] & in2[146];
    assign P[67] = in[146] ^ in2[146];
    assign G[68] = in[145] & in2[145];
    assign P[68] = in[145] ^ in2[145];
    assign G[69] = in[144] & in2[144];
    assign P[69] = in[144] ^ in2[144];
    assign G[70] = in[143] & in2[143];
    assign P[70] = in[143] ^ in2[143];
    assign G[71] = in[142] & in2[142];
    assign P[71] = in[142] ^ in2[142];
    assign G[72] = in[141] & in2[141];
    assign P[72] = in[141] ^ in2[141];
    assign G[73] = in[140] & in2[140];
    assign P[73] = in[140] ^ in2[140];
    assign G[74] = in[139] & in2[139];
    assign P[74] = in[139] ^ in2[139];
    assign G[75] = in[138] & in2[138];
    assign P[75] = in[138] ^ in2[138];
    assign G[76] = in[137] & in2[137];
    assign P[76] = in[137] ^ in2[137];
    assign G[77] = in[136] & in2[136];
    assign P[77] = in[136] ^ in2[136];
    assign G[78] = in[135] & in2[135];
    assign P[78] = in[135] ^ in2[135];
    assign G[79] = in[134] & in2[134];
    assign P[79] = in[134] ^ in2[134];
    assign G[80] = in[133] & in2[133];
    assign P[80] = in[133] ^ in2[133];
    assign G[81] = in[132] & in2[132];
    assign P[81] = in[132] ^ in2[132];
    assign G[82] = in[131] & in2[131];
    assign P[82] = in[131] ^ in2[131];
    assign G[83] = in[130] & in2[130];
    assign P[83] = in[130] ^ in2[130];
    assign G[84] = in[129] & in2[129];
    assign P[84] = in[129] ^ in2[129];
    assign G[85] = in[128] & in2[128];
    assign P[85] = in[128] ^ in2[128];
    assign G[86] = in[127] & in2[127];
    assign P[86] = in[127] ^ in2[127];
    assign G[87] = in[126] & in2[126];
    assign P[87] = in[126] ^ in2[126];
    assign G[88] = in[125] & in2[125];
    assign P[88] = in[125] ^ in2[125];
    assign G[89] = in[124] & in2[124];
    assign P[89] = in[124] ^ in2[124];
    assign G[90] = in[123] & in2[123];
    assign P[90] = in[123] ^ in2[123];
    assign G[91] = in[122] & in2[122];
    assign P[91] = in[122] ^ in2[122];
    assign G[92] = in[121] & in2[121];
    assign P[92] = in[121] ^ in2[121];
    assign G[93] = in[120] & in2[120];
    assign P[93] = in[120] ^ in2[120];
    assign G[94] = in[119] & in2[119];
    assign P[94] = in[119] ^ in2[119];
    assign G[95] = in[118] & in2[118];
    assign P[95] = in[118] ^ in2[118];
    assign G[96] = in[117] & in2[117];
    assign P[96] = in[117] ^ in2[117];
    assign G[97] = in[116] & in2[116];
    assign P[97] = in[116] ^ in2[116];
    assign G[98] = in[115] & in2[115];
    assign P[98] = in[115] ^ in2[115];
    assign G[99] = in[114] & in2[114];
    assign P[99] = in[114] ^ in2[114];
    assign G[100] = in[113] & in2[113];
    assign P[100] = in[113] ^ in2[113];
    assign G[101] = in[112] & in2[112];
    assign P[101] = in[112] ^ in2[112];
    assign G[102] = in[111] & in2[111];
    assign P[102] = in[111] ^ in2[111];
    assign G[103] = in[110] & in2[110];
    assign P[103] = in[110] ^ in2[110];
    assign G[104] = in[109] & in2[109];
    assign P[104] = in[109] ^ in2[109];
    assign G[105] = in[108] & in2[108];
    assign P[105] = in[108] ^ in2[108];
    assign G[106] = in[107] & in2[107];
    assign P[106] = in[107] ^ in2[107];
    assign G[107] = in[106] & in2[106];
    assign P[107] = in[106] ^ in2[106];
    assign G[108] = in[105] & in2[105];
    assign P[108] = in[105] ^ in2[105];
    assign G[109] = in[104] & in2[104];
    assign P[109] = in[104] ^ in2[104];
    assign G[110] = in[103] & in2[103];
    assign P[110] = in[103] ^ in2[103];
    assign G[111] = in[102] & in2[102];
    assign P[111] = in[102] ^ in2[102];
    assign G[112] = in[101] & in2[101];
    assign P[112] = in[101] ^ in2[101];
    assign G[113] = in[100] & in2[100];
    assign P[113] = in[100] ^ in2[100];
    assign G[114] = in[99] & in2[99];
    assign P[114] = in[99] ^ in2[99];
    assign G[115] = in[98] & in2[98];
    assign P[115] = in[98] ^ in2[98];
    assign G[116] = in[97] & in2[97];
    assign P[116] = in[97] ^ in2[97];
    assign G[117] = in[96] & in2[96];
    assign P[117] = in[96] ^ in2[96];
    assign G[118] = in[95] & in2[95];
    assign P[118] = in[95] ^ in2[95];
    assign G[119] = in[94] & in2[94];
    assign P[119] = in[94] ^ in2[94];
    assign G[120] = in[93] & in2[93];
    assign P[120] = in[93] ^ in2[93];
    assign G[121] = in[92] & in2[92];
    assign P[121] = in[92] ^ in2[92];
    assign G[122] = in[91] & in2[91];
    assign P[122] = in[91] ^ in2[91];
    assign G[123] = in[90] & in2[90];
    assign P[123] = in[90] ^ in2[90];
    assign G[124] = in[89] & in2[89];
    assign P[124] = in[89] ^ in2[89];
    assign G[125] = in[88] & in2[88];
    assign P[125] = in[88] ^ in2[88];
    assign G[126] = in[87] & in2[87];
    assign P[126] = in[87] ^ in2[87];
    assign G[127] = in[86] & in2[86];
    assign P[127] = in[86] ^ in2[86];
    assign G[128] = in[85] & in2[85];
    assign P[128] = in[85] ^ in2[85];
    assign G[129] = in[84] & in2[84];
    assign P[129] = in[84] ^ in2[84];
    assign G[130] = in[83] & in2[83];
    assign P[130] = in[83] ^ in2[83];
    assign G[131] = in[82] & in2[82];
    assign P[131] = in[82] ^ in2[82];
    assign G[132] = in[81] & in2[81];
    assign P[132] = in[81] ^ in2[81];
    assign G[133] = in[80] & in2[80];
    assign P[133] = in[80] ^ in2[80];
    assign G[134] = in[79] & in2[79];
    assign P[134] = in[79] ^ in2[79];
    assign G[135] = in[78] & in2[78];
    assign P[135] = in[78] ^ in2[78];
    assign G[136] = in[77] & in2[77];
    assign P[136] = in[77] ^ in2[77];
    assign G[137] = in[76] & in2[76];
    assign P[137] = in[76] ^ in2[76];
    assign G[138] = in[75] & in2[75];
    assign P[138] = in[75] ^ in2[75];
    assign G[139] = in[74] & in2[74];
    assign P[139] = in[74] ^ in2[74];
    assign G[140] = in[73] & in2[73];
    assign P[140] = in[73] ^ in2[73];
    assign G[141] = in[72] & in2[72];
    assign P[141] = in[72] ^ in2[72];
    assign G[142] = in[71] & in2[71];
    assign P[142] = in[71] ^ in2[71];
    assign G[143] = in[70] & in2[70];
    assign P[143] = in[70] ^ in2[70];
    assign G[144] = in[69] & in2[69];
    assign P[144] = in[69] ^ in2[69];
    assign G[145] = in[68] & in2[68];
    assign P[145] = in[68] ^ in2[68];
    assign G[146] = in[67] & in2[67];
    assign P[146] = in[67] ^ in2[67];
    assign G[147] = in[66] & in2[66];
    assign P[147] = in[66] ^ in2[66];
    assign G[148] = in[65] & in2[65];
    assign P[148] = in[65] ^ in2[65];
    assign G[149] = in[64] & in2[64];
    assign P[149] = in[64] ^ in2[64];
    assign G[150] = in[63] & in2[63];
    assign P[150] = in[63] ^ in2[63];
    assign G[151] = in[62] & in2[62];
    assign P[151] = in[62] ^ in2[62];
    assign G[152] = in[61] & in2[61];
    assign P[152] = in[61] ^ in2[61];
    assign G[153] = in[60] & in2[60];
    assign P[153] = in[60] ^ in2[60];
    assign G[154] = in[59] & in2[59];
    assign P[154] = in[59] ^ in2[59];
    assign G[155] = in[58] & in2[58];
    assign P[155] = in[58] ^ in2[58];
    assign G[156] = in[57] & in2[57];
    assign P[156] = in[57] ^ in2[57];
    assign G[157] = in[56] & in2[56];
    assign P[157] = in[56] ^ in2[56];
    assign G[158] = in[55] & in2[55];
    assign P[158] = in[55] ^ in2[55];
    assign G[159] = in[54] & in2[54];
    assign P[159] = in[54] ^ in2[54];
    assign G[160] = in[53] & in2[53];
    assign P[160] = in[53] ^ in2[53];
    assign G[161] = in[52] & in2[52];
    assign P[161] = in[52] ^ in2[52];
    assign G[162] = in[51] & in2[51];
    assign P[162] = in[51] ^ in2[51];
    assign G[163] = in[50] & in2[50];
    assign P[163] = in[50] ^ in2[50];
    assign G[164] = in[49] & in2[49];
    assign P[164] = in[49] ^ in2[49];
    assign G[165] = in[48] & in2[48];
    assign P[165] = in[48] ^ in2[48];
    assign G[166] = in[47] & in2[47];
    assign P[166] = in[47] ^ in2[47];
    assign G[167] = in[46] & in2[46];
    assign P[167] = in[46] ^ in2[46];
    assign G[168] = in[45] & in2[45];
    assign P[168] = in[45] ^ in2[45];
    assign G[169] = in[44] & in2[44];
    assign P[169] = in[44] ^ in2[44];
    assign G[170] = in[43] & in2[43];
    assign P[170] = in[43] ^ in2[43];
    assign G[171] = in[42] & in2[42];
    assign P[171] = in[42] ^ in2[42];
    assign G[172] = in[41] & in2[41];
    assign P[172] = in[41] ^ in2[41];
    assign G[173] = in[40] & in2[40];
    assign P[173] = in[40] ^ in2[40];
    assign G[174] = in[39] & in2[39];
    assign P[174] = in[39] ^ in2[39];
    assign G[175] = in[38] & in2[38];
    assign P[175] = in[38] ^ in2[38];
    assign G[176] = in[37] & in2[37];
    assign P[176] = in[37] ^ in2[37];
    assign G[177] = in[36] & in2[36];
    assign P[177] = in[36] ^ in2[36];
    assign G[178] = in[35] & in2[35];
    assign P[178] = in[35] ^ in2[35];
    assign G[179] = in[34] & in2[34];
    assign P[179] = in[34] ^ in2[34];
    assign G[180] = in[33] & in2[33];
    assign P[180] = in[33] ^ in2[33];
    assign G[181] = in[32] & in2[32];
    assign P[181] = in[32] ^ in2[32];
    assign G[182] = in[31] & in2[31];
    assign P[182] = in[31] ^ in2[31];
    assign G[183] = in[30] & in2[30];
    assign P[183] = in[30] ^ in2[30];
    assign G[184] = in[29] & in2[29];
    assign P[184] = in[29] ^ in2[29];
    assign G[185] = in[28] & in2[28];
    assign P[185] = in[28] ^ in2[28];
    assign G[186] = in[27] & in2[27];
    assign P[186] = in[27] ^ in2[27];
    assign G[187] = in[26] & in2[26];
    assign P[187] = in[26] ^ in2[26];
    assign G[188] = in[25] & in2[25];
    assign P[188] = in[25] ^ in2[25];
    assign G[189] = in[24] & in2[24];
    assign P[189] = in[24] ^ in2[24];
    assign G[190] = in[23] & in2[23];
    assign P[190] = in[23] ^ in2[23];
    assign G[191] = in[22] & in2[22];
    assign P[191] = in[22] ^ in2[22];
    assign G[192] = in[21] & in2[21];
    assign P[192] = in[21] ^ in2[21];
    assign G[193] = in[20] & in2[20];
    assign P[193] = in[20] ^ in2[20];
    assign G[194] = in[19] & in2[19];
    assign P[194] = in[19] ^ in2[19];
    assign G[195] = in[18] & in2[18];
    assign P[195] = in[18] ^ in2[18];
    assign G[196] = in[17] & in2[17];
    assign P[196] = in[17] ^ in2[17];
    assign G[197] = in[16] & in2[16];
    assign P[197] = in[16] ^ in2[16];
    assign G[198] = in[15] & in2[15];
    assign P[198] = in[15] ^ in2[15];
    assign G[199] = in[14] & in2[14];
    assign P[199] = in[14] ^ in2[14];
    assign G[200] = in[13] & in2[13];
    assign P[200] = in[13] ^ in2[13];
    assign G[201] = in[12] & in2[12];
    assign P[201] = in[12] ^ in2[12];
    assign G[202] = in[11] & in2[11];
    assign P[202] = in[11] ^ in2[11];
    assign G[203] = in[10] & in2[10];
    assign P[203] = in[10] ^ in2[10];
    assign G[204] = in[9] & in2[9];
    assign P[204] = in[9] ^ in2[9];
    assign G[205] = in[8] & in2[8];
    assign P[205] = in[8] ^ in2[8];
    assign G[206] = in[7] & in2[7];
    assign P[206] = in[7] ^ in2[7];
    assign G[207] = in[6] & in2[6];
    assign P[207] = in[6] ^ in2[6];
    assign G[208] = in[5] & in2[5];
    assign P[208] = in[5] ^ in2[5];
    assign G[209] = in[4] & in2[4];
    assign P[209] = in[4] ^ in2[4];
    assign G[210] = in[3] & in2[3];
    assign P[210] = in[3] ^ in2[3];
    assign G[211] = in[2] & in2[2];
    assign P[211] = in[2] ^ in2[2];
    assign G[212] = in[1] & in2[1];
    assign P[212] = in[1] ^ in2[1];
    assign G[213] = in[0] & in2[0];
    assign P[213] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign C[213] = G[212] | (P[212] & C[212]);
    assign cout = G[213] | (P[213] & C[213]);
    assign sum = P ^ C;
endmodule

module CLA213(output [212:0] sum, output cout, input [212:0] in1, input [212:0] in2;

    wire[212:0] G;
    wire[212:0] C;
    wire[212:0] P;

    assign G[0] = in[212] & in2[212];
    assign P[0] = in[212] ^ in2[212];
    assign G[1] = in[211] & in2[211];
    assign P[1] = in[211] ^ in2[211];
    assign G[2] = in[210] & in2[210];
    assign P[2] = in[210] ^ in2[210];
    assign G[3] = in[209] & in2[209];
    assign P[3] = in[209] ^ in2[209];
    assign G[4] = in[208] & in2[208];
    assign P[4] = in[208] ^ in2[208];
    assign G[5] = in[207] & in2[207];
    assign P[5] = in[207] ^ in2[207];
    assign G[6] = in[206] & in2[206];
    assign P[6] = in[206] ^ in2[206];
    assign G[7] = in[205] & in2[205];
    assign P[7] = in[205] ^ in2[205];
    assign G[8] = in[204] & in2[204];
    assign P[8] = in[204] ^ in2[204];
    assign G[9] = in[203] & in2[203];
    assign P[9] = in[203] ^ in2[203];
    assign G[10] = in[202] & in2[202];
    assign P[10] = in[202] ^ in2[202];
    assign G[11] = in[201] & in2[201];
    assign P[11] = in[201] ^ in2[201];
    assign G[12] = in[200] & in2[200];
    assign P[12] = in[200] ^ in2[200];
    assign G[13] = in[199] & in2[199];
    assign P[13] = in[199] ^ in2[199];
    assign G[14] = in[198] & in2[198];
    assign P[14] = in[198] ^ in2[198];
    assign G[15] = in[197] & in2[197];
    assign P[15] = in[197] ^ in2[197];
    assign G[16] = in[196] & in2[196];
    assign P[16] = in[196] ^ in2[196];
    assign G[17] = in[195] & in2[195];
    assign P[17] = in[195] ^ in2[195];
    assign G[18] = in[194] & in2[194];
    assign P[18] = in[194] ^ in2[194];
    assign G[19] = in[193] & in2[193];
    assign P[19] = in[193] ^ in2[193];
    assign G[20] = in[192] & in2[192];
    assign P[20] = in[192] ^ in2[192];
    assign G[21] = in[191] & in2[191];
    assign P[21] = in[191] ^ in2[191];
    assign G[22] = in[190] & in2[190];
    assign P[22] = in[190] ^ in2[190];
    assign G[23] = in[189] & in2[189];
    assign P[23] = in[189] ^ in2[189];
    assign G[24] = in[188] & in2[188];
    assign P[24] = in[188] ^ in2[188];
    assign G[25] = in[187] & in2[187];
    assign P[25] = in[187] ^ in2[187];
    assign G[26] = in[186] & in2[186];
    assign P[26] = in[186] ^ in2[186];
    assign G[27] = in[185] & in2[185];
    assign P[27] = in[185] ^ in2[185];
    assign G[28] = in[184] & in2[184];
    assign P[28] = in[184] ^ in2[184];
    assign G[29] = in[183] & in2[183];
    assign P[29] = in[183] ^ in2[183];
    assign G[30] = in[182] & in2[182];
    assign P[30] = in[182] ^ in2[182];
    assign G[31] = in[181] & in2[181];
    assign P[31] = in[181] ^ in2[181];
    assign G[32] = in[180] & in2[180];
    assign P[32] = in[180] ^ in2[180];
    assign G[33] = in[179] & in2[179];
    assign P[33] = in[179] ^ in2[179];
    assign G[34] = in[178] & in2[178];
    assign P[34] = in[178] ^ in2[178];
    assign G[35] = in[177] & in2[177];
    assign P[35] = in[177] ^ in2[177];
    assign G[36] = in[176] & in2[176];
    assign P[36] = in[176] ^ in2[176];
    assign G[37] = in[175] & in2[175];
    assign P[37] = in[175] ^ in2[175];
    assign G[38] = in[174] & in2[174];
    assign P[38] = in[174] ^ in2[174];
    assign G[39] = in[173] & in2[173];
    assign P[39] = in[173] ^ in2[173];
    assign G[40] = in[172] & in2[172];
    assign P[40] = in[172] ^ in2[172];
    assign G[41] = in[171] & in2[171];
    assign P[41] = in[171] ^ in2[171];
    assign G[42] = in[170] & in2[170];
    assign P[42] = in[170] ^ in2[170];
    assign G[43] = in[169] & in2[169];
    assign P[43] = in[169] ^ in2[169];
    assign G[44] = in[168] & in2[168];
    assign P[44] = in[168] ^ in2[168];
    assign G[45] = in[167] & in2[167];
    assign P[45] = in[167] ^ in2[167];
    assign G[46] = in[166] & in2[166];
    assign P[46] = in[166] ^ in2[166];
    assign G[47] = in[165] & in2[165];
    assign P[47] = in[165] ^ in2[165];
    assign G[48] = in[164] & in2[164];
    assign P[48] = in[164] ^ in2[164];
    assign G[49] = in[163] & in2[163];
    assign P[49] = in[163] ^ in2[163];
    assign G[50] = in[162] & in2[162];
    assign P[50] = in[162] ^ in2[162];
    assign G[51] = in[161] & in2[161];
    assign P[51] = in[161] ^ in2[161];
    assign G[52] = in[160] & in2[160];
    assign P[52] = in[160] ^ in2[160];
    assign G[53] = in[159] & in2[159];
    assign P[53] = in[159] ^ in2[159];
    assign G[54] = in[158] & in2[158];
    assign P[54] = in[158] ^ in2[158];
    assign G[55] = in[157] & in2[157];
    assign P[55] = in[157] ^ in2[157];
    assign G[56] = in[156] & in2[156];
    assign P[56] = in[156] ^ in2[156];
    assign G[57] = in[155] & in2[155];
    assign P[57] = in[155] ^ in2[155];
    assign G[58] = in[154] & in2[154];
    assign P[58] = in[154] ^ in2[154];
    assign G[59] = in[153] & in2[153];
    assign P[59] = in[153] ^ in2[153];
    assign G[60] = in[152] & in2[152];
    assign P[60] = in[152] ^ in2[152];
    assign G[61] = in[151] & in2[151];
    assign P[61] = in[151] ^ in2[151];
    assign G[62] = in[150] & in2[150];
    assign P[62] = in[150] ^ in2[150];
    assign G[63] = in[149] & in2[149];
    assign P[63] = in[149] ^ in2[149];
    assign G[64] = in[148] & in2[148];
    assign P[64] = in[148] ^ in2[148];
    assign G[65] = in[147] & in2[147];
    assign P[65] = in[147] ^ in2[147];
    assign G[66] = in[146] & in2[146];
    assign P[66] = in[146] ^ in2[146];
    assign G[67] = in[145] & in2[145];
    assign P[67] = in[145] ^ in2[145];
    assign G[68] = in[144] & in2[144];
    assign P[68] = in[144] ^ in2[144];
    assign G[69] = in[143] & in2[143];
    assign P[69] = in[143] ^ in2[143];
    assign G[70] = in[142] & in2[142];
    assign P[70] = in[142] ^ in2[142];
    assign G[71] = in[141] & in2[141];
    assign P[71] = in[141] ^ in2[141];
    assign G[72] = in[140] & in2[140];
    assign P[72] = in[140] ^ in2[140];
    assign G[73] = in[139] & in2[139];
    assign P[73] = in[139] ^ in2[139];
    assign G[74] = in[138] & in2[138];
    assign P[74] = in[138] ^ in2[138];
    assign G[75] = in[137] & in2[137];
    assign P[75] = in[137] ^ in2[137];
    assign G[76] = in[136] & in2[136];
    assign P[76] = in[136] ^ in2[136];
    assign G[77] = in[135] & in2[135];
    assign P[77] = in[135] ^ in2[135];
    assign G[78] = in[134] & in2[134];
    assign P[78] = in[134] ^ in2[134];
    assign G[79] = in[133] & in2[133];
    assign P[79] = in[133] ^ in2[133];
    assign G[80] = in[132] & in2[132];
    assign P[80] = in[132] ^ in2[132];
    assign G[81] = in[131] & in2[131];
    assign P[81] = in[131] ^ in2[131];
    assign G[82] = in[130] & in2[130];
    assign P[82] = in[130] ^ in2[130];
    assign G[83] = in[129] & in2[129];
    assign P[83] = in[129] ^ in2[129];
    assign G[84] = in[128] & in2[128];
    assign P[84] = in[128] ^ in2[128];
    assign G[85] = in[127] & in2[127];
    assign P[85] = in[127] ^ in2[127];
    assign G[86] = in[126] & in2[126];
    assign P[86] = in[126] ^ in2[126];
    assign G[87] = in[125] & in2[125];
    assign P[87] = in[125] ^ in2[125];
    assign G[88] = in[124] & in2[124];
    assign P[88] = in[124] ^ in2[124];
    assign G[89] = in[123] & in2[123];
    assign P[89] = in[123] ^ in2[123];
    assign G[90] = in[122] & in2[122];
    assign P[90] = in[122] ^ in2[122];
    assign G[91] = in[121] & in2[121];
    assign P[91] = in[121] ^ in2[121];
    assign G[92] = in[120] & in2[120];
    assign P[92] = in[120] ^ in2[120];
    assign G[93] = in[119] & in2[119];
    assign P[93] = in[119] ^ in2[119];
    assign G[94] = in[118] & in2[118];
    assign P[94] = in[118] ^ in2[118];
    assign G[95] = in[117] & in2[117];
    assign P[95] = in[117] ^ in2[117];
    assign G[96] = in[116] & in2[116];
    assign P[96] = in[116] ^ in2[116];
    assign G[97] = in[115] & in2[115];
    assign P[97] = in[115] ^ in2[115];
    assign G[98] = in[114] & in2[114];
    assign P[98] = in[114] ^ in2[114];
    assign G[99] = in[113] & in2[113];
    assign P[99] = in[113] ^ in2[113];
    assign G[100] = in[112] & in2[112];
    assign P[100] = in[112] ^ in2[112];
    assign G[101] = in[111] & in2[111];
    assign P[101] = in[111] ^ in2[111];
    assign G[102] = in[110] & in2[110];
    assign P[102] = in[110] ^ in2[110];
    assign G[103] = in[109] & in2[109];
    assign P[103] = in[109] ^ in2[109];
    assign G[104] = in[108] & in2[108];
    assign P[104] = in[108] ^ in2[108];
    assign G[105] = in[107] & in2[107];
    assign P[105] = in[107] ^ in2[107];
    assign G[106] = in[106] & in2[106];
    assign P[106] = in[106] ^ in2[106];
    assign G[107] = in[105] & in2[105];
    assign P[107] = in[105] ^ in2[105];
    assign G[108] = in[104] & in2[104];
    assign P[108] = in[104] ^ in2[104];
    assign G[109] = in[103] & in2[103];
    assign P[109] = in[103] ^ in2[103];
    assign G[110] = in[102] & in2[102];
    assign P[110] = in[102] ^ in2[102];
    assign G[111] = in[101] & in2[101];
    assign P[111] = in[101] ^ in2[101];
    assign G[112] = in[100] & in2[100];
    assign P[112] = in[100] ^ in2[100];
    assign G[113] = in[99] & in2[99];
    assign P[113] = in[99] ^ in2[99];
    assign G[114] = in[98] & in2[98];
    assign P[114] = in[98] ^ in2[98];
    assign G[115] = in[97] & in2[97];
    assign P[115] = in[97] ^ in2[97];
    assign G[116] = in[96] & in2[96];
    assign P[116] = in[96] ^ in2[96];
    assign G[117] = in[95] & in2[95];
    assign P[117] = in[95] ^ in2[95];
    assign G[118] = in[94] & in2[94];
    assign P[118] = in[94] ^ in2[94];
    assign G[119] = in[93] & in2[93];
    assign P[119] = in[93] ^ in2[93];
    assign G[120] = in[92] & in2[92];
    assign P[120] = in[92] ^ in2[92];
    assign G[121] = in[91] & in2[91];
    assign P[121] = in[91] ^ in2[91];
    assign G[122] = in[90] & in2[90];
    assign P[122] = in[90] ^ in2[90];
    assign G[123] = in[89] & in2[89];
    assign P[123] = in[89] ^ in2[89];
    assign G[124] = in[88] & in2[88];
    assign P[124] = in[88] ^ in2[88];
    assign G[125] = in[87] & in2[87];
    assign P[125] = in[87] ^ in2[87];
    assign G[126] = in[86] & in2[86];
    assign P[126] = in[86] ^ in2[86];
    assign G[127] = in[85] & in2[85];
    assign P[127] = in[85] ^ in2[85];
    assign G[128] = in[84] & in2[84];
    assign P[128] = in[84] ^ in2[84];
    assign G[129] = in[83] & in2[83];
    assign P[129] = in[83] ^ in2[83];
    assign G[130] = in[82] & in2[82];
    assign P[130] = in[82] ^ in2[82];
    assign G[131] = in[81] & in2[81];
    assign P[131] = in[81] ^ in2[81];
    assign G[132] = in[80] & in2[80];
    assign P[132] = in[80] ^ in2[80];
    assign G[133] = in[79] & in2[79];
    assign P[133] = in[79] ^ in2[79];
    assign G[134] = in[78] & in2[78];
    assign P[134] = in[78] ^ in2[78];
    assign G[135] = in[77] & in2[77];
    assign P[135] = in[77] ^ in2[77];
    assign G[136] = in[76] & in2[76];
    assign P[136] = in[76] ^ in2[76];
    assign G[137] = in[75] & in2[75];
    assign P[137] = in[75] ^ in2[75];
    assign G[138] = in[74] & in2[74];
    assign P[138] = in[74] ^ in2[74];
    assign G[139] = in[73] & in2[73];
    assign P[139] = in[73] ^ in2[73];
    assign G[140] = in[72] & in2[72];
    assign P[140] = in[72] ^ in2[72];
    assign G[141] = in[71] & in2[71];
    assign P[141] = in[71] ^ in2[71];
    assign G[142] = in[70] & in2[70];
    assign P[142] = in[70] ^ in2[70];
    assign G[143] = in[69] & in2[69];
    assign P[143] = in[69] ^ in2[69];
    assign G[144] = in[68] & in2[68];
    assign P[144] = in[68] ^ in2[68];
    assign G[145] = in[67] & in2[67];
    assign P[145] = in[67] ^ in2[67];
    assign G[146] = in[66] & in2[66];
    assign P[146] = in[66] ^ in2[66];
    assign G[147] = in[65] & in2[65];
    assign P[147] = in[65] ^ in2[65];
    assign G[148] = in[64] & in2[64];
    assign P[148] = in[64] ^ in2[64];
    assign G[149] = in[63] & in2[63];
    assign P[149] = in[63] ^ in2[63];
    assign G[150] = in[62] & in2[62];
    assign P[150] = in[62] ^ in2[62];
    assign G[151] = in[61] & in2[61];
    assign P[151] = in[61] ^ in2[61];
    assign G[152] = in[60] & in2[60];
    assign P[152] = in[60] ^ in2[60];
    assign G[153] = in[59] & in2[59];
    assign P[153] = in[59] ^ in2[59];
    assign G[154] = in[58] & in2[58];
    assign P[154] = in[58] ^ in2[58];
    assign G[155] = in[57] & in2[57];
    assign P[155] = in[57] ^ in2[57];
    assign G[156] = in[56] & in2[56];
    assign P[156] = in[56] ^ in2[56];
    assign G[157] = in[55] & in2[55];
    assign P[157] = in[55] ^ in2[55];
    assign G[158] = in[54] & in2[54];
    assign P[158] = in[54] ^ in2[54];
    assign G[159] = in[53] & in2[53];
    assign P[159] = in[53] ^ in2[53];
    assign G[160] = in[52] & in2[52];
    assign P[160] = in[52] ^ in2[52];
    assign G[161] = in[51] & in2[51];
    assign P[161] = in[51] ^ in2[51];
    assign G[162] = in[50] & in2[50];
    assign P[162] = in[50] ^ in2[50];
    assign G[163] = in[49] & in2[49];
    assign P[163] = in[49] ^ in2[49];
    assign G[164] = in[48] & in2[48];
    assign P[164] = in[48] ^ in2[48];
    assign G[165] = in[47] & in2[47];
    assign P[165] = in[47] ^ in2[47];
    assign G[166] = in[46] & in2[46];
    assign P[166] = in[46] ^ in2[46];
    assign G[167] = in[45] & in2[45];
    assign P[167] = in[45] ^ in2[45];
    assign G[168] = in[44] & in2[44];
    assign P[168] = in[44] ^ in2[44];
    assign G[169] = in[43] & in2[43];
    assign P[169] = in[43] ^ in2[43];
    assign G[170] = in[42] & in2[42];
    assign P[170] = in[42] ^ in2[42];
    assign G[171] = in[41] & in2[41];
    assign P[171] = in[41] ^ in2[41];
    assign G[172] = in[40] & in2[40];
    assign P[172] = in[40] ^ in2[40];
    assign G[173] = in[39] & in2[39];
    assign P[173] = in[39] ^ in2[39];
    assign G[174] = in[38] & in2[38];
    assign P[174] = in[38] ^ in2[38];
    assign G[175] = in[37] & in2[37];
    assign P[175] = in[37] ^ in2[37];
    assign G[176] = in[36] & in2[36];
    assign P[176] = in[36] ^ in2[36];
    assign G[177] = in[35] & in2[35];
    assign P[177] = in[35] ^ in2[35];
    assign G[178] = in[34] & in2[34];
    assign P[178] = in[34] ^ in2[34];
    assign G[179] = in[33] & in2[33];
    assign P[179] = in[33] ^ in2[33];
    assign G[180] = in[32] & in2[32];
    assign P[180] = in[32] ^ in2[32];
    assign G[181] = in[31] & in2[31];
    assign P[181] = in[31] ^ in2[31];
    assign G[182] = in[30] & in2[30];
    assign P[182] = in[30] ^ in2[30];
    assign G[183] = in[29] & in2[29];
    assign P[183] = in[29] ^ in2[29];
    assign G[184] = in[28] & in2[28];
    assign P[184] = in[28] ^ in2[28];
    assign G[185] = in[27] & in2[27];
    assign P[185] = in[27] ^ in2[27];
    assign G[186] = in[26] & in2[26];
    assign P[186] = in[26] ^ in2[26];
    assign G[187] = in[25] & in2[25];
    assign P[187] = in[25] ^ in2[25];
    assign G[188] = in[24] & in2[24];
    assign P[188] = in[24] ^ in2[24];
    assign G[189] = in[23] & in2[23];
    assign P[189] = in[23] ^ in2[23];
    assign G[190] = in[22] & in2[22];
    assign P[190] = in[22] ^ in2[22];
    assign G[191] = in[21] & in2[21];
    assign P[191] = in[21] ^ in2[21];
    assign G[192] = in[20] & in2[20];
    assign P[192] = in[20] ^ in2[20];
    assign G[193] = in[19] & in2[19];
    assign P[193] = in[19] ^ in2[19];
    assign G[194] = in[18] & in2[18];
    assign P[194] = in[18] ^ in2[18];
    assign G[195] = in[17] & in2[17];
    assign P[195] = in[17] ^ in2[17];
    assign G[196] = in[16] & in2[16];
    assign P[196] = in[16] ^ in2[16];
    assign G[197] = in[15] & in2[15];
    assign P[197] = in[15] ^ in2[15];
    assign G[198] = in[14] & in2[14];
    assign P[198] = in[14] ^ in2[14];
    assign G[199] = in[13] & in2[13];
    assign P[199] = in[13] ^ in2[13];
    assign G[200] = in[12] & in2[12];
    assign P[200] = in[12] ^ in2[12];
    assign G[201] = in[11] & in2[11];
    assign P[201] = in[11] ^ in2[11];
    assign G[202] = in[10] & in2[10];
    assign P[202] = in[10] ^ in2[10];
    assign G[203] = in[9] & in2[9];
    assign P[203] = in[9] ^ in2[9];
    assign G[204] = in[8] & in2[8];
    assign P[204] = in[8] ^ in2[8];
    assign G[205] = in[7] & in2[7];
    assign P[205] = in[7] ^ in2[7];
    assign G[206] = in[6] & in2[6];
    assign P[206] = in[6] ^ in2[6];
    assign G[207] = in[5] & in2[5];
    assign P[207] = in[5] ^ in2[5];
    assign G[208] = in[4] & in2[4];
    assign P[208] = in[4] ^ in2[4];
    assign G[209] = in[3] & in2[3];
    assign P[209] = in[3] ^ in2[3];
    assign G[210] = in[2] & in2[2];
    assign P[210] = in[2] ^ in2[2];
    assign G[211] = in[1] & in2[1];
    assign P[211] = in[1] ^ in2[1];
    assign G[212] = in[0] & in2[0];
    assign P[212] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign C[212] = G[211] | (P[211] & C[211]);
    assign cout = G[212] | (P[212] & C[212]);
    assign sum = P ^ C;
endmodule

module CLA212(output [211:0] sum, output cout, input [211:0] in1, input [211:0] in2;

    wire[211:0] G;
    wire[211:0] C;
    wire[211:0] P;

    assign G[0] = in[211] & in2[211];
    assign P[0] = in[211] ^ in2[211];
    assign G[1] = in[210] & in2[210];
    assign P[1] = in[210] ^ in2[210];
    assign G[2] = in[209] & in2[209];
    assign P[2] = in[209] ^ in2[209];
    assign G[3] = in[208] & in2[208];
    assign P[3] = in[208] ^ in2[208];
    assign G[4] = in[207] & in2[207];
    assign P[4] = in[207] ^ in2[207];
    assign G[5] = in[206] & in2[206];
    assign P[5] = in[206] ^ in2[206];
    assign G[6] = in[205] & in2[205];
    assign P[6] = in[205] ^ in2[205];
    assign G[7] = in[204] & in2[204];
    assign P[7] = in[204] ^ in2[204];
    assign G[8] = in[203] & in2[203];
    assign P[8] = in[203] ^ in2[203];
    assign G[9] = in[202] & in2[202];
    assign P[9] = in[202] ^ in2[202];
    assign G[10] = in[201] & in2[201];
    assign P[10] = in[201] ^ in2[201];
    assign G[11] = in[200] & in2[200];
    assign P[11] = in[200] ^ in2[200];
    assign G[12] = in[199] & in2[199];
    assign P[12] = in[199] ^ in2[199];
    assign G[13] = in[198] & in2[198];
    assign P[13] = in[198] ^ in2[198];
    assign G[14] = in[197] & in2[197];
    assign P[14] = in[197] ^ in2[197];
    assign G[15] = in[196] & in2[196];
    assign P[15] = in[196] ^ in2[196];
    assign G[16] = in[195] & in2[195];
    assign P[16] = in[195] ^ in2[195];
    assign G[17] = in[194] & in2[194];
    assign P[17] = in[194] ^ in2[194];
    assign G[18] = in[193] & in2[193];
    assign P[18] = in[193] ^ in2[193];
    assign G[19] = in[192] & in2[192];
    assign P[19] = in[192] ^ in2[192];
    assign G[20] = in[191] & in2[191];
    assign P[20] = in[191] ^ in2[191];
    assign G[21] = in[190] & in2[190];
    assign P[21] = in[190] ^ in2[190];
    assign G[22] = in[189] & in2[189];
    assign P[22] = in[189] ^ in2[189];
    assign G[23] = in[188] & in2[188];
    assign P[23] = in[188] ^ in2[188];
    assign G[24] = in[187] & in2[187];
    assign P[24] = in[187] ^ in2[187];
    assign G[25] = in[186] & in2[186];
    assign P[25] = in[186] ^ in2[186];
    assign G[26] = in[185] & in2[185];
    assign P[26] = in[185] ^ in2[185];
    assign G[27] = in[184] & in2[184];
    assign P[27] = in[184] ^ in2[184];
    assign G[28] = in[183] & in2[183];
    assign P[28] = in[183] ^ in2[183];
    assign G[29] = in[182] & in2[182];
    assign P[29] = in[182] ^ in2[182];
    assign G[30] = in[181] & in2[181];
    assign P[30] = in[181] ^ in2[181];
    assign G[31] = in[180] & in2[180];
    assign P[31] = in[180] ^ in2[180];
    assign G[32] = in[179] & in2[179];
    assign P[32] = in[179] ^ in2[179];
    assign G[33] = in[178] & in2[178];
    assign P[33] = in[178] ^ in2[178];
    assign G[34] = in[177] & in2[177];
    assign P[34] = in[177] ^ in2[177];
    assign G[35] = in[176] & in2[176];
    assign P[35] = in[176] ^ in2[176];
    assign G[36] = in[175] & in2[175];
    assign P[36] = in[175] ^ in2[175];
    assign G[37] = in[174] & in2[174];
    assign P[37] = in[174] ^ in2[174];
    assign G[38] = in[173] & in2[173];
    assign P[38] = in[173] ^ in2[173];
    assign G[39] = in[172] & in2[172];
    assign P[39] = in[172] ^ in2[172];
    assign G[40] = in[171] & in2[171];
    assign P[40] = in[171] ^ in2[171];
    assign G[41] = in[170] & in2[170];
    assign P[41] = in[170] ^ in2[170];
    assign G[42] = in[169] & in2[169];
    assign P[42] = in[169] ^ in2[169];
    assign G[43] = in[168] & in2[168];
    assign P[43] = in[168] ^ in2[168];
    assign G[44] = in[167] & in2[167];
    assign P[44] = in[167] ^ in2[167];
    assign G[45] = in[166] & in2[166];
    assign P[45] = in[166] ^ in2[166];
    assign G[46] = in[165] & in2[165];
    assign P[46] = in[165] ^ in2[165];
    assign G[47] = in[164] & in2[164];
    assign P[47] = in[164] ^ in2[164];
    assign G[48] = in[163] & in2[163];
    assign P[48] = in[163] ^ in2[163];
    assign G[49] = in[162] & in2[162];
    assign P[49] = in[162] ^ in2[162];
    assign G[50] = in[161] & in2[161];
    assign P[50] = in[161] ^ in2[161];
    assign G[51] = in[160] & in2[160];
    assign P[51] = in[160] ^ in2[160];
    assign G[52] = in[159] & in2[159];
    assign P[52] = in[159] ^ in2[159];
    assign G[53] = in[158] & in2[158];
    assign P[53] = in[158] ^ in2[158];
    assign G[54] = in[157] & in2[157];
    assign P[54] = in[157] ^ in2[157];
    assign G[55] = in[156] & in2[156];
    assign P[55] = in[156] ^ in2[156];
    assign G[56] = in[155] & in2[155];
    assign P[56] = in[155] ^ in2[155];
    assign G[57] = in[154] & in2[154];
    assign P[57] = in[154] ^ in2[154];
    assign G[58] = in[153] & in2[153];
    assign P[58] = in[153] ^ in2[153];
    assign G[59] = in[152] & in2[152];
    assign P[59] = in[152] ^ in2[152];
    assign G[60] = in[151] & in2[151];
    assign P[60] = in[151] ^ in2[151];
    assign G[61] = in[150] & in2[150];
    assign P[61] = in[150] ^ in2[150];
    assign G[62] = in[149] & in2[149];
    assign P[62] = in[149] ^ in2[149];
    assign G[63] = in[148] & in2[148];
    assign P[63] = in[148] ^ in2[148];
    assign G[64] = in[147] & in2[147];
    assign P[64] = in[147] ^ in2[147];
    assign G[65] = in[146] & in2[146];
    assign P[65] = in[146] ^ in2[146];
    assign G[66] = in[145] & in2[145];
    assign P[66] = in[145] ^ in2[145];
    assign G[67] = in[144] & in2[144];
    assign P[67] = in[144] ^ in2[144];
    assign G[68] = in[143] & in2[143];
    assign P[68] = in[143] ^ in2[143];
    assign G[69] = in[142] & in2[142];
    assign P[69] = in[142] ^ in2[142];
    assign G[70] = in[141] & in2[141];
    assign P[70] = in[141] ^ in2[141];
    assign G[71] = in[140] & in2[140];
    assign P[71] = in[140] ^ in2[140];
    assign G[72] = in[139] & in2[139];
    assign P[72] = in[139] ^ in2[139];
    assign G[73] = in[138] & in2[138];
    assign P[73] = in[138] ^ in2[138];
    assign G[74] = in[137] & in2[137];
    assign P[74] = in[137] ^ in2[137];
    assign G[75] = in[136] & in2[136];
    assign P[75] = in[136] ^ in2[136];
    assign G[76] = in[135] & in2[135];
    assign P[76] = in[135] ^ in2[135];
    assign G[77] = in[134] & in2[134];
    assign P[77] = in[134] ^ in2[134];
    assign G[78] = in[133] & in2[133];
    assign P[78] = in[133] ^ in2[133];
    assign G[79] = in[132] & in2[132];
    assign P[79] = in[132] ^ in2[132];
    assign G[80] = in[131] & in2[131];
    assign P[80] = in[131] ^ in2[131];
    assign G[81] = in[130] & in2[130];
    assign P[81] = in[130] ^ in2[130];
    assign G[82] = in[129] & in2[129];
    assign P[82] = in[129] ^ in2[129];
    assign G[83] = in[128] & in2[128];
    assign P[83] = in[128] ^ in2[128];
    assign G[84] = in[127] & in2[127];
    assign P[84] = in[127] ^ in2[127];
    assign G[85] = in[126] & in2[126];
    assign P[85] = in[126] ^ in2[126];
    assign G[86] = in[125] & in2[125];
    assign P[86] = in[125] ^ in2[125];
    assign G[87] = in[124] & in2[124];
    assign P[87] = in[124] ^ in2[124];
    assign G[88] = in[123] & in2[123];
    assign P[88] = in[123] ^ in2[123];
    assign G[89] = in[122] & in2[122];
    assign P[89] = in[122] ^ in2[122];
    assign G[90] = in[121] & in2[121];
    assign P[90] = in[121] ^ in2[121];
    assign G[91] = in[120] & in2[120];
    assign P[91] = in[120] ^ in2[120];
    assign G[92] = in[119] & in2[119];
    assign P[92] = in[119] ^ in2[119];
    assign G[93] = in[118] & in2[118];
    assign P[93] = in[118] ^ in2[118];
    assign G[94] = in[117] & in2[117];
    assign P[94] = in[117] ^ in2[117];
    assign G[95] = in[116] & in2[116];
    assign P[95] = in[116] ^ in2[116];
    assign G[96] = in[115] & in2[115];
    assign P[96] = in[115] ^ in2[115];
    assign G[97] = in[114] & in2[114];
    assign P[97] = in[114] ^ in2[114];
    assign G[98] = in[113] & in2[113];
    assign P[98] = in[113] ^ in2[113];
    assign G[99] = in[112] & in2[112];
    assign P[99] = in[112] ^ in2[112];
    assign G[100] = in[111] & in2[111];
    assign P[100] = in[111] ^ in2[111];
    assign G[101] = in[110] & in2[110];
    assign P[101] = in[110] ^ in2[110];
    assign G[102] = in[109] & in2[109];
    assign P[102] = in[109] ^ in2[109];
    assign G[103] = in[108] & in2[108];
    assign P[103] = in[108] ^ in2[108];
    assign G[104] = in[107] & in2[107];
    assign P[104] = in[107] ^ in2[107];
    assign G[105] = in[106] & in2[106];
    assign P[105] = in[106] ^ in2[106];
    assign G[106] = in[105] & in2[105];
    assign P[106] = in[105] ^ in2[105];
    assign G[107] = in[104] & in2[104];
    assign P[107] = in[104] ^ in2[104];
    assign G[108] = in[103] & in2[103];
    assign P[108] = in[103] ^ in2[103];
    assign G[109] = in[102] & in2[102];
    assign P[109] = in[102] ^ in2[102];
    assign G[110] = in[101] & in2[101];
    assign P[110] = in[101] ^ in2[101];
    assign G[111] = in[100] & in2[100];
    assign P[111] = in[100] ^ in2[100];
    assign G[112] = in[99] & in2[99];
    assign P[112] = in[99] ^ in2[99];
    assign G[113] = in[98] & in2[98];
    assign P[113] = in[98] ^ in2[98];
    assign G[114] = in[97] & in2[97];
    assign P[114] = in[97] ^ in2[97];
    assign G[115] = in[96] & in2[96];
    assign P[115] = in[96] ^ in2[96];
    assign G[116] = in[95] & in2[95];
    assign P[116] = in[95] ^ in2[95];
    assign G[117] = in[94] & in2[94];
    assign P[117] = in[94] ^ in2[94];
    assign G[118] = in[93] & in2[93];
    assign P[118] = in[93] ^ in2[93];
    assign G[119] = in[92] & in2[92];
    assign P[119] = in[92] ^ in2[92];
    assign G[120] = in[91] & in2[91];
    assign P[120] = in[91] ^ in2[91];
    assign G[121] = in[90] & in2[90];
    assign P[121] = in[90] ^ in2[90];
    assign G[122] = in[89] & in2[89];
    assign P[122] = in[89] ^ in2[89];
    assign G[123] = in[88] & in2[88];
    assign P[123] = in[88] ^ in2[88];
    assign G[124] = in[87] & in2[87];
    assign P[124] = in[87] ^ in2[87];
    assign G[125] = in[86] & in2[86];
    assign P[125] = in[86] ^ in2[86];
    assign G[126] = in[85] & in2[85];
    assign P[126] = in[85] ^ in2[85];
    assign G[127] = in[84] & in2[84];
    assign P[127] = in[84] ^ in2[84];
    assign G[128] = in[83] & in2[83];
    assign P[128] = in[83] ^ in2[83];
    assign G[129] = in[82] & in2[82];
    assign P[129] = in[82] ^ in2[82];
    assign G[130] = in[81] & in2[81];
    assign P[130] = in[81] ^ in2[81];
    assign G[131] = in[80] & in2[80];
    assign P[131] = in[80] ^ in2[80];
    assign G[132] = in[79] & in2[79];
    assign P[132] = in[79] ^ in2[79];
    assign G[133] = in[78] & in2[78];
    assign P[133] = in[78] ^ in2[78];
    assign G[134] = in[77] & in2[77];
    assign P[134] = in[77] ^ in2[77];
    assign G[135] = in[76] & in2[76];
    assign P[135] = in[76] ^ in2[76];
    assign G[136] = in[75] & in2[75];
    assign P[136] = in[75] ^ in2[75];
    assign G[137] = in[74] & in2[74];
    assign P[137] = in[74] ^ in2[74];
    assign G[138] = in[73] & in2[73];
    assign P[138] = in[73] ^ in2[73];
    assign G[139] = in[72] & in2[72];
    assign P[139] = in[72] ^ in2[72];
    assign G[140] = in[71] & in2[71];
    assign P[140] = in[71] ^ in2[71];
    assign G[141] = in[70] & in2[70];
    assign P[141] = in[70] ^ in2[70];
    assign G[142] = in[69] & in2[69];
    assign P[142] = in[69] ^ in2[69];
    assign G[143] = in[68] & in2[68];
    assign P[143] = in[68] ^ in2[68];
    assign G[144] = in[67] & in2[67];
    assign P[144] = in[67] ^ in2[67];
    assign G[145] = in[66] & in2[66];
    assign P[145] = in[66] ^ in2[66];
    assign G[146] = in[65] & in2[65];
    assign P[146] = in[65] ^ in2[65];
    assign G[147] = in[64] & in2[64];
    assign P[147] = in[64] ^ in2[64];
    assign G[148] = in[63] & in2[63];
    assign P[148] = in[63] ^ in2[63];
    assign G[149] = in[62] & in2[62];
    assign P[149] = in[62] ^ in2[62];
    assign G[150] = in[61] & in2[61];
    assign P[150] = in[61] ^ in2[61];
    assign G[151] = in[60] & in2[60];
    assign P[151] = in[60] ^ in2[60];
    assign G[152] = in[59] & in2[59];
    assign P[152] = in[59] ^ in2[59];
    assign G[153] = in[58] & in2[58];
    assign P[153] = in[58] ^ in2[58];
    assign G[154] = in[57] & in2[57];
    assign P[154] = in[57] ^ in2[57];
    assign G[155] = in[56] & in2[56];
    assign P[155] = in[56] ^ in2[56];
    assign G[156] = in[55] & in2[55];
    assign P[156] = in[55] ^ in2[55];
    assign G[157] = in[54] & in2[54];
    assign P[157] = in[54] ^ in2[54];
    assign G[158] = in[53] & in2[53];
    assign P[158] = in[53] ^ in2[53];
    assign G[159] = in[52] & in2[52];
    assign P[159] = in[52] ^ in2[52];
    assign G[160] = in[51] & in2[51];
    assign P[160] = in[51] ^ in2[51];
    assign G[161] = in[50] & in2[50];
    assign P[161] = in[50] ^ in2[50];
    assign G[162] = in[49] & in2[49];
    assign P[162] = in[49] ^ in2[49];
    assign G[163] = in[48] & in2[48];
    assign P[163] = in[48] ^ in2[48];
    assign G[164] = in[47] & in2[47];
    assign P[164] = in[47] ^ in2[47];
    assign G[165] = in[46] & in2[46];
    assign P[165] = in[46] ^ in2[46];
    assign G[166] = in[45] & in2[45];
    assign P[166] = in[45] ^ in2[45];
    assign G[167] = in[44] & in2[44];
    assign P[167] = in[44] ^ in2[44];
    assign G[168] = in[43] & in2[43];
    assign P[168] = in[43] ^ in2[43];
    assign G[169] = in[42] & in2[42];
    assign P[169] = in[42] ^ in2[42];
    assign G[170] = in[41] & in2[41];
    assign P[170] = in[41] ^ in2[41];
    assign G[171] = in[40] & in2[40];
    assign P[171] = in[40] ^ in2[40];
    assign G[172] = in[39] & in2[39];
    assign P[172] = in[39] ^ in2[39];
    assign G[173] = in[38] & in2[38];
    assign P[173] = in[38] ^ in2[38];
    assign G[174] = in[37] & in2[37];
    assign P[174] = in[37] ^ in2[37];
    assign G[175] = in[36] & in2[36];
    assign P[175] = in[36] ^ in2[36];
    assign G[176] = in[35] & in2[35];
    assign P[176] = in[35] ^ in2[35];
    assign G[177] = in[34] & in2[34];
    assign P[177] = in[34] ^ in2[34];
    assign G[178] = in[33] & in2[33];
    assign P[178] = in[33] ^ in2[33];
    assign G[179] = in[32] & in2[32];
    assign P[179] = in[32] ^ in2[32];
    assign G[180] = in[31] & in2[31];
    assign P[180] = in[31] ^ in2[31];
    assign G[181] = in[30] & in2[30];
    assign P[181] = in[30] ^ in2[30];
    assign G[182] = in[29] & in2[29];
    assign P[182] = in[29] ^ in2[29];
    assign G[183] = in[28] & in2[28];
    assign P[183] = in[28] ^ in2[28];
    assign G[184] = in[27] & in2[27];
    assign P[184] = in[27] ^ in2[27];
    assign G[185] = in[26] & in2[26];
    assign P[185] = in[26] ^ in2[26];
    assign G[186] = in[25] & in2[25];
    assign P[186] = in[25] ^ in2[25];
    assign G[187] = in[24] & in2[24];
    assign P[187] = in[24] ^ in2[24];
    assign G[188] = in[23] & in2[23];
    assign P[188] = in[23] ^ in2[23];
    assign G[189] = in[22] & in2[22];
    assign P[189] = in[22] ^ in2[22];
    assign G[190] = in[21] & in2[21];
    assign P[190] = in[21] ^ in2[21];
    assign G[191] = in[20] & in2[20];
    assign P[191] = in[20] ^ in2[20];
    assign G[192] = in[19] & in2[19];
    assign P[192] = in[19] ^ in2[19];
    assign G[193] = in[18] & in2[18];
    assign P[193] = in[18] ^ in2[18];
    assign G[194] = in[17] & in2[17];
    assign P[194] = in[17] ^ in2[17];
    assign G[195] = in[16] & in2[16];
    assign P[195] = in[16] ^ in2[16];
    assign G[196] = in[15] & in2[15];
    assign P[196] = in[15] ^ in2[15];
    assign G[197] = in[14] & in2[14];
    assign P[197] = in[14] ^ in2[14];
    assign G[198] = in[13] & in2[13];
    assign P[198] = in[13] ^ in2[13];
    assign G[199] = in[12] & in2[12];
    assign P[199] = in[12] ^ in2[12];
    assign G[200] = in[11] & in2[11];
    assign P[200] = in[11] ^ in2[11];
    assign G[201] = in[10] & in2[10];
    assign P[201] = in[10] ^ in2[10];
    assign G[202] = in[9] & in2[9];
    assign P[202] = in[9] ^ in2[9];
    assign G[203] = in[8] & in2[8];
    assign P[203] = in[8] ^ in2[8];
    assign G[204] = in[7] & in2[7];
    assign P[204] = in[7] ^ in2[7];
    assign G[205] = in[6] & in2[6];
    assign P[205] = in[6] ^ in2[6];
    assign G[206] = in[5] & in2[5];
    assign P[206] = in[5] ^ in2[5];
    assign G[207] = in[4] & in2[4];
    assign P[207] = in[4] ^ in2[4];
    assign G[208] = in[3] & in2[3];
    assign P[208] = in[3] ^ in2[3];
    assign G[209] = in[2] & in2[2];
    assign P[209] = in[2] ^ in2[2];
    assign G[210] = in[1] & in2[1];
    assign P[210] = in[1] ^ in2[1];
    assign G[211] = in[0] & in2[0];
    assign P[211] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign C[211] = G[210] | (P[210] & C[210]);
    assign cout = G[211] | (P[211] & C[211]);
    assign sum = P ^ C;
endmodule

module CLA211(output [210:0] sum, output cout, input [210:0] in1, input [210:0] in2;

    wire[210:0] G;
    wire[210:0] C;
    wire[210:0] P;

    assign G[0] = in[210] & in2[210];
    assign P[0] = in[210] ^ in2[210];
    assign G[1] = in[209] & in2[209];
    assign P[1] = in[209] ^ in2[209];
    assign G[2] = in[208] & in2[208];
    assign P[2] = in[208] ^ in2[208];
    assign G[3] = in[207] & in2[207];
    assign P[3] = in[207] ^ in2[207];
    assign G[4] = in[206] & in2[206];
    assign P[4] = in[206] ^ in2[206];
    assign G[5] = in[205] & in2[205];
    assign P[5] = in[205] ^ in2[205];
    assign G[6] = in[204] & in2[204];
    assign P[6] = in[204] ^ in2[204];
    assign G[7] = in[203] & in2[203];
    assign P[7] = in[203] ^ in2[203];
    assign G[8] = in[202] & in2[202];
    assign P[8] = in[202] ^ in2[202];
    assign G[9] = in[201] & in2[201];
    assign P[9] = in[201] ^ in2[201];
    assign G[10] = in[200] & in2[200];
    assign P[10] = in[200] ^ in2[200];
    assign G[11] = in[199] & in2[199];
    assign P[11] = in[199] ^ in2[199];
    assign G[12] = in[198] & in2[198];
    assign P[12] = in[198] ^ in2[198];
    assign G[13] = in[197] & in2[197];
    assign P[13] = in[197] ^ in2[197];
    assign G[14] = in[196] & in2[196];
    assign P[14] = in[196] ^ in2[196];
    assign G[15] = in[195] & in2[195];
    assign P[15] = in[195] ^ in2[195];
    assign G[16] = in[194] & in2[194];
    assign P[16] = in[194] ^ in2[194];
    assign G[17] = in[193] & in2[193];
    assign P[17] = in[193] ^ in2[193];
    assign G[18] = in[192] & in2[192];
    assign P[18] = in[192] ^ in2[192];
    assign G[19] = in[191] & in2[191];
    assign P[19] = in[191] ^ in2[191];
    assign G[20] = in[190] & in2[190];
    assign P[20] = in[190] ^ in2[190];
    assign G[21] = in[189] & in2[189];
    assign P[21] = in[189] ^ in2[189];
    assign G[22] = in[188] & in2[188];
    assign P[22] = in[188] ^ in2[188];
    assign G[23] = in[187] & in2[187];
    assign P[23] = in[187] ^ in2[187];
    assign G[24] = in[186] & in2[186];
    assign P[24] = in[186] ^ in2[186];
    assign G[25] = in[185] & in2[185];
    assign P[25] = in[185] ^ in2[185];
    assign G[26] = in[184] & in2[184];
    assign P[26] = in[184] ^ in2[184];
    assign G[27] = in[183] & in2[183];
    assign P[27] = in[183] ^ in2[183];
    assign G[28] = in[182] & in2[182];
    assign P[28] = in[182] ^ in2[182];
    assign G[29] = in[181] & in2[181];
    assign P[29] = in[181] ^ in2[181];
    assign G[30] = in[180] & in2[180];
    assign P[30] = in[180] ^ in2[180];
    assign G[31] = in[179] & in2[179];
    assign P[31] = in[179] ^ in2[179];
    assign G[32] = in[178] & in2[178];
    assign P[32] = in[178] ^ in2[178];
    assign G[33] = in[177] & in2[177];
    assign P[33] = in[177] ^ in2[177];
    assign G[34] = in[176] & in2[176];
    assign P[34] = in[176] ^ in2[176];
    assign G[35] = in[175] & in2[175];
    assign P[35] = in[175] ^ in2[175];
    assign G[36] = in[174] & in2[174];
    assign P[36] = in[174] ^ in2[174];
    assign G[37] = in[173] & in2[173];
    assign P[37] = in[173] ^ in2[173];
    assign G[38] = in[172] & in2[172];
    assign P[38] = in[172] ^ in2[172];
    assign G[39] = in[171] & in2[171];
    assign P[39] = in[171] ^ in2[171];
    assign G[40] = in[170] & in2[170];
    assign P[40] = in[170] ^ in2[170];
    assign G[41] = in[169] & in2[169];
    assign P[41] = in[169] ^ in2[169];
    assign G[42] = in[168] & in2[168];
    assign P[42] = in[168] ^ in2[168];
    assign G[43] = in[167] & in2[167];
    assign P[43] = in[167] ^ in2[167];
    assign G[44] = in[166] & in2[166];
    assign P[44] = in[166] ^ in2[166];
    assign G[45] = in[165] & in2[165];
    assign P[45] = in[165] ^ in2[165];
    assign G[46] = in[164] & in2[164];
    assign P[46] = in[164] ^ in2[164];
    assign G[47] = in[163] & in2[163];
    assign P[47] = in[163] ^ in2[163];
    assign G[48] = in[162] & in2[162];
    assign P[48] = in[162] ^ in2[162];
    assign G[49] = in[161] & in2[161];
    assign P[49] = in[161] ^ in2[161];
    assign G[50] = in[160] & in2[160];
    assign P[50] = in[160] ^ in2[160];
    assign G[51] = in[159] & in2[159];
    assign P[51] = in[159] ^ in2[159];
    assign G[52] = in[158] & in2[158];
    assign P[52] = in[158] ^ in2[158];
    assign G[53] = in[157] & in2[157];
    assign P[53] = in[157] ^ in2[157];
    assign G[54] = in[156] & in2[156];
    assign P[54] = in[156] ^ in2[156];
    assign G[55] = in[155] & in2[155];
    assign P[55] = in[155] ^ in2[155];
    assign G[56] = in[154] & in2[154];
    assign P[56] = in[154] ^ in2[154];
    assign G[57] = in[153] & in2[153];
    assign P[57] = in[153] ^ in2[153];
    assign G[58] = in[152] & in2[152];
    assign P[58] = in[152] ^ in2[152];
    assign G[59] = in[151] & in2[151];
    assign P[59] = in[151] ^ in2[151];
    assign G[60] = in[150] & in2[150];
    assign P[60] = in[150] ^ in2[150];
    assign G[61] = in[149] & in2[149];
    assign P[61] = in[149] ^ in2[149];
    assign G[62] = in[148] & in2[148];
    assign P[62] = in[148] ^ in2[148];
    assign G[63] = in[147] & in2[147];
    assign P[63] = in[147] ^ in2[147];
    assign G[64] = in[146] & in2[146];
    assign P[64] = in[146] ^ in2[146];
    assign G[65] = in[145] & in2[145];
    assign P[65] = in[145] ^ in2[145];
    assign G[66] = in[144] & in2[144];
    assign P[66] = in[144] ^ in2[144];
    assign G[67] = in[143] & in2[143];
    assign P[67] = in[143] ^ in2[143];
    assign G[68] = in[142] & in2[142];
    assign P[68] = in[142] ^ in2[142];
    assign G[69] = in[141] & in2[141];
    assign P[69] = in[141] ^ in2[141];
    assign G[70] = in[140] & in2[140];
    assign P[70] = in[140] ^ in2[140];
    assign G[71] = in[139] & in2[139];
    assign P[71] = in[139] ^ in2[139];
    assign G[72] = in[138] & in2[138];
    assign P[72] = in[138] ^ in2[138];
    assign G[73] = in[137] & in2[137];
    assign P[73] = in[137] ^ in2[137];
    assign G[74] = in[136] & in2[136];
    assign P[74] = in[136] ^ in2[136];
    assign G[75] = in[135] & in2[135];
    assign P[75] = in[135] ^ in2[135];
    assign G[76] = in[134] & in2[134];
    assign P[76] = in[134] ^ in2[134];
    assign G[77] = in[133] & in2[133];
    assign P[77] = in[133] ^ in2[133];
    assign G[78] = in[132] & in2[132];
    assign P[78] = in[132] ^ in2[132];
    assign G[79] = in[131] & in2[131];
    assign P[79] = in[131] ^ in2[131];
    assign G[80] = in[130] & in2[130];
    assign P[80] = in[130] ^ in2[130];
    assign G[81] = in[129] & in2[129];
    assign P[81] = in[129] ^ in2[129];
    assign G[82] = in[128] & in2[128];
    assign P[82] = in[128] ^ in2[128];
    assign G[83] = in[127] & in2[127];
    assign P[83] = in[127] ^ in2[127];
    assign G[84] = in[126] & in2[126];
    assign P[84] = in[126] ^ in2[126];
    assign G[85] = in[125] & in2[125];
    assign P[85] = in[125] ^ in2[125];
    assign G[86] = in[124] & in2[124];
    assign P[86] = in[124] ^ in2[124];
    assign G[87] = in[123] & in2[123];
    assign P[87] = in[123] ^ in2[123];
    assign G[88] = in[122] & in2[122];
    assign P[88] = in[122] ^ in2[122];
    assign G[89] = in[121] & in2[121];
    assign P[89] = in[121] ^ in2[121];
    assign G[90] = in[120] & in2[120];
    assign P[90] = in[120] ^ in2[120];
    assign G[91] = in[119] & in2[119];
    assign P[91] = in[119] ^ in2[119];
    assign G[92] = in[118] & in2[118];
    assign P[92] = in[118] ^ in2[118];
    assign G[93] = in[117] & in2[117];
    assign P[93] = in[117] ^ in2[117];
    assign G[94] = in[116] & in2[116];
    assign P[94] = in[116] ^ in2[116];
    assign G[95] = in[115] & in2[115];
    assign P[95] = in[115] ^ in2[115];
    assign G[96] = in[114] & in2[114];
    assign P[96] = in[114] ^ in2[114];
    assign G[97] = in[113] & in2[113];
    assign P[97] = in[113] ^ in2[113];
    assign G[98] = in[112] & in2[112];
    assign P[98] = in[112] ^ in2[112];
    assign G[99] = in[111] & in2[111];
    assign P[99] = in[111] ^ in2[111];
    assign G[100] = in[110] & in2[110];
    assign P[100] = in[110] ^ in2[110];
    assign G[101] = in[109] & in2[109];
    assign P[101] = in[109] ^ in2[109];
    assign G[102] = in[108] & in2[108];
    assign P[102] = in[108] ^ in2[108];
    assign G[103] = in[107] & in2[107];
    assign P[103] = in[107] ^ in2[107];
    assign G[104] = in[106] & in2[106];
    assign P[104] = in[106] ^ in2[106];
    assign G[105] = in[105] & in2[105];
    assign P[105] = in[105] ^ in2[105];
    assign G[106] = in[104] & in2[104];
    assign P[106] = in[104] ^ in2[104];
    assign G[107] = in[103] & in2[103];
    assign P[107] = in[103] ^ in2[103];
    assign G[108] = in[102] & in2[102];
    assign P[108] = in[102] ^ in2[102];
    assign G[109] = in[101] & in2[101];
    assign P[109] = in[101] ^ in2[101];
    assign G[110] = in[100] & in2[100];
    assign P[110] = in[100] ^ in2[100];
    assign G[111] = in[99] & in2[99];
    assign P[111] = in[99] ^ in2[99];
    assign G[112] = in[98] & in2[98];
    assign P[112] = in[98] ^ in2[98];
    assign G[113] = in[97] & in2[97];
    assign P[113] = in[97] ^ in2[97];
    assign G[114] = in[96] & in2[96];
    assign P[114] = in[96] ^ in2[96];
    assign G[115] = in[95] & in2[95];
    assign P[115] = in[95] ^ in2[95];
    assign G[116] = in[94] & in2[94];
    assign P[116] = in[94] ^ in2[94];
    assign G[117] = in[93] & in2[93];
    assign P[117] = in[93] ^ in2[93];
    assign G[118] = in[92] & in2[92];
    assign P[118] = in[92] ^ in2[92];
    assign G[119] = in[91] & in2[91];
    assign P[119] = in[91] ^ in2[91];
    assign G[120] = in[90] & in2[90];
    assign P[120] = in[90] ^ in2[90];
    assign G[121] = in[89] & in2[89];
    assign P[121] = in[89] ^ in2[89];
    assign G[122] = in[88] & in2[88];
    assign P[122] = in[88] ^ in2[88];
    assign G[123] = in[87] & in2[87];
    assign P[123] = in[87] ^ in2[87];
    assign G[124] = in[86] & in2[86];
    assign P[124] = in[86] ^ in2[86];
    assign G[125] = in[85] & in2[85];
    assign P[125] = in[85] ^ in2[85];
    assign G[126] = in[84] & in2[84];
    assign P[126] = in[84] ^ in2[84];
    assign G[127] = in[83] & in2[83];
    assign P[127] = in[83] ^ in2[83];
    assign G[128] = in[82] & in2[82];
    assign P[128] = in[82] ^ in2[82];
    assign G[129] = in[81] & in2[81];
    assign P[129] = in[81] ^ in2[81];
    assign G[130] = in[80] & in2[80];
    assign P[130] = in[80] ^ in2[80];
    assign G[131] = in[79] & in2[79];
    assign P[131] = in[79] ^ in2[79];
    assign G[132] = in[78] & in2[78];
    assign P[132] = in[78] ^ in2[78];
    assign G[133] = in[77] & in2[77];
    assign P[133] = in[77] ^ in2[77];
    assign G[134] = in[76] & in2[76];
    assign P[134] = in[76] ^ in2[76];
    assign G[135] = in[75] & in2[75];
    assign P[135] = in[75] ^ in2[75];
    assign G[136] = in[74] & in2[74];
    assign P[136] = in[74] ^ in2[74];
    assign G[137] = in[73] & in2[73];
    assign P[137] = in[73] ^ in2[73];
    assign G[138] = in[72] & in2[72];
    assign P[138] = in[72] ^ in2[72];
    assign G[139] = in[71] & in2[71];
    assign P[139] = in[71] ^ in2[71];
    assign G[140] = in[70] & in2[70];
    assign P[140] = in[70] ^ in2[70];
    assign G[141] = in[69] & in2[69];
    assign P[141] = in[69] ^ in2[69];
    assign G[142] = in[68] & in2[68];
    assign P[142] = in[68] ^ in2[68];
    assign G[143] = in[67] & in2[67];
    assign P[143] = in[67] ^ in2[67];
    assign G[144] = in[66] & in2[66];
    assign P[144] = in[66] ^ in2[66];
    assign G[145] = in[65] & in2[65];
    assign P[145] = in[65] ^ in2[65];
    assign G[146] = in[64] & in2[64];
    assign P[146] = in[64] ^ in2[64];
    assign G[147] = in[63] & in2[63];
    assign P[147] = in[63] ^ in2[63];
    assign G[148] = in[62] & in2[62];
    assign P[148] = in[62] ^ in2[62];
    assign G[149] = in[61] & in2[61];
    assign P[149] = in[61] ^ in2[61];
    assign G[150] = in[60] & in2[60];
    assign P[150] = in[60] ^ in2[60];
    assign G[151] = in[59] & in2[59];
    assign P[151] = in[59] ^ in2[59];
    assign G[152] = in[58] & in2[58];
    assign P[152] = in[58] ^ in2[58];
    assign G[153] = in[57] & in2[57];
    assign P[153] = in[57] ^ in2[57];
    assign G[154] = in[56] & in2[56];
    assign P[154] = in[56] ^ in2[56];
    assign G[155] = in[55] & in2[55];
    assign P[155] = in[55] ^ in2[55];
    assign G[156] = in[54] & in2[54];
    assign P[156] = in[54] ^ in2[54];
    assign G[157] = in[53] & in2[53];
    assign P[157] = in[53] ^ in2[53];
    assign G[158] = in[52] & in2[52];
    assign P[158] = in[52] ^ in2[52];
    assign G[159] = in[51] & in2[51];
    assign P[159] = in[51] ^ in2[51];
    assign G[160] = in[50] & in2[50];
    assign P[160] = in[50] ^ in2[50];
    assign G[161] = in[49] & in2[49];
    assign P[161] = in[49] ^ in2[49];
    assign G[162] = in[48] & in2[48];
    assign P[162] = in[48] ^ in2[48];
    assign G[163] = in[47] & in2[47];
    assign P[163] = in[47] ^ in2[47];
    assign G[164] = in[46] & in2[46];
    assign P[164] = in[46] ^ in2[46];
    assign G[165] = in[45] & in2[45];
    assign P[165] = in[45] ^ in2[45];
    assign G[166] = in[44] & in2[44];
    assign P[166] = in[44] ^ in2[44];
    assign G[167] = in[43] & in2[43];
    assign P[167] = in[43] ^ in2[43];
    assign G[168] = in[42] & in2[42];
    assign P[168] = in[42] ^ in2[42];
    assign G[169] = in[41] & in2[41];
    assign P[169] = in[41] ^ in2[41];
    assign G[170] = in[40] & in2[40];
    assign P[170] = in[40] ^ in2[40];
    assign G[171] = in[39] & in2[39];
    assign P[171] = in[39] ^ in2[39];
    assign G[172] = in[38] & in2[38];
    assign P[172] = in[38] ^ in2[38];
    assign G[173] = in[37] & in2[37];
    assign P[173] = in[37] ^ in2[37];
    assign G[174] = in[36] & in2[36];
    assign P[174] = in[36] ^ in2[36];
    assign G[175] = in[35] & in2[35];
    assign P[175] = in[35] ^ in2[35];
    assign G[176] = in[34] & in2[34];
    assign P[176] = in[34] ^ in2[34];
    assign G[177] = in[33] & in2[33];
    assign P[177] = in[33] ^ in2[33];
    assign G[178] = in[32] & in2[32];
    assign P[178] = in[32] ^ in2[32];
    assign G[179] = in[31] & in2[31];
    assign P[179] = in[31] ^ in2[31];
    assign G[180] = in[30] & in2[30];
    assign P[180] = in[30] ^ in2[30];
    assign G[181] = in[29] & in2[29];
    assign P[181] = in[29] ^ in2[29];
    assign G[182] = in[28] & in2[28];
    assign P[182] = in[28] ^ in2[28];
    assign G[183] = in[27] & in2[27];
    assign P[183] = in[27] ^ in2[27];
    assign G[184] = in[26] & in2[26];
    assign P[184] = in[26] ^ in2[26];
    assign G[185] = in[25] & in2[25];
    assign P[185] = in[25] ^ in2[25];
    assign G[186] = in[24] & in2[24];
    assign P[186] = in[24] ^ in2[24];
    assign G[187] = in[23] & in2[23];
    assign P[187] = in[23] ^ in2[23];
    assign G[188] = in[22] & in2[22];
    assign P[188] = in[22] ^ in2[22];
    assign G[189] = in[21] & in2[21];
    assign P[189] = in[21] ^ in2[21];
    assign G[190] = in[20] & in2[20];
    assign P[190] = in[20] ^ in2[20];
    assign G[191] = in[19] & in2[19];
    assign P[191] = in[19] ^ in2[19];
    assign G[192] = in[18] & in2[18];
    assign P[192] = in[18] ^ in2[18];
    assign G[193] = in[17] & in2[17];
    assign P[193] = in[17] ^ in2[17];
    assign G[194] = in[16] & in2[16];
    assign P[194] = in[16] ^ in2[16];
    assign G[195] = in[15] & in2[15];
    assign P[195] = in[15] ^ in2[15];
    assign G[196] = in[14] & in2[14];
    assign P[196] = in[14] ^ in2[14];
    assign G[197] = in[13] & in2[13];
    assign P[197] = in[13] ^ in2[13];
    assign G[198] = in[12] & in2[12];
    assign P[198] = in[12] ^ in2[12];
    assign G[199] = in[11] & in2[11];
    assign P[199] = in[11] ^ in2[11];
    assign G[200] = in[10] & in2[10];
    assign P[200] = in[10] ^ in2[10];
    assign G[201] = in[9] & in2[9];
    assign P[201] = in[9] ^ in2[9];
    assign G[202] = in[8] & in2[8];
    assign P[202] = in[8] ^ in2[8];
    assign G[203] = in[7] & in2[7];
    assign P[203] = in[7] ^ in2[7];
    assign G[204] = in[6] & in2[6];
    assign P[204] = in[6] ^ in2[6];
    assign G[205] = in[5] & in2[5];
    assign P[205] = in[5] ^ in2[5];
    assign G[206] = in[4] & in2[4];
    assign P[206] = in[4] ^ in2[4];
    assign G[207] = in[3] & in2[3];
    assign P[207] = in[3] ^ in2[3];
    assign G[208] = in[2] & in2[2];
    assign P[208] = in[2] ^ in2[2];
    assign G[209] = in[1] & in2[1];
    assign P[209] = in[1] ^ in2[1];
    assign G[210] = in[0] & in2[0];
    assign P[210] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign C[210] = G[209] | (P[209] & C[209]);
    assign cout = G[210] | (P[210] & C[210]);
    assign sum = P ^ C;
endmodule

module CLA210(output [209:0] sum, output cout, input [209:0] in1, input [209:0] in2;

    wire[209:0] G;
    wire[209:0] C;
    wire[209:0] P;

    assign G[0] = in[209] & in2[209];
    assign P[0] = in[209] ^ in2[209];
    assign G[1] = in[208] & in2[208];
    assign P[1] = in[208] ^ in2[208];
    assign G[2] = in[207] & in2[207];
    assign P[2] = in[207] ^ in2[207];
    assign G[3] = in[206] & in2[206];
    assign P[3] = in[206] ^ in2[206];
    assign G[4] = in[205] & in2[205];
    assign P[4] = in[205] ^ in2[205];
    assign G[5] = in[204] & in2[204];
    assign P[5] = in[204] ^ in2[204];
    assign G[6] = in[203] & in2[203];
    assign P[6] = in[203] ^ in2[203];
    assign G[7] = in[202] & in2[202];
    assign P[7] = in[202] ^ in2[202];
    assign G[8] = in[201] & in2[201];
    assign P[8] = in[201] ^ in2[201];
    assign G[9] = in[200] & in2[200];
    assign P[9] = in[200] ^ in2[200];
    assign G[10] = in[199] & in2[199];
    assign P[10] = in[199] ^ in2[199];
    assign G[11] = in[198] & in2[198];
    assign P[11] = in[198] ^ in2[198];
    assign G[12] = in[197] & in2[197];
    assign P[12] = in[197] ^ in2[197];
    assign G[13] = in[196] & in2[196];
    assign P[13] = in[196] ^ in2[196];
    assign G[14] = in[195] & in2[195];
    assign P[14] = in[195] ^ in2[195];
    assign G[15] = in[194] & in2[194];
    assign P[15] = in[194] ^ in2[194];
    assign G[16] = in[193] & in2[193];
    assign P[16] = in[193] ^ in2[193];
    assign G[17] = in[192] & in2[192];
    assign P[17] = in[192] ^ in2[192];
    assign G[18] = in[191] & in2[191];
    assign P[18] = in[191] ^ in2[191];
    assign G[19] = in[190] & in2[190];
    assign P[19] = in[190] ^ in2[190];
    assign G[20] = in[189] & in2[189];
    assign P[20] = in[189] ^ in2[189];
    assign G[21] = in[188] & in2[188];
    assign P[21] = in[188] ^ in2[188];
    assign G[22] = in[187] & in2[187];
    assign P[22] = in[187] ^ in2[187];
    assign G[23] = in[186] & in2[186];
    assign P[23] = in[186] ^ in2[186];
    assign G[24] = in[185] & in2[185];
    assign P[24] = in[185] ^ in2[185];
    assign G[25] = in[184] & in2[184];
    assign P[25] = in[184] ^ in2[184];
    assign G[26] = in[183] & in2[183];
    assign P[26] = in[183] ^ in2[183];
    assign G[27] = in[182] & in2[182];
    assign P[27] = in[182] ^ in2[182];
    assign G[28] = in[181] & in2[181];
    assign P[28] = in[181] ^ in2[181];
    assign G[29] = in[180] & in2[180];
    assign P[29] = in[180] ^ in2[180];
    assign G[30] = in[179] & in2[179];
    assign P[30] = in[179] ^ in2[179];
    assign G[31] = in[178] & in2[178];
    assign P[31] = in[178] ^ in2[178];
    assign G[32] = in[177] & in2[177];
    assign P[32] = in[177] ^ in2[177];
    assign G[33] = in[176] & in2[176];
    assign P[33] = in[176] ^ in2[176];
    assign G[34] = in[175] & in2[175];
    assign P[34] = in[175] ^ in2[175];
    assign G[35] = in[174] & in2[174];
    assign P[35] = in[174] ^ in2[174];
    assign G[36] = in[173] & in2[173];
    assign P[36] = in[173] ^ in2[173];
    assign G[37] = in[172] & in2[172];
    assign P[37] = in[172] ^ in2[172];
    assign G[38] = in[171] & in2[171];
    assign P[38] = in[171] ^ in2[171];
    assign G[39] = in[170] & in2[170];
    assign P[39] = in[170] ^ in2[170];
    assign G[40] = in[169] & in2[169];
    assign P[40] = in[169] ^ in2[169];
    assign G[41] = in[168] & in2[168];
    assign P[41] = in[168] ^ in2[168];
    assign G[42] = in[167] & in2[167];
    assign P[42] = in[167] ^ in2[167];
    assign G[43] = in[166] & in2[166];
    assign P[43] = in[166] ^ in2[166];
    assign G[44] = in[165] & in2[165];
    assign P[44] = in[165] ^ in2[165];
    assign G[45] = in[164] & in2[164];
    assign P[45] = in[164] ^ in2[164];
    assign G[46] = in[163] & in2[163];
    assign P[46] = in[163] ^ in2[163];
    assign G[47] = in[162] & in2[162];
    assign P[47] = in[162] ^ in2[162];
    assign G[48] = in[161] & in2[161];
    assign P[48] = in[161] ^ in2[161];
    assign G[49] = in[160] & in2[160];
    assign P[49] = in[160] ^ in2[160];
    assign G[50] = in[159] & in2[159];
    assign P[50] = in[159] ^ in2[159];
    assign G[51] = in[158] & in2[158];
    assign P[51] = in[158] ^ in2[158];
    assign G[52] = in[157] & in2[157];
    assign P[52] = in[157] ^ in2[157];
    assign G[53] = in[156] & in2[156];
    assign P[53] = in[156] ^ in2[156];
    assign G[54] = in[155] & in2[155];
    assign P[54] = in[155] ^ in2[155];
    assign G[55] = in[154] & in2[154];
    assign P[55] = in[154] ^ in2[154];
    assign G[56] = in[153] & in2[153];
    assign P[56] = in[153] ^ in2[153];
    assign G[57] = in[152] & in2[152];
    assign P[57] = in[152] ^ in2[152];
    assign G[58] = in[151] & in2[151];
    assign P[58] = in[151] ^ in2[151];
    assign G[59] = in[150] & in2[150];
    assign P[59] = in[150] ^ in2[150];
    assign G[60] = in[149] & in2[149];
    assign P[60] = in[149] ^ in2[149];
    assign G[61] = in[148] & in2[148];
    assign P[61] = in[148] ^ in2[148];
    assign G[62] = in[147] & in2[147];
    assign P[62] = in[147] ^ in2[147];
    assign G[63] = in[146] & in2[146];
    assign P[63] = in[146] ^ in2[146];
    assign G[64] = in[145] & in2[145];
    assign P[64] = in[145] ^ in2[145];
    assign G[65] = in[144] & in2[144];
    assign P[65] = in[144] ^ in2[144];
    assign G[66] = in[143] & in2[143];
    assign P[66] = in[143] ^ in2[143];
    assign G[67] = in[142] & in2[142];
    assign P[67] = in[142] ^ in2[142];
    assign G[68] = in[141] & in2[141];
    assign P[68] = in[141] ^ in2[141];
    assign G[69] = in[140] & in2[140];
    assign P[69] = in[140] ^ in2[140];
    assign G[70] = in[139] & in2[139];
    assign P[70] = in[139] ^ in2[139];
    assign G[71] = in[138] & in2[138];
    assign P[71] = in[138] ^ in2[138];
    assign G[72] = in[137] & in2[137];
    assign P[72] = in[137] ^ in2[137];
    assign G[73] = in[136] & in2[136];
    assign P[73] = in[136] ^ in2[136];
    assign G[74] = in[135] & in2[135];
    assign P[74] = in[135] ^ in2[135];
    assign G[75] = in[134] & in2[134];
    assign P[75] = in[134] ^ in2[134];
    assign G[76] = in[133] & in2[133];
    assign P[76] = in[133] ^ in2[133];
    assign G[77] = in[132] & in2[132];
    assign P[77] = in[132] ^ in2[132];
    assign G[78] = in[131] & in2[131];
    assign P[78] = in[131] ^ in2[131];
    assign G[79] = in[130] & in2[130];
    assign P[79] = in[130] ^ in2[130];
    assign G[80] = in[129] & in2[129];
    assign P[80] = in[129] ^ in2[129];
    assign G[81] = in[128] & in2[128];
    assign P[81] = in[128] ^ in2[128];
    assign G[82] = in[127] & in2[127];
    assign P[82] = in[127] ^ in2[127];
    assign G[83] = in[126] & in2[126];
    assign P[83] = in[126] ^ in2[126];
    assign G[84] = in[125] & in2[125];
    assign P[84] = in[125] ^ in2[125];
    assign G[85] = in[124] & in2[124];
    assign P[85] = in[124] ^ in2[124];
    assign G[86] = in[123] & in2[123];
    assign P[86] = in[123] ^ in2[123];
    assign G[87] = in[122] & in2[122];
    assign P[87] = in[122] ^ in2[122];
    assign G[88] = in[121] & in2[121];
    assign P[88] = in[121] ^ in2[121];
    assign G[89] = in[120] & in2[120];
    assign P[89] = in[120] ^ in2[120];
    assign G[90] = in[119] & in2[119];
    assign P[90] = in[119] ^ in2[119];
    assign G[91] = in[118] & in2[118];
    assign P[91] = in[118] ^ in2[118];
    assign G[92] = in[117] & in2[117];
    assign P[92] = in[117] ^ in2[117];
    assign G[93] = in[116] & in2[116];
    assign P[93] = in[116] ^ in2[116];
    assign G[94] = in[115] & in2[115];
    assign P[94] = in[115] ^ in2[115];
    assign G[95] = in[114] & in2[114];
    assign P[95] = in[114] ^ in2[114];
    assign G[96] = in[113] & in2[113];
    assign P[96] = in[113] ^ in2[113];
    assign G[97] = in[112] & in2[112];
    assign P[97] = in[112] ^ in2[112];
    assign G[98] = in[111] & in2[111];
    assign P[98] = in[111] ^ in2[111];
    assign G[99] = in[110] & in2[110];
    assign P[99] = in[110] ^ in2[110];
    assign G[100] = in[109] & in2[109];
    assign P[100] = in[109] ^ in2[109];
    assign G[101] = in[108] & in2[108];
    assign P[101] = in[108] ^ in2[108];
    assign G[102] = in[107] & in2[107];
    assign P[102] = in[107] ^ in2[107];
    assign G[103] = in[106] & in2[106];
    assign P[103] = in[106] ^ in2[106];
    assign G[104] = in[105] & in2[105];
    assign P[104] = in[105] ^ in2[105];
    assign G[105] = in[104] & in2[104];
    assign P[105] = in[104] ^ in2[104];
    assign G[106] = in[103] & in2[103];
    assign P[106] = in[103] ^ in2[103];
    assign G[107] = in[102] & in2[102];
    assign P[107] = in[102] ^ in2[102];
    assign G[108] = in[101] & in2[101];
    assign P[108] = in[101] ^ in2[101];
    assign G[109] = in[100] & in2[100];
    assign P[109] = in[100] ^ in2[100];
    assign G[110] = in[99] & in2[99];
    assign P[110] = in[99] ^ in2[99];
    assign G[111] = in[98] & in2[98];
    assign P[111] = in[98] ^ in2[98];
    assign G[112] = in[97] & in2[97];
    assign P[112] = in[97] ^ in2[97];
    assign G[113] = in[96] & in2[96];
    assign P[113] = in[96] ^ in2[96];
    assign G[114] = in[95] & in2[95];
    assign P[114] = in[95] ^ in2[95];
    assign G[115] = in[94] & in2[94];
    assign P[115] = in[94] ^ in2[94];
    assign G[116] = in[93] & in2[93];
    assign P[116] = in[93] ^ in2[93];
    assign G[117] = in[92] & in2[92];
    assign P[117] = in[92] ^ in2[92];
    assign G[118] = in[91] & in2[91];
    assign P[118] = in[91] ^ in2[91];
    assign G[119] = in[90] & in2[90];
    assign P[119] = in[90] ^ in2[90];
    assign G[120] = in[89] & in2[89];
    assign P[120] = in[89] ^ in2[89];
    assign G[121] = in[88] & in2[88];
    assign P[121] = in[88] ^ in2[88];
    assign G[122] = in[87] & in2[87];
    assign P[122] = in[87] ^ in2[87];
    assign G[123] = in[86] & in2[86];
    assign P[123] = in[86] ^ in2[86];
    assign G[124] = in[85] & in2[85];
    assign P[124] = in[85] ^ in2[85];
    assign G[125] = in[84] & in2[84];
    assign P[125] = in[84] ^ in2[84];
    assign G[126] = in[83] & in2[83];
    assign P[126] = in[83] ^ in2[83];
    assign G[127] = in[82] & in2[82];
    assign P[127] = in[82] ^ in2[82];
    assign G[128] = in[81] & in2[81];
    assign P[128] = in[81] ^ in2[81];
    assign G[129] = in[80] & in2[80];
    assign P[129] = in[80] ^ in2[80];
    assign G[130] = in[79] & in2[79];
    assign P[130] = in[79] ^ in2[79];
    assign G[131] = in[78] & in2[78];
    assign P[131] = in[78] ^ in2[78];
    assign G[132] = in[77] & in2[77];
    assign P[132] = in[77] ^ in2[77];
    assign G[133] = in[76] & in2[76];
    assign P[133] = in[76] ^ in2[76];
    assign G[134] = in[75] & in2[75];
    assign P[134] = in[75] ^ in2[75];
    assign G[135] = in[74] & in2[74];
    assign P[135] = in[74] ^ in2[74];
    assign G[136] = in[73] & in2[73];
    assign P[136] = in[73] ^ in2[73];
    assign G[137] = in[72] & in2[72];
    assign P[137] = in[72] ^ in2[72];
    assign G[138] = in[71] & in2[71];
    assign P[138] = in[71] ^ in2[71];
    assign G[139] = in[70] & in2[70];
    assign P[139] = in[70] ^ in2[70];
    assign G[140] = in[69] & in2[69];
    assign P[140] = in[69] ^ in2[69];
    assign G[141] = in[68] & in2[68];
    assign P[141] = in[68] ^ in2[68];
    assign G[142] = in[67] & in2[67];
    assign P[142] = in[67] ^ in2[67];
    assign G[143] = in[66] & in2[66];
    assign P[143] = in[66] ^ in2[66];
    assign G[144] = in[65] & in2[65];
    assign P[144] = in[65] ^ in2[65];
    assign G[145] = in[64] & in2[64];
    assign P[145] = in[64] ^ in2[64];
    assign G[146] = in[63] & in2[63];
    assign P[146] = in[63] ^ in2[63];
    assign G[147] = in[62] & in2[62];
    assign P[147] = in[62] ^ in2[62];
    assign G[148] = in[61] & in2[61];
    assign P[148] = in[61] ^ in2[61];
    assign G[149] = in[60] & in2[60];
    assign P[149] = in[60] ^ in2[60];
    assign G[150] = in[59] & in2[59];
    assign P[150] = in[59] ^ in2[59];
    assign G[151] = in[58] & in2[58];
    assign P[151] = in[58] ^ in2[58];
    assign G[152] = in[57] & in2[57];
    assign P[152] = in[57] ^ in2[57];
    assign G[153] = in[56] & in2[56];
    assign P[153] = in[56] ^ in2[56];
    assign G[154] = in[55] & in2[55];
    assign P[154] = in[55] ^ in2[55];
    assign G[155] = in[54] & in2[54];
    assign P[155] = in[54] ^ in2[54];
    assign G[156] = in[53] & in2[53];
    assign P[156] = in[53] ^ in2[53];
    assign G[157] = in[52] & in2[52];
    assign P[157] = in[52] ^ in2[52];
    assign G[158] = in[51] & in2[51];
    assign P[158] = in[51] ^ in2[51];
    assign G[159] = in[50] & in2[50];
    assign P[159] = in[50] ^ in2[50];
    assign G[160] = in[49] & in2[49];
    assign P[160] = in[49] ^ in2[49];
    assign G[161] = in[48] & in2[48];
    assign P[161] = in[48] ^ in2[48];
    assign G[162] = in[47] & in2[47];
    assign P[162] = in[47] ^ in2[47];
    assign G[163] = in[46] & in2[46];
    assign P[163] = in[46] ^ in2[46];
    assign G[164] = in[45] & in2[45];
    assign P[164] = in[45] ^ in2[45];
    assign G[165] = in[44] & in2[44];
    assign P[165] = in[44] ^ in2[44];
    assign G[166] = in[43] & in2[43];
    assign P[166] = in[43] ^ in2[43];
    assign G[167] = in[42] & in2[42];
    assign P[167] = in[42] ^ in2[42];
    assign G[168] = in[41] & in2[41];
    assign P[168] = in[41] ^ in2[41];
    assign G[169] = in[40] & in2[40];
    assign P[169] = in[40] ^ in2[40];
    assign G[170] = in[39] & in2[39];
    assign P[170] = in[39] ^ in2[39];
    assign G[171] = in[38] & in2[38];
    assign P[171] = in[38] ^ in2[38];
    assign G[172] = in[37] & in2[37];
    assign P[172] = in[37] ^ in2[37];
    assign G[173] = in[36] & in2[36];
    assign P[173] = in[36] ^ in2[36];
    assign G[174] = in[35] & in2[35];
    assign P[174] = in[35] ^ in2[35];
    assign G[175] = in[34] & in2[34];
    assign P[175] = in[34] ^ in2[34];
    assign G[176] = in[33] & in2[33];
    assign P[176] = in[33] ^ in2[33];
    assign G[177] = in[32] & in2[32];
    assign P[177] = in[32] ^ in2[32];
    assign G[178] = in[31] & in2[31];
    assign P[178] = in[31] ^ in2[31];
    assign G[179] = in[30] & in2[30];
    assign P[179] = in[30] ^ in2[30];
    assign G[180] = in[29] & in2[29];
    assign P[180] = in[29] ^ in2[29];
    assign G[181] = in[28] & in2[28];
    assign P[181] = in[28] ^ in2[28];
    assign G[182] = in[27] & in2[27];
    assign P[182] = in[27] ^ in2[27];
    assign G[183] = in[26] & in2[26];
    assign P[183] = in[26] ^ in2[26];
    assign G[184] = in[25] & in2[25];
    assign P[184] = in[25] ^ in2[25];
    assign G[185] = in[24] & in2[24];
    assign P[185] = in[24] ^ in2[24];
    assign G[186] = in[23] & in2[23];
    assign P[186] = in[23] ^ in2[23];
    assign G[187] = in[22] & in2[22];
    assign P[187] = in[22] ^ in2[22];
    assign G[188] = in[21] & in2[21];
    assign P[188] = in[21] ^ in2[21];
    assign G[189] = in[20] & in2[20];
    assign P[189] = in[20] ^ in2[20];
    assign G[190] = in[19] & in2[19];
    assign P[190] = in[19] ^ in2[19];
    assign G[191] = in[18] & in2[18];
    assign P[191] = in[18] ^ in2[18];
    assign G[192] = in[17] & in2[17];
    assign P[192] = in[17] ^ in2[17];
    assign G[193] = in[16] & in2[16];
    assign P[193] = in[16] ^ in2[16];
    assign G[194] = in[15] & in2[15];
    assign P[194] = in[15] ^ in2[15];
    assign G[195] = in[14] & in2[14];
    assign P[195] = in[14] ^ in2[14];
    assign G[196] = in[13] & in2[13];
    assign P[196] = in[13] ^ in2[13];
    assign G[197] = in[12] & in2[12];
    assign P[197] = in[12] ^ in2[12];
    assign G[198] = in[11] & in2[11];
    assign P[198] = in[11] ^ in2[11];
    assign G[199] = in[10] & in2[10];
    assign P[199] = in[10] ^ in2[10];
    assign G[200] = in[9] & in2[9];
    assign P[200] = in[9] ^ in2[9];
    assign G[201] = in[8] & in2[8];
    assign P[201] = in[8] ^ in2[8];
    assign G[202] = in[7] & in2[7];
    assign P[202] = in[7] ^ in2[7];
    assign G[203] = in[6] & in2[6];
    assign P[203] = in[6] ^ in2[6];
    assign G[204] = in[5] & in2[5];
    assign P[204] = in[5] ^ in2[5];
    assign G[205] = in[4] & in2[4];
    assign P[205] = in[4] ^ in2[4];
    assign G[206] = in[3] & in2[3];
    assign P[206] = in[3] ^ in2[3];
    assign G[207] = in[2] & in2[2];
    assign P[207] = in[2] ^ in2[2];
    assign G[208] = in[1] & in2[1];
    assign P[208] = in[1] ^ in2[1];
    assign G[209] = in[0] & in2[0];
    assign P[209] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign C[209] = G[208] | (P[208] & C[208]);
    assign cout = G[209] | (P[209] & C[209]);
    assign sum = P ^ C;
endmodule

module CLA209(output [208:0] sum, output cout, input [208:0] in1, input [208:0] in2;

    wire[208:0] G;
    wire[208:0] C;
    wire[208:0] P;

    assign G[0] = in[208] & in2[208];
    assign P[0] = in[208] ^ in2[208];
    assign G[1] = in[207] & in2[207];
    assign P[1] = in[207] ^ in2[207];
    assign G[2] = in[206] & in2[206];
    assign P[2] = in[206] ^ in2[206];
    assign G[3] = in[205] & in2[205];
    assign P[3] = in[205] ^ in2[205];
    assign G[4] = in[204] & in2[204];
    assign P[4] = in[204] ^ in2[204];
    assign G[5] = in[203] & in2[203];
    assign P[5] = in[203] ^ in2[203];
    assign G[6] = in[202] & in2[202];
    assign P[6] = in[202] ^ in2[202];
    assign G[7] = in[201] & in2[201];
    assign P[7] = in[201] ^ in2[201];
    assign G[8] = in[200] & in2[200];
    assign P[8] = in[200] ^ in2[200];
    assign G[9] = in[199] & in2[199];
    assign P[9] = in[199] ^ in2[199];
    assign G[10] = in[198] & in2[198];
    assign P[10] = in[198] ^ in2[198];
    assign G[11] = in[197] & in2[197];
    assign P[11] = in[197] ^ in2[197];
    assign G[12] = in[196] & in2[196];
    assign P[12] = in[196] ^ in2[196];
    assign G[13] = in[195] & in2[195];
    assign P[13] = in[195] ^ in2[195];
    assign G[14] = in[194] & in2[194];
    assign P[14] = in[194] ^ in2[194];
    assign G[15] = in[193] & in2[193];
    assign P[15] = in[193] ^ in2[193];
    assign G[16] = in[192] & in2[192];
    assign P[16] = in[192] ^ in2[192];
    assign G[17] = in[191] & in2[191];
    assign P[17] = in[191] ^ in2[191];
    assign G[18] = in[190] & in2[190];
    assign P[18] = in[190] ^ in2[190];
    assign G[19] = in[189] & in2[189];
    assign P[19] = in[189] ^ in2[189];
    assign G[20] = in[188] & in2[188];
    assign P[20] = in[188] ^ in2[188];
    assign G[21] = in[187] & in2[187];
    assign P[21] = in[187] ^ in2[187];
    assign G[22] = in[186] & in2[186];
    assign P[22] = in[186] ^ in2[186];
    assign G[23] = in[185] & in2[185];
    assign P[23] = in[185] ^ in2[185];
    assign G[24] = in[184] & in2[184];
    assign P[24] = in[184] ^ in2[184];
    assign G[25] = in[183] & in2[183];
    assign P[25] = in[183] ^ in2[183];
    assign G[26] = in[182] & in2[182];
    assign P[26] = in[182] ^ in2[182];
    assign G[27] = in[181] & in2[181];
    assign P[27] = in[181] ^ in2[181];
    assign G[28] = in[180] & in2[180];
    assign P[28] = in[180] ^ in2[180];
    assign G[29] = in[179] & in2[179];
    assign P[29] = in[179] ^ in2[179];
    assign G[30] = in[178] & in2[178];
    assign P[30] = in[178] ^ in2[178];
    assign G[31] = in[177] & in2[177];
    assign P[31] = in[177] ^ in2[177];
    assign G[32] = in[176] & in2[176];
    assign P[32] = in[176] ^ in2[176];
    assign G[33] = in[175] & in2[175];
    assign P[33] = in[175] ^ in2[175];
    assign G[34] = in[174] & in2[174];
    assign P[34] = in[174] ^ in2[174];
    assign G[35] = in[173] & in2[173];
    assign P[35] = in[173] ^ in2[173];
    assign G[36] = in[172] & in2[172];
    assign P[36] = in[172] ^ in2[172];
    assign G[37] = in[171] & in2[171];
    assign P[37] = in[171] ^ in2[171];
    assign G[38] = in[170] & in2[170];
    assign P[38] = in[170] ^ in2[170];
    assign G[39] = in[169] & in2[169];
    assign P[39] = in[169] ^ in2[169];
    assign G[40] = in[168] & in2[168];
    assign P[40] = in[168] ^ in2[168];
    assign G[41] = in[167] & in2[167];
    assign P[41] = in[167] ^ in2[167];
    assign G[42] = in[166] & in2[166];
    assign P[42] = in[166] ^ in2[166];
    assign G[43] = in[165] & in2[165];
    assign P[43] = in[165] ^ in2[165];
    assign G[44] = in[164] & in2[164];
    assign P[44] = in[164] ^ in2[164];
    assign G[45] = in[163] & in2[163];
    assign P[45] = in[163] ^ in2[163];
    assign G[46] = in[162] & in2[162];
    assign P[46] = in[162] ^ in2[162];
    assign G[47] = in[161] & in2[161];
    assign P[47] = in[161] ^ in2[161];
    assign G[48] = in[160] & in2[160];
    assign P[48] = in[160] ^ in2[160];
    assign G[49] = in[159] & in2[159];
    assign P[49] = in[159] ^ in2[159];
    assign G[50] = in[158] & in2[158];
    assign P[50] = in[158] ^ in2[158];
    assign G[51] = in[157] & in2[157];
    assign P[51] = in[157] ^ in2[157];
    assign G[52] = in[156] & in2[156];
    assign P[52] = in[156] ^ in2[156];
    assign G[53] = in[155] & in2[155];
    assign P[53] = in[155] ^ in2[155];
    assign G[54] = in[154] & in2[154];
    assign P[54] = in[154] ^ in2[154];
    assign G[55] = in[153] & in2[153];
    assign P[55] = in[153] ^ in2[153];
    assign G[56] = in[152] & in2[152];
    assign P[56] = in[152] ^ in2[152];
    assign G[57] = in[151] & in2[151];
    assign P[57] = in[151] ^ in2[151];
    assign G[58] = in[150] & in2[150];
    assign P[58] = in[150] ^ in2[150];
    assign G[59] = in[149] & in2[149];
    assign P[59] = in[149] ^ in2[149];
    assign G[60] = in[148] & in2[148];
    assign P[60] = in[148] ^ in2[148];
    assign G[61] = in[147] & in2[147];
    assign P[61] = in[147] ^ in2[147];
    assign G[62] = in[146] & in2[146];
    assign P[62] = in[146] ^ in2[146];
    assign G[63] = in[145] & in2[145];
    assign P[63] = in[145] ^ in2[145];
    assign G[64] = in[144] & in2[144];
    assign P[64] = in[144] ^ in2[144];
    assign G[65] = in[143] & in2[143];
    assign P[65] = in[143] ^ in2[143];
    assign G[66] = in[142] & in2[142];
    assign P[66] = in[142] ^ in2[142];
    assign G[67] = in[141] & in2[141];
    assign P[67] = in[141] ^ in2[141];
    assign G[68] = in[140] & in2[140];
    assign P[68] = in[140] ^ in2[140];
    assign G[69] = in[139] & in2[139];
    assign P[69] = in[139] ^ in2[139];
    assign G[70] = in[138] & in2[138];
    assign P[70] = in[138] ^ in2[138];
    assign G[71] = in[137] & in2[137];
    assign P[71] = in[137] ^ in2[137];
    assign G[72] = in[136] & in2[136];
    assign P[72] = in[136] ^ in2[136];
    assign G[73] = in[135] & in2[135];
    assign P[73] = in[135] ^ in2[135];
    assign G[74] = in[134] & in2[134];
    assign P[74] = in[134] ^ in2[134];
    assign G[75] = in[133] & in2[133];
    assign P[75] = in[133] ^ in2[133];
    assign G[76] = in[132] & in2[132];
    assign P[76] = in[132] ^ in2[132];
    assign G[77] = in[131] & in2[131];
    assign P[77] = in[131] ^ in2[131];
    assign G[78] = in[130] & in2[130];
    assign P[78] = in[130] ^ in2[130];
    assign G[79] = in[129] & in2[129];
    assign P[79] = in[129] ^ in2[129];
    assign G[80] = in[128] & in2[128];
    assign P[80] = in[128] ^ in2[128];
    assign G[81] = in[127] & in2[127];
    assign P[81] = in[127] ^ in2[127];
    assign G[82] = in[126] & in2[126];
    assign P[82] = in[126] ^ in2[126];
    assign G[83] = in[125] & in2[125];
    assign P[83] = in[125] ^ in2[125];
    assign G[84] = in[124] & in2[124];
    assign P[84] = in[124] ^ in2[124];
    assign G[85] = in[123] & in2[123];
    assign P[85] = in[123] ^ in2[123];
    assign G[86] = in[122] & in2[122];
    assign P[86] = in[122] ^ in2[122];
    assign G[87] = in[121] & in2[121];
    assign P[87] = in[121] ^ in2[121];
    assign G[88] = in[120] & in2[120];
    assign P[88] = in[120] ^ in2[120];
    assign G[89] = in[119] & in2[119];
    assign P[89] = in[119] ^ in2[119];
    assign G[90] = in[118] & in2[118];
    assign P[90] = in[118] ^ in2[118];
    assign G[91] = in[117] & in2[117];
    assign P[91] = in[117] ^ in2[117];
    assign G[92] = in[116] & in2[116];
    assign P[92] = in[116] ^ in2[116];
    assign G[93] = in[115] & in2[115];
    assign P[93] = in[115] ^ in2[115];
    assign G[94] = in[114] & in2[114];
    assign P[94] = in[114] ^ in2[114];
    assign G[95] = in[113] & in2[113];
    assign P[95] = in[113] ^ in2[113];
    assign G[96] = in[112] & in2[112];
    assign P[96] = in[112] ^ in2[112];
    assign G[97] = in[111] & in2[111];
    assign P[97] = in[111] ^ in2[111];
    assign G[98] = in[110] & in2[110];
    assign P[98] = in[110] ^ in2[110];
    assign G[99] = in[109] & in2[109];
    assign P[99] = in[109] ^ in2[109];
    assign G[100] = in[108] & in2[108];
    assign P[100] = in[108] ^ in2[108];
    assign G[101] = in[107] & in2[107];
    assign P[101] = in[107] ^ in2[107];
    assign G[102] = in[106] & in2[106];
    assign P[102] = in[106] ^ in2[106];
    assign G[103] = in[105] & in2[105];
    assign P[103] = in[105] ^ in2[105];
    assign G[104] = in[104] & in2[104];
    assign P[104] = in[104] ^ in2[104];
    assign G[105] = in[103] & in2[103];
    assign P[105] = in[103] ^ in2[103];
    assign G[106] = in[102] & in2[102];
    assign P[106] = in[102] ^ in2[102];
    assign G[107] = in[101] & in2[101];
    assign P[107] = in[101] ^ in2[101];
    assign G[108] = in[100] & in2[100];
    assign P[108] = in[100] ^ in2[100];
    assign G[109] = in[99] & in2[99];
    assign P[109] = in[99] ^ in2[99];
    assign G[110] = in[98] & in2[98];
    assign P[110] = in[98] ^ in2[98];
    assign G[111] = in[97] & in2[97];
    assign P[111] = in[97] ^ in2[97];
    assign G[112] = in[96] & in2[96];
    assign P[112] = in[96] ^ in2[96];
    assign G[113] = in[95] & in2[95];
    assign P[113] = in[95] ^ in2[95];
    assign G[114] = in[94] & in2[94];
    assign P[114] = in[94] ^ in2[94];
    assign G[115] = in[93] & in2[93];
    assign P[115] = in[93] ^ in2[93];
    assign G[116] = in[92] & in2[92];
    assign P[116] = in[92] ^ in2[92];
    assign G[117] = in[91] & in2[91];
    assign P[117] = in[91] ^ in2[91];
    assign G[118] = in[90] & in2[90];
    assign P[118] = in[90] ^ in2[90];
    assign G[119] = in[89] & in2[89];
    assign P[119] = in[89] ^ in2[89];
    assign G[120] = in[88] & in2[88];
    assign P[120] = in[88] ^ in2[88];
    assign G[121] = in[87] & in2[87];
    assign P[121] = in[87] ^ in2[87];
    assign G[122] = in[86] & in2[86];
    assign P[122] = in[86] ^ in2[86];
    assign G[123] = in[85] & in2[85];
    assign P[123] = in[85] ^ in2[85];
    assign G[124] = in[84] & in2[84];
    assign P[124] = in[84] ^ in2[84];
    assign G[125] = in[83] & in2[83];
    assign P[125] = in[83] ^ in2[83];
    assign G[126] = in[82] & in2[82];
    assign P[126] = in[82] ^ in2[82];
    assign G[127] = in[81] & in2[81];
    assign P[127] = in[81] ^ in2[81];
    assign G[128] = in[80] & in2[80];
    assign P[128] = in[80] ^ in2[80];
    assign G[129] = in[79] & in2[79];
    assign P[129] = in[79] ^ in2[79];
    assign G[130] = in[78] & in2[78];
    assign P[130] = in[78] ^ in2[78];
    assign G[131] = in[77] & in2[77];
    assign P[131] = in[77] ^ in2[77];
    assign G[132] = in[76] & in2[76];
    assign P[132] = in[76] ^ in2[76];
    assign G[133] = in[75] & in2[75];
    assign P[133] = in[75] ^ in2[75];
    assign G[134] = in[74] & in2[74];
    assign P[134] = in[74] ^ in2[74];
    assign G[135] = in[73] & in2[73];
    assign P[135] = in[73] ^ in2[73];
    assign G[136] = in[72] & in2[72];
    assign P[136] = in[72] ^ in2[72];
    assign G[137] = in[71] & in2[71];
    assign P[137] = in[71] ^ in2[71];
    assign G[138] = in[70] & in2[70];
    assign P[138] = in[70] ^ in2[70];
    assign G[139] = in[69] & in2[69];
    assign P[139] = in[69] ^ in2[69];
    assign G[140] = in[68] & in2[68];
    assign P[140] = in[68] ^ in2[68];
    assign G[141] = in[67] & in2[67];
    assign P[141] = in[67] ^ in2[67];
    assign G[142] = in[66] & in2[66];
    assign P[142] = in[66] ^ in2[66];
    assign G[143] = in[65] & in2[65];
    assign P[143] = in[65] ^ in2[65];
    assign G[144] = in[64] & in2[64];
    assign P[144] = in[64] ^ in2[64];
    assign G[145] = in[63] & in2[63];
    assign P[145] = in[63] ^ in2[63];
    assign G[146] = in[62] & in2[62];
    assign P[146] = in[62] ^ in2[62];
    assign G[147] = in[61] & in2[61];
    assign P[147] = in[61] ^ in2[61];
    assign G[148] = in[60] & in2[60];
    assign P[148] = in[60] ^ in2[60];
    assign G[149] = in[59] & in2[59];
    assign P[149] = in[59] ^ in2[59];
    assign G[150] = in[58] & in2[58];
    assign P[150] = in[58] ^ in2[58];
    assign G[151] = in[57] & in2[57];
    assign P[151] = in[57] ^ in2[57];
    assign G[152] = in[56] & in2[56];
    assign P[152] = in[56] ^ in2[56];
    assign G[153] = in[55] & in2[55];
    assign P[153] = in[55] ^ in2[55];
    assign G[154] = in[54] & in2[54];
    assign P[154] = in[54] ^ in2[54];
    assign G[155] = in[53] & in2[53];
    assign P[155] = in[53] ^ in2[53];
    assign G[156] = in[52] & in2[52];
    assign P[156] = in[52] ^ in2[52];
    assign G[157] = in[51] & in2[51];
    assign P[157] = in[51] ^ in2[51];
    assign G[158] = in[50] & in2[50];
    assign P[158] = in[50] ^ in2[50];
    assign G[159] = in[49] & in2[49];
    assign P[159] = in[49] ^ in2[49];
    assign G[160] = in[48] & in2[48];
    assign P[160] = in[48] ^ in2[48];
    assign G[161] = in[47] & in2[47];
    assign P[161] = in[47] ^ in2[47];
    assign G[162] = in[46] & in2[46];
    assign P[162] = in[46] ^ in2[46];
    assign G[163] = in[45] & in2[45];
    assign P[163] = in[45] ^ in2[45];
    assign G[164] = in[44] & in2[44];
    assign P[164] = in[44] ^ in2[44];
    assign G[165] = in[43] & in2[43];
    assign P[165] = in[43] ^ in2[43];
    assign G[166] = in[42] & in2[42];
    assign P[166] = in[42] ^ in2[42];
    assign G[167] = in[41] & in2[41];
    assign P[167] = in[41] ^ in2[41];
    assign G[168] = in[40] & in2[40];
    assign P[168] = in[40] ^ in2[40];
    assign G[169] = in[39] & in2[39];
    assign P[169] = in[39] ^ in2[39];
    assign G[170] = in[38] & in2[38];
    assign P[170] = in[38] ^ in2[38];
    assign G[171] = in[37] & in2[37];
    assign P[171] = in[37] ^ in2[37];
    assign G[172] = in[36] & in2[36];
    assign P[172] = in[36] ^ in2[36];
    assign G[173] = in[35] & in2[35];
    assign P[173] = in[35] ^ in2[35];
    assign G[174] = in[34] & in2[34];
    assign P[174] = in[34] ^ in2[34];
    assign G[175] = in[33] & in2[33];
    assign P[175] = in[33] ^ in2[33];
    assign G[176] = in[32] & in2[32];
    assign P[176] = in[32] ^ in2[32];
    assign G[177] = in[31] & in2[31];
    assign P[177] = in[31] ^ in2[31];
    assign G[178] = in[30] & in2[30];
    assign P[178] = in[30] ^ in2[30];
    assign G[179] = in[29] & in2[29];
    assign P[179] = in[29] ^ in2[29];
    assign G[180] = in[28] & in2[28];
    assign P[180] = in[28] ^ in2[28];
    assign G[181] = in[27] & in2[27];
    assign P[181] = in[27] ^ in2[27];
    assign G[182] = in[26] & in2[26];
    assign P[182] = in[26] ^ in2[26];
    assign G[183] = in[25] & in2[25];
    assign P[183] = in[25] ^ in2[25];
    assign G[184] = in[24] & in2[24];
    assign P[184] = in[24] ^ in2[24];
    assign G[185] = in[23] & in2[23];
    assign P[185] = in[23] ^ in2[23];
    assign G[186] = in[22] & in2[22];
    assign P[186] = in[22] ^ in2[22];
    assign G[187] = in[21] & in2[21];
    assign P[187] = in[21] ^ in2[21];
    assign G[188] = in[20] & in2[20];
    assign P[188] = in[20] ^ in2[20];
    assign G[189] = in[19] & in2[19];
    assign P[189] = in[19] ^ in2[19];
    assign G[190] = in[18] & in2[18];
    assign P[190] = in[18] ^ in2[18];
    assign G[191] = in[17] & in2[17];
    assign P[191] = in[17] ^ in2[17];
    assign G[192] = in[16] & in2[16];
    assign P[192] = in[16] ^ in2[16];
    assign G[193] = in[15] & in2[15];
    assign P[193] = in[15] ^ in2[15];
    assign G[194] = in[14] & in2[14];
    assign P[194] = in[14] ^ in2[14];
    assign G[195] = in[13] & in2[13];
    assign P[195] = in[13] ^ in2[13];
    assign G[196] = in[12] & in2[12];
    assign P[196] = in[12] ^ in2[12];
    assign G[197] = in[11] & in2[11];
    assign P[197] = in[11] ^ in2[11];
    assign G[198] = in[10] & in2[10];
    assign P[198] = in[10] ^ in2[10];
    assign G[199] = in[9] & in2[9];
    assign P[199] = in[9] ^ in2[9];
    assign G[200] = in[8] & in2[8];
    assign P[200] = in[8] ^ in2[8];
    assign G[201] = in[7] & in2[7];
    assign P[201] = in[7] ^ in2[7];
    assign G[202] = in[6] & in2[6];
    assign P[202] = in[6] ^ in2[6];
    assign G[203] = in[5] & in2[5];
    assign P[203] = in[5] ^ in2[5];
    assign G[204] = in[4] & in2[4];
    assign P[204] = in[4] ^ in2[4];
    assign G[205] = in[3] & in2[3];
    assign P[205] = in[3] ^ in2[3];
    assign G[206] = in[2] & in2[2];
    assign P[206] = in[2] ^ in2[2];
    assign G[207] = in[1] & in2[1];
    assign P[207] = in[1] ^ in2[1];
    assign G[208] = in[0] & in2[0];
    assign P[208] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign C[208] = G[207] | (P[207] & C[207]);
    assign cout = G[208] | (P[208] & C[208]);
    assign sum = P ^ C;
endmodule

module CLA208(output [207:0] sum, output cout, input [207:0] in1, input [207:0] in2;

    wire[207:0] G;
    wire[207:0] C;
    wire[207:0] P;

    assign G[0] = in[207] & in2[207];
    assign P[0] = in[207] ^ in2[207];
    assign G[1] = in[206] & in2[206];
    assign P[1] = in[206] ^ in2[206];
    assign G[2] = in[205] & in2[205];
    assign P[2] = in[205] ^ in2[205];
    assign G[3] = in[204] & in2[204];
    assign P[3] = in[204] ^ in2[204];
    assign G[4] = in[203] & in2[203];
    assign P[4] = in[203] ^ in2[203];
    assign G[5] = in[202] & in2[202];
    assign P[5] = in[202] ^ in2[202];
    assign G[6] = in[201] & in2[201];
    assign P[6] = in[201] ^ in2[201];
    assign G[7] = in[200] & in2[200];
    assign P[7] = in[200] ^ in2[200];
    assign G[8] = in[199] & in2[199];
    assign P[8] = in[199] ^ in2[199];
    assign G[9] = in[198] & in2[198];
    assign P[9] = in[198] ^ in2[198];
    assign G[10] = in[197] & in2[197];
    assign P[10] = in[197] ^ in2[197];
    assign G[11] = in[196] & in2[196];
    assign P[11] = in[196] ^ in2[196];
    assign G[12] = in[195] & in2[195];
    assign P[12] = in[195] ^ in2[195];
    assign G[13] = in[194] & in2[194];
    assign P[13] = in[194] ^ in2[194];
    assign G[14] = in[193] & in2[193];
    assign P[14] = in[193] ^ in2[193];
    assign G[15] = in[192] & in2[192];
    assign P[15] = in[192] ^ in2[192];
    assign G[16] = in[191] & in2[191];
    assign P[16] = in[191] ^ in2[191];
    assign G[17] = in[190] & in2[190];
    assign P[17] = in[190] ^ in2[190];
    assign G[18] = in[189] & in2[189];
    assign P[18] = in[189] ^ in2[189];
    assign G[19] = in[188] & in2[188];
    assign P[19] = in[188] ^ in2[188];
    assign G[20] = in[187] & in2[187];
    assign P[20] = in[187] ^ in2[187];
    assign G[21] = in[186] & in2[186];
    assign P[21] = in[186] ^ in2[186];
    assign G[22] = in[185] & in2[185];
    assign P[22] = in[185] ^ in2[185];
    assign G[23] = in[184] & in2[184];
    assign P[23] = in[184] ^ in2[184];
    assign G[24] = in[183] & in2[183];
    assign P[24] = in[183] ^ in2[183];
    assign G[25] = in[182] & in2[182];
    assign P[25] = in[182] ^ in2[182];
    assign G[26] = in[181] & in2[181];
    assign P[26] = in[181] ^ in2[181];
    assign G[27] = in[180] & in2[180];
    assign P[27] = in[180] ^ in2[180];
    assign G[28] = in[179] & in2[179];
    assign P[28] = in[179] ^ in2[179];
    assign G[29] = in[178] & in2[178];
    assign P[29] = in[178] ^ in2[178];
    assign G[30] = in[177] & in2[177];
    assign P[30] = in[177] ^ in2[177];
    assign G[31] = in[176] & in2[176];
    assign P[31] = in[176] ^ in2[176];
    assign G[32] = in[175] & in2[175];
    assign P[32] = in[175] ^ in2[175];
    assign G[33] = in[174] & in2[174];
    assign P[33] = in[174] ^ in2[174];
    assign G[34] = in[173] & in2[173];
    assign P[34] = in[173] ^ in2[173];
    assign G[35] = in[172] & in2[172];
    assign P[35] = in[172] ^ in2[172];
    assign G[36] = in[171] & in2[171];
    assign P[36] = in[171] ^ in2[171];
    assign G[37] = in[170] & in2[170];
    assign P[37] = in[170] ^ in2[170];
    assign G[38] = in[169] & in2[169];
    assign P[38] = in[169] ^ in2[169];
    assign G[39] = in[168] & in2[168];
    assign P[39] = in[168] ^ in2[168];
    assign G[40] = in[167] & in2[167];
    assign P[40] = in[167] ^ in2[167];
    assign G[41] = in[166] & in2[166];
    assign P[41] = in[166] ^ in2[166];
    assign G[42] = in[165] & in2[165];
    assign P[42] = in[165] ^ in2[165];
    assign G[43] = in[164] & in2[164];
    assign P[43] = in[164] ^ in2[164];
    assign G[44] = in[163] & in2[163];
    assign P[44] = in[163] ^ in2[163];
    assign G[45] = in[162] & in2[162];
    assign P[45] = in[162] ^ in2[162];
    assign G[46] = in[161] & in2[161];
    assign P[46] = in[161] ^ in2[161];
    assign G[47] = in[160] & in2[160];
    assign P[47] = in[160] ^ in2[160];
    assign G[48] = in[159] & in2[159];
    assign P[48] = in[159] ^ in2[159];
    assign G[49] = in[158] & in2[158];
    assign P[49] = in[158] ^ in2[158];
    assign G[50] = in[157] & in2[157];
    assign P[50] = in[157] ^ in2[157];
    assign G[51] = in[156] & in2[156];
    assign P[51] = in[156] ^ in2[156];
    assign G[52] = in[155] & in2[155];
    assign P[52] = in[155] ^ in2[155];
    assign G[53] = in[154] & in2[154];
    assign P[53] = in[154] ^ in2[154];
    assign G[54] = in[153] & in2[153];
    assign P[54] = in[153] ^ in2[153];
    assign G[55] = in[152] & in2[152];
    assign P[55] = in[152] ^ in2[152];
    assign G[56] = in[151] & in2[151];
    assign P[56] = in[151] ^ in2[151];
    assign G[57] = in[150] & in2[150];
    assign P[57] = in[150] ^ in2[150];
    assign G[58] = in[149] & in2[149];
    assign P[58] = in[149] ^ in2[149];
    assign G[59] = in[148] & in2[148];
    assign P[59] = in[148] ^ in2[148];
    assign G[60] = in[147] & in2[147];
    assign P[60] = in[147] ^ in2[147];
    assign G[61] = in[146] & in2[146];
    assign P[61] = in[146] ^ in2[146];
    assign G[62] = in[145] & in2[145];
    assign P[62] = in[145] ^ in2[145];
    assign G[63] = in[144] & in2[144];
    assign P[63] = in[144] ^ in2[144];
    assign G[64] = in[143] & in2[143];
    assign P[64] = in[143] ^ in2[143];
    assign G[65] = in[142] & in2[142];
    assign P[65] = in[142] ^ in2[142];
    assign G[66] = in[141] & in2[141];
    assign P[66] = in[141] ^ in2[141];
    assign G[67] = in[140] & in2[140];
    assign P[67] = in[140] ^ in2[140];
    assign G[68] = in[139] & in2[139];
    assign P[68] = in[139] ^ in2[139];
    assign G[69] = in[138] & in2[138];
    assign P[69] = in[138] ^ in2[138];
    assign G[70] = in[137] & in2[137];
    assign P[70] = in[137] ^ in2[137];
    assign G[71] = in[136] & in2[136];
    assign P[71] = in[136] ^ in2[136];
    assign G[72] = in[135] & in2[135];
    assign P[72] = in[135] ^ in2[135];
    assign G[73] = in[134] & in2[134];
    assign P[73] = in[134] ^ in2[134];
    assign G[74] = in[133] & in2[133];
    assign P[74] = in[133] ^ in2[133];
    assign G[75] = in[132] & in2[132];
    assign P[75] = in[132] ^ in2[132];
    assign G[76] = in[131] & in2[131];
    assign P[76] = in[131] ^ in2[131];
    assign G[77] = in[130] & in2[130];
    assign P[77] = in[130] ^ in2[130];
    assign G[78] = in[129] & in2[129];
    assign P[78] = in[129] ^ in2[129];
    assign G[79] = in[128] & in2[128];
    assign P[79] = in[128] ^ in2[128];
    assign G[80] = in[127] & in2[127];
    assign P[80] = in[127] ^ in2[127];
    assign G[81] = in[126] & in2[126];
    assign P[81] = in[126] ^ in2[126];
    assign G[82] = in[125] & in2[125];
    assign P[82] = in[125] ^ in2[125];
    assign G[83] = in[124] & in2[124];
    assign P[83] = in[124] ^ in2[124];
    assign G[84] = in[123] & in2[123];
    assign P[84] = in[123] ^ in2[123];
    assign G[85] = in[122] & in2[122];
    assign P[85] = in[122] ^ in2[122];
    assign G[86] = in[121] & in2[121];
    assign P[86] = in[121] ^ in2[121];
    assign G[87] = in[120] & in2[120];
    assign P[87] = in[120] ^ in2[120];
    assign G[88] = in[119] & in2[119];
    assign P[88] = in[119] ^ in2[119];
    assign G[89] = in[118] & in2[118];
    assign P[89] = in[118] ^ in2[118];
    assign G[90] = in[117] & in2[117];
    assign P[90] = in[117] ^ in2[117];
    assign G[91] = in[116] & in2[116];
    assign P[91] = in[116] ^ in2[116];
    assign G[92] = in[115] & in2[115];
    assign P[92] = in[115] ^ in2[115];
    assign G[93] = in[114] & in2[114];
    assign P[93] = in[114] ^ in2[114];
    assign G[94] = in[113] & in2[113];
    assign P[94] = in[113] ^ in2[113];
    assign G[95] = in[112] & in2[112];
    assign P[95] = in[112] ^ in2[112];
    assign G[96] = in[111] & in2[111];
    assign P[96] = in[111] ^ in2[111];
    assign G[97] = in[110] & in2[110];
    assign P[97] = in[110] ^ in2[110];
    assign G[98] = in[109] & in2[109];
    assign P[98] = in[109] ^ in2[109];
    assign G[99] = in[108] & in2[108];
    assign P[99] = in[108] ^ in2[108];
    assign G[100] = in[107] & in2[107];
    assign P[100] = in[107] ^ in2[107];
    assign G[101] = in[106] & in2[106];
    assign P[101] = in[106] ^ in2[106];
    assign G[102] = in[105] & in2[105];
    assign P[102] = in[105] ^ in2[105];
    assign G[103] = in[104] & in2[104];
    assign P[103] = in[104] ^ in2[104];
    assign G[104] = in[103] & in2[103];
    assign P[104] = in[103] ^ in2[103];
    assign G[105] = in[102] & in2[102];
    assign P[105] = in[102] ^ in2[102];
    assign G[106] = in[101] & in2[101];
    assign P[106] = in[101] ^ in2[101];
    assign G[107] = in[100] & in2[100];
    assign P[107] = in[100] ^ in2[100];
    assign G[108] = in[99] & in2[99];
    assign P[108] = in[99] ^ in2[99];
    assign G[109] = in[98] & in2[98];
    assign P[109] = in[98] ^ in2[98];
    assign G[110] = in[97] & in2[97];
    assign P[110] = in[97] ^ in2[97];
    assign G[111] = in[96] & in2[96];
    assign P[111] = in[96] ^ in2[96];
    assign G[112] = in[95] & in2[95];
    assign P[112] = in[95] ^ in2[95];
    assign G[113] = in[94] & in2[94];
    assign P[113] = in[94] ^ in2[94];
    assign G[114] = in[93] & in2[93];
    assign P[114] = in[93] ^ in2[93];
    assign G[115] = in[92] & in2[92];
    assign P[115] = in[92] ^ in2[92];
    assign G[116] = in[91] & in2[91];
    assign P[116] = in[91] ^ in2[91];
    assign G[117] = in[90] & in2[90];
    assign P[117] = in[90] ^ in2[90];
    assign G[118] = in[89] & in2[89];
    assign P[118] = in[89] ^ in2[89];
    assign G[119] = in[88] & in2[88];
    assign P[119] = in[88] ^ in2[88];
    assign G[120] = in[87] & in2[87];
    assign P[120] = in[87] ^ in2[87];
    assign G[121] = in[86] & in2[86];
    assign P[121] = in[86] ^ in2[86];
    assign G[122] = in[85] & in2[85];
    assign P[122] = in[85] ^ in2[85];
    assign G[123] = in[84] & in2[84];
    assign P[123] = in[84] ^ in2[84];
    assign G[124] = in[83] & in2[83];
    assign P[124] = in[83] ^ in2[83];
    assign G[125] = in[82] & in2[82];
    assign P[125] = in[82] ^ in2[82];
    assign G[126] = in[81] & in2[81];
    assign P[126] = in[81] ^ in2[81];
    assign G[127] = in[80] & in2[80];
    assign P[127] = in[80] ^ in2[80];
    assign G[128] = in[79] & in2[79];
    assign P[128] = in[79] ^ in2[79];
    assign G[129] = in[78] & in2[78];
    assign P[129] = in[78] ^ in2[78];
    assign G[130] = in[77] & in2[77];
    assign P[130] = in[77] ^ in2[77];
    assign G[131] = in[76] & in2[76];
    assign P[131] = in[76] ^ in2[76];
    assign G[132] = in[75] & in2[75];
    assign P[132] = in[75] ^ in2[75];
    assign G[133] = in[74] & in2[74];
    assign P[133] = in[74] ^ in2[74];
    assign G[134] = in[73] & in2[73];
    assign P[134] = in[73] ^ in2[73];
    assign G[135] = in[72] & in2[72];
    assign P[135] = in[72] ^ in2[72];
    assign G[136] = in[71] & in2[71];
    assign P[136] = in[71] ^ in2[71];
    assign G[137] = in[70] & in2[70];
    assign P[137] = in[70] ^ in2[70];
    assign G[138] = in[69] & in2[69];
    assign P[138] = in[69] ^ in2[69];
    assign G[139] = in[68] & in2[68];
    assign P[139] = in[68] ^ in2[68];
    assign G[140] = in[67] & in2[67];
    assign P[140] = in[67] ^ in2[67];
    assign G[141] = in[66] & in2[66];
    assign P[141] = in[66] ^ in2[66];
    assign G[142] = in[65] & in2[65];
    assign P[142] = in[65] ^ in2[65];
    assign G[143] = in[64] & in2[64];
    assign P[143] = in[64] ^ in2[64];
    assign G[144] = in[63] & in2[63];
    assign P[144] = in[63] ^ in2[63];
    assign G[145] = in[62] & in2[62];
    assign P[145] = in[62] ^ in2[62];
    assign G[146] = in[61] & in2[61];
    assign P[146] = in[61] ^ in2[61];
    assign G[147] = in[60] & in2[60];
    assign P[147] = in[60] ^ in2[60];
    assign G[148] = in[59] & in2[59];
    assign P[148] = in[59] ^ in2[59];
    assign G[149] = in[58] & in2[58];
    assign P[149] = in[58] ^ in2[58];
    assign G[150] = in[57] & in2[57];
    assign P[150] = in[57] ^ in2[57];
    assign G[151] = in[56] & in2[56];
    assign P[151] = in[56] ^ in2[56];
    assign G[152] = in[55] & in2[55];
    assign P[152] = in[55] ^ in2[55];
    assign G[153] = in[54] & in2[54];
    assign P[153] = in[54] ^ in2[54];
    assign G[154] = in[53] & in2[53];
    assign P[154] = in[53] ^ in2[53];
    assign G[155] = in[52] & in2[52];
    assign P[155] = in[52] ^ in2[52];
    assign G[156] = in[51] & in2[51];
    assign P[156] = in[51] ^ in2[51];
    assign G[157] = in[50] & in2[50];
    assign P[157] = in[50] ^ in2[50];
    assign G[158] = in[49] & in2[49];
    assign P[158] = in[49] ^ in2[49];
    assign G[159] = in[48] & in2[48];
    assign P[159] = in[48] ^ in2[48];
    assign G[160] = in[47] & in2[47];
    assign P[160] = in[47] ^ in2[47];
    assign G[161] = in[46] & in2[46];
    assign P[161] = in[46] ^ in2[46];
    assign G[162] = in[45] & in2[45];
    assign P[162] = in[45] ^ in2[45];
    assign G[163] = in[44] & in2[44];
    assign P[163] = in[44] ^ in2[44];
    assign G[164] = in[43] & in2[43];
    assign P[164] = in[43] ^ in2[43];
    assign G[165] = in[42] & in2[42];
    assign P[165] = in[42] ^ in2[42];
    assign G[166] = in[41] & in2[41];
    assign P[166] = in[41] ^ in2[41];
    assign G[167] = in[40] & in2[40];
    assign P[167] = in[40] ^ in2[40];
    assign G[168] = in[39] & in2[39];
    assign P[168] = in[39] ^ in2[39];
    assign G[169] = in[38] & in2[38];
    assign P[169] = in[38] ^ in2[38];
    assign G[170] = in[37] & in2[37];
    assign P[170] = in[37] ^ in2[37];
    assign G[171] = in[36] & in2[36];
    assign P[171] = in[36] ^ in2[36];
    assign G[172] = in[35] & in2[35];
    assign P[172] = in[35] ^ in2[35];
    assign G[173] = in[34] & in2[34];
    assign P[173] = in[34] ^ in2[34];
    assign G[174] = in[33] & in2[33];
    assign P[174] = in[33] ^ in2[33];
    assign G[175] = in[32] & in2[32];
    assign P[175] = in[32] ^ in2[32];
    assign G[176] = in[31] & in2[31];
    assign P[176] = in[31] ^ in2[31];
    assign G[177] = in[30] & in2[30];
    assign P[177] = in[30] ^ in2[30];
    assign G[178] = in[29] & in2[29];
    assign P[178] = in[29] ^ in2[29];
    assign G[179] = in[28] & in2[28];
    assign P[179] = in[28] ^ in2[28];
    assign G[180] = in[27] & in2[27];
    assign P[180] = in[27] ^ in2[27];
    assign G[181] = in[26] & in2[26];
    assign P[181] = in[26] ^ in2[26];
    assign G[182] = in[25] & in2[25];
    assign P[182] = in[25] ^ in2[25];
    assign G[183] = in[24] & in2[24];
    assign P[183] = in[24] ^ in2[24];
    assign G[184] = in[23] & in2[23];
    assign P[184] = in[23] ^ in2[23];
    assign G[185] = in[22] & in2[22];
    assign P[185] = in[22] ^ in2[22];
    assign G[186] = in[21] & in2[21];
    assign P[186] = in[21] ^ in2[21];
    assign G[187] = in[20] & in2[20];
    assign P[187] = in[20] ^ in2[20];
    assign G[188] = in[19] & in2[19];
    assign P[188] = in[19] ^ in2[19];
    assign G[189] = in[18] & in2[18];
    assign P[189] = in[18] ^ in2[18];
    assign G[190] = in[17] & in2[17];
    assign P[190] = in[17] ^ in2[17];
    assign G[191] = in[16] & in2[16];
    assign P[191] = in[16] ^ in2[16];
    assign G[192] = in[15] & in2[15];
    assign P[192] = in[15] ^ in2[15];
    assign G[193] = in[14] & in2[14];
    assign P[193] = in[14] ^ in2[14];
    assign G[194] = in[13] & in2[13];
    assign P[194] = in[13] ^ in2[13];
    assign G[195] = in[12] & in2[12];
    assign P[195] = in[12] ^ in2[12];
    assign G[196] = in[11] & in2[11];
    assign P[196] = in[11] ^ in2[11];
    assign G[197] = in[10] & in2[10];
    assign P[197] = in[10] ^ in2[10];
    assign G[198] = in[9] & in2[9];
    assign P[198] = in[9] ^ in2[9];
    assign G[199] = in[8] & in2[8];
    assign P[199] = in[8] ^ in2[8];
    assign G[200] = in[7] & in2[7];
    assign P[200] = in[7] ^ in2[7];
    assign G[201] = in[6] & in2[6];
    assign P[201] = in[6] ^ in2[6];
    assign G[202] = in[5] & in2[5];
    assign P[202] = in[5] ^ in2[5];
    assign G[203] = in[4] & in2[4];
    assign P[203] = in[4] ^ in2[4];
    assign G[204] = in[3] & in2[3];
    assign P[204] = in[3] ^ in2[3];
    assign G[205] = in[2] & in2[2];
    assign P[205] = in[2] ^ in2[2];
    assign G[206] = in[1] & in2[1];
    assign P[206] = in[1] ^ in2[1];
    assign G[207] = in[0] & in2[0];
    assign P[207] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign C[207] = G[206] | (P[206] & C[206]);
    assign cout = G[207] | (P[207] & C[207]);
    assign sum = P ^ C;
endmodule

module CLA207(output [206:0] sum, output cout, input [206:0] in1, input [206:0] in2;

    wire[206:0] G;
    wire[206:0] C;
    wire[206:0] P;

    assign G[0] = in[206] & in2[206];
    assign P[0] = in[206] ^ in2[206];
    assign G[1] = in[205] & in2[205];
    assign P[1] = in[205] ^ in2[205];
    assign G[2] = in[204] & in2[204];
    assign P[2] = in[204] ^ in2[204];
    assign G[3] = in[203] & in2[203];
    assign P[3] = in[203] ^ in2[203];
    assign G[4] = in[202] & in2[202];
    assign P[4] = in[202] ^ in2[202];
    assign G[5] = in[201] & in2[201];
    assign P[5] = in[201] ^ in2[201];
    assign G[6] = in[200] & in2[200];
    assign P[6] = in[200] ^ in2[200];
    assign G[7] = in[199] & in2[199];
    assign P[7] = in[199] ^ in2[199];
    assign G[8] = in[198] & in2[198];
    assign P[8] = in[198] ^ in2[198];
    assign G[9] = in[197] & in2[197];
    assign P[9] = in[197] ^ in2[197];
    assign G[10] = in[196] & in2[196];
    assign P[10] = in[196] ^ in2[196];
    assign G[11] = in[195] & in2[195];
    assign P[11] = in[195] ^ in2[195];
    assign G[12] = in[194] & in2[194];
    assign P[12] = in[194] ^ in2[194];
    assign G[13] = in[193] & in2[193];
    assign P[13] = in[193] ^ in2[193];
    assign G[14] = in[192] & in2[192];
    assign P[14] = in[192] ^ in2[192];
    assign G[15] = in[191] & in2[191];
    assign P[15] = in[191] ^ in2[191];
    assign G[16] = in[190] & in2[190];
    assign P[16] = in[190] ^ in2[190];
    assign G[17] = in[189] & in2[189];
    assign P[17] = in[189] ^ in2[189];
    assign G[18] = in[188] & in2[188];
    assign P[18] = in[188] ^ in2[188];
    assign G[19] = in[187] & in2[187];
    assign P[19] = in[187] ^ in2[187];
    assign G[20] = in[186] & in2[186];
    assign P[20] = in[186] ^ in2[186];
    assign G[21] = in[185] & in2[185];
    assign P[21] = in[185] ^ in2[185];
    assign G[22] = in[184] & in2[184];
    assign P[22] = in[184] ^ in2[184];
    assign G[23] = in[183] & in2[183];
    assign P[23] = in[183] ^ in2[183];
    assign G[24] = in[182] & in2[182];
    assign P[24] = in[182] ^ in2[182];
    assign G[25] = in[181] & in2[181];
    assign P[25] = in[181] ^ in2[181];
    assign G[26] = in[180] & in2[180];
    assign P[26] = in[180] ^ in2[180];
    assign G[27] = in[179] & in2[179];
    assign P[27] = in[179] ^ in2[179];
    assign G[28] = in[178] & in2[178];
    assign P[28] = in[178] ^ in2[178];
    assign G[29] = in[177] & in2[177];
    assign P[29] = in[177] ^ in2[177];
    assign G[30] = in[176] & in2[176];
    assign P[30] = in[176] ^ in2[176];
    assign G[31] = in[175] & in2[175];
    assign P[31] = in[175] ^ in2[175];
    assign G[32] = in[174] & in2[174];
    assign P[32] = in[174] ^ in2[174];
    assign G[33] = in[173] & in2[173];
    assign P[33] = in[173] ^ in2[173];
    assign G[34] = in[172] & in2[172];
    assign P[34] = in[172] ^ in2[172];
    assign G[35] = in[171] & in2[171];
    assign P[35] = in[171] ^ in2[171];
    assign G[36] = in[170] & in2[170];
    assign P[36] = in[170] ^ in2[170];
    assign G[37] = in[169] & in2[169];
    assign P[37] = in[169] ^ in2[169];
    assign G[38] = in[168] & in2[168];
    assign P[38] = in[168] ^ in2[168];
    assign G[39] = in[167] & in2[167];
    assign P[39] = in[167] ^ in2[167];
    assign G[40] = in[166] & in2[166];
    assign P[40] = in[166] ^ in2[166];
    assign G[41] = in[165] & in2[165];
    assign P[41] = in[165] ^ in2[165];
    assign G[42] = in[164] & in2[164];
    assign P[42] = in[164] ^ in2[164];
    assign G[43] = in[163] & in2[163];
    assign P[43] = in[163] ^ in2[163];
    assign G[44] = in[162] & in2[162];
    assign P[44] = in[162] ^ in2[162];
    assign G[45] = in[161] & in2[161];
    assign P[45] = in[161] ^ in2[161];
    assign G[46] = in[160] & in2[160];
    assign P[46] = in[160] ^ in2[160];
    assign G[47] = in[159] & in2[159];
    assign P[47] = in[159] ^ in2[159];
    assign G[48] = in[158] & in2[158];
    assign P[48] = in[158] ^ in2[158];
    assign G[49] = in[157] & in2[157];
    assign P[49] = in[157] ^ in2[157];
    assign G[50] = in[156] & in2[156];
    assign P[50] = in[156] ^ in2[156];
    assign G[51] = in[155] & in2[155];
    assign P[51] = in[155] ^ in2[155];
    assign G[52] = in[154] & in2[154];
    assign P[52] = in[154] ^ in2[154];
    assign G[53] = in[153] & in2[153];
    assign P[53] = in[153] ^ in2[153];
    assign G[54] = in[152] & in2[152];
    assign P[54] = in[152] ^ in2[152];
    assign G[55] = in[151] & in2[151];
    assign P[55] = in[151] ^ in2[151];
    assign G[56] = in[150] & in2[150];
    assign P[56] = in[150] ^ in2[150];
    assign G[57] = in[149] & in2[149];
    assign P[57] = in[149] ^ in2[149];
    assign G[58] = in[148] & in2[148];
    assign P[58] = in[148] ^ in2[148];
    assign G[59] = in[147] & in2[147];
    assign P[59] = in[147] ^ in2[147];
    assign G[60] = in[146] & in2[146];
    assign P[60] = in[146] ^ in2[146];
    assign G[61] = in[145] & in2[145];
    assign P[61] = in[145] ^ in2[145];
    assign G[62] = in[144] & in2[144];
    assign P[62] = in[144] ^ in2[144];
    assign G[63] = in[143] & in2[143];
    assign P[63] = in[143] ^ in2[143];
    assign G[64] = in[142] & in2[142];
    assign P[64] = in[142] ^ in2[142];
    assign G[65] = in[141] & in2[141];
    assign P[65] = in[141] ^ in2[141];
    assign G[66] = in[140] & in2[140];
    assign P[66] = in[140] ^ in2[140];
    assign G[67] = in[139] & in2[139];
    assign P[67] = in[139] ^ in2[139];
    assign G[68] = in[138] & in2[138];
    assign P[68] = in[138] ^ in2[138];
    assign G[69] = in[137] & in2[137];
    assign P[69] = in[137] ^ in2[137];
    assign G[70] = in[136] & in2[136];
    assign P[70] = in[136] ^ in2[136];
    assign G[71] = in[135] & in2[135];
    assign P[71] = in[135] ^ in2[135];
    assign G[72] = in[134] & in2[134];
    assign P[72] = in[134] ^ in2[134];
    assign G[73] = in[133] & in2[133];
    assign P[73] = in[133] ^ in2[133];
    assign G[74] = in[132] & in2[132];
    assign P[74] = in[132] ^ in2[132];
    assign G[75] = in[131] & in2[131];
    assign P[75] = in[131] ^ in2[131];
    assign G[76] = in[130] & in2[130];
    assign P[76] = in[130] ^ in2[130];
    assign G[77] = in[129] & in2[129];
    assign P[77] = in[129] ^ in2[129];
    assign G[78] = in[128] & in2[128];
    assign P[78] = in[128] ^ in2[128];
    assign G[79] = in[127] & in2[127];
    assign P[79] = in[127] ^ in2[127];
    assign G[80] = in[126] & in2[126];
    assign P[80] = in[126] ^ in2[126];
    assign G[81] = in[125] & in2[125];
    assign P[81] = in[125] ^ in2[125];
    assign G[82] = in[124] & in2[124];
    assign P[82] = in[124] ^ in2[124];
    assign G[83] = in[123] & in2[123];
    assign P[83] = in[123] ^ in2[123];
    assign G[84] = in[122] & in2[122];
    assign P[84] = in[122] ^ in2[122];
    assign G[85] = in[121] & in2[121];
    assign P[85] = in[121] ^ in2[121];
    assign G[86] = in[120] & in2[120];
    assign P[86] = in[120] ^ in2[120];
    assign G[87] = in[119] & in2[119];
    assign P[87] = in[119] ^ in2[119];
    assign G[88] = in[118] & in2[118];
    assign P[88] = in[118] ^ in2[118];
    assign G[89] = in[117] & in2[117];
    assign P[89] = in[117] ^ in2[117];
    assign G[90] = in[116] & in2[116];
    assign P[90] = in[116] ^ in2[116];
    assign G[91] = in[115] & in2[115];
    assign P[91] = in[115] ^ in2[115];
    assign G[92] = in[114] & in2[114];
    assign P[92] = in[114] ^ in2[114];
    assign G[93] = in[113] & in2[113];
    assign P[93] = in[113] ^ in2[113];
    assign G[94] = in[112] & in2[112];
    assign P[94] = in[112] ^ in2[112];
    assign G[95] = in[111] & in2[111];
    assign P[95] = in[111] ^ in2[111];
    assign G[96] = in[110] & in2[110];
    assign P[96] = in[110] ^ in2[110];
    assign G[97] = in[109] & in2[109];
    assign P[97] = in[109] ^ in2[109];
    assign G[98] = in[108] & in2[108];
    assign P[98] = in[108] ^ in2[108];
    assign G[99] = in[107] & in2[107];
    assign P[99] = in[107] ^ in2[107];
    assign G[100] = in[106] & in2[106];
    assign P[100] = in[106] ^ in2[106];
    assign G[101] = in[105] & in2[105];
    assign P[101] = in[105] ^ in2[105];
    assign G[102] = in[104] & in2[104];
    assign P[102] = in[104] ^ in2[104];
    assign G[103] = in[103] & in2[103];
    assign P[103] = in[103] ^ in2[103];
    assign G[104] = in[102] & in2[102];
    assign P[104] = in[102] ^ in2[102];
    assign G[105] = in[101] & in2[101];
    assign P[105] = in[101] ^ in2[101];
    assign G[106] = in[100] & in2[100];
    assign P[106] = in[100] ^ in2[100];
    assign G[107] = in[99] & in2[99];
    assign P[107] = in[99] ^ in2[99];
    assign G[108] = in[98] & in2[98];
    assign P[108] = in[98] ^ in2[98];
    assign G[109] = in[97] & in2[97];
    assign P[109] = in[97] ^ in2[97];
    assign G[110] = in[96] & in2[96];
    assign P[110] = in[96] ^ in2[96];
    assign G[111] = in[95] & in2[95];
    assign P[111] = in[95] ^ in2[95];
    assign G[112] = in[94] & in2[94];
    assign P[112] = in[94] ^ in2[94];
    assign G[113] = in[93] & in2[93];
    assign P[113] = in[93] ^ in2[93];
    assign G[114] = in[92] & in2[92];
    assign P[114] = in[92] ^ in2[92];
    assign G[115] = in[91] & in2[91];
    assign P[115] = in[91] ^ in2[91];
    assign G[116] = in[90] & in2[90];
    assign P[116] = in[90] ^ in2[90];
    assign G[117] = in[89] & in2[89];
    assign P[117] = in[89] ^ in2[89];
    assign G[118] = in[88] & in2[88];
    assign P[118] = in[88] ^ in2[88];
    assign G[119] = in[87] & in2[87];
    assign P[119] = in[87] ^ in2[87];
    assign G[120] = in[86] & in2[86];
    assign P[120] = in[86] ^ in2[86];
    assign G[121] = in[85] & in2[85];
    assign P[121] = in[85] ^ in2[85];
    assign G[122] = in[84] & in2[84];
    assign P[122] = in[84] ^ in2[84];
    assign G[123] = in[83] & in2[83];
    assign P[123] = in[83] ^ in2[83];
    assign G[124] = in[82] & in2[82];
    assign P[124] = in[82] ^ in2[82];
    assign G[125] = in[81] & in2[81];
    assign P[125] = in[81] ^ in2[81];
    assign G[126] = in[80] & in2[80];
    assign P[126] = in[80] ^ in2[80];
    assign G[127] = in[79] & in2[79];
    assign P[127] = in[79] ^ in2[79];
    assign G[128] = in[78] & in2[78];
    assign P[128] = in[78] ^ in2[78];
    assign G[129] = in[77] & in2[77];
    assign P[129] = in[77] ^ in2[77];
    assign G[130] = in[76] & in2[76];
    assign P[130] = in[76] ^ in2[76];
    assign G[131] = in[75] & in2[75];
    assign P[131] = in[75] ^ in2[75];
    assign G[132] = in[74] & in2[74];
    assign P[132] = in[74] ^ in2[74];
    assign G[133] = in[73] & in2[73];
    assign P[133] = in[73] ^ in2[73];
    assign G[134] = in[72] & in2[72];
    assign P[134] = in[72] ^ in2[72];
    assign G[135] = in[71] & in2[71];
    assign P[135] = in[71] ^ in2[71];
    assign G[136] = in[70] & in2[70];
    assign P[136] = in[70] ^ in2[70];
    assign G[137] = in[69] & in2[69];
    assign P[137] = in[69] ^ in2[69];
    assign G[138] = in[68] & in2[68];
    assign P[138] = in[68] ^ in2[68];
    assign G[139] = in[67] & in2[67];
    assign P[139] = in[67] ^ in2[67];
    assign G[140] = in[66] & in2[66];
    assign P[140] = in[66] ^ in2[66];
    assign G[141] = in[65] & in2[65];
    assign P[141] = in[65] ^ in2[65];
    assign G[142] = in[64] & in2[64];
    assign P[142] = in[64] ^ in2[64];
    assign G[143] = in[63] & in2[63];
    assign P[143] = in[63] ^ in2[63];
    assign G[144] = in[62] & in2[62];
    assign P[144] = in[62] ^ in2[62];
    assign G[145] = in[61] & in2[61];
    assign P[145] = in[61] ^ in2[61];
    assign G[146] = in[60] & in2[60];
    assign P[146] = in[60] ^ in2[60];
    assign G[147] = in[59] & in2[59];
    assign P[147] = in[59] ^ in2[59];
    assign G[148] = in[58] & in2[58];
    assign P[148] = in[58] ^ in2[58];
    assign G[149] = in[57] & in2[57];
    assign P[149] = in[57] ^ in2[57];
    assign G[150] = in[56] & in2[56];
    assign P[150] = in[56] ^ in2[56];
    assign G[151] = in[55] & in2[55];
    assign P[151] = in[55] ^ in2[55];
    assign G[152] = in[54] & in2[54];
    assign P[152] = in[54] ^ in2[54];
    assign G[153] = in[53] & in2[53];
    assign P[153] = in[53] ^ in2[53];
    assign G[154] = in[52] & in2[52];
    assign P[154] = in[52] ^ in2[52];
    assign G[155] = in[51] & in2[51];
    assign P[155] = in[51] ^ in2[51];
    assign G[156] = in[50] & in2[50];
    assign P[156] = in[50] ^ in2[50];
    assign G[157] = in[49] & in2[49];
    assign P[157] = in[49] ^ in2[49];
    assign G[158] = in[48] & in2[48];
    assign P[158] = in[48] ^ in2[48];
    assign G[159] = in[47] & in2[47];
    assign P[159] = in[47] ^ in2[47];
    assign G[160] = in[46] & in2[46];
    assign P[160] = in[46] ^ in2[46];
    assign G[161] = in[45] & in2[45];
    assign P[161] = in[45] ^ in2[45];
    assign G[162] = in[44] & in2[44];
    assign P[162] = in[44] ^ in2[44];
    assign G[163] = in[43] & in2[43];
    assign P[163] = in[43] ^ in2[43];
    assign G[164] = in[42] & in2[42];
    assign P[164] = in[42] ^ in2[42];
    assign G[165] = in[41] & in2[41];
    assign P[165] = in[41] ^ in2[41];
    assign G[166] = in[40] & in2[40];
    assign P[166] = in[40] ^ in2[40];
    assign G[167] = in[39] & in2[39];
    assign P[167] = in[39] ^ in2[39];
    assign G[168] = in[38] & in2[38];
    assign P[168] = in[38] ^ in2[38];
    assign G[169] = in[37] & in2[37];
    assign P[169] = in[37] ^ in2[37];
    assign G[170] = in[36] & in2[36];
    assign P[170] = in[36] ^ in2[36];
    assign G[171] = in[35] & in2[35];
    assign P[171] = in[35] ^ in2[35];
    assign G[172] = in[34] & in2[34];
    assign P[172] = in[34] ^ in2[34];
    assign G[173] = in[33] & in2[33];
    assign P[173] = in[33] ^ in2[33];
    assign G[174] = in[32] & in2[32];
    assign P[174] = in[32] ^ in2[32];
    assign G[175] = in[31] & in2[31];
    assign P[175] = in[31] ^ in2[31];
    assign G[176] = in[30] & in2[30];
    assign P[176] = in[30] ^ in2[30];
    assign G[177] = in[29] & in2[29];
    assign P[177] = in[29] ^ in2[29];
    assign G[178] = in[28] & in2[28];
    assign P[178] = in[28] ^ in2[28];
    assign G[179] = in[27] & in2[27];
    assign P[179] = in[27] ^ in2[27];
    assign G[180] = in[26] & in2[26];
    assign P[180] = in[26] ^ in2[26];
    assign G[181] = in[25] & in2[25];
    assign P[181] = in[25] ^ in2[25];
    assign G[182] = in[24] & in2[24];
    assign P[182] = in[24] ^ in2[24];
    assign G[183] = in[23] & in2[23];
    assign P[183] = in[23] ^ in2[23];
    assign G[184] = in[22] & in2[22];
    assign P[184] = in[22] ^ in2[22];
    assign G[185] = in[21] & in2[21];
    assign P[185] = in[21] ^ in2[21];
    assign G[186] = in[20] & in2[20];
    assign P[186] = in[20] ^ in2[20];
    assign G[187] = in[19] & in2[19];
    assign P[187] = in[19] ^ in2[19];
    assign G[188] = in[18] & in2[18];
    assign P[188] = in[18] ^ in2[18];
    assign G[189] = in[17] & in2[17];
    assign P[189] = in[17] ^ in2[17];
    assign G[190] = in[16] & in2[16];
    assign P[190] = in[16] ^ in2[16];
    assign G[191] = in[15] & in2[15];
    assign P[191] = in[15] ^ in2[15];
    assign G[192] = in[14] & in2[14];
    assign P[192] = in[14] ^ in2[14];
    assign G[193] = in[13] & in2[13];
    assign P[193] = in[13] ^ in2[13];
    assign G[194] = in[12] & in2[12];
    assign P[194] = in[12] ^ in2[12];
    assign G[195] = in[11] & in2[11];
    assign P[195] = in[11] ^ in2[11];
    assign G[196] = in[10] & in2[10];
    assign P[196] = in[10] ^ in2[10];
    assign G[197] = in[9] & in2[9];
    assign P[197] = in[9] ^ in2[9];
    assign G[198] = in[8] & in2[8];
    assign P[198] = in[8] ^ in2[8];
    assign G[199] = in[7] & in2[7];
    assign P[199] = in[7] ^ in2[7];
    assign G[200] = in[6] & in2[6];
    assign P[200] = in[6] ^ in2[6];
    assign G[201] = in[5] & in2[5];
    assign P[201] = in[5] ^ in2[5];
    assign G[202] = in[4] & in2[4];
    assign P[202] = in[4] ^ in2[4];
    assign G[203] = in[3] & in2[3];
    assign P[203] = in[3] ^ in2[3];
    assign G[204] = in[2] & in2[2];
    assign P[204] = in[2] ^ in2[2];
    assign G[205] = in[1] & in2[1];
    assign P[205] = in[1] ^ in2[1];
    assign G[206] = in[0] & in2[0];
    assign P[206] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign C[206] = G[205] | (P[205] & C[205]);
    assign cout = G[206] | (P[206] & C[206]);
    assign sum = P ^ C;
endmodule

module CLA206(output [205:0] sum, output cout, input [205:0] in1, input [205:0] in2;

    wire[205:0] G;
    wire[205:0] C;
    wire[205:0] P;

    assign G[0] = in[205] & in2[205];
    assign P[0] = in[205] ^ in2[205];
    assign G[1] = in[204] & in2[204];
    assign P[1] = in[204] ^ in2[204];
    assign G[2] = in[203] & in2[203];
    assign P[2] = in[203] ^ in2[203];
    assign G[3] = in[202] & in2[202];
    assign P[3] = in[202] ^ in2[202];
    assign G[4] = in[201] & in2[201];
    assign P[4] = in[201] ^ in2[201];
    assign G[5] = in[200] & in2[200];
    assign P[5] = in[200] ^ in2[200];
    assign G[6] = in[199] & in2[199];
    assign P[6] = in[199] ^ in2[199];
    assign G[7] = in[198] & in2[198];
    assign P[7] = in[198] ^ in2[198];
    assign G[8] = in[197] & in2[197];
    assign P[8] = in[197] ^ in2[197];
    assign G[9] = in[196] & in2[196];
    assign P[9] = in[196] ^ in2[196];
    assign G[10] = in[195] & in2[195];
    assign P[10] = in[195] ^ in2[195];
    assign G[11] = in[194] & in2[194];
    assign P[11] = in[194] ^ in2[194];
    assign G[12] = in[193] & in2[193];
    assign P[12] = in[193] ^ in2[193];
    assign G[13] = in[192] & in2[192];
    assign P[13] = in[192] ^ in2[192];
    assign G[14] = in[191] & in2[191];
    assign P[14] = in[191] ^ in2[191];
    assign G[15] = in[190] & in2[190];
    assign P[15] = in[190] ^ in2[190];
    assign G[16] = in[189] & in2[189];
    assign P[16] = in[189] ^ in2[189];
    assign G[17] = in[188] & in2[188];
    assign P[17] = in[188] ^ in2[188];
    assign G[18] = in[187] & in2[187];
    assign P[18] = in[187] ^ in2[187];
    assign G[19] = in[186] & in2[186];
    assign P[19] = in[186] ^ in2[186];
    assign G[20] = in[185] & in2[185];
    assign P[20] = in[185] ^ in2[185];
    assign G[21] = in[184] & in2[184];
    assign P[21] = in[184] ^ in2[184];
    assign G[22] = in[183] & in2[183];
    assign P[22] = in[183] ^ in2[183];
    assign G[23] = in[182] & in2[182];
    assign P[23] = in[182] ^ in2[182];
    assign G[24] = in[181] & in2[181];
    assign P[24] = in[181] ^ in2[181];
    assign G[25] = in[180] & in2[180];
    assign P[25] = in[180] ^ in2[180];
    assign G[26] = in[179] & in2[179];
    assign P[26] = in[179] ^ in2[179];
    assign G[27] = in[178] & in2[178];
    assign P[27] = in[178] ^ in2[178];
    assign G[28] = in[177] & in2[177];
    assign P[28] = in[177] ^ in2[177];
    assign G[29] = in[176] & in2[176];
    assign P[29] = in[176] ^ in2[176];
    assign G[30] = in[175] & in2[175];
    assign P[30] = in[175] ^ in2[175];
    assign G[31] = in[174] & in2[174];
    assign P[31] = in[174] ^ in2[174];
    assign G[32] = in[173] & in2[173];
    assign P[32] = in[173] ^ in2[173];
    assign G[33] = in[172] & in2[172];
    assign P[33] = in[172] ^ in2[172];
    assign G[34] = in[171] & in2[171];
    assign P[34] = in[171] ^ in2[171];
    assign G[35] = in[170] & in2[170];
    assign P[35] = in[170] ^ in2[170];
    assign G[36] = in[169] & in2[169];
    assign P[36] = in[169] ^ in2[169];
    assign G[37] = in[168] & in2[168];
    assign P[37] = in[168] ^ in2[168];
    assign G[38] = in[167] & in2[167];
    assign P[38] = in[167] ^ in2[167];
    assign G[39] = in[166] & in2[166];
    assign P[39] = in[166] ^ in2[166];
    assign G[40] = in[165] & in2[165];
    assign P[40] = in[165] ^ in2[165];
    assign G[41] = in[164] & in2[164];
    assign P[41] = in[164] ^ in2[164];
    assign G[42] = in[163] & in2[163];
    assign P[42] = in[163] ^ in2[163];
    assign G[43] = in[162] & in2[162];
    assign P[43] = in[162] ^ in2[162];
    assign G[44] = in[161] & in2[161];
    assign P[44] = in[161] ^ in2[161];
    assign G[45] = in[160] & in2[160];
    assign P[45] = in[160] ^ in2[160];
    assign G[46] = in[159] & in2[159];
    assign P[46] = in[159] ^ in2[159];
    assign G[47] = in[158] & in2[158];
    assign P[47] = in[158] ^ in2[158];
    assign G[48] = in[157] & in2[157];
    assign P[48] = in[157] ^ in2[157];
    assign G[49] = in[156] & in2[156];
    assign P[49] = in[156] ^ in2[156];
    assign G[50] = in[155] & in2[155];
    assign P[50] = in[155] ^ in2[155];
    assign G[51] = in[154] & in2[154];
    assign P[51] = in[154] ^ in2[154];
    assign G[52] = in[153] & in2[153];
    assign P[52] = in[153] ^ in2[153];
    assign G[53] = in[152] & in2[152];
    assign P[53] = in[152] ^ in2[152];
    assign G[54] = in[151] & in2[151];
    assign P[54] = in[151] ^ in2[151];
    assign G[55] = in[150] & in2[150];
    assign P[55] = in[150] ^ in2[150];
    assign G[56] = in[149] & in2[149];
    assign P[56] = in[149] ^ in2[149];
    assign G[57] = in[148] & in2[148];
    assign P[57] = in[148] ^ in2[148];
    assign G[58] = in[147] & in2[147];
    assign P[58] = in[147] ^ in2[147];
    assign G[59] = in[146] & in2[146];
    assign P[59] = in[146] ^ in2[146];
    assign G[60] = in[145] & in2[145];
    assign P[60] = in[145] ^ in2[145];
    assign G[61] = in[144] & in2[144];
    assign P[61] = in[144] ^ in2[144];
    assign G[62] = in[143] & in2[143];
    assign P[62] = in[143] ^ in2[143];
    assign G[63] = in[142] & in2[142];
    assign P[63] = in[142] ^ in2[142];
    assign G[64] = in[141] & in2[141];
    assign P[64] = in[141] ^ in2[141];
    assign G[65] = in[140] & in2[140];
    assign P[65] = in[140] ^ in2[140];
    assign G[66] = in[139] & in2[139];
    assign P[66] = in[139] ^ in2[139];
    assign G[67] = in[138] & in2[138];
    assign P[67] = in[138] ^ in2[138];
    assign G[68] = in[137] & in2[137];
    assign P[68] = in[137] ^ in2[137];
    assign G[69] = in[136] & in2[136];
    assign P[69] = in[136] ^ in2[136];
    assign G[70] = in[135] & in2[135];
    assign P[70] = in[135] ^ in2[135];
    assign G[71] = in[134] & in2[134];
    assign P[71] = in[134] ^ in2[134];
    assign G[72] = in[133] & in2[133];
    assign P[72] = in[133] ^ in2[133];
    assign G[73] = in[132] & in2[132];
    assign P[73] = in[132] ^ in2[132];
    assign G[74] = in[131] & in2[131];
    assign P[74] = in[131] ^ in2[131];
    assign G[75] = in[130] & in2[130];
    assign P[75] = in[130] ^ in2[130];
    assign G[76] = in[129] & in2[129];
    assign P[76] = in[129] ^ in2[129];
    assign G[77] = in[128] & in2[128];
    assign P[77] = in[128] ^ in2[128];
    assign G[78] = in[127] & in2[127];
    assign P[78] = in[127] ^ in2[127];
    assign G[79] = in[126] & in2[126];
    assign P[79] = in[126] ^ in2[126];
    assign G[80] = in[125] & in2[125];
    assign P[80] = in[125] ^ in2[125];
    assign G[81] = in[124] & in2[124];
    assign P[81] = in[124] ^ in2[124];
    assign G[82] = in[123] & in2[123];
    assign P[82] = in[123] ^ in2[123];
    assign G[83] = in[122] & in2[122];
    assign P[83] = in[122] ^ in2[122];
    assign G[84] = in[121] & in2[121];
    assign P[84] = in[121] ^ in2[121];
    assign G[85] = in[120] & in2[120];
    assign P[85] = in[120] ^ in2[120];
    assign G[86] = in[119] & in2[119];
    assign P[86] = in[119] ^ in2[119];
    assign G[87] = in[118] & in2[118];
    assign P[87] = in[118] ^ in2[118];
    assign G[88] = in[117] & in2[117];
    assign P[88] = in[117] ^ in2[117];
    assign G[89] = in[116] & in2[116];
    assign P[89] = in[116] ^ in2[116];
    assign G[90] = in[115] & in2[115];
    assign P[90] = in[115] ^ in2[115];
    assign G[91] = in[114] & in2[114];
    assign P[91] = in[114] ^ in2[114];
    assign G[92] = in[113] & in2[113];
    assign P[92] = in[113] ^ in2[113];
    assign G[93] = in[112] & in2[112];
    assign P[93] = in[112] ^ in2[112];
    assign G[94] = in[111] & in2[111];
    assign P[94] = in[111] ^ in2[111];
    assign G[95] = in[110] & in2[110];
    assign P[95] = in[110] ^ in2[110];
    assign G[96] = in[109] & in2[109];
    assign P[96] = in[109] ^ in2[109];
    assign G[97] = in[108] & in2[108];
    assign P[97] = in[108] ^ in2[108];
    assign G[98] = in[107] & in2[107];
    assign P[98] = in[107] ^ in2[107];
    assign G[99] = in[106] & in2[106];
    assign P[99] = in[106] ^ in2[106];
    assign G[100] = in[105] & in2[105];
    assign P[100] = in[105] ^ in2[105];
    assign G[101] = in[104] & in2[104];
    assign P[101] = in[104] ^ in2[104];
    assign G[102] = in[103] & in2[103];
    assign P[102] = in[103] ^ in2[103];
    assign G[103] = in[102] & in2[102];
    assign P[103] = in[102] ^ in2[102];
    assign G[104] = in[101] & in2[101];
    assign P[104] = in[101] ^ in2[101];
    assign G[105] = in[100] & in2[100];
    assign P[105] = in[100] ^ in2[100];
    assign G[106] = in[99] & in2[99];
    assign P[106] = in[99] ^ in2[99];
    assign G[107] = in[98] & in2[98];
    assign P[107] = in[98] ^ in2[98];
    assign G[108] = in[97] & in2[97];
    assign P[108] = in[97] ^ in2[97];
    assign G[109] = in[96] & in2[96];
    assign P[109] = in[96] ^ in2[96];
    assign G[110] = in[95] & in2[95];
    assign P[110] = in[95] ^ in2[95];
    assign G[111] = in[94] & in2[94];
    assign P[111] = in[94] ^ in2[94];
    assign G[112] = in[93] & in2[93];
    assign P[112] = in[93] ^ in2[93];
    assign G[113] = in[92] & in2[92];
    assign P[113] = in[92] ^ in2[92];
    assign G[114] = in[91] & in2[91];
    assign P[114] = in[91] ^ in2[91];
    assign G[115] = in[90] & in2[90];
    assign P[115] = in[90] ^ in2[90];
    assign G[116] = in[89] & in2[89];
    assign P[116] = in[89] ^ in2[89];
    assign G[117] = in[88] & in2[88];
    assign P[117] = in[88] ^ in2[88];
    assign G[118] = in[87] & in2[87];
    assign P[118] = in[87] ^ in2[87];
    assign G[119] = in[86] & in2[86];
    assign P[119] = in[86] ^ in2[86];
    assign G[120] = in[85] & in2[85];
    assign P[120] = in[85] ^ in2[85];
    assign G[121] = in[84] & in2[84];
    assign P[121] = in[84] ^ in2[84];
    assign G[122] = in[83] & in2[83];
    assign P[122] = in[83] ^ in2[83];
    assign G[123] = in[82] & in2[82];
    assign P[123] = in[82] ^ in2[82];
    assign G[124] = in[81] & in2[81];
    assign P[124] = in[81] ^ in2[81];
    assign G[125] = in[80] & in2[80];
    assign P[125] = in[80] ^ in2[80];
    assign G[126] = in[79] & in2[79];
    assign P[126] = in[79] ^ in2[79];
    assign G[127] = in[78] & in2[78];
    assign P[127] = in[78] ^ in2[78];
    assign G[128] = in[77] & in2[77];
    assign P[128] = in[77] ^ in2[77];
    assign G[129] = in[76] & in2[76];
    assign P[129] = in[76] ^ in2[76];
    assign G[130] = in[75] & in2[75];
    assign P[130] = in[75] ^ in2[75];
    assign G[131] = in[74] & in2[74];
    assign P[131] = in[74] ^ in2[74];
    assign G[132] = in[73] & in2[73];
    assign P[132] = in[73] ^ in2[73];
    assign G[133] = in[72] & in2[72];
    assign P[133] = in[72] ^ in2[72];
    assign G[134] = in[71] & in2[71];
    assign P[134] = in[71] ^ in2[71];
    assign G[135] = in[70] & in2[70];
    assign P[135] = in[70] ^ in2[70];
    assign G[136] = in[69] & in2[69];
    assign P[136] = in[69] ^ in2[69];
    assign G[137] = in[68] & in2[68];
    assign P[137] = in[68] ^ in2[68];
    assign G[138] = in[67] & in2[67];
    assign P[138] = in[67] ^ in2[67];
    assign G[139] = in[66] & in2[66];
    assign P[139] = in[66] ^ in2[66];
    assign G[140] = in[65] & in2[65];
    assign P[140] = in[65] ^ in2[65];
    assign G[141] = in[64] & in2[64];
    assign P[141] = in[64] ^ in2[64];
    assign G[142] = in[63] & in2[63];
    assign P[142] = in[63] ^ in2[63];
    assign G[143] = in[62] & in2[62];
    assign P[143] = in[62] ^ in2[62];
    assign G[144] = in[61] & in2[61];
    assign P[144] = in[61] ^ in2[61];
    assign G[145] = in[60] & in2[60];
    assign P[145] = in[60] ^ in2[60];
    assign G[146] = in[59] & in2[59];
    assign P[146] = in[59] ^ in2[59];
    assign G[147] = in[58] & in2[58];
    assign P[147] = in[58] ^ in2[58];
    assign G[148] = in[57] & in2[57];
    assign P[148] = in[57] ^ in2[57];
    assign G[149] = in[56] & in2[56];
    assign P[149] = in[56] ^ in2[56];
    assign G[150] = in[55] & in2[55];
    assign P[150] = in[55] ^ in2[55];
    assign G[151] = in[54] & in2[54];
    assign P[151] = in[54] ^ in2[54];
    assign G[152] = in[53] & in2[53];
    assign P[152] = in[53] ^ in2[53];
    assign G[153] = in[52] & in2[52];
    assign P[153] = in[52] ^ in2[52];
    assign G[154] = in[51] & in2[51];
    assign P[154] = in[51] ^ in2[51];
    assign G[155] = in[50] & in2[50];
    assign P[155] = in[50] ^ in2[50];
    assign G[156] = in[49] & in2[49];
    assign P[156] = in[49] ^ in2[49];
    assign G[157] = in[48] & in2[48];
    assign P[157] = in[48] ^ in2[48];
    assign G[158] = in[47] & in2[47];
    assign P[158] = in[47] ^ in2[47];
    assign G[159] = in[46] & in2[46];
    assign P[159] = in[46] ^ in2[46];
    assign G[160] = in[45] & in2[45];
    assign P[160] = in[45] ^ in2[45];
    assign G[161] = in[44] & in2[44];
    assign P[161] = in[44] ^ in2[44];
    assign G[162] = in[43] & in2[43];
    assign P[162] = in[43] ^ in2[43];
    assign G[163] = in[42] & in2[42];
    assign P[163] = in[42] ^ in2[42];
    assign G[164] = in[41] & in2[41];
    assign P[164] = in[41] ^ in2[41];
    assign G[165] = in[40] & in2[40];
    assign P[165] = in[40] ^ in2[40];
    assign G[166] = in[39] & in2[39];
    assign P[166] = in[39] ^ in2[39];
    assign G[167] = in[38] & in2[38];
    assign P[167] = in[38] ^ in2[38];
    assign G[168] = in[37] & in2[37];
    assign P[168] = in[37] ^ in2[37];
    assign G[169] = in[36] & in2[36];
    assign P[169] = in[36] ^ in2[36];
    assign G[170] = in[35] & in2[35];
    assign P[170] = in[35] ^ in2[35];
    assign G[171] = in[34] & in2[34];
    assign P[171] = in[34] ^ in2[34];
    assign G[172] = in[33] & in2[33];
    assign P[172] = in[33] ^ in2[33];
    assign G[173] = in[32] & in2[32];
    assign P[173] = in[32] ^ in2[32];
    assign G[174] = in[31] & in2[31];
    assign P[174] = in[31] ^ in2[31];
    assign G[175] = in[30] & in2[30];
    assign P[175] = in[30] ^ in2[30];
    assign G[176] = in[29] & in2[29];
    assign P[176] = in[29] ^ in2[29];
    assign G[177] = in[28] & in2[28];
    assign P[177] = in[28] ^ in2[28];
    assign G[178] = in[27] & in2[27];
    assign P[178] = in[27] ^ in2[27];
    assign G[179] = in[26] & in2[26];
    assign P[179] = in[26] ^ in2[26];
    assign G[180] = in[25] & in2[25];
    assign P[180] = in[25] ^ in2[25];
    assign G[181] = in[24] & in2[24];
    assign P[181] = in[24] ^ in2[24];
    assign G[182] = in[23] & in2[23];
    assign P[182] = in[23] ^ in2[23];
    assign G[183] = in[22] & in2[22];
    assign P[183] = in[22] ^ in2[22];
    assign G[184] = in[21] & in2[21];
    assign P[184] = in[21] ^ in2[21];
    assign G[185] = in[20] & in2[20];
    assign P[185] = in[20] ^ in2[20];
    assign G[186] = in[19] & in2[19];
    assign P[186] = in[19] ^ in2[19];
    assign G[187] = in[18] & in2[18];
    assign P[187] = in[18] ^ in2[18];
    assign G[188] = in[17] & in2[17];
    assign P[188] = in[17] ^ in2[17];
    assign G[189] = in[16] & in2[16];
    assign P[189] = in[16] ^ in2[16];
    assign G[190] = in[15] & in2[15];
    assign P[190] = in[15] ^ in2[15];
    assign G[191] = in[14] & in2[14];
    assign P[191] = in[14] ^ in2[14];
    assign G[192] = in[13] & in2[13];
    assign P[192] = in[13] ^ in2[13];
    assign G[193] = in[12] & in2[12];
    assign P[193] = in[12] ^ in2[12];
    assign G[194] = in[11] & in2[11];
    assign P[194] = in[11] ^ in2[11];
    assign G[195] = in[10] & in2[10];
    assign P[195] = in[10] ^ in2[10];
    assign G[196] = in[9] & in2[9];
    assign P[196] = in[9] ^ in2[9];
    assign G[197] = in[8] & in2[8];
    assign P[197] = in[8] ^ in2[8];
    assign G[198] = in[7] & in2[7];
    assign P[198] = in[7] ^ in2[7];
    assign G[199] = in[6] & in2[6];
    assign P[199] = in[6] ^ in2[6];
    assign G[200] = in[5] & in2[5];
    assign P[200] = in[5] ^ in2[5];
    assign G[201] = in[4] & in2[4];
    assign P[201] = in[4] ^ in2[4];
    assign G[202] = in[3] & in2[3];
    assign P[202] = in[3] ^ in2[3];
    assign G[203] = in[2] & in2[2];
    assign P[203] = in[2] ^ in2[2];
    assign G[204] = in[1] & in2[1];
    assign P[204] = in[1] ^ in2[1];
    assign G[205] = in[0] & in2[0];
    assign P[205] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign C[205] = G[204] | (P[204] & C[204]);
    assign cout = G[205] | (P[205] & C[205]);
    assign sum = P ^ C;
endmodule

module CLA205(output [204:0] sum, output cout, input [204:0] in1, input [204:0] in2;

    wire[204:0] G;
    wire[204:0] C;
    wire[204:0] P;

    assign G[0] = in[204] & in2[204];
    assign P[0] = in[204] ^ in2[204];
    assign G[1] = in[203] & in2[203];
    assign P[1] = in[203] ^ in2[203];
    assign G[2] = in[202] & in2[202];
    assign P[2] = in[202] ^ in2[202];
    assign G[3] = in[201] & in2[201];
    assign P[3] = in[201] ^ in2[201];
    assign G[4] = in[200] & in2[200];
    assign P[4] = in[200] ^ in2[200];
    assign G[5] = in[199] & in2[199];
    assign P[5] = in[199] ^ in2[199];
    assign G[6] = in[198] & in2[198];
    assign P[6] = in[198] ^ in2[198];
    assign G[7] = in[197] & in2[197];
    assign P[7] = in[197] ^ in2[197];
    assign G[8] = in[196] & in2[196];
    assign P[8] = in[196] ^ in2[196];
    assign G[9] = in[195] & in2[195];
    assign P[9] = in[195] ^ in2[195];
    assign G[10] = in[194] & in2[194];
    assign P[10] = in[194] ^ in2[194];
    assign G[11] = in[193] & in2[193];
    assign P[11] = in[193] ^ in2[193];
    assign G[12] = in[192] & in2[192];
    assign P[12] = in[192] ^ in2[192];
    assign G[13] = in[191] & in2[191];
    assign P[13] = in[191] ^ in2[191];
    assign G[14] = in[190] & in2[190];
    assign P[14] = in[190] ^ in2[190];
    assign G[15] = in[189] & in2[189];
    assign P[15] = in[189] ^ in2[189];
    assign G[16] = in[188] & in2[188];
    assign P[16] = in[188] ^ in2[188];
    assign G[17] = in[187] & in2[187];
    assign P[17] = in[187] ^ in2[187];
    assign G[18] = in[186] & in2[186];
    assign P[18] = in[186] ^ in2[186];
    assign G[19] = in[185] & in2[185];
    assign P[19] = in[185] ^ in2[185];
    assign G[20] = in[184] & in2[184];
    assign P[20] = in[184] ^ in2[184];
    assign G[21] = in[183] & in2[183];
    assign P[21] = in[183] ^ in2[183];
    assign G[22] = in[182] & in2[182];
    assign P[22] = in[182] ^ in2[182];
    assign G[23] = in[181] & in2[181];
    assign P[23] = in[181] ^ in2[181];
    assign G[24] = in[180] & in2[180];
    assign P[24] = in[180] ^ in2[180];
    assign G[25] = in[179] & in2[179];
    assign P[25] = in[179] ^ in2[179];
    assign G[26] = in[178] & in2[178];
    assign P[26] = in[178] ^ in2[178];
    assign G[27] = in[177] & in2[177];
    assign P[27] = in[177] ^ in2[177];
    assign G[28] = in[176] & in2[176];
    assign P[28] = in[176] ^ in2[176];
    assign G[29] = in[175] & in2[175];
    assign P[29] = in[175] ^ in2[175];
    assign G[30] = in[174] & in2[174];
    assign P[30] = in[174] ^ in2[174];
    assign G[31] = in[173] & in2[173];
    assign P[31] = in[173] ^ in2[173];
    assign G[32] = in[172] & in2[172];
    assign P[32] = in[172] ^ in2[172];
    assign G[33] = in[171] & in2[171];
    assign P[33] = in[171] ^ in2[171];
    assign G[34] = in[170] & in2[170];
    assign P[34] = in[170] ^ in2[170];
    assign G[35] = in[169] & in2[169];
    assign P[35] = in[169] ^ in2[169];
    assign G[36] = in[168] & in2[168];
    assign P[36] = in[168] ^ in2[168];
    assign G[37] = in[167] & in2[167];
    assign P[37] = in[167] ^ in2[167];
    assign G[38] = in[166] & in2[166];
    assign P[38] = in[166] ^ in2[166];
    assign G[39] = in[165] & in2[165];
    assign P[39] = in[165] ^ in2[165];
    assign G[40] = in[164] & in2[164];
    assign P[40] = in[164] ^ in2[164];
    assign G[41] = in[163] & in2[163];
    assign P[41] = in[163] ^ in2[163];
    assign G[42] = in[162] & in2[162];
    assign P[42] = in[162] ^ in2[162];
    assign G[43] = in[161] & in2[161];
    assign P[43] = in[161] ^ in2[161];
    assign G[44] = in[160] & in2[160];
    assign P[44] = in[160] ^ in2[160];
    assign G[45] = in[159] & in2[159];
    assign P[45] = in[159] ^ in2[159];
    assign G[46] = in[158] & in2[158];
    assign P[46] = in[158] ^ in2[158];
    assign G[47] = in[157] & in2[157];
    assign P[47] = in[157] ^ in2[157];
    assign G[48] = in[156] & in2[156];
    assign P[48] = in[156] ^ in2[156];
    assign G[49] = in[155] & in2[155];
    assign P[49] = in[155] ^ in2[155];
    assign G[50] = in[154] & in2[154];
    assign P[50] = in[154] ^ in2[154];
    assign G[51] = in[153] & in2[153];
    assign P[51] = in[153] ^ in2[153];
    assign G[52] = in[152] & in2[152];
    assign P[52] = in[152] ^ in2[152];
    assign G[53] = in[151] & in2[151];
    assign P[53] = in[151] ^ in2[151];
    assign G[54] = in[150] & in2[150];
    assign P[54] = in[150] ^ in2[150];
    assign G[55] = in[149] & in2[149];
    assign P[55] = in[149] ^ in2[149];
    assign G[56] = in[148] & in2[148];
    assign P[56] = in[148] ^ in2[148];
    assign G[57] = in[147] & in2[147];
    assign P[57] = in[147] ^ in2[147];
    assign G[58] = in[146] & in2[146];
    assign P[58] = in[146] ^ in2[146];
    assign G[59] = in[145] & in2[145];
    assign P[59] = in[145] ^ in2[145];
    assign G[60] = in[144] & in2[144];
    assign P[60] = in[144] ^ in2[144];
    assign G[61] = in[143] & in2[143];
    assign P[61] = in[143] ^ in2[143];
    assign G[62] = in[142] & in2[142];
    assign P[62] = in[142] ^ in2[142];
    assign G[63] = in[141] & in2[141];
    assign P[63] = in[141] ^ in2[141];
    assign G[64] = in[140] & in2[140];
    assign P[64] = in[140] ^ in2[140];
    assign G[65] = in[139] & in2[139];
    assign P[65] = in[139] ^ in2[139];
    assign G[66] = in[138] & in2[138];
    assign P[66] = in[138] ^ in2[138];
    assign G[67] = in[137] & in2[137];
    assign P[67] = in[137] ^ in2[137];
    assign G[68] = in[136] & in2[136];
    assign P[68] = in[136] ^ in2[136];
    assign G[69] = in[135] & in2[135];
    assign P[69] = in[135] ^ in2[135];
    assign G[70] = in[134] & in2[134];
    assign P[70] = in[134] ^ in2[134];
    assign G[71] = in[133] & in2[133];
    assign P[71] = in[133] ^ in2[133];
    assign G[72] = in[132] & in2[132];
    assign P[72] = in[132] ^ in2[132];
    assign G[73] = in[131] & in2[131];
    assign P[73] = in[131] ^ in2[131];
    assign G[74] = in[130] & in2[130];
    assign P[74] = in[130] ^ in2[130];
    assign G[75] = in[129] & in2[129];
    assign P[75] = in[129] ^ in2[129];
    assign G[76] = in[128] & in2[128];
    assign P[76] = in[128] ^ in2[128];
    assign G[77] = in[127] & in2[127];
    assign P[77] = in[127] ^ in2[127];
    assign G[78] = in[126] & in2[126];
    assign P[78] = in[126] ^ in2[126];
    assign G[79] = in[125] & in2[125];
    assign P[79] = in[125] ^ in2[125];
    assign G[80] = in[124] & in2[124];
    assign P[80] = in[124] ^ in2[124];
    assign G[81] = in[123] & in2[123];
    assign P[81] = in[123] ^ in2[123];
    assign G[82] = in[122] & in2[122];
    assign P[82] = in[122] ^ in2[122];
    assign G[83] = in[121] & in2[121];
    assign P[83] = in[121] ^ in2[121];
    assign G[84] = in[120] & in2[120];
    assign P[84] = in[120] ^ in2[120];
    assign G[85] = in[119] & in2[119];
    assign P[85] = in[119] ^ in2[119];
    assign G[86] = in[118] & in2[118];
    assign P[86] = in[118] ^ in2[118];
    assign G[87] = in[117] & in2[117];
    assign P[87] = in[117] ^ in2[117];
    assign G[88] = in[116] & in2[116];
    assign P[88] = in[116] ^ in2[116];
    assign G[89] = in[115] & in2[115];
    assign P[89] = in[115] ^ in2[115];
    assign G[90] = in[114] & in2[114];
    assign P[90] = in[114] ^ in2[114];
    assign G[91] = in[113] & in2[113];
    assign P[91] = in[113] ^ in2[113];
    assign G[92] = in[112] & in2[112];
    assign P[92] = in[112] ^ in2[112];
    assign G[93] = in[111] & in2[111];
    assign P[93] = in[111] ^ in2[111];
    assign G[94] = in[110] & in2[110];
    assign P[94] = in[110] ^ in2[110];
    assign G[95] = in[109] & in2[109];
    assign P[95] = in[109] ^ in2[109];
    assign G[96] = in[108] & in2[108];
    assign P[96] = in[108] ^ in2[108];
    assign G[97] = in[107] & in2[107];
    assign P[97] = in[107] ^ in2[107];
    assign G[98] = in[106] & in2[106];
    assign P[98] = in[106] ^ in2[106];
    assign G[99] = in[105] & in2[105];
    assign P[99] = in[105] ^ in2[105];
    assign G[100] = in[104] & in2[104];
    assign P[100] = in[104] ^ in2[104];
    assign G[101] = in[103] & in2[103];
    assign P[101] = in[103] ^ in2[103];
    assign G[102] = in[102] & in2[102];
    assign P[102] = in[102] ^ in2[102];
    assign G[103] = in[101] & in2[101];
    assign P[103] = in[101] ^ in2[101];
    assign G[104] = in[100] & in2[100];
    assign P[104] = in[100] ^ in2[100];
    assign G[105] = in[99] & in2[99];
    assign P[105] = in[99] ^ in2[99];
    assign G[106] = in[98] & in2[98];
    assign P[106] = in[98] ^ in2[98];
    assign G[107] = in[97] & in2[97];
    assign P[107] = in[97] ^ in2[97];
    assign G[108] = in[96] & in2[96];
    assign P[108] = in[96] ^ in2[96];
    assign G[109] = in[95] & in2[95];
    assign P[109] = in[95] ^ in2[95];
    assign G[110] = in[94] & in2[94];
    assign P[110] = in[94] ^ in2[94];
    assign G[111] = in[93] & in2[93];
    assign P[111] = in[93] ^ in2[93];
    assign G[112] = in[92] & in2[92];
    assign P[112] = in[92] ^ in2[92];
    assign G[113] = in[91] & in2[91];
    assign P[113] = in[91] ^ in2[91];
    assign G[114] = in[90] & in2[90];
    assign P[114] = in[90] ^ in2[90];
    assign G[115] = in[89] & in2[89];
    assign P[115] = in[89] ^ in2[89];
    assign G[116] = in[88] & in2[88];
    assign P[116] = in[88] ^ in2[88];
    assign G[117] = in[87] & in2[87];
    assign P[117] = in[87] ^ in2[87];
    assign G[118] = in[86] & in2[86];
    assign P[118] = in[86] ^ in2[86];
    assign G[119] = in[85] & in2[85];
    assign P[119] = in[85] ^ in2[85];
    assign G[120] = in[84] & in2[84];
    assign P[120] = in[84] ^ in2[84];
    assign G[121] = in[83] & in2[83];
    assign P[121] = in[83] ^ in2[83];
    assign G[122] = in[82] & in2[82];
    assign P[122] = in[82] ^ in2[82];
    assign G[123] = in[81] & in2[81];
    assign P[123] = in[81] ^ in2[81];
    assign G[124] = in[80] & in2[80];
    assign P[124] = in[80] ^ in2[80];
    assign G[125] = in[79] & in2[79];
    assign P[125] = in[79] ^ in2[79];
    assign G[126] = in[78] & in2[78];
    assign P[126] = in[78] ^ in2[78];
    assign G[127] = in[77] & in2[77];
    assign P[127] = in[77] ^ in2[77];
    assign G[128] = in[76] & in2[76];
    assign P[128] = in[76] ^ in2[76];
    assign G[129] = in[75] & in2[75];
    assign P[129] = in[75] ^ in2[75];
    assign G[130] = in[74] & in2[74];
    assign P[130] = in[74] ^ in2[74];
    assign G[131] = in[73] & in2[73];
    assign P[131] = in[73] ^ in2[73];
    assign G[132] = in[72] & in2[72];
    assign P[132] = in[72] ^ in2[72];
    assign G[133] = in[71] & in2[71];
    assign P[133] = in[71] ^ in2[71];
    assign G[134] = in[70] & in2[70];
    assign P[134] = in[70] ^ in2[70];
    assign G[135] = in[69] & in2[69];
    assign P[135] = in[69] ^ in2[69];
    assign G[136] = in[68] & in2[68];
    assign P[136] = in[68] ^ in2[68];
    assign G[137] = in[67] & in2[67];
    assign P[137] = in[67] ^ in2[67];
    assign G[138] = in[66] & in2[66];
    assign P[138] = in[66] ^ in2[66];
    assign G[139] = in[65] & in2[65];
    assign P[139] = in[65] ^ in2[65];
    assign G[140] = in[64] & in2[64];
    assign P[140] = in[64] ^ in2[64];
    assign G[141] = in[63] & in2[63];
    assign P[141] = in[63] ^ in2[63];
    assign G[142] = in[62] & in2[62];
    assign P[142] = in[62] ^ in2[62];
    assign G[143] = in[61] & in2[61];
    assign P[143] = in[61] ^ in2[61];
    assign G[144] = in[60] & in2[60];
    assign P[144] = in[60] ^ in2[60];
    assign G[145] = in[59] & in2[59];
    assign P[145] = in[59] ^ in2[59];
    assign G[146] = in[58] & in2[58];
    assign P[146] = in[58] ^ in2[58];
    assign G[147] = in[57] & in2[57];
    assign P[147] = in[57] ^ in2[57];
    assign G[148] = in[56] & in2[56];
    assign P[148] = in[56] ^ in2[56];
    assign G[149] = in[55] & in2[55];
    assign P[149] = in[55] ^ in2[55];
    assign G[150] = in[54] & in2[54];
    assign P[150] = in[54] ^ in2[54];
    assign G[151] = in[53] & in2[53];
    assign P[151] = in[53] ^ in2[53];
    assign G[152] = in[52] & in2[52];
    assign P[152] = in[52] ^ in2[52];
    assign G[153] = in[51] & in2[51];
    assign P[153] = in[51] ^ in2[51];
    assign G[154] = in[50] & in2[50];
    assign P[154] = in[50] ^ in2[50];
    assign G[155] = in[49] & in2[49];
    assign P[155] = in[49] ^ in2[49];
    assign G[156] = in[48] & in2[48];
    assign P[156] = in[48] ^ in2[48];
    assign G[157] = in[47] & in2[47];
    assign P[157] = in[47] ^ in2[47];
    assign G[158] = in[46] & in2[46];
    assign P[158] = in[46] ^ in2[46];
    assign G[159] = in[45] & in2[45];
    assign P[159] = in[45] ^ in2[45];
    assign G[160] = in[44] & in2[44];
    assign P[160] = in[44] ^ in2[44];
    assign G[161] = in[43] & in2[43];
    assign P[161] = in[43] ^ in2[43];
    assign G[162] = in[42] & in2[42];
    assign P[162] = in[42] ^ in2[42];
    assign G[163] = in[41] & in2[41];
    assign P[163] = in[41] ^ in2[41];
    assign G[164] = in[40] & in2[40];
    assign P[164] = in[40] ^ in2[40];
    assign G[165] = in[39] & in2[39];
    assign P[165] = in[39] ^ in2[39];
    assign G[166] = in[38] & in2[38];
    assign P[166] = in[38] ^ in2[38];
    assign G[167] = in[37] & in2[37];
    assign P[167] = in[37] ^ in2[37];
    assign G[168] = in[36] & in2[36];
    assign P[168] = in[36] ^ in2[36];
    assign G[169] = in[35] & in2[35];
    assign P[169] = in[35] ^ in2[35];
    assign G[170] = in[34] & in2[34];
    assign P[170] = in[34] ^ in2[34];
    assign G[171] = in[33] & in2[33];
    assign P[171] = in[33] ^ in2[33];
    assign G[172] = in[32] & in2[32];
    assign P[172] = in[32] ^ in2[32];
    assign G[173] = in[31] & in2[31];
    assign P[173] = in[31] ^ in2[31];
    assign G[174] = in[30] & in2[30];
    assign P[174] = in[30] ^ in2[30];
    assign G[175] = in[29] & in2[29];
    assign P[175] = in[29] ^ in2[29];
    assign G[176] = in[28] & in2[28];
    assign P[176] = in[28] ^ in2[28];
    assign G[177] = in[27] & in2[27];
    assign P[177] = in[27] ^ in2[27];
    assign G[178] = in[26] & in2[26];
    assign P[178] = in[26] ^ in2[26];
    assign G[179] = in[25] & in2[25];
    assign P[179] = in[25] ^ in2[25];
    assign G[180] = in[24] & in2[24];
    assign P[180] = in[24] ^ in2[24];
    assign G[181] = in[23] & in2[23];
    assign P[181] = in[23] ^ in2[23];
    assign G[182] = in[22] & in2[22];
    assign P[182] = in[22] ^ in2[22];
    assign G[183] = in[21] & in2[21];
    assign P[183] = in[21] ^ in2[21];
    assign G[184] = in[20] & in2[20];
    assign P[184] = in[20] ^ in2[20];
    assign G[185] = in[19] & in2[19];
    assign P[185] = in[19] ^ in2[19];
    assign G[186] = in[18] & in2[18];
    assign P[186] = in[18] ^ in2[18];
    assign G[187] = in[17] & in2[17];
    assign P[187] = in[17] ^ in2[17];
    assign G[188] = in[16] & in2[16];
    assign P[188] = in[16] ^ in2[16];
    assign G[189] = in[15] & in2[15];
    assign P[189] = in[15] ^ in2[15];
    assign G[190] = in[14] & in2[14];
    assign P[190] = in[14] ^ in2[14];
    assign G[191] = in[13] & in2[13];
    assign P[191] = in[13] ^ in2[13];
    assign G[192] = in[12] & in2[12];
    assign P[192] = in[12] ^ in2[12];
    assign G[193] = in[11] & in2[11];
    assign P[193] = in[11] ^ in2[11];
    assign G[194] = in[10] & in2[10];
    assign P[194] = in[10] ^ in2[10];
    assign G[195] = in[9] & in2[9];
    assign P[195] = in[9] ^ in2[9];
    assign G[196] = in[8] & in2[8];
    assign P[196] = in[8] ^ in2[8];
    assign G[197] = in[7] & in2[7];
    assign P[197] = in[7] ^ in2[7];
    assign G[198] = in[6] & in2[6];
    assign P[198] = in[6] ^ in2[6];
    assign G[199] = in[5] & in2[5];
    assign P[199] = in[5] ^ in2[5];
    assign G[200] = in[4] & in2[4];
    assign P[200] = in[4] ^ in2[4];
    assign G[201] = in[3] & in2[3];
    assign P[201] = in[3] ^ in2[3];
    assign G[202] = in[2] & in2[2];
    assign P[202] = in[2] ^ in2[2];
    assign G[203] = in[1] & in2[1];
    assign P[203] = in[1] ^ in2[1];
    assign G[204] = in[0] & in2[0];
    assign P[204] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign C[204] = G[203] | (P[203] & C[203]);
    assign cout = G[204] | (P[204] & C[204]);
    assign sum = P ^ C;
endmodule

module CLA204(output [203:0] sum, output cout, input [203:0] in1, input [203:0] in2;

    wire[203:0] G;
    wire[203:0] C;
    wire[203:0] P;

    assign G[0] = in[203] & in2[203];
    assign P[0] = in[203] ^ in2[203];
    assign G[1] = in[202] & in2[202];
    assign P[1] = in[202] ^ in2[202];
    assign G[2] = in[201] & in2[201];
    assign P[2] = in[201] ^ in2[201];
    assign G[3] = in[200] & in2[200];
    assign P[3] = in[200] ^ in2[200];
    assign G[4] = in[199] & in2[199];
    assign P[4] = in[199] ^ in2[199];
    assign G[5] = in[198] & in2[198];
    assign P[5] = in[198] ^ in2[198];
    assign G[6] = in[197] & in2[197];
    assign P[6] = in[197] ^ in2[197];
    assign G[7] = in[196] & in2[196];
    assign P[7] = in[196] ^ in2[196];
    assign G[8] = in[195] & in2[195];
    assign P[8] = in[195] ^ in2[195];
    assign G[9] = in[194] & in2[194];
    assign P[9] = in[194] ^ in2[194];
    assign G[10] = in[193] & in2[193];
    assign P[10] = in[193] ^ in2[193];
    assign G[11] = in[192] & in2[192];
    assign P[11] = in[192] ^ in2[192];
    assign G[12] = in[191] & in2[191];
    assign P[12] = in[191] ^ in2[191];
    assign G[13] = in[190] & in2[190];
    assign P[13] = in[190] ^ in2[190];
    assign G[14] = in[189] & in2[189];
    assign P[14] = in[189] ^ in2[189];
    assign G[15] = in[188] & in2[188];
    assign P[15] = in[188] ^ in2[188];
    assign G[16] = in[187] & in2[187];
    assign P[16] = in[187] ^ in2[187];
    assign G[17] = in[186] & in2[186];
    assign P[17] = in[186] ^ in2[186];
    assign G[18] = in[185] & in2[185];
    assign P[18] = in[185] ^ in2[185];
    assign G[19] = in[184] & in2[184];
    assign P[19] = in[184] ^ in2[184];
    assign G[20] = in[183] & in2[183];
    assign P[20] = in[183] ^ in2[183];
    assign G[21] = in[182] & in2[182];
    assign P[21] = in[182] ^ in2[182];
    assign G[22] = in[181] & in2[181];
    assign P[22] = in[181] ^ in2[181];
    assign G[23] = in[180] & in2[180];
    assign P[23] = in[180] ^ in2[180];
    assign G[24] = in[179] & in2[179];
    assign P[24] = in[179] ^ in2[179];
    assign G[25] = in[178] & in2[178];
    assign P[25] = in[178] ^ in2[178];
    assign G[26] = in[177] & in2[177];
    assign P[26] = in[177] ^ in2[177];
    assign G[27] = in[176] & in2[176];
    assign P[27] = in[176] ^ in2[176];
    assign G[28] = in[175] & in2[175];
    assign P[28] = in[175] ^ in2[175];
    assign G[29] = in[174] & in2[174];
    assign P[29] = in[174] ^ in2[174];
    assign G[30] = in[173] & in2[173];
    assign P[30] = in[173] ^ in2[173];
    assign G[31] = in[172] & in2[172];
    assign P[31] = in[172] ^ in2[172];
    assign G[32] = in[171] & in2[171];
    assign P[32] = in[171] ^ in2[171];
    assign G[33] = in[170] & in2[170];
    assign P[33] = in[170] ^ in2[170];
    assign G[34] = in[169] & in2[169];
    assign P[34] = in[169] ^ in2[169];
    assign G[35] = in[168] & in2[168];
    assign P[35] = in[168] ^ in2[168];
    assign G[36] = in[167] & in2[167];
    assign P[36] = in[167] ^ in2[167];
    assign G[37] = in[166] & in2[166];
    assign P[37] = in[166] ^ in2[166];
    assign G[38] = in[165] & in2[165];
    assign P[38] = in[165] ^ in2[165];
    assign G[39] = in[164] & in2[164];
    assign P[39] = in[164] ^ in2[164];
    assign G[40] = in[163] & in2[163];
    assign P[40] = in[163] ^ in2[163];
    assign G[41] = in[162] & in2[162];
    assign P[41] = in[162] ^ in2[162];
    assign G[42] = in[161] & in2[161];
    assign P[42] = in[161] ^ in2[161];
    assign G[43] = in[160] & in2[160];
    assign P[43] = in[160] ^ in2[160];
    assign G[44] = in[159] & in2[159];
    assign P[44] = in[159] ^ in2[159];
    assign G[45] = in[158] & in2[158];
    assign P[45] = in[158] ^ in2[158];
    assign G[46] = in[157] & in2[157];
    assign P[46] = in[157] ^ in2[157];
    assign G[47] = in[156] & in2[156];
    assign P[47] = in[156] ^ in2[156];
    assign G[48] = in[155] & in2[155];
    assign P[48] = in[155] ^ in2[155];
    assign G[49] = in[154] & in2[154];
    assign P[49] = in[154] ^ in2[154];
    assign G[50] = in[153] & in2[153];
    assign P[50] = in[153] ^ in2[153];
    assign G[51] = in[152] & in2[152];
    assign P[51] = in[152] ^ in2[152];
    assign G[52] = in[151] & in2[151];
    assign P[52] = in[151] ^ in2[151];
    assign G[53] = in[150] & in2[150];
    assign P[53] = in[150] ^ in2[150];
    assign G[54] = in[149] & in2[149];
    assign P[54] = in[149] ^ in2[149];
    assign G[55] = in[148] & in2[148];
    assign P[55] = in[148] ^ in2[148];
    assign G[56] = in[147] & in2[147];
    assign P[56] = in[147] ^ in2[147];
    assign G[57] = in[146] & in2[146];
    assign P[57] = in[146] ^ in2[146];
    assign G[58] = in[145] & in2[145];
    assign P[58] = in[145] ^ in2[145];
    assign G[59] = in[144] & in2[144];
    assign P[59] = in[144] ^ in2[144];
    assign G[60] = in[143] & in2[143];
    assign P[60] = in[143] ^ in2[143];
    assign G[61] = in[142] & in2[142];
    assign P[61] = in[142] ^ in2[142];
    assign G[62] = in[141] & in2[141];
    assign P[62] = in[141] ^ in2[141];
    assign G[63] = in[140] & in2[140];
    assign P[63] = in[140] ^ in2[140];
    assign G[64] = in[139] & in2[139];
    assign P[64] = in[139] ^ in2[139];
    assign G[65] = in[138] & in2[138];
    assign P[65] = in[138] ^ in2[138];
    assign G[66] = in[137] & in2[137];
    assign P[66] = in[137] ^ in2[137];
    assign G[67] = in[136] & in2[136];
    assign P[67] = in[136] ^ in2[136];
    assign G[68] = in[135] & in2[135];
    assign P[68] = in[135] ^ in2[135];
    assign G[69] = in[134] & in2[134];
    assign P[69] = in[134] ^ in2[134];
    assign G[70] = in[133] & in2[133];
    assign P[70] = in[133] ^ in2[133];
    assign G[71] = in[132] & in2[132];
    assign P[71] = in[132] ^ in2[132];
    assign G[72] = in[131] & in2[131];
    assign P[72] = in[131] ^ in2[131];
    assign G[73] = in[130] & in2[130];
    assign P[73] = in[130] ^ in2[130];
    assign G[74] = in[129] & in2[129];
    assign P[74] = in[129] ^ in2[129];
    assign G[75] = in[128] & in2[128];
    assign P[75] = in[128] ^ in2[128];
    assign G[76] = in[127] & in2[127];
    assign P[76] = in[127] ^ in2[127];
    assign G[77] = in[126] & in2[126];
    assign P[77] = in[126] ^ in2[126];
    assign G[78] = in[125] & in2[125];
    assign P[78] = in[125] ^ in2[125];
    assign G[79] = in[124] & in2[124];
    assign P[79] = in[124] ^ in2[124];
    assign G[80] = in[123] & in2[123];
    assign P[80] = in[123] ^ in2[123];
    assign G[81] = in[122] & in2[122];
    assign P[81] = in[122] ^ in2[122];
    assign G[82] = in[121] & in2[121];
    assign P[82] = in[121] ^ in2[121];
    assign G[83] = in[120] & in2[120];
    assign P[83] = in[120] ^ in2[120];
    assign G[84] = in[119] & in2[119];
    assign P[84] = in[119] ^ in2[119];
    assign G[85] = in[118] & in2[118];
    assign P[85] = in[118] ^ in2[118];
    assign G[86] = in[117] & in2[117];
    assign P[86] = in[117] ^ in2[117];
    assign G[87] = in[116] & in2[116];
    assign P[87] = in[116] ^ in2[116];
    assign G[88] = in[115] & in2[115];
    assign P[88] = in[115] ^ in2[115];
    assign G[89] = in[114] & in2[114];
    assign P[89] = in[114] ^ in2[114];
    assign G[90] = in[113] & in2[113];
    assign P[90] = in[113] ^ in2[113];
    assign G[91] = in[112] & in2[112];
    assign P[91] = in[112] ^ in2[112];
    assign G[92] = in[111] & in2[111];
    assign P[92] = in[111] ^ in2[111];
    assign G[93] = in[110] & in2[110];
    assign P[93] = in[110] ^ in2[110];
    assign G[94] = in[109] & in2[109];
    assign P[94] = in[109] ^ in2[109];
    assign G[95] = in[108] & in2[108];
    assign P[95] = in[108] ^ in2[108];
    assign G[96] = in[107] & in2[107];
    assign P[96] = in[107] ^ in2[107];
    assign G[97] = in[106] & in2[106];
    assign P[97] = in[106] ^ in2[106];
    assign G[98] = in[105] & in2[105];
    assign P[98] = in[105] ^ in2[105];
    assign G[99] = in[104] & in2[104];
    assign P[99] = in[104] ^ in2[104];
    assign G[100] = in[103] & in2[103];
    assign P[100] = in[103] ^ in2[103];
    assign G[101] = in[102] & in2[102];
    assign P[101] = in[102] ^ in2[102];
    assign G[102] = in[101] & in2[101];
    assign P[102] = in[101] ^ in2[101];
    assign G[103] = in[100] & in2[100];
    assign P[103] = in[100] ^ in2[100];
    assign G[104] = in[99] & in2[99];
    assign P[104] = in[99] ^ in2[99];
    assign G[105] = in[98] & in2[98];
    assign P[105] = in[98] ^ in2[98];
    assign G[106] = in[97] & in2[97];
    assign P[106] = in[97] ^ in2[97];
    assign G[107] = in[96] & in2[96];
    assign P[107] = in[96] ^ in2[96];
    assign G[108] = in[95] & in2[95];
    assign P[108] = in[95] ^ in2[95];
    assign G[109] = in[94] & in2[94];
    assign P[109] = in[94] ^ in2[94];
    assign G[110] = in[93] & in2[93];
    assign P[110] = in[93] ^ in2[93];
    assign G[111] = in[92] & in2[92];
    assign P[111] = in[92] ^ in2[92];
    assign G[112] = in[91] & in2[91];
    assign P[112] = in[91] ^ in2[91];
    assign G[113] = in[90] & in2[90];
    assign P[113] = in[90] ^ in2[90];
    assign G[114] = in[89] & in2[89];
    assign P[114] = in[89] ^ in2[89];
    assign G[115] = in[88] & in2[88];
    assign P[115] = in[88] ^ in2[88];
    assign G[116] = in[87] & in2[87];
    assign P[116] = in[87] ^ in2[87];
    assign G[117] = in[86] & in2[86];
    assign P[117] = in[86] ^ in2[86];
    assign G[118] = in[85] & in2[85];
    assign P[118] = in[85] ^ in2[85];
    assign G[119] = in[84] & in2[84];
    assign P[119] = in[84] ^ in2[84];
    assign G[120] = in[83] & in2[83];
    assign P[120] = in[83] ^ in2[83];
    assign G[121] = in[82] & in2[82];
    assign P[121] = in[82] ^ in2[82];
    assign G[122] = in[81] & in2[81];
    assign P[122] = in[81] ^ in2[81];
    assign G[123] = in[80] & in2[80];
    assign P[123] = in[80] ^ in2[80];
    assign G[124] = in[79] & in2[79];
    assign P[124] = in[79] ^ in2[79];
    assign G[125] = in[78] & in2[78];
    assign P[125] = in[78] ^ in2[78];
    assign G[126] = in[77] & in2[77];
    assign P[126] = in[77] ^ in2[77];
    assign G[127] = in[76] & in2[76];
    assign P[127] = in[76] ^ in2[76];
    assign G[128] = in[75] & in2[75];
    assign P[128] = in[75] ^ in2[75];
    assign G[129] = in[74] & in2[74];
    assign P[129] = in[74] ^ in2[74];
    assign G[130] = in[73] & in2[73];
    assign P[130] = in[73] ^ in2[73];
    assign G[131] = in[72] & in2[72];
    assign P[131] = in[72] ^ in2[72];
    assign G[132] = in[71] & in2[71];
    assign P[132] = in[71] ^ in2[71];
    assign G[133] = in[70] & in2[70];
    assign P[133] = in[70] ^ in2[70];
    assign G[134] = in[69] & in2[69];
    assign P[134] = in[69] ^ in2[69];
    assign G[135] = in[68] & in2[68];
    assign P[135] = in[68] ^ in2[68];
    assign G[136] = in[67] & in2[67];
    assign P[136] = in[67] ^ in2[67];
    assign G[137] = in[66] & in2[66];
    assign P[137] = in[66] ^ in2[66];
    assign G[138] = in[65] & in2[65];
    assign P[138] = in[65] ^ in2[65];
    assign G[139] = in[64] & in2[64];
    assign P[139] = in[64] ^ in2[64];
    assign G[140] = in[63] & in2[63];
    assign P[140] = in[63] ^ in2[63];
    assign G[141] = in[62] & in2[62];
    assign P[141] = in[62] ^ in2[62];
    assign G[142] = in[61] & in2[61];
    assign P[142] = in[61] ^ in2[61];
    assign G[143] = in[60] & in2[60];
    assign P[143] = in[60] ^ in2[60];
    assign G[144] = in[59] & in2[59];
    assign P[144] = in[59] ^ in2[59];
    assign G[145] = in[58] & in2[58];
    assign P[145] = in[58] ^ in2[58];
    assign G[146] = in[57] & in2[57];
    assign P[146] = in[57] ^ in2[57];
    assign G[147] = in[56] & in2[56];
    assign P[147] = in[56] ^ in2[56];
    assign G[148] = in[55] & in2[55];
    assign P[148] = in[55] ^ in2[55];
    assign G[149] = in[54] & in2[54];
    assign P[149] = in[54] ^ in2[54];
    assign G[150] = in[53] & in2[53];
    assign P[150] = in[53] ^ in2[53];
    assign G[151] = in[52] & in2[52];
    assign P[151] = in[52] ^ in2[52];
    assign G[152] = in[51] & in2[51];
    assign P[152] = in[51] ^ in2[51];
    assign G[153] = in[50] & in2[50];
    assign P[153] = in[50] ^ in2[50];
    assign G[154] = in[49] & in2[49];
    assign P[154] = in[49] ^ in2[49];
    assign G[155] = in[48] & in2[48];
    assign P[155] = in[48] ^ in2[48];
    assign G[156] = in[47] & in2[47];
    assign P[156] = in[47] ^ in2[47];
    assign G[157] = in[46] & in2[46];
    assign P[157] = in[46] ^ in2[46];
    assign G[158] = in[45] & in2[45];
    assign P[158] = in[45] ^ in2[45];
    assign G[159] = in[44] & in2[44];
    assign P[159] = in[44] ^ in2[44];
    assign G[160] = in[43] & in2[43];
    assign P[160] = in[43] ^ in2[43];
    assign G[161] = in[42] & in2[42];
    assign P[161] = in[42] ^ in2[42];
    assign G[162] = in[41] & in2[41];
    assign P[162] = in[41] ^ in2[41];
    assign G[163] = in[40] & in2[40];
    assign P[163] = in[40] ^ in2[40];
    assign G[164] = in[39] & in2[39];
    assign P[164] = in[39] ^ in2[39];
    assign G[165] = in[38] & in2[38];
    assign P[165] = in[38] ^ in2[38];
    assign G[166] = in[37] & in2[37];
    assign P[166] = in[37] ^ in2[37];
    assign G[167] = in[36] & in2[36];
    assign P[167] = in[36] ^ in2[36];
    assign G[168] = in[35] & in2[35];
    assign P[168] = in[35] ^ in2[35];
    assign G[169] = in[34] & in2[34];
    assign P[169] = in[34] ^ in2[34];
    assign G[170] = in[33] & in2[33];
    assign P[170] = in[33] ^ in2[33];
    assign G[171] = in[32] & in2[32];
    assign P[171] = in[32] ^ in2[32];
    assign G[172] = in[31] & in2[31];
    assign P[172] = in[31] ^ in2[31];
    assign G[173] = in[30] & in2[30];
    assign P[173] = in[30] ^ in2[30];
    assign G[174] = in[29] & in2[29];
    assign P[174] = in[29] ^ in2[29];
    assign G[175] = in[28] & in2[28];
    assign P[175] = in[28] ^ in2[28];
    assign G[176] = in[27] & in2[27];
    assign P[176] = in[27] ^ in2[27];
    assign G[177] = in[26] & in2[26];
    assign P[177] = in[26] ^ in2[26];
    assign G[178] = in[25] & in2[25];
    assign P[178] = in[25] ^ in2[25];
    assign G[179] = in[24] & in2[24];
    assign P[179] = in[24] ^ in2[24];
    assign G[180] = in[23] & in2[23];
    assign P[180] = in[23] ^ in2[23];
    assign G[181] = in[22] & in2[22];
    assign P[181] = in[22] ^ in2[22];
    assign G[182] = in[21] & in2[21];
    assign P[182] = in[21] ^ in2[21];
    assign G[183] = in[20] & in2[20];
    assign P[183] = in[20] ^ in2[20];
    assign G[184] = in[19] & in2[19];
    assign P[184] = in[19] ^ in2[19];
    assign G[185] = in[18] & in2[18];
    assign P[185] = in[18] ^ in2[18];
    assign G[186] = in[17] & in2[17];
    assign P[186] = in[17] ^ in2[17];
    assign G[187] = in[16] & in2[16];
    assign P[187] = in[16] ^ in2[16];
    assign G[188] = in[15] & in2[15];
    assign P[188] = in[15] ^ in2[15];
    assign G[189] = in[14] & in2[14];
    assign P[189] = in[14] ^ in2[14];
    assign G[190] = in[13] & in2[13];
    assign P[190] = in[13] ^ in2[13];
    assign G[191] = in[12] & in2[12];
    assign P[191] = in[12] ^ in2[12];
    assign G[192] = in[11] & in2[11];
    assign P[192] = in[11] ^ in2[11];
    assign G[193] = in[10] & in2[10];
    assign P[193] = in[10] ^ in2[10];
    assign G[194] = in[9] & in2[9];
    assign P[194] = in[9] ^ in2[9];
    assign G[195] = in[8] & in2[8];
    assign P[195] = in[8] ^ in2[8];
    assign G[196] = in[7] & in2[7];
    assign P[196] = in[7] ^ in2[7];
    assign G[197] = in[6] & in2[6];
    assign P[197] = in[6] ^ in2[6];
    assign G[198] = in[5] & in2[5];
    assign P[198] = in[5] ^ in2[5];
    assign G[199] = in[4] & in2[4];
    assign P[199] = in[4] ^ in2[4];
    assign G[200] = in[3] & in2[3];
    assign P[200] = in[3] ^ in2[3];
    assign G[201] = in[2] & in2[2];
    assign P[201] = in[2] ^ in2[2];
    assign G[202] = in[1] & in2[1];
    assign P[202] = in[1] ^ in2[1];
    assign G[203] = in[0] & in2[0];
    assign P[203] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign C[203] = G[202] | (P[202] & C[202]);
    assign cout = G[203] | (P[203] & C[203]);
    assign sum = P ^ C;
endmodule

module CLA203(output [202:0] sum, output cout, input [202:0] in1, input [202:0] in2;

    wire[202:0] G;
    wire[202:0] C;
    wire[202:0] P;

    assign G[0] = in[202] & in2[202];
    assign P[0] = in[202] ^ in2[202];
    assign G[1] = in[201] & in2[201];
    assign P[1] = in[201] ^ in2[201];
    assign G[2] = in[200] & in2[200];
    assign P[2] = in[200] ^ in2[200];
    assign G[3] = in[199] & in2[199];
    assign P[3] = in[199] ^ in2[199];
    assign G[4] = in[198] & in2[198];
    assign P[4] = in[198] ^ in2[198];
    assign G[5] = in[197] & in2[197];
    assign P[5] = in[197] ^ in2[197];
    assign G[6] = in[196] & in2[196];
    assign P[6] = in[196] ^ in2[196];
    assign G[7] = in[195] & in2[195];
    assign P[7] = in[195] ^ in2[195];
    assign G[8] = in[194] & in2[194];
    assign P[8] = in[194] ^ in2[194];
    assign G[9] = in[193] & in2[193];
    assign P[9] = in[193] ^ in2[193];
    assign G[10] = in[192] & in2[192];
    assign P[10] = in[192] ^ in2[192];
    assign G[11] = in[191] & in2[191];
    assign P[11] = in[191] ^ in2[191];
    assign G[12] = in[190] & in2[190];
    assign P[12] = in[190] ^ in2[190];
    assign G[13] = in[189] & in2[189];
    assign P[13] = in[189] ^ in2[189];
    assign G[14] = in[188] & in2[188];
    assign P[14] = in[188] ^ in2[188];
    assign G[15] = in[187] & in2[187];
    assign P[15] = in[187] ^ in2[187];
    assign G[16] = in[186] & in2[186];
    assign P[16] = in[186] ^ in2[186];
    assign G[17] = in[185] & in2[185];
    assign P[17] = in[185] ^ in2[185];
    assign G[18] = in[184] & in2[184];
    assign P[18] = in[184] ^ in2[184];
    assign G[19] = in[183] & in2[183];
    assign P[19] = in[183] ^ in2[183];
    assign G[20] = in[182] & in2[182];
    assign P[20] = in[182] ^ in2[182];
    assign G[21] = in[181] & in2[181];
    assign P[21] = in[181] ^ in2[181];
    assign G[22] = in[180] & in2[180];
    assign P[22] = in[180] ^ in2[180];
    assign G[23] = in[179] & in2[179];
    assign P[23] = in[179] ^ in2[179];
    assign G[24] = in[178] & in2[178];
    assign P[24] = in[178] ^ in2[178];
    assign G[25] = in[177] & in2[177];
    assign P[25] = in[177] ^ in2[177];
    assign G[26] = in[176] & in2[176];
    assign P[26] = in[176] ^ in2[176];
    assign G[27] = in[175] & in2[175];
    assign P[27] = in[175] ^ in2[175];
    assign G[28] = in[174] & in2[174];
    assign P[28] = in[174] ^ in2[174];
    assign G[29] = in[173] & in2[173];
    assign P[29] = in[173] ^ in2[173];
    assign G[30] = in[172] & in2[172];
    assign P[30] = in[172] ^ in2[172];
    assign G[31] = in[171] & in2[171];
    assign P[31] = in[171] ^ in2[171];
    assign G[32] = in[170] & in2[170];
    assign P[32] = in[170] ^ in2[170];
    assign G[33] = in[169] & in2[169];
    assign P[33] = in[169] ^ in2[169];
    assign G[34] = in[168] & in2[168];
    assign P[34] = in[168] ^ in2[168];
    assign G[35] = in[167] & in2[167];
    assign P[35] = in[167] ^ in2[167];
    assign G[36] = in[166] & in2[166];
    assign P[36] = in[166] ^ in2[166];
    assign G[37] = in[165] & in2[165];
    assign P[37] = in[165] ^ in2[165];
    assign G[38] = in[164] & in2[164];
    assign P[38] = in[164] ^ in2[164];
    assign G[39] = in[163] & in2[163];
    assign P[39] = in[163] ^ in2[163];
    assign G[40] = in[162] & in2[162];
    assign P[40] = in[162] ^ in2[162];
    assign G[41] = in[161] & in2[161];
    assign P[41] = in[161] ^ in2[161];
    assign G[42] = in[160] & in2[160];
    assign P[42] = in[160] ^ in2[160];
    assign G[43] = in[159] & in2[159];
    assign P[43] = in[159] ^ in2[159];
    assign G[44] = in[158] & in2[158];
    assign P[44] = in[158] ^ in2[158];
    assign G[45] = in[157] & in2[157];
    assign P[45] = in[157] ^ in2[157];
    assign G[46] = in[156] & in2[156];
    assign P[46] = in[156] ^ in2[156];
    assign G[47] = in[155] & in2[155];
    assign P[47] = in[155] ^ in2[155];
    assign G[48] = in[154] & in2[154];
    assign P[48] = in[154] ^ in2[154];
    assign G[49] = in[153] & in2[153];
    assign P[49] = in[153] ^ in2[153];
    assign G[50] = in[152] & in2[152];
    assign P[50] = in[152] ^ in2[152];
    assign G[51] = in[151] & in2[151];
    assign P[51] = in[151] ^ in2[151];
    assign G[52] = in[150] & in2[150];
    assign P[52] = in[150] ^ in2[150];
    assign G[53] = in[149] & in2[149];
    assign P[53] = in[149] ^ in2[149];
    assign G[54] = in[148] & in2[148];
    assign P[54] = in[148] ^ in2[148];
    assign G[55] = in[147] & in2[147];
    assign P[55] = in[147] ^ in2[147];
    assign G[56] = in[146] & in2[146];
    assign P[56] = in[146] ^ in2[146];
    assign G[57] = in[145] & in2[145];
    assign P[57] = in[145] ^ in2[145];
    assign G[58] = in[144] & in2[144];
    assign P[58] = in[144] ^ in2[144];
    assign G[59] = in[143] & in2[143];
    assign P[59] = in[143] ^ in2[143];
    assign G[60] = in[142] & in2[142];
    assign P[60] = in[142] ^ in2[142];
    assign G[61] = in[141] & in2[141];
    assign P[61] = in[141] ^ in2[141];
    assign G[62] = in[140] & in2[140];
    assign P[62] = in[140] ^ in2[140];
    assign G[63] = in[139] & in2[139];
    assign P[63] = in[139] ^ in2[139];
    assign G[64] = in[138] & in2[138];
    assign P[64] = in[138] ^ in2[138];
    assign G[65] = in[137] & in2[137];
    assign P[65] = in[137] ^ in2[137];
    assign G[66] = in[136] & in2[136];
    assign P[66] = in[136] ^ in2[136];
    assign G[67] = in[135] & in2[135];
    assign P[67] = in[135] ^ in2[135];
    assign G[68] = in[134] & in2[134];
    assign P[68] = in[134] ^ in2[134];
    assign G[69] = in[133] & in2[133];
    assign P[69] = in[133] ^ in2[133];
    assign G[70] = in[132] & in2[132];
    assign P[70] = in[132] ^ in2[132];
    assign G[71] = in[131] & in2[131];
    assign P[71] = in[131] ^ in2[131];
    assign G[72] = in[130] & in2[130];
    assign P[72] = in[130] ^ in2[130];
    assign G[73] = in[129] & in2[129];
    assign P[73] = in[129] ^ in2[129];
    assign G[74] = in[128] & in2[128];
    assign P[74] = in[128] ^ in2[128];
    assign G[75] = in[127] & in2[127];
    assign P[75] = in[127] ^ in2[127];
    assign G[76] = in[126] & in2[126];
    assign P[76] = in[126] ^ in2[126];
    assign G[77] = in[125] & in2[125];
    assign P[77] = in[125] ^ in2[125];
    assign G[78] = in[124] & in2[124];
    assign P[78] = in[124] ^ in2[124];
    assign G[79] = in[123] & in2[123];
    assign P[79] = in[123] ^ in2[123];
    assign G[80] = in[122] & in2[122];
    assign P[80] = in[122] ^ in2[122];
    assign G[81] = in[121] & in2[121];
    assign P[81] = in[121] ^ in2[121];
    assign G[82] = in[120] & in2[120];
    assign P[82] = in[120] ^ in2[120];
    assign G[83] = in[119] & in2[119];
    assign P[83] = in[119] ^ in2[119];
    assign G[84] = in[118] & in2[118];
    assign P[84] = in[118] ^ in2[118];
    assign G[85] = in[117] & in2[117];
    assign P[85] = in[117] ^ in2[117];
    assign G[86] = in[116] & in2[116];
    assign P[86] = in[116] ^ in2[116];
    assign G[87] = in[115] & in2[115];
    assign P[87] = in[115] ^ in2[115];
    assign G[88] = in[114] & in2[114];
    assign P[88] = in[114] ^ in2[114];
    assign G[89] = in[113] & in2[113];
    assign P[89] = in[113] ^ in2[113];
    assign G[90] = in[112] & in2[112];
    assign P[90] = in[112] ^ in2[112];
    assign G[91] = in[111] & in2[111];
    assign P[91] = in[111] ^ in2[111];
    assign G[92] = in[110] & in2[110];
    assign P[92] = in[110] ^ in2[110];
    assign G[93] = in[109] & in2[109];
    assign P[93] = in[109] ^ in2[109];
    assign G[94] = in[108] & in2[108];
    assign P[94] = in[108] ^ in2[108];
    assign G[95] = in[107] & in2[107];
    assign P[95] = in[107] ^ in2[107];
    assign G[96] = in[106] & in2[106];
    assign P[96] = in[106] ^ in2[106];
    assign G[97] = in[105] & in2[105];
    assign P[97] = in[105] ^ in2[105];
    assign G[98] = in[104] & in2[104];
    assign P[98] = in[104] ^ in2[104];
    assign G[99] = in[103] & in2[103];
    assign P[99] = in[103] ^ in2[103];
    assign G[100] = in[102] & in2[102];
    assign P[100] = in[102] ^ in2[102];
    assign G[101] = in[101] & in2[101];
    assign P[101] = in[101] ^ in2[101];
    assign G[102] = in[100] & in2[100];
    assign P[102] = in[100] ^ in2[100];
    assign G[103] = in[99] & in2[99];
    assign P[103] = in[99] ^ in2[99];
    assign G[104] = in[98] & in2[98];
    assign P[104] = in[98] ^ in2[98];
    assign G[105] = in[97] & in2[97];
    assign P[105] = in[97] ^ in2[97];
    assign G[106] = in[96] & in2[96];
    assign P[106] = in[96] ^ in2[96];
    assign G[107] = in[95] & in2[95];
    assign P[107] = in[95] ^ in2[95];
    assign G[108] = in[94] & in2[94];
    assign P[108] = in[94] ^ in2[94];
    assign G[109] = in[93] & in2[93];
    assign P[109] = in[93] ^ in2[93];
    assign G[110] = in[92] & in2[92];
    assign P[110] = in[92] ^ in2[92];
    assign G[111] = in[91] & in2[91];
    assign P[111] = in[91] ^ in2[91];
    assign G[112] = in[90] & in2[90];
    assign P[112] = in[90] ^ in2[90];
    assign G[113] = in[89] & in2[89];
    assign P[113] = in[89] ^ in2[89];
    assign G[114] = in[88] & in2[88];
    assign P[114] = in[88] ^ in2[88];
    assign G[115] = in[87] & in2[87];
    assign P[115] = in[87] ^ in2[87];
    assign G[116] = in[86] & in2[86];
    assign P[116] = in[86] ^ in2[86];
    assign G[117] = in[85] & in2[85];
    assign P[117] = in[85] ^ in2[85];
    assign G[118] = in[84] & in2[84];
    assign P[118] = in[84] ^ in2[84];
    assign G[119] = in[83] & in2[83];
    assign P[119] = in[83] ^ in2[83];
    assign G[120] = in[82] & in2[82];
    assign P[120] = in[82] ^ in2[82];
    assign G[121] = in[81] & in2[81];
    assign P[121] = in[81] ^ in2[81];
    assign G[122] = in[80] & in2[80];
    assign P[122] = in[80] ^ in2[80];
    assign G[123] = in[79] & in2[79];
    assign P[123] = in[79] ^ in2[79];
    assign G[124] = in[78] & in2[78];
    assign P[124] = in[78] ^ in2[78];
    assign G[125] = in[77] & in2[77];
    assign P[125] = in[77] ^ in2[77];
    assign G[126] = in[76] & in2[76];
    assign P[126] = in[76] ^ in2[76];
    assign G[127] = in[75] & in2[75];
    assign P[127] = in[75] ^ in2[75];
    assign G[128] = in[74] & in2[74];
    assign P[128] = in[74] ^ in2[74];
    assign G[129] = in[73] & in2[73];
    assign P[129] = in[73] ^ in2[73];
    assign G[130] = in[72] & in2[72];
    assign P[130] = in[72] ^ in2[72];
    assign G[131] = in[71] & in2[71];
    assign P[131] = in[71] ^ in2[71];
    assign G[132] = in[70] & in2[70];
    assign P[132] = in[70] ^ in2[70];
    assign G[133] = in[69] & in2[69];
    assign P[133] = in[69] ^ in2[69];
    assign G[134] = in[68] & in2[68];
    assign P[134] = in[68] ^ in2[68];
    assign G[135] = in[67] & in2[67];
    assign P[135] = in[67] ^ in2[67];
    assign G[136] = in[66] & in2[66];
    assign P[136] = in[66] ^ in2[66];
    assign G[137] = in[65] & in2[65];
    assign P[137] = in[65] ^ in2[65];
    assign G[138] = in[64] & in2[64];
    assign P[138] = in[64] ^ in2[64];
    assign G[139] = in[63] & in2[63];
    assign P[139] = in[63] ^ in2[63];
    assign G[140] = in[62] & in2[62];
    assign P[140] = in[62] ^ in2[62];
    assign G[141] = in[61] & in2[61];
    assign P[141] = in[61] ^ in2[61];
    assign G[142] = in[60] & in2[60];
    assign P[142] = in[60] ^ in2[60];
    assign G[143] = in[59] & in2[59];
    assign P[143] = in[59] ^ in2[59];
    assign G[144] = in[58] & in2[58];
    assign P[144] = in[58] ^ in2[58];
    assign G[145] = in[57] & in2[57];
    assign P[145] = in[57] ^ in2[57];
    assign G[146] = in[56] & in2[56];
    assign P[146] = in[56] ^ in2[56];
    assign G[147] = in[55] & in2[55];
    assign P[147] = in[55] ^ in2[55];
    assign G[148] = in[54] & in2[54];
    assign P[148] = in[54] ^ in2[54];
    assign G[149] = in[53] & in2[53];
    assign P[149] = in[53] ^ in2[53];
    assign G[150] = in[52] & in2[52];
    assign P[150] = in[52] ^ in2[52];
    assign G[151] = in[51] & in2[51];
    assign P[151] = in[51] ^ in2[51];
    assign G[152] = in[50] & in2[50];
    assign P[152] = in[50] ^ in2[50];
    assign G[153] = in[49] & in2[49];
    assign P[153] = in[49] ^ in2[49];
    assign G[154] = in[48] & in2[48];
    assign P[154] = in[48] ^ in2[48];
    assign G[155] = in[47] & in2[47];
    assign P[155] = in[47] ^ in2[47];
    assign G[156] = in[46] & in2[46];
    assign P[156] = in[46] ^ in2[46];
    assign G[157] = in[45] & in2[45];
    assign P[157] = in[45] ^ in2[45];
    assign G[158] = in[44] & in2[44];
    assign P[158] = in[44] ^ in2[44];
    assign G[159] = in[43] & in2[43];
    assign P[159] = in[43] ^ in2[43];
    assign G[160] = in[42] & in2[42];
    assign P[160] = in[42] ^ in2[42];
    assign G[161] = in[41] & in2[41];
    assign P[161] = in[41] ^ in2[41];
    assign G[162] = in[40] & in2[40];
    assign P[162] = in[40] ^ in2[40];
    assign G[163] = in[39] & in2[39];
    assign P[163] = in[39] ^ in2[39];
    assign G[164] = in[38] & in2[38];
    assign P[164] = in[38] ^ in2[38];
    assign G[165] = in[37] & in2[37];
    assign P[165] = in[37] ^ in2[37];
    assign G[166] = in[36] & in2[36];
    assign P[166] = in[36] ^ in2[36];
    assign G[167] = in[35] & in2[35];
    assign P[167] = in[35] ^ in2[35];
    assign G[168] = in[34] & in2[34];
    assign P[168] = in[34] ^ in2[34];
    assign G[169] = in[33] & in2[33];
    assign P[169] = in[33] ^ in2[33];
    assign G[170] = in[32] & in2[32];
    assign P[170] = in[32] ^ in2[32];
    assign G[171] = in[31] & in2[31];
    assign P[171] = in[31] ^ in2[31];
    assign G[172] = in[30] & in2[30];
    assign P[172] = in[30] ^ in2[30];
    assign G[173] = in[29] & in2[29];
    assign P[173] = in[29] ^ in2[29];
    assign G[174] = in[28] & in2[28];
    assign P[174] = in[28] ^ in2[28];
    assign G[175] = in[27] & in2[27];
    assign P[175] = in[27] ^ in2[27];
    assign G[176] = in[26] & in2[26];
    assign P[176] = in[26] ^ in2[26];
    assign G[177] = in[25] & in2[25];
    assign P[177] = in[25] ^ in2[25];
    assign G[178] = in[24] & in2[24];
    assign P[178] = in[24] ^ in2[24];
    assign G[179] = in[23] & in2[23];
    assign P[179] = in[23] ^ in2[23];
    assign G[180] = in[22] & in2[22];
    assign P[180] = in[22] ^ in2[22];
    assign G[181] = in[21] & in2[21];
    assign P[181] = in[21] ^ in2[21];
    assign G[182] = in[20] & in2[20];
    assign P[182] = in[20] ^ in2[20];
    assign G[183] = in[19] & in2[19];
    assign P[183] = in[19] ^ in2[19];
    assign G[184] = in[18] & in2[18];
    assign P[184] = in[18] ^ in2[18];
    assign G[185] = in[17] & in2[17];
    assign P[185] = in[17] ^ in2[17];
    assign G[186] = in[16] & in2[16];
    assign P[186] = in[16] ^ in2[16];
    assign G[187] = in[15] & in2[15];
    assign P[187] = in[15] ^ in2[15];
    assign G[188] = in[14] & in2[14];
    assign P[188] = in[14] ^ in2[14];
    assign G[189] = in[13] & in2[13];
    assign P[189] = in[13] ^ in2[13];
    assign G[190] = in[12] & in2[12];
    assign P[190] = in[12] ^ in2[12];
    assign G[191] = in[11] & in2[11];
    assign P[191] = in[11] ^ in2[11];
    assign G[192] = in[10] & in2[10];
    assign P[192] = in[10] ^ in2[10];
    assign G[193] = in[9] & in2[9];
    assign P[193] = in[9] ^ in2[9];
    assign G[194] = in[8] & in2[8];
    assign P[194] = in[8] ^ in2[8];
    assign G[195] = in[7] & in2[7];
    assign P[195] = in[7] ^ in2[7];
    assign G[196] = in[6] & in2[6];
    assign P[196] = in[6] ^ in2[6];
    assign G[197] = in[5] & in2[5];
    assign P[197] = in[5] ^ in2[5];
    assign G[198] = in[4] & in2[4];
    assign P[198] = in[4] ^ in2[4];
    assign G[199] = in[3] & in2[3];
    assign P[199] = in[3] ^ in2[3];
    assign G[200] = in[2] & in2[2];
    assign P[200] = in[2] ^ in2[2];
    assign G[201] = in[1] & in2[1];
    assign P[201] = in[1] ^ in2[1];
    assign G[202] = in[0] & in2[0];
    assign P[202] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign C[202] = G[201] | (P[201] & C[201]);
    assign cout = G[202] | (P[202] & C[202]);
    assign sum = P ^ C;
endmodule

module CLA202(output [201:0] sum, output cout, input [201:0] in1, input [201:0] in2;

    wire[201:0] G;
    wire[201:0] C;
    wire[201:0] P;

    assign G[0] = in[201] & in2[201];
    assign P[0] = in[201] ^ in2[201];
    assign G[1] = in[200] & in2[200];
    assign P[1] = in[200] ^ in2[200];
    assign G[2] = in[199] & in2[199];
    assign P[2] = in[199] ^ in2[199];
    assign G[3] = in[198] & in2[198];
    assign P[3] = in[198] ^ in2[198];
    assign G[4] = in[197] & in2[197];
    assign P[4] = in[197] ^ in2[197];
    assign G[5] = in[196] & in2[196];
    assign P[5] = in[196] ^ in2[196];
    assign G[6] = in[195] & in2[195];
    assign P[6] = in[195] ^ in2[195];
    assign G[7] = in[194] & in2[194];
    assign P[7] = in[194] ^ in2[194];
    assign G[8] = in[193] & in2[193];
    assign P[8] = in[193] ^ in2[193];
    assign G[9] = in[192] & in2[192];
    assign P[9] = in[192] ^ in2[192];
    assign G[10] = in[191] & in2[191];
    assign P[10] = in[191] ^ in2[191];
    assign G[11] = in[190] & in2[190];
    assign P[11] = in[190] ^ in2[190];
    assign G[12] = in[189] & in2[189];
    assign P[12] = in[189] ^ in2[189];
    assign G[13] = in[188] & in2[188];
    assign P[13] = in[188] ^ in2[188];
    assign G[14] = in[187] & in2[187];
    assign P[14] = in[187] ^ in2[187];
    assign G[15] = in[186] & in2[186];
    assign P[15] = in[186] ^ in2[186];
    assign G[16] = in[185] & in2[185];
    assign P[16] = in[185] ^ in2[185];
    assign G[17] = in[184] & in2[184];
    assign P[17] = in[184] ^ in2[184];
    assign G[18] = in[183] & in2[183];
    assign P[18] = in[183] ^ in2[183];
    assign G[19] = in[182] & in2[182];
    assign P[19] = in[182] ^ in2[182];
    assign G[20] = in[181] & in2[181];
    assign P[20] = in[181] ^ in2[181];
    assign G[21] = in[180] & in2[180];
    assign P[21] = in[180] ^ in2[180];
    assign G[22] = in[179] & in2[179];
    assign P[22] = in[179] ^ in2[179];
    assign G[23] = in[178] & in2[178];
    assign P[23] = in[178] ^ in2[178];
    assign G[24] = in[177] & in2[177];
    assign P[24] = in[177] ^ in2[177];
    assign G[25] = in[176] & in2[176];
    assign P[25] = in[176] ^ in2[176];
    assign G[26] = in[175] & in2[175];
    assign P[26] = in[175] ^ in2[175];
    assign G[27] = in[174] & in2[174];
    assign P[27] = in[174] ^ in2[174];
    assign G[28] = in[173] & in2[173];
    assign P[28] = in[173] ^ in2[173];
    assign G[29] = in[172] & in2[172];
    assign P[29] = in[172] ^ in2[172];
    assign G[30] = in[171] & in2[171];
    assign P[30] = in[171] ^ in2[171];
    assign G[31] = in[170] & in2[170];
    assign P[31] = in[170] ^ in2[170];
    assign G[32] = in[169] & in2[169];
    assign P[32] = in[169] ^ in2[169];
    assign G[33] = in[168] & in2[168];
    assign P[33] = in[168] ^ in2[168];
    assign G[34] = in[167] & in2[167];
    assign P[34] = in[167] ^ in2[167];
    assign G[35] = in[166] & in2[166];
    assign P[35] = in[166] ^ in2[166];
    assign G[36] = in[165] & in2[165];
    assign P[36] = in[165] ^ in2[165];
    assign G[37] = in[164] & in2[164];
    assign P[37] = in[164] ^ in2[164];
    assign G[38] = in[163] & in2[163];
    assign P[38] = in[163] ^ in2[163];
    assign G[39] = in[162] & in2[162];
    assign P[39] = in[162] ^ in2[162];
    assign G[40] = in[161] & in2[161];
    assign P[40] = in[161] ^ in2[161];
    assign G[41] = in[160] & in2[160];
    assign P[41] = in[160] ^ in2[160];
    assign G[42] = in[159] & in2[159];
    assign P[42] = in[159] ^ in2[159];
    assign G[43] = in[158] & in2[158];
    assign P[43] = in[158] ^ in2[158];
    assign G[44] = in[157] & in2[157];
    assign P[44] = in[157] ^ in2[157];
    assign G[45] = in[156] & in2[156];
    assign P[45] = in[156] ^ in2[156];
    assign G[46] = in[155] & in2[155];
    assign P[46] = in[155] ^ in2[155];
    assign G[47] = in[154] & in2[154];
    assign P[47] = in[154] ^ in2[154];
    assign G[48] = in[153] & in2[153];
    assign P[48] = in[153] ^ in2[153];
    assign G[49] = in[152] & in2[152];
    assign P[49] = in[152] ^ in2[152];
    assign G[50] = in[151] & in2[151];
    assign P[50] = in[151] ^ in2[151];
    assign G[51] = in[150] & in2[150];
    assign P[51] = in[150] ^ in2[150];
    assign G[52] = in[149] & in2[149];
    assign P[52] = in[149] ^ in2[149];
    assign G[53] = in[148] & in2[148];
    assign P[53] = in[148] ^ in2[148];
    assign G[54] = in[147] & in2[147];
    assign P[54] = in[147] ^ in2[147];
    assign G[55] = in[146] & in2[146];
    assign P[55] = in[146] ^ in2[146];
    assign G[56] = in[145] & in2[145];
    assign P[56] = in[145] ^ in2[145];
    assign G[57] = in[144] & in2[144];
    assign P[57] = in[144] ^ in2[144];
    assign G[58] = in[143] & in2[143];
    assign P[58] = in[143] ^ in2[143];
    assign G[59] = in[142] & in2[142];
    assign P[59] = in[142] ^ in2[142];
    assign G[60] = in[141] & in2[141];
    assign P[60] = in[141] ^ in2[141];
    assign G[61] = in[140] & in2[140];
    assign P[61] = in[140] ^ in2[140];
    assign G[62] = in[139] & in2[139];
    assign P[62] = in[139] ^ in2[139];
    assign G[63] = in[138] & in2[138];
    assign P[63] = in[138] ^ in2[138];
    assign G[64] = in[137] & in2[137];
    assign P[64] = in[137] ^ in2[137];
    assign G[65] = in[136] & in2[136];
    assign P[65] = in[136] ^ in2[136];
    assign G[66] = in[135] & in2[135];
    assign P[66] = in[135] ^ in2[135];
    assign G[67] = in[134] & in2[134];
    assign P[67] = in[134] ^ in2[134];
    assign G[68] = in[133] & in2[133];
    assign P[68] = in[133] ^ in2[133];
    assign G[69] = in[132] & in2[132];
    assign P[69] = in[132] ^ in2[132];
    assign G[70] = in[131] & in2[131];
    assign P[70] = in[131] ^ in2[131];
    assign G[71] = in[130] & in2[130];
    assign P[71] = in[130] ^ in2[130];
    assign G[72] = in[129] & in2[129];
    assign P[72] = in[129] ^ in2[129];
    assign G[73] = in[128] & in2[128];
    assign P[73] = in[128] ^ in2[128];
    assign G[74] = in[127] & in2[127];
    assign P[74] = in[127] ^ in2[127];
    assign G[75] = in[126] & in2[126];
    assign P[75] = in[126] ^ in2[126];
    assign G[76] = in[125] & in2[125];
    assign P[76] = in[125] ^ in2[125];
    assign G[77] = in[124] & in2[124];
    assign P[77] = in[124] ^ in2[124];
    assign G[78] = in[123] & in2[123];
    assign P[78] = in[123] ^ in2[123];
    assign G[79] = in[122] & in2[122];
    assign P[79] = in[122] ^ in2[122];
    assign G[80] = in[121] & in2[121];
    assign P[80] = in[121] ^ in2[121];
    assign G[81] = in[120] & in2[120];
    assign P[81] = in[120] ^ in2[120];
    assign G[82] = in[119] & in2[119];
    assign P[82] = in[119] ^ in2[119];
    assign G[83] = in[118] & in2[118];
    assign P[83] = in[118] ^ in2[118];
    assign G[84] = in[117] & in2[117];
    assign P[84] = in[117] ^ in2[117];
    assign G[85] = in[116] & in2[116];
    assign P[85] = in[116] ^ in2[116];
    assign G[86] = in[115] & in2[115];
    assign P[86] = in[115] ^ in2[115];
    assign G[87] = in[114] & in2[114];
    assign P[87] = in[114] ^ in2[114];
    assign G[88] = in[113] & in2[113];
    assign P[88] = in[113] ^ in2[113];
    assign G[89] = in[112] & in2[112];
    assign P[89] = in[112] ^ in2[112];
    assign G[90] = in[111] & in2[111];
    assign P[90] = in[111] ^ in2[111];
    assign G[91] = in[110] & in2[110];
    assign P[91] = in[110] ^ in2[110];
    assign G[92] = in[109] & in2[109];
    assign P[92] = in[109] ^ in2[109];
    assign G[93] = in[108] & in2[108];
    assign P[93] = in[108] ^ in2[108];
    assign G[94] = in[107] & in2[107];
    assign P[94] = in[107] ^ in2[107];
    assign G[95] = in[106] & in2[106];
    assign P[95] = in[106] ^ in2[106];
    assign G[96] = in[105] & in2[105];
    assign P[96] = in[105] ^ in2[105];
    assign G[97] = in[104] & in2[104];
    assign P[97] = in[104] ^ in2[104];
    assign G[98] = in[103] & in2[103];
    assign P[98] = in[103] ^ in2[103];
    assign G[99] = in[102] & in2[102];
    assign P[99] = in[102] ^ in2[102];
    assign G[100] = in[101] & in2[101];
    assign P[100] = in[101] ^ in2[101];
    assign G[101] = in[100] & in2[100];
    assign P[101] = in[100] ^ in2[100];
    assign G[102] = in[99] & in2[99];
    assign P[102] = in[99] ^ in2[99];
    assign G[103] = in[98] & in2[98];
    assign P[103] = in[98] ^ in2[98];
    assign G[104] = in[97] & in2[97];
    assign P[104] = in[97] ^ in2[97];
    assign G[105] = in[96] & in2[96];
    assign P[105] = in[96] ^ in2[96];
    assign G[106] = in[95] & in2[95];
    assign P[106] = in[95] ^ in2[95];
    assign G[107] = in[94] & in2[94];
    assign P[107] = in[94] ^ in2[94];
    assign G[108] = in[93] & in2[93];
    assign P[108] = in[93] ^ in2[93];
    assign G[109] = in[92] & in2[92];
    assign P[109] = in[92] ^ in2[92];
    assign G[110] = in[91] & in2[91];
    assign P[110] = in[91] ^ in2[91];
    assign G[111] = in[90] & in2[90];
    assign P[111] = in[90] ^ in2[90];
    assign G[112] = in[89] & in2[89];
    assign P[112] = in[89] ^ in2[89];
    assign G[113] = in[88] & in2[88];
    assign P[113] = in[88] ^ in2[88];
    assign G[114] = in[87] & in2[87];
    assign P[114] = in[87] ^ in2[87];
    assign G[115] = in[86] & in2[86];
    assign P[115] = in[86] ^ in2[86];
    assign G[116] = in[85] & in2[85];
    assign P[116] = in[85] ^ in2[85];
    assign G[117] = in[84] & in2[84];
    assign P[117] = in[84] ^ in2[84];
    assign G[118] = in[83] & in2[83];
    assign P[118] = in[83] ^ in2[83];
    assign G[119] = in[82] & in2[82];
    assign P[119] = in[82] ^ in2[82];
    assign G[120] = in[81] & in2[81];
    assign P[120] = in[81] ^ in2[81];
    assign G[121] = in[80] & in2[80];
    assign P[121] = in[80] ^ in2[80];
    assign G[122] = in[79] & in2[79];
    assign P[122] = in[79] ^ in2[79];
    assign G[123] = in[78] & in2[78];
    assign P[123] = in[78] ^ in2[78];
    assign G[124] = in[77] & in2[77];
    assign P[124] = in[77] ^ in2[77];
    assign G[125] = in[76] & in2[76];
    assign P[125] = in[76] ^ in2[76];
    assign G[126] = in[75] & in2[75];
    assign P[126] = in[75] ^ in2[75];
    assign G[127] = in[74] & in2[74];
    assign P[127] = in[74] ^ in2[74];
    assign G[128] = in[73] & in2[73];
    assign P[128] = in[73] ^ in2[73];
    assign G[129] = in[72] & in2[72];
    assign P[129] = in[72] ^ in2[72];
    assign G[130] = in[71] & in2[71];
    assign P[130] = in[71] ^ in2[71];
    assign G[131] = in[70] & in2[70];
    assign P[131] = in[70] ^ in2[70];
    assign G[132] = in[69] & in2[69];
    assign P[132] = in[69] ^ in2[69];
    assign G[133] = in[68] & in2[68];
    assign P[133] = in[68] ^ in2[68];
    assign G[134] = in[67] & in2[67];
    assign P[134] = in[67] ^ in2[67];
    assign G[135] = in[66] & in2[66];
    assign P[135] = in[66] ^ in2[66];
    assign G[136] = in[65] & in2[65];
    assign P[136] = in[65] ^ in2[65];
    assign G[137] = in[64] & in2[64];
    assign P[137] = in[64] ^ in2[64];
    assign G[138] = in[63] & in2[63];
    assign P[138] = in[63] ^ in2[63];
    assign G[139] = in[62] & in2[62];
    assign P[139] = in[62] ^ in2[62];
    assign G[140] = in[61] & in2[61];
    assign P[140] = in[61] ^ in2[61];
    assign G[141] = in[60] & in2[60];
    assign P[141] = in[60] ^ in2[60];
    assign G[142] = in[59] & in2[59];
    assign P[142] = in[59] ^ in2[59];
    assign G[143] = in[58] & in2[58];
    assign P[143] = in[58] ^ in2[58];
    assign G[144] = in[57] & in2[57];
    assign P[144] = in[57] ^ in2[57];
    assign G[145] = in[56] & in2[56];
    assign P[145] = in[56] ^ in2[56];
    assign G[146] = in[55] & in2[55];
    assign P[146] = in[55] ^ in2[55];
    assign G[147] = in[54] & in2[54];
    assign P[147] = in[54] ^ in2[54];
    assign G[148] = in[53] & in2[53];
    assign P[148] = in[53] ^ in2[53];
    assign G[149] = in[52] & in2[52];
    assign P[149] = in[52] ^ in2[52];
    assign G[150] = in[51] & in2[51];
    assign P[150] = in[51] ^ in2[51];
    assign G[151] = in[50] & in2[50];
    assign P[151] = in[50] ^ in2[50];
    assign G[152] = in[49] & in2[49];
    assign P[152] = in[49] ^ in2[49];
    assign G[153] = in[48] & in2[48];
    assign P[153] = in[48] ^ in2[48];
    assign G[154] = in[47] & in2[47];
    assign P[154] = in[47] ^ in2[47];
    assign G[155] = in[46] & in2[46];
    assign P[155] = in[46] ^ in2[46];
    assign G[156] = in[45] & in2[45];
    assign P[156] = in[45] ^ in2[45];
    assign G[157] = in[44] & in2[44];
    assign P[157] = in[44] ^ in2[44];
    assign G[158] = in[43] & in2[43];
    assign P[158] = in[43] ^ in2[43];
    assign G[159] = in[42] & in2[42];
    assign P[159] = in[42] ^ in2[42];
    assign G[160] = in[41] & in2[41];
    assign P[160] = in[41] ^ in2[41];
    assign G[161] = in[40] & in2[40];
    assign P[161] = in[40] ^ in2[40];
    assign G[162] = in[39] & in2[39];
    assign P[162] = in[39] ^ in2[39];
    assign G[163] = in[38] & in2[38];
    assign P[163] = in[38] ^ in2[38];
    assign G[164] = in[37] & in2[37];
    assign P[164] = in[37] ^ in2[37];
    assign G[165] = in[36] & in2[36];
    assign P[165] = in[36] ^ in2[36];
    assign G[166] = in[35] & in2[35];
    assign P[166] = in[35] ^ in2[35];
    assign G[167] = in[34] & in2[34];
    assign P[167] = in[34] ^ in2[34];
    assign G[168] = in[33] & in2[33];
    assign P[168] = in[33] ^ in2[33];
    assign G[169] = in[32] & in2[32];
    assign P[169] = in[32] ^ in2[32];
    assign G[170] = in[31] & in2[31];
    assign P[170] = in[31] ^ in2[31];
    assign G[171] = in[30] & in2[30];
    assign P[171] = in[30] ^ in2[30];
    assign G[172] = in[29] & in2[29];
    assign P[172] = in[29] ^ in2[29];
    assign G[173] = in[28] & in2[28];
    assign P[173] = in[28] ^ in2[28];
    assign G[174] = in[27] & in2[27];
    assign P[174] = in[27] ^ in2[27];
    assign G[175] = in[26] & in2[26];
    assign P[175] = in[26] ^ in2[26];
    assign G[176] = in[25] & in2[25];
    assign P[176] = in[25] ^ in2[25];
    assign G[177] = in[24] & in2[24];
    assign P[177] = in[24] ^ in2[24];
    assign G[178] = in[23] & in2[23];
    assign P[178] = in[23] ^ in2[23];
    assign G[179] = in[22] & in2[22];
    assign P[179] = in[22] ^ in2[22];
    assign G[180] = in[21] & in2[21];
    assign P[180] = in[21] ^ in2[21];
    assign G[181] = in[20] & in2[20];
    assign P[181] = in[20] ^ in2[20];
    assign G[182] = in[19] & in2[19];
    assign P[182] = in[19] ^ in2[19];
    assign G[183] = in[18] & in2[18];
    assign P[183] = in[18] ^ in2[18];
    assign G[184] = in[17] & in2[17];
    assign P[184] = in[17] ^ in2[17];
    assign G[185] = in[16] & in2[16];
    assign P[185] = in[16] ^ in2[16];
    assign G[186] = in[15] & in2[15];
    assign P[186] = in[15] ^ in2[15];
    assign G[187] = in[14] & in2[14];
    assign P[187] = in[14] ^ in2[14];
    assign G[188] = in[13] & in2[13];
    assign P[188] = in[13] ^ in2[13];
    assign G[189] = in[12] & in2[12];
    assign P[189] = in[12] ^ in2[12];
    assign G[190] = in[11] & in2[11];
    assign P[190] = in[11] ^ in2[11];
    assign G[191] = in[10] & in2[10];
    assign P[191] = in[10] ^ in2[10];
    assign G[192] = in[9] & in2[9];
    assign P[192] = in[9] ^ in2[9];
    assign G[193] = in[8] & in2[8];
    assign P[193] = in[8] ^ in2[8];
    assign G[194] = in[7] & in2[7];
    assign P[194] = in[7] ^ in2[7];
    assign G[195] = in[6] & in2[6];
    assign P[195] = in[6] ^ in2[6];
    assign G[196] = in[5] & in2[5];
    assign P[196] = in[5] ^ in2[5];
    assign G[197] = in[4] & in2[4];
    assign P[197] = in[4] ^ in2[4];
    assign G[198] = in[3] & in2[3];
    assign P[198] = in[3] ^ in2[3];
    assign G[199] = in[2] & in2[2];
    assign P[199] = in[2] ^ in2[2];
    assign G[200] = in[1] & in2[1];
    assign P[200] = in[1] ^ in2[1];
    assign G[201] = in[0] & in2[0];
    assign P[201] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign C[201] = G[200] | (P[200] & C[200]);
    assign cout = G[201] | (P[201] & C[201]);
    assign sum = P ^ C;
endmodule

module CLA201(output [200:0] sum, output cout, input [200:0] in1, input [200:0] in2;

    wire[200:0] G;
    wire[200:0] C;
    wire[200:0] P;

    assign G[0] = in[200] & in2[200];
    assign P[0] = in[200] ^ in2[200];
    assign G[1] = in[199] & in2[199];
    assign P[1] = in[199] ^ in2[199];
    assign G[2] = in[198] & in2[198];
    assign P[2] = in[198] ^ in2[198];
    assign G[3] = in[197] & in2[197];
    assign P[3] = in[197] ^ in2[197];
    assign G[4] = in[196] & in2[196];
    assign P[4] = in[196] ^ in2[196];
    assign G[5] = in[195] & in2[195];
    assign P[5] = in[195] ^ in2[195];
    assign G[6] = in[194] & in2[194];
    assign P[6] = in[194] ^ in2[194];
    assign G[7] = in[193] & in2[193];
    assign P[7] = in[193] ^ in2[193];
    assign G[8] = in[192] & in2[192];
    assign P[8] = in[192] ^ in2[192];
    assign G[9] = in[191] & in2[191];
    assign P[9] = in[191] ^ in2[191];
    assign G[10] = in[190] & in2[190];
    assign P[10] = in[190] ^ in2[190];
    assign G[11] = in[189] & in2[189];
    assign P[11] = in[189] ^ in2[189];
    assign G[12] = in[188] & in2[188];
    assign P[12] = in[188] ^ in2[188];
    assign G[13] = in[187] & in2[187];
    assign P[13] = in[187] ^ in2[187];
    assign G[14] = in[186] & in2[186];
    assign P[14] = in[186] ^ in2[186];
    assign G[15] = in[185] & in2[185];
    assign P[15] = in[185] ^ in2[185];
    assign G[16] = in[184] & in2[184];
    assign P[16] = in[184] ^ in2[184];
    assign G[17] = in[183] & in2[183];
    assign P[17] = in[183] ^ in2[183];
    assign G[18] = in[182] & in2[182];
    assign P[18] = in[182] ^ in2[182];
    assign G[19] = in[181] & in2[181];
    assign P[19] = in[181] ^ in2[181];
    assign G[20] = in[180] & in2[180];
    assign P[20] = in[180] ^ in2[180];
    assign G[21] = in[179] & in2[179];
    assign P[21] = in[179] ^ in2[179];
    assign G[22] = in[178] & in2[178];
    assign P[22] = in[178] ^ in2[178];
    assign G[23] = in[177] & in2[177];
    assign P[23] = in[177] ^ in2[177];
    assign G[24] = in[176] & in2[176];
    assign P[24] = in[176] ^ in2[176];
    assign G[25] = in[175] & in2[175];
    assign P[25] = in[175] ^ in2[175];
    assign G[26] = in[174] & in2[174];
    assign P[26] = in[174] ^ in2[174];
    assign G[27] = in[173] & in2[173];
    assign P[27] = in[173] ^ in2[173];
    assign G[28] = in[172] & in2[172];
    assign P[28] = in[172] ^ in2[172];
    assign G[29] = in[171] & in2[171];
    assign P[29] = in[171] ^ in2[171];
    assign G[30] = in[170] & in2[170];
    assign P[30] = in[170] ^ in2[170];
    assign G[31] = in[169] & in2[169];
    assign P[31] = in[169] ^ in2[169];
    assign G[32] = in[168] & in2[168];
    assign P[32] = in[168] ^ in2[168];
    assign G[33] = in[167] & in2[167];
    assign P[33] = in[167] ^ in2[167];
    assign G[34] = in[166] & in2[166];
    assign P[34] = in[166] ^ in2[166];
    assign G[35] = in[165] & in2[165];
    assign P[35] = in[165] ^ in2[165];
    assign G[36] = in[164] & in2[164];
    assign P[36] = in[164] ^ in2[164];
    assign G[37] = in[163] & in2[163];
    assign P[37] = in[163] ^ in2[163];
    assign G[38] = in[162] & in2[162];
    assign P[38] = in[162] ^ in2[162];
    assign G[39] = in[161] & in2[161];
    assign P[39] = in[161] ^ in2[161];
    assign G[40] = in[160] & in2[160];
    assign P[40] = in[160] ^ in2[160];
    assign G[41] = in[159] & in2[159];
    assign P[41] = in[159] ^ in2[159];
    assign G[42] = in[158] & in2[158];
    assign P[42] = in[158] ^ in2[158];
    assign G[43] = in[157] & in2[157];
    assign P[43] = in[157] ^ in2[157];
    assign G[44] = in[156] & in2[156];
    assign P[44] = in[156] ^ in2[156];
    assign G[45] = in[155] & in2[155];
    assign P[45] = in[155] ^ in2[155];
    assign G[46] = in[154] & in2[154];
    assign P[46] = in[154] ^ in2[154];
    assign G[47] = in[153] & in2[153];
    assign P[47] = in[153] ^ in2[153];
    assign G[48] = in[152] & in2[152];
    assign P[48] = in[152] ^ in2[152];
    assign G[49] = in[151] & in2[151];
    assign P[49] = in[151] ^ in2[151];
    assign G[50] = in[150] & in2[150];
    assign P[50] = in[150] ^ in2[150];
    assign G[51] = in[149] & in2[149];
    assign P[51] = in[149] ^ in2[149];
    assign G[52] = in[148] & in2[148];
    assign P[52] = in[148] ^ in2[148];
    assign G[53] = in[147] & in2[147];
    assign P[53] = in[147] ^ in2[147];
    assign G[54] = in[146] & in2[146];
    assign P[54] = in[146] ^ in2[146];
    assign G[55] = in[145] & in2[145];
    assign P[55] = in[145] ^ in2[145];
    assign G[56] = in[144] & in2[144];
    assign P[56] = in[144] ^ in2[144];
    assign G[57] = in[143] & in2[143];
    assign P[57] = in[143] ^ in2[143];
    assign G[58] = in[142] & in2[142];
    assign P[58] = in[142] ^ in2[142];
    assign G[59] = in[141] & in2[141];
    assign P[59] = in[141] ^ in2[141];
    assign G[60] = in[140] & in2[140];
    assign P[60] = in[140] ^ in2[140];
    assign G[61] = in[139] & in2[139];
    assign P[61] = in[139] ^ in2[139];
    assign G[62] = in[138] & in2[138];
    assign P[62] = in[138] ^ in2[138];
    assign G[63] = in[137] & in2[137];
    assign P[63] = in[137] ^ in2[137];
    assign G[64] = in[136] & in2[136];
    assign P[64] = in[136] ^ in2[136];
    assign G[65] = in[135] & in2[135];
    assign P[65] = in[135] ^ in2[135];
    assign G[66] = in[134] & in2[134];
    assign P[66] = in[134] ^ in2[134];
    assign G[67] = in[133] & in2[133];
    assign P[67] = in[133] ^ in2[133];
    assign G[68] = in[132] & in2[132];
    assign P[68] = in[132] ^ in2[132];
    assign G[69] = in[131] & in2[131];
    assign P[69] = in[131] ^ in2[131];
    assign G[70] = in[130] & in2[130];
    assign P[70] = in[130] ^ in2[130];
    assign G[71] = in[129] & in2[129];
    assign P[71] = in[129] ^ in2[129];
    assign G[72] = in[128] & in2[128];
    assign P[72] = in[128] ^ in2[128];
    assign G[73] = in[127] & in2[127];
    assign P[73] = in[127] ^ in2[127];
    assign G[74] = in[126] & in2[126];
    assign P[74] = in[126] ^ in2[126];
    assign G[75] = in[125] & in2[125];
    assign P[75] = in[125] ^ in2[125];
    assign G[76] = in[124] & in2[124];
    assign P[76] = in[124] ^ in2[124];
    assign G[77] = in[123] & in2[123];
    assign P[77] = in[123] ^ in2[123];
    assign G[78] = in[122] & in2[122];
    assign P[78] = in[122] ^ in2[122];
    assign G[79] = in[121] & in2[121];
    assign P[79] = in[121] ^ in2[121];
    assign G[80] = in[120] & in2[120];
    assign P[80] = in[120] ^ in2[120];
    assign G[81] = in[119] & in2[119];
    assign P[81] = in[119] ^ in2[119];
    assign G[82] = in[118] & in2[118];
    assign P[82] = in[118] ^ in2[118];
    assign G[83] = in[117] & in2[117];
    assign P[83] = in[117] ^ in2[117];
    assign G[84] = in[116] & in2[116];
    assign P[84] = in[116] ^ in2[116];
    assign G[85] = in[115] & in2[115];
    assign P[85] = in[115] ^ in2[115];
    assign G[86] = in[114] & in2[114];
    assign P[86] = in[114] ^ in2[114];
    assign G[87] = in[113] & in2[113];
    assign P[87] = in[113] ^ in2[113];
    assign G[88] = in[112] & in2[112];
    assign P[88] = in[112] ^ in2[112];
    assign G[89] = in[111] & in2[111];
    assign P[89] = in[111] ^ in2[111];
    assign G[90] = in[110] & in2[110];
    assign P[90] = in[110] ^ in2[110];
    assign G[91] = in[109] & in2[109];
    assign P[91] = in[109] ^ in2[109];
    assign G[92] = in[108] & in2[108];
    assign P[92] = in[108] ^ in2[108];
    assign G[93] = in[107] & in2[107];
    assign P[93] = in[107] ^ in2[107];
    assign G[94] = in[106] & in2[106];
    assign P[94] = in[106] ^ in2[106];
    assign G[95] = in[105] & in2[105];
    assign P[95] = in[105] ^ in2[105];
    assign G[96] = in[104] & in2[104];
    assign P[96] = in[104] ^ in2[104];
    assign G[97] = in[103] & in2[103];
    assign P[97] = in[103] ^ in2[103];
    assign G[98] = in[102] & in2[102];
    assign P[98] = in[102] ^ in2[102];
    assign G[99] = in[101] & in2[101];
    assign P[99] = in[101] ^ in2[101];
    assign G[100] = in[100] & in2[100];
    assign P[100] = in[100] ^ in2[100];
    assign G[101] = in[99] & in2[99];
    assign P[101] = in[99] ^ in2[99];
    assign G[102] = in[98] & in2[98];
    assign P[102] = in[98] ^ in2[98];
    assign G[103] = in[97] & in2[97];
    assign P[103] = in[97] ^ in2[97];
    assign G[104] = in[96] & in2[96];
    assign P[104] = in[96] ^ in2[96];
    assign G[105] = in[95] & in2[95];
    assign P[105] = in[95] ^ in2[95];
    assign G[106] = in[94] & in2[94];
    assign P[106] = in[94] ^ in2[94];
    assign G[107] = in[93] & in2[93];
    assign P[107] = in[93] ^ in2[93];
    assign G[108] = in[92] & in2[92];
    assign P[108] = in[92] ^ in2[92];
    assign G[109] = in[91] & in2[91];
    assign P[109] = in[91] ^ in2[91];
    assign G[110] = in[90] & in2[90];
    assign P[110] = in[90] ^ in2[90];
    assign G[111] = in[89] & in2[89];
    assign P[111] = in[89] ^ in2[89];
    assign G[112] = in[88] & in2[88];
    assign P[112] = in[88] ^ in2[88];
    assign G[113] = in[87] & in2[87];
    assign P[113] = in[87] ^ in2[87];
    assign G[114] = in[86] & in2[86];
    assign P[114] = in[86] ^ in2[86];
    assign G[115] = in[85] & in2[85];
    assign P[115] = in[85] ^ in2[85];
    assign G[116] = in[84] & in2[84];
    assign P[116] = in[84] ^ in2[84];
    assign G[117] = in[83] & in2[83];
    assign P[117] = in[83] ^ in2[83];
    assign G[118] = in[82] & in2[82];
    assign P[118] = in[82] ^ in2[82];
    assign G[119] = in[81] & in2[81];
    assign P[119] = in[81] ^ in2[81];
    assign G[120] = in[80] & in2[80];
    assign P[120] = in[80] ^ in2[80];
    assign G[121] = in[79] & in2[79];
    assign P[121] = in[79] ^ in2[79];
    assign G[122] = in[78] & in2[78];
    assign P[122] = in[78] ^ in2[78];
    assign G[123] = in[77] & in2[77];
    assign P[123] = in[77] ^ in2[77];
    assign G[124] = in[76] & in2[76];
    assign P[124] = in[76] ^ in2[76];
    assign G[125] = in[75] & in2[75];
    assign P[125] = in[75] ^ in2[75];
    assign G[126] = in[74] & in2[74];
    assign P[126] = in[74] ^ in2[74];
    assign G[127] = in[73] & in2[73];
    assign P[127] = in[73] ^ in2[73];
    assign G[128] = in[72] & in2[72];
    assign P[128] = in[72] ^ in2[72];
    assign G[129] = in[71] & in2[71];
    assign P[129] = in[71] ^ in2[71];
    assign G[130] = in[70] & in2[70];
    assign P[130] = in[70] ^ in2[70];
    assign G[131] = in[69] & in2[69];
    assign P[131] = in[69] ^ in2[69];
    assign G[132] = in[68] & in2[68];
    assign P[132] = in[68] ^ in2[68];
    assign G[133] = in[67] & in2[67];
    assign P[133] = in[67] ^ in2[67];
    assign G[134] = in[66] & in2[66];
    assign P[134] = in[66] ^ in2[66];
    assign G[135] = in[65] & in2[65];
    assign P[135] = in[65] ^ in2[65];
    assign G[136] = in[64] & in2[64];
    assign P[136] = in[64] ^ in2[64];
    assign G[137] = in[63] & in2[63];
    assign P[137] = in[63] ^ in2[63];
    assign G[138] = in[62] & in2[62];
    assign P[138] = in[62] ^ in2[62];
    assign G[139] = in[61] & in2[61];
    assign P[139] = in[61] ^ in2[61];
    assign G[140] = in[60] & in2[60];
    assign P[140] = in[60] ^ in2[60];
    assign G[141] = in[59] & in2[59];
    assign P[141] = in[59] ^ in2[59];
    assign G[142] = in[58] & in2[58];
    assign P[142] = in[58] ^ in2[58];
    assign G[143] = in[57] & in2[57];
    assign P[143] = in[57] ^ in2[57];
    assign G[144] = in[56] & in2[56];
    assign P[144] = in[56] ^ in2[56];
    assign G[145] = in[55] & in2[55];
    assign P[145] = in[55] ^ in2[55];
    assign G[146] = in[54] & in2[54];
    assign P[146] = in[54] ^ in2[54];
    assign G[147] = in[53] & in2[53];
    assign P[147] = in[53] ^ in2[53];
    assign G[148] = in[52] & in2[52];
    assign P[148] = in[52] ^ in2[52];
    assign G[149] = in[51] & in2[51];
    assign P[149] = in[51] ^ in2[51];
    assign G[150] = in[50] & in2[50];
    assign P[150] = in[50] ^ in2[50];
    assign G[151] = in[49] & in2[49];
    assign P[151] = in[49] ^ in2[49];
    assign G[152] = in[48] & in2[48];
    assign P[152] = in[48] ^ in2[48];
    assign G[153] = in[47] & in2[47];
    assign P[153] = in[47] ^ in2[47];
    assign G[154] = in[46] & in2[46];
    assign P[154] = in[46] ^ in2[46];
    assign G[155] = in[45] & in2[45];
    assign P[155] = in[45] ^ in2[45];
    assign G[156] = in[44] & in2[44];
    assign P[156] = in[44] ^ in2[44];
    assign G[157] = in[43] & in2[43];
    assign P[157] = in[43] ^ in2[43];
    assign G[158] = in[42] & in2[42];
    assign P[158] = in[42] ^ in2[42];
    assign G[159] = in[41] & in2[41];
    assign P[159] = in[41] ^ in2[41];
    assign G[160] = in[40] & in2[40];
    assign P[160] = in[40] ^ in2[40];
    assign G[161] = in[39] & in2[39];
    assign P[161] = in[39] ^ in2[39];
    assign G[162] = in[38] & in2[38];
    assign P[162] = in[38] ^ in2[38];
    assign G[163] = in[37] & in2[37];
    assign P[163] = in[37] ^ in2[37];
    assign G[164] = in[36] & in2[36];
    assign P[164] = in[36] ^ in2[36];
    assign G[165] = in[35] & in2[35];
    assign P[165] = in[35] ^ in2[35];
    assign G[166] = in[34] & in2[34];
    assign P[166] = in[34] ^ in2[34];
    assign G[167] = in[33] & in2[33];
    assign P[167] = in[33] ^ in2[33];
    assign G[168] = in[32] & in2[32];
    assign P[168] = in[32] ^ in2[32];
    assign G[169] = in[31] & in2[31];
    assign P[169] = in[31] ^ in2[31];
    assign G[170] = in[30] & in2[30];
    assign P[170] = in[30] ^ in2[30];
    assign G[171] = in[29] & in2[29];
    assign P[171] = in[29] ^ in2[29];
    assign G[172] = in[28] & in2[28];
    assign P[172] = in[28] ^ in2[28];
    assign G[173] = in[27] & in2[27];
    assign P[173] = in[27] ^ in2[27];
    assign G[174] = in[26] & in2[26];
    assign P[174] = in[26] ^ in2[26];
    assign G[175] = in[25] & in2[25];
    assign P[175] = in[25] ^ in2[25];
    assign G[176] = in[24] & in2[24];
    assign P[176] = in[24] ^ in2[24];
    assign G[177] = in[23] & in2[23];
    assign P[177] = in[23] ^ in2[23];
    assign G[178] = in[22] & in2[22];
    assign P[178] = in[22] ^ in2[22];
    assign G[179] = in[21] & in2[21];
    assign P[179] = in[21] ^ in2[21];
    assign G[180] = in[20] & in2[20];
    assign P[180] = in[20] ^ in2[20];
    assign G[181] = in[19] & in2[19];
    assign P[181] = in[19] ^ in2[19];
    assign G[182] = in[18] & in2[18];
    assign P[182] = in[18] ^ in2[18];
    assign G[183] = in[17] & in2[17];
    assign P[183] = in[17] ^ in2[17];
    assign G[184] = in[16] & in2[16];
    assign P[184] = in[16] ^ in2[16];
    assign G[185] = in[15] & in2[15];
    assign P[185] = in[15] ^ in2[15];
    assign G[186] = in[14] & in2[14];
    assign P[186] = in[14] ^ in2[14];
    assign G[187] = in[13] & in2[13];
    assign P[187] = in[13] ^ in2[13];
    assign G[188] = in[12] & in2[12];
    assign P[188] = in[12] ^ in2[12];
    assign G[189] = in[11] & in2[11];
    assign P[189] = in[11] ^ in2[11];
    assign G[190] = in[10] & in2[10];
    assign P[190] = in[10] ^ in2[10];
    assign G[191] = in[9] & in2[9];
    assign P[191] = in[9] ^ in2[9];
    assign G[192] = in[8] & in2[8];
    assign P[192] = in[8] ^ in2[8];
    assign G[193] = in[7] & in2[7];
    assign P[193] = in[7] ^ in2[7];
    assign G[194] = in[6] & in2[6];
    assign P[194] = in[6] ^ in2[6];
    assign G[195] = in[5] & in2[5];
    assign P[195] = in[5] ^ in2[5];
    assign G[196] = in[4] & in2[4];
    assign P[196] = in[4] ^ in2[4];
    assign G[197] = in[3] & in2[3];
    assign P[197] = in[3] ^ in2[3];
    assign G[198] = in[2] & in2[2];
    assign P[198] = in[2] ^ in2[2];
    assign G[199] = in[1] & in2[1];
    assign P[199] = in[1] ^ in2[1];
    assign G[200] = in[0] & in2[0];
    assign P[200] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign C[200] = G[199] | (P[199] & C[199]);
    assign cout = G[200] | (P[200] & C[200]);
    assign sum = P ^ C;
endmodule

module CLA200(output [199:0] sum, output cout, input [199:0] in1, input [199:0] in2;

    wire[199:0] G;
    wire[199:0] C;
    wire[199:0] P;

    assign G[0] = in[199] & in2[199];
    assign P[0] = in[199] ^ in2[199];
    assign G[1] = in[198] & in2[198];
    assign P[1] = in[198] ^ in2[198];
    assign G[2] = in[197] & in2[197];
    assign P[2] = in[197] ^ in2[197];
    assign G[3] = in[196] & in2[196];
    assign P[3] = in[196] ^ in2[196];
    assign G[4] = in[195] & in2[195];
    assign P[4] = in[195] ^ in2[195];
    assign G[5] = in[194] & in2[194];
    assign P[5] = in[194] ^ in2[194];
    assign G[6] = in[193] & in2[193];
    assign P[6] = in[193] ^ in2[193];
    assign G[7] = in[192] & in2[192];
    assign P[7] = in[192] ^ in2[192];
    assign G[8] = in[191] & in2[191];
    assign P[8] = in[191] ^ in2[191];
    assign G[9] = in[190] & in2[190];
    assign P[9] = in[190] ^ in2[190];
    assign G[10] = in[189] & in2[189];
    assign P[10] = in[189] ^ in2[189];
    assign G[11] = in[188] & in2[188];
    assign P[11] = in[188] ^ in2[188];
    assign G[12] = in[187] & in2[187];
    assign P[12] = in[187] ^ in2[187];
    assign G[13] = in[186] & in2[186];
    assign P[13] = in[186] ^ in2[186];
    assign G[14] = in[185] & in2[185];
    assign P[14] = in[185] ^ in2[185];
    assign G[15] = in[184] & in2[184];
    assign P[15] = in[184] ^ in2[184];
    assign G[16] = in[183] & in2[183];
    assign P[16] = in[183] ^ in2[183];
    assign G[17] = in[182] & in2[182];
    assign P[17] = in[182] ^ in2[182];
    assign G[18] = in[181] & in2[181];
    assign P[18] = in[181] ^ in2[181];
    assign G[19] = in[180] & in2[180];
    assign P[19] = in[180] ^ in2[180];
    assign G[20] = in[179] & in2[179];
    assign P[20] = in[179] ^ in2[179];
    assign G[21] = in[178] & in2[178];
    assign P[21] = in[178] ^ in2[178];
    assign G[22] = in[177] & in2[177];
    assign P[22] = in[177] ^ in2[177];
    assign G[23] = in[176] & in2[176];
    assign P[23] = in[176] ^ in2[176];
    assign G[24] = in[175] & in2[175];
    assign P[24] = in[175] ^ in2[175];
    assign G[25] = in[174] & in2[174];
    assign P[25] = in[174] ^ in2[174];
    assign G[26] = in[173] & in2[173];
    assign P[26] = in[173] ^ in2[173];
    assign G[27] = in[172] & in2[172];
    assign P[27] = in[172] ^ in2[172];
    assign G[28] = in[171] & in2[171];
    assign P[28] = in[171] ^ in2[171];
    assign G[29] = in[170] & in2[170];
    assign P[29] = in[170] ^ in2[170];
    assign G[30] = in[169] & in2[169];
    assign P[30] = in[169] ^ in2[169];
    assign G[31] = in[168] & in2[168];
    assign P[31] = in[168] ^ in2[168];
    assign G[32] = in[167] & in2[167];
    assign P[32] = in[167] ^ in2[167];
    assign G[33] = in[166] & in2[166];
    assign P[33] = in[166] ^ in2[166];
    assign G[34] = in[165] & in2[165];
    assign P[34] = in[165] ^ in2[165];
    assign G[35] = in[164] & in2[164];
    assign P[35] = in[164] ^ in2[164];
    assign G[36] = in[163] & in2[163];
    assign P[36] = in[163] ^ in2[163];
    assign G[37] = in[162] & in2[162];
    assign P[37] = in[162] ^ in2[162];
    assign G[38] = in[161] & in2[161];
    assign P[38] = in[161] ^ in2[161];
    assign G[39] = in[160] & in2[160];
    assign P[39] = in[160] ^ in2[160];
    assign G[40] = in[159] & in2[159];
    assign P[40] = in[159] ^ in2[159];
    assign G[41] = in[158] & in2[158];
    assign P[41] = in[158] ^ in2[158];
    assign G[42] = in[157] & in2[157];
    assign P[42] = in[157] ^ in2[157];
    assign G[43] = in[156] & in2[156];
    assign P[43] = in[156] ^ in2[156];
    assign G[44] = in[155] & in2[155];
    assign P[44] = in[155] ^ in2[155];
    assign G[45] = in[154] & in2[154];
    assign P[45] = in[154] ^ in2[154];
    assign G[46] = in[153] & in2[153];
    assign P[46] = in[153] ^ in2[153];
    assign G[47] = in[152] & in2[152];
    assign P[47] = in[152] ^ in2[152];
    assign G[48] = in[151] & in2[151];
    assign P[48] = in[151] ^ in2[151];
    assign G[49] = in[150] & in2[150];
    assign P[49] = in[150] ^ in2[150];
    assign G[50] = in[149] & in2[149];
    assign P[50] = in[149] ^ in2[149];
    assign G[51] = in[148] & in2[148];
    assign P[51] = in[148] ^ in2[148];
    assign G[52] = in[147] & in2[147];
    assign P[52] = in[147] ^ in2[147];
    assign G[53] = in[146] & in2[146];
    assign P[53] = in[146] ^ in2[146];
    assign G[54] = in[145] & in2[145];
    assign P[54] = in[145] ^ in2[145];
    assign G[55] = in[144] & in2[144];
    assign P[55] = in[144] ^ in2[144];
    assign G[56] = in[143] & in2[143];
    assign P[56] = in[143] ^ in2[143];
    assign G[57] = in[142] & in2[142];
    assign P[57] = in[142] ^ in2[142];
    assign G[58] = in[141] & in2[141];
    assign P[58] = in[141] ^ in2[141];
    assign G[59] = in[140] & in2[140];
    assign P[59] = in[140] ^ in2[140];
    assign G[60] = in[139] & in2[139];
    assign P[60] = in[139] ^ in2[139];
    assign G[61] = in[138] & in2[138];
    assign P[61] = in[138] ^ in2[138];
    assign G[62] = in[137] & in2[137];
    assign P[62] = in[137] ^ in2[137];
    assign G[63] = in[136] & in2[136];
    assign P[63] = in[136] ^ in2[136];
    assign G[64] = in[135] & in2[135];
    assign P[64] = in[135] ^ in2[135];
    assign G[65] = in[134] & in2[134];
    assign P[65] = in[134] ^ in2[134];
    assign G[66] = in[133] & in2[133];
    assign P[66] = in[133] ^ in2[133];
    assign G[67] = in[132] & in2[132];
    assign P[67] = in[132] ^ in2[132];
    assign G[68] = in[131] & in2[131];
    assign P[68] = in[131] ^ in2[131];
    assign G[69] = in[130] & in2[130];
    assign P[69] = in[130] ^ in2[130];
    assign G[70] = in[129] & in2[129];
    assign P[70] = in[129] ^ in2[129];
    assign G[71] = in[128] & in2[128];
    assign P[71] = in[128] ^ in2[128];
    assign G[72] = in[127] & in2[127];
    assign P[72] = in[127] ^ in2[127];
    assign G[73] = in[126] & in2[126];
    assign P[73] = in[126] ^ in2[126];
    assign G[74] = in[125] & in2[125];
    assign P[74] = in[125] ^ in2[125];
    assign G[75] = in[124] & in2[124];
    assign P[75] = in[124] ^ in2[124];
    assign G[76] = in[123] & in2[123];
    assign P[76] = in[123] ^ in2[123];
    assign G[77] = in[122] & in2[122];
    assign P[77] = in[122] ^ in2[122];
    assign G[78] = in[121] & in2[121];
    assign P[78] = in[121] ^ in2[121];
    assign G[79] = in[120] & in2[120];
    assign P[79] = in[120] ^ in2[120];
    assign G[80] = in[119] & in2[119];
    assign P[80] = in[119] ^ in2[119];
    assign G[81] = in[118] & in2[118];
    assign P[81] = in[118] ^ in2[118];
    assign G[82] = in[117] & in2[117];
    assign P[82] = in[117] ^ in2[117];
    assign G[83] = in[116] & in2[116];
    assign P[83] = in[116] ^ in2[116];
    assign G[84] = in[115] & in2[115];
    assign P[84] = in[115] ^ in2[115];
    assign G[85] = in[114] & in2[114];
    assign P[85] = in[114] ^ in2[114];
    assign G[86] = in[113] & in2[113];
    assign P[86] = in[113] ^ in2[113];
    assign G[87] = in[112] & in2[112];
    assign P[87] = in[112] ^ in2[112];
    assign G[88] = in[111] & in2[111];
    assign P[88] = in[111] ^ in2[111];
    assign G[89] = in[110] & in2[110];
    assign P[89] = in[110] ^ in2[110];
    assign G[90] = in[109] & in2[109];
    assign P[90] = in[109] ^ in2[109];
    assign G[91] = in[108] & in2[108];
    assign P[91] = in[108] ^ in2[108];
    assign G[92] = in[107] & in2[107];
    assign P[92] = in[107] ^ in2[107];
    assign G[93] = in[106] & in2[106];
    assign P[93] = in[106] ^ in2[106];
    assign G[94] = in[105] & in2[105];
    assign P[94] = in[105] ^ in2[105];
    assign G[95] = in[104] & in2[104];
    assign P[95] = in[104] ^ in2[104];
    assign G[96] = in[103] & in2[103];
    assign P[96] = in[103] ^ in2[103];
    assign G[97] = in[102] & in2[102];
    assign P[97] = in[102] ^ in2[102];
    assign G[98] = in[101] & in2[101];
    assign P[98] = in[101] ^ in2[101];
    assign G[99] = in[100] & in2[100];
    assign P[99] = in[100] ^ in2[100];
    assign G[100] = in[99] & in2[99];
    assign P[100] = in[99] ^ in2[99];
    assign G[101] = in[98] & in2[98];
    assign P[101] = in[98] ^ in2[98];
    assign G[102] = in[97] & in2[97];
    assign P[102] = in[97] ^ in2[97];
    assign G[103] = in[96] & in2[96];
    assign P[103] = in[96] ^ in2[96];
    assign G[104] = in[95] & in2[95];
    assign P[104] = in[95] ^ in2[95];
    assign G[105] = in[94] & in2[94];
    assign P[105] = in[94] ^ in2[94];
    assign G[106] = in[93] & in2[93];
    assign P[106] = in[93] ^ in2[93];
    assign G[107] = in[92] & in2[92];
    assign P[107] = in[92] ^ in2[92];
    assign G[108] = in[91] & in2[91];
    assign P[108] = in[91] ^ in2[91];
    assign G[109] = in[90] & in2[90];
    assign P[109] = in[90] ^ in2[90];
    assign G[110] = in[89] & in2[89];
    assign P[110] = in[89] ^ in2[89];
    assign G[111] = in[88] & in2[88];
    assign P[111] = in[88] ^ in2[88];
    assign G[112] = in[87] & in2[87];
    assign P[112] = in[87] ^ in2[87];
    assign G[113] = in[86] & in2[86];
    assign P[113] = in[86] ^ in2[86];
    assign G[114] = in[85] & in2[85];
    assign P[114] = in[85] ^ in2[85];
    assign G[115] = in[84] & in2[84];
    assign P[115] = in[84] ^ in2[84];
    assign G[116] = in[83] & in2[83];
    assign P[116] = in[83] ^ in2[83];
    assign G[117] = in[82] & in2[82];
    assign P[117] = in[82] ^ in2[82];
    assign G[118] = in[81] & in2[81];
    assign P[118] = in[81] ^ in2[81];
    assign G[119] = in[80] & in2[80];
    assign P[119] = in[80] ^ in2[80];
    assign G[120] = in[79] & in2[79];
    assign P[120] = in[79] ^ in2[79];
    assign G[121] = in[78] & in2[78];
    assign P[121] = in[78] ^ in2[78];
    assign G[122] = in[77] & in2[77];
    assign P[122] = in[77] ^ in2[77];
    assign G[123] = in[76] & in2[76];
    assign P[123] = in[76] ^ in2[76];
    assign G[124] = in[75] & in2[75];
    assign P[124] = in[75] ^ in2[75];
    assign G[125] = in[74] & in2[74];
    assign P[125] = in[74] ^ in2[74];
    assign G[126] = in[73] & in2[73];
    assign P[126] = in[73] ^ in2[73];
    assign G[127] = in[72] & in2[72];
    assign P[127] = in[72] ^ in2[72];
    assign G[128] = in[71] & in2[71];
    assign P[128] = in[71] ^ in2[71];
    assign G[129] = in[70] & in2[70];
    assign P[129] = in[70] ^ in2[70];
    assign G[130] = in[69] & in2[69];
    assign P[130] = in[69] ^ in2[69];
    assign G[131] = in[68] & in2[68];
    assign P[131] = in[68] ^ in2[68];
    assign G[132] = in[67] & in2[67];
    assign P[132] = in[67] ^ in2[67];
    assign G[133] = in[66] & in2[66];
    assign P[133] = in[66] ^ in2[66];
    assign G[134] = in[65] & in2[65];
    assign P[134] = in[65] ^ in2[65];
    assign G[135] = in[64] & in2[64];
    assign P[135] = in[64] ^ in2[64];
    assign G[136] = in[63] & in2[63];
    assign P[136] = in[63] ^ in2[63];
    assign G[137] = in[62] & in2[62];
    assign P[137] = in[62] ^ in2[62];
    assign G[138] = in[61] & in2[61];
    assign P[138] = in[61] ^ in2[61];
    assign G[139] = in[60] & in2[60];
    assign P[139] = in[60] ^ in2[60];
    assign G[140] = in[59] & in2[59];
    assign P[140] = in[59] ^ in2[59];
    assign G[141] = in[58] & in2[58];
    assign P[141] = in[58] ^ in2[58];
    assign G[142] = in[57] & in2[57];
    assign P[142] = in[57] ^ in2[57];
    assign G[143] = in[56] & in2[56];
    assign P[143] = in[56] ^ in2[56];
    assign G[144] = in[55] & in2[55];
    assign P[144] = in[55] ^ in2[55];
    assign G[145] = in[54] & in2[54];
    assign P[145] = in[54] ^ in2[54];
    assign G[146] = in[53] & in2[53];
    assign P[146] = in[53] ^ in2[53];
    assign G[147] = in[52] & in2[52];
    assign P[147] = in[52] ^ in2[52];
    assign G[148] = in[51] & in2[51];
    assign P[148] = in[51] ^ in2[51];
    assign G[149] = in[50] & in2[50];
    assign P[149] = in[50] ^ in2[50];
    assign G[150] = in[49] & in2[49];
    assign P[150] = in[49] ^ in2[49];
    assign G[151] = in[48] & in2[48];
    assign P[151] = in[48] ^ in2[48];
    assign G[152] = in[47] & in2[47];
    assign P[152] = in[47] ^ in2[47];
    assign G[153] = in[46] & in2[46];
    assign P[153] = in[46] ^ in2[46];
    assign G[154] = in[45] & in2[45];
    assign P[154] = in[45] ^ in2[45];
    assign G[155] = in[44] & in2[44];
    assign P[155] = in[44] ^ in2[44];
    assign G[156] = in[43] & in2[43];
    assign P[156] = in[43] ^ in2[43];
    assign G[157] = in[42] & in2[42];
    assign P[157] = in[42] ^ in2[42];
    assign G[158] = in[41] & in2[41];
    assign P[158] = in[41] ^ in2[41];
    assign G[159] = in[40] & in2[40];
    assign P[159] = in[40] ^ in2[40];
    assign G[160] = in[39] & in2[39];
    assign P[160] = in[39] ^ in2[39];
    assign G[161] = in[38] & in2[38];
    assign P[161] = in[38] ^ in2[38];
    assign G[162] = in[37] & in2[37];
    assign P[162] = in[37] ^ in2[37];
    assign G[163] = in[36] & in2[36];
    assign P[163] = in[36] ^ in2[36];
    assign G[164] = in[35] & in2[35];
    assign P[164] = in[35] ^ in2[35];
    assign G[165] = in[34] & in2[34];
    assign P[165] = in[34] ^ in2[34];
    assign G[166] = in[33] & in2[33];
    assign P[166] = in[33] ^ in2[33];
    assign G[167] = in[32] & in2[32];
    assign P[167] = in[32] ^ in2[32];
    assign G[168] = in[31] & in2[31];
    assign P[168] = in[31] ^ in2[31];
    assign G[169] = in[30] & in2[30];
    assign P[169] = in[30] ^ in2[30];
    assign G[170] = in[29] & in2[29];
    assign P[170] = in[29] ^ in2[29];
    assign G[171] = in[28] & in2[28];
    assign P[171] = in[28] ^ in2[28];
    assign G[172] = in[27] & in2[27];
    assign P[172] = in[27] ^ in2[27];
    assign G[173] = in[26] & in2[26];
    assign P[173] = in[26] ^ in2[26];
    assign G[174] = in[25] & in2[25];
    assign P[174] = in[25] ^ in2[25];
    assign G[175] = in[24] & in2[24];
    assign P[175] = in[24] ^ in2[24];
    assign G[176] = in[23] & in2[23];
    assign P[176] = in[23] ^ in2[23];
    assign G[177] = in[22] & in2[22];
    assign P[177] = in[22] ^ in2[22];
    assign G[178] = in[21] & in2[21];
    assign P[178] = in[21] ^ in2[21];
    assign G[179] = in[20] & in2[20];
    assign P[179] = in[20] ^ in2[20];
    assign G[180] = in[19] & in2[19];
    assign P[180] = in[19] ^ in2[19];
    assign G[181] = in[18] & in2[18];
    assign P[181] = in[18] ^ in2[18];
    assign G[182] = in[17] & in2[17];
    assign P[182] = in[17] ^ in2[17];
    assign G[183] = in[16] & in2[16];
    assign P[183] = in[16] ^ in2[16];
    assign G[184] = in[15] & in2[15];
    assign P[184] = in[15] ^ in2[15];
    assign G[185] = in[14] & in2[14];
    assign P[185] = in[14] ^ in2[14];
    assign G[186] = in[13] & in2[13];
    assign P[186] = in[13] ^ in2[13];
    assign G[187] = in[12] & in2[12];
    assign P[187] = in[12] ^ in2[12];
    assign G[188] = in[11] & in2[11];
    assign P[188] = in[11] ^ in2[11];
    assign G[189] = in[10] & in2[10];
    assign P[189] = in[10] ^ in2[10];
    assign G[190] = in[9] & in2[9];
    assign P[190] = in[9] ^ in2[9];
    assign G[191] = in[8] & in2[8];
    assign P[191] = in[8] ^ in2[8];
    assign G[192] = in[7] & in2[7];
    assign P[192] = in[7] ^ in2[7];
    assign G[193] = in[6] & in2[6];
    assign P[193] = in[6] ^ in2[6];
    assign G[194] = in[5] & in2[5];
    assign P[194] = in[5] ^ in2[5];
    assign G[195] = in[4] & in2[4];
    assign P[195] = in[4] ^ in2[4];
    assign G[196] = in[3] & in2[3];
    assign P[196] = in[3] ^ in2[3];
    assign G[197] = in[2] & in2[2];
    assign P[197] = in[2] ^ in2[2];
    assign G[198] = in[1] & in2[1];
    assign P[198] = in[1] ^ in2[1];
    assign G[199] = in[0] & in2[0];
    assign P[199] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign C[199] = G[198] | (P[198] & C[198]);
    assign cout = G[199] | (P[199] & C[199]);
    assign sum = P ^ C;
endmodule

module CLA199(output [198:0] sum, output cout, input [198:0] in1, input [198:0] in2;

    wire[198:0] G;
    wire[198:0] C;
    wire[198:0] P;

    assign G[0] = in[198] & in2[198];
    assign P[0] = in[198] ^ in2[198];
    assign G[1] = in[197] & in2[197];
    assign P[1] = in[197] ^ in2[197];
    assign G[2] = in[196] & in2[196];
    assign P[2] = in[196] ^ in2[196];
    assign G[3] = in[195] & in2[195];
    assign P[3] = in[195] ^ in2[195];
    assign G[4] = in[194] & in2[194];
    assign P[4] = in[194] ^ in2[194];
    assign G[5] = in[193] & in2[193];
    assign P[5] = in[193] ^ in2[193];
    assign G[6] = in[192] & in2[192];
    assign P[6] = in[192] ^ in2[192];
    assign G[7] = in[191] & in2[191];
    assign P[7] = in[191] ^ in2[191];
    assign G[8] = in[190] & in2[190];
    assign P[8] = in[190] ^ in2[190];
    assign G[9] = in[189] & in2[189];
    assign P[9] = in[189] ^ in2[189];
    assign G[10] = in[188] & in2[188];
    assign P[10] = in[188] ^ in2[188];
    assign G[11] = in[187] & in2[187];
    assign P[11] = in[187] ^ in2[187];
    assign G[12] = in[186] & in2[186];
    assign P[12] = in[186] ^ in2[186];
    assign G[13] = in[185] & in2[185];
    assign P[13] = in[185] ^ in2[185];
    assign G[14] = in[184] & in2[184];
    assign P[14] = in[184] ^ in2[184];
    assign G[15] = in[183] & in2[183];
    assign P[15] = in[183] ^ in2[183];
    assign G[16] = in[182] & in2[182];
    assign P[16] = in[182] ^ in2[182];
    assign G[17] = in[181] & in2[181];
    assign P[17] = in[181] ^ in2[181];
    assign G[18] = in[180] & in2[180];
    assign P[18] = in[180] ^ in2[180];
    assign G[19] = in[179] & in2[179];
    assign P[19] = in[179] ^ in2[179];
    assign G[20] = in[178] & in2[178];
    assign P[20] = in[178] ^ in2[178];
    assign G[21] = in[177] & in2[177];
    assign P[21] = in[177] ^ in2[177];
    assign G[22] = in[176] & in2[176];
    assign P[22] = in[176] ^ in2[176];
    assign G[23] = in[175] & in2[175];
    assign P[23] = in[175] ^ in2[175];
    assign G[24] = in[174] & in2[174];
    assign P[24] = in[174] ^ in2[174];
    assign G[25] = in[173] & in2[173];
    assign P[25] = in[173] ^ in2[173];
    assign G[26] = in[172] & in2[172];
    assign P[26] = in[172] ^ in2[172];
    assign G[27] = in[171] & in2[171];
    assign P[27] = in[171] ^ in2[171];
    assign G[28] = in[170] & in2[170];
    assign P[28] = in[170] ^ in2[170];
    assign G[29] = in[169] & in2[169];
    assign P[29] = in[169] ^ in2[169];
    assign G[30] = in[168] & in2[168];
    assign P[30] = in[168] ^ in2[168];
    assign G[31] = in[167] & in2[167];
    assign P[31] = in[167] ^ in2[167];
    assign G[32] = in[166] & in2[166];
    assign P[32] = in[166] ^ in2[166];
    assign G[33] = in[165] & in2[165];
    assign P[33] = in[165] ^ in2[165];
    assign G[34] = in[164] & in2[164];
    assign P[34] = in[164] ^ in2[164];
    assign G[35] = in[163] & in2[163];
    assign P[35] = in[163] ^ in2[163];
    assign G[36] = in[162] & in2[162];
    assign P[36] = in[162] ^ in2[162];
    assign G[37] = in[161] & in2[161];
    assign P[37] = in[161] ^ in2[161];
    assign G[38] = in[160] & in2[160];
    assign P[38] = in[160] ^ in2[160];
    assign G[39] = in[159] & in2[159];
    assign P[39] = in[159] ^ in2[159];
    assign G[40] = in[158] & in2[158];
    assign P[40] = in[158] ^ in2[158];
    assign G[41] = in[157] & in2[157];
    assign P[41] = in[157] ^ in2[157];
    assign G[42] = in[156] & in2[156];
    assign P[42] = in[156] ^ in2[156];
    assign G[43] = in[155] & in2[155];
    assign P[43] = in[155] ^ in2[155];
    assign G[44] = in[154] & in2[154];
    assign P[44] = in[154] ^ in2[154];
    assign G[45] = in[153] & in2[153];
    assign P[45] = in[153] ^ in2[153];
    assign G[46] = in[152] & in2[152];
    assign P[46] = in[152] ^ in2[152];
    assign G[47] = in[151] & in2[151];
    assign P[47] = in[151] ^ in2[151];
    assign G[48] = in[150] & in2[150];
    assign P[48] = in[150] ^ in2[150];
    assign G[49] = in[149] & in2[149];
    assign P[49] = in[149] ^ in2[149];
    assign G[50] = in[148] & in2[148];
    assign P[50] = in[148] ^ in2[148];
    assign G[51] = in[147] & in2[147];
    assign P[51] = in[147] ^ in2[147];
    assign G[52] = in[146] & in2[146];
    assign P[52] = in[146] ^ in2[146];
    assign G[53] = in[145] & in2[145];
    assign P[53] = in[145] ^ in2[145];
    assign G[54] = in[144] & in2[144];
    assign P[54] = in[144] ^ in2[144];
    assign G[55] = in[143] & in2[143];
    assign P[55] = in[143] ^ in2[143];
    assign G[56] = in[142] & in2[142];
    assign P[56] = in[142] ^ in2[142];
    assign G[57] = in[141] & in2[141];
    assign P[57] = in[141] ^ in2[141];
    assign G[58] = in[140] & in2[140];
    assign P[58] = in[140] ^ in2[140];
    assign G[59] = in[139] & in2[139];
    assign P[59] = in[139] ^ in2[139];
    assign G[60] = in[138] & in2[138];
    assign P[60] = in[138] ^ in2[138];
    assign G[61] = in[137] & in2[137];
    assign P[61] = in[137] ^ in2[137];
    assign G[62] = in[136] & in2[136];
    assign P[62] = in[136] ^ in2[136];
    assign G[63] = in[135] & in2[135];
    assign P[63] = in[135] ^ in2[135];
    assign G[64] = in[134] & in2[134];
    assign P[64] = in[134] ^ in2[134];
    assign G[65] = in[133] & in2[133];
    assign P[65] = in[133] ^ in2[133];
    assign G[66] = in[132] & in2[132];
    assign P[66] = in[132] ^ in2[132];
    assign G[67] = in[131] & in2[131];
    assign P[67] = in[131] ^ in2[131];
    assign G[68] = in[130] & in2[130];
    assign P[68] = in[130] ^ in2[130];
    assign G[69] = in[129] & in2[129];
    assign P[69] = in[129] ^ in2[129];
    assign G[70] = in[128] & in2[128];
    assign P[70] = in[128] ^ in2[128];
    assign G[71] = in[127] & in2[127];
    assign P[71] = in[127] ^ in2[127];
    assign G[72] = in[126] & in2[126];
    assign P[72] = in[126] ^ in2[126];
    assign G[73] = in[125] & in2[125];
    assign P[73] = in[125] ^ in2[125];
    assign G[74] = in[124] & in2[124];
    assign P[74] = in[124] ^ in2[124];
    assign G[75] = in[123] & in2[123];
    assign P[75] = in[123] ^ in2[123];
    assign G[76] = in[122] & in2[122];
    assign P[76] = in[122] ^ in2[122];
    assign G[77] = in[121] & in2[121];
    assign P[77] = in[121] ^ in2[121];
    assign G[78] = in[120] & in2[120];
    assign P[78] = in[120] ^ in2[120];
    assign G[79] = in[119] & in2[119];
    assign P[79] = in[119] ^ in2[119];
    assign G[80] = in[118] & in2[118];
    assign P[80] = in[118] ^ in2[118];
    assign G[81] = in[117] & in2[117];
    assign P[81] = in[117] ^ in2[117];
    assign G[82] = in[116] & in2[116];
    assign P[82] = in[116] ^ in2[116];
    assign G[83] = in[115] & in2[115];
    assign P[83] = in[115] ^ in2[115];
    assign G[84] = in[114] & in2[114];
    assign P[84] = in[114] ^ in2[114];
    assign G[85] = in[113] & in2[113];
    assign P[85] = in[113] ^ in2[113];
    assign G[86] = in[112] & in2[112];
    assign P[86] = in[112] ^ in2[112];
    assign G[87] = in[111] & in2[111];
    assign P[87] = in[111] ^ in2[111];
    assign G[88] = in[110] & in2[110];
    assign P[88] = in[110] ^ in2[110];
    assign G[89] = in[109] & in2[109];
    assign P[89] = in[109] ^ in2[109];
    assign G[90] = in[108] & in2[108];
    assign P[90] = in[108] ^ in2[108];
    assign G[91] = in[107] & in2[107];
    assign P[91] = in[107] ^ in2[107];
    assign G[92] = in[106] & in2[106];
    assign P[92] = in[106] ^ in2[106];
    assign G[93] = in[105] & in2[105];
    assign P[93] = in[105] ^ in2[105];
    assign G[94] = in[104] & in2[104];
    assign P[94] = in[104] ^ in2[104];
    assign G[95] = in[103] & in2[103];
    assign P[95] = in[103] ^ in2[103];
    assign G[96] = in[102] & in2[102];
    assign P[96] = in[102] ^ in2[102];
    assign G[97] = in[101] & in2[101];
    assign P[97] = in[101] ^ in2[101];
    assign G[98] = in[100] & in2[100];
    assign P[98] = in[100] ^ in2[100];
    assign G[99] = in[99] & in2[99];
    assign P[99] = in[99] ^ in2[99];
    assign G[100] = in[98] & in2[98];
    assign P[100] = in[98] ^ in2[98];
    assign G[101] = in[97] & in2[97];
    assign P[101] = in[97] ^ in2[97];
    assign G[102] = in[96] & in2[96];
    assign P[102] = in[96] ^ in2[96];
    assign G[103] = in[95] & in2[95];
    assign P[103] = in[95] ^ in2[95];
    assign G[104] = in[94] & in2[94];
    assign P[104] = in[94] ^ in2[94];
    assign G[105] = in[93] & in2[93];
    assign P[105] = in[93] ^ in2[93];
    assign G[106] = in[92] & in2[92];
    assign P[106] = in[92] ^ in2[92];
    assign G[107] = in[91] & in2[91];
    assign P[107] = in[91] ^ in2[91];
    assign G[108] = in[90] & in2[90];
    assign P[108] = in[90] ^ in2[90];
    assign G[109] = in[89] & in2[89];
    assign P[109] = in[89] ^ in2[89];
    assign G[110] = in[88] & in2[88];
    assign P[110] = in[88] ^ in2[88];
    assign G[111] = in[87] & in2[87];
    assign P[111] = in[87] ^ in2[87];
    assign G[112] = in[86] & in2[86];
    assign P[112] = in[86] ^ in2[86];
    assign G[113] = in[85] & in2[85];
    assign P[113] = in[85] ^ in2[85];
    assign G[114] = in[84] & in2[84];
    assign P[114] = in[84] ^ in2[84];
    assign G[115] = in[83] & in2[83];
    assign P[115] = in[83] ^ in2[83];
    assign G[116] = in[82] & in2[82];
    assign P[116] = in[82] ^ in2[82];
    assign G[117] = in[81] & in2[81];
    assign P[117] = in[81] ^ in2[81];
    assign G[118] = in[80] & in2[80];
    assign P[118] = in[80] ^ in2[80];
    assign G[119] = in[79] & in2[79];
    assign P[119] = in[79] ^ in2[79];
    assign G[120] = in[78] & in2[78];
    assign P[120] = in[78] ^ in2[78];
    assign G[121] = in[77] & in2[77];
    assign P[121] = in[77] ^ in2[77];
    assign G[122] = in[76] & in2[76];
    assign P[122] = in[76] ^ in2[76];
    assign G[123] = in[75] & in2[75];
    assign P[123] = in[75] ^ in2[75];
    assign G[124] = in[74] & in2[74];
    assign P[124] = in[74] ^ in2[74];
    assign G[125] = in[73] & in2[73];
    assign P[125] = in[73] ^ in2[73];
    assign G[126] = in[72] & in2[72];
    assign P[126] = in[72] ^ in2[72];
    assign G[127] = in[71] & in2[71];
    assign P[127] = in[71] ^ in2[71];
    assign G[128] = in[70] & in2[70];
    assign P[128] = in[70] ^ in2[70];
    assign G[129] = in[69] & in2[69];
    assign P[129] = in[69] ^ in2[69];
    assign G[130] = in[68] & in2[68];
    assign P[130] = in[68] ^ in2[68];
    assign G[131] = in[67] & in2[67];
    assign P[131] = in[67] ^ in2[67];
    assign G[132] = in[66] & in2[66];
    assign P[132] = in[66] ^ in2[66];
    assign G[133] = in[65] & in2[65];
    assign P[133] = in[65] ^ in2[65];
    assign G[134] = in[64] & in2[64];
    assign P[134] = in[64] ^ in2[64];
    assign G[135] = in[63] & in2[63];
    assign P[135] = in[63] ^ in2[63];
    assign G[136] = in[62] & in2[62];
    assign P[136] = in[62] ^ in2[62];
    assign G[137] = in[61] & in2[61];
    assign P[137] = in[61] ^ in2[61];
    assign G[138] = in[60] & in2[60];
    assign P[138] = in[60] ^ in2[60];
    assign G[139] = in[59] & in2[59];
    assign P[139] = in[59] ^ in2[59];
    assign G[140] = in[58] & in2[58];
    assign P[140] = in[58] ^ in2[58];
    assign G[141] = in[57] & in2[57];
    assign P[141] = in[57] ^ in2[57];
    assign G[142] = in[56] & in2[56];
    assign P[142] = in[56] ^ in2[56];
    assign G[143] = in[55] & in2[55];
    assign P[143] = in[55] ^ in2[55];
    assign G[144] = in[54] & in2[54];
    assign P[144] = in[54] ^ in2[54];
    assign G[145] = in[53] & in2[53];
    assign P[145] = in[53] ^ in2[53];
    assign G[146] = in[52] & in2[52];
    assign P[146] = in[52] ^ in2[52];
    assign G[147] = in[51] & in2[51];
    assign P[147] = in[51] ^ in2[51];
    assign G[148] = in[50] & in2[50];
    assign P[148] = in[50] ^ in2[50];
    assign G[149] = in[49] & in2[49];
    assign P[149] = in[49] ^ in2[49];
    assign G[150] = in[48] & in2[48];
    assign P[150] = in[48] ^ in2[48];
    assign G[151] = in[47] & in2[47];
    assign P[151] = in[47] ^ in2[47];
    assign G[152] = in[46] & in2[46];
    assign P[152] = in[46] ^ in2[46];
    assign G[153] = in[45] & in2[45];
    assign P[153] = in[45] ^ in2[45];
    assign G[154] = in[44] & in2[44];
    assign P[154] = in[44] ^ in2[44];
    assign G[155] = in[43] & in2[43];
    assign P[155] = in[43] ^ in2[43];
    assign G[156] = in[42] & in2[42];
    assign P[156] = in[42] ^ in2[42];
    assign G[157] = in[41] & in2[41];
    assign P[157] = in[41] ^ in2[41];
    assign G[158] = in[40] & in2[40];
    assign P[158] = in[40] ^ in2[40];
    assign G[159] = in[39] & in2[39];
    assign P[159] = in[39] ^ in2[39];
    assign G[160] = in[38] & in2[38];
    assign P[160] = in[38] ^ in2[38];
    assign G[161] = in[37] & in2[37];
    assign P[161] = in[37] ^ in2[37];
    assign G[162] = in[36] & in2[36];
    assign P[162] = in[36] ^ in2[36];
    assign G[163] = in[35] & in2[35];
    assign P[163] = in[35] ^ in2[35];
    assign G[164] = in[34] & in2[34];
    assign P[164] = in[34] ^ in2[34];
    assign G[165] = in[33] & in2[33];
    assign P[165] = in[33] ^ in2[33];
    assign G[166] = in[32] & in2[32];
    assign P[166] = in[32] ^ in2[32];
    assign G[167] = in[31] & in2[31];
    assign P[167] = in[31] ^ in2[31];
    assign G[168] = in[30] & in2[30];
    assign P[168] = in[30] ^ in2[30];
    assign G[169] = in[29] & in2[29];
    assign P[169] = in[29] ^ in2[29];
    assign G[170] = in[28] & in2[28];
    assign P[170] = in[28] ^ in2[28];
    assign G[171] = in[27] & in2[27];
    assign P[171] = in[27] ^ in2[27];
    assign G[172] = in[26] & in2[26];
    assign P[172] = in[26] ^ in2[26];
    assign G[173] = in[25] & in2[25];
    assign P[173] = in[25] ^ in2[25];
    assign G[174] = in[24] & in2[24];
    assign P[174] = in[24] ^ in2[24];
    assign G[175] = in[23] & in2[23];
    assign P[175] = in[23] ^ in2[23];
    assign G[176] = in[22] & in2[22];
    assign P[176] = in[22] ^ in2[22];
    assign G[177] = in[21] & in2[21];
    assign P[177] = in[21] ^ in2[21];
    assign G[178] = in[20] & in2[20];
    assign P[178] = in[20] ^ in2[20];
    assign G[179] = in[19] & in2[19];
    assign P[179] = in[19] ^ in2[19];
    assign G[180] = in[18] & in2[18];
    assign P[180] = in[18] ^ in2[18];
    assign G[181] = in[17] & in2[17];
    assign P[181] = in[17] ^ in2[17];
    assign G[182] = in[16] & in2[16];
    assign P[182] = in[16] ^ in2[16];
    assign G[183] = in[15] & in2[15];
    assign P[183] = in[15] ^ in2[15];
    assign G[184] = in[14] & in2[14];
    assign P[184] = in[14] ^ in2[14];
    assign G[185] = in[13] & in2[13];
    assign P[185] = in[13] ^ in2[13];
    assign G[186] = in[12] & in2[12];
    assign P[186] = in[12] ^ in2[12];
    assign G[187] = in[11] & in2[11];
    assign P[187] = in[11] ^ in2[11];
    assign G[188] = in[10] & in2[10];
    assign P[188] = in[10] ^ in2[10];
    assign G[189] = in[9] & in2[9];
    assign P[189] = in[9] ^ in2[9];
    assign G[190] = in[8] & in2[8];
    assign P[190] = in[8] ^ in2[8];
    assign G[191] = in[7] & in2[7];
    assign P[191] = in[7] ^ in2[7];
    assign G[192] = in[6] & in2[6];
    assign P[192] = in[6] ^ in2[6];
    assign G[193] = in[5] & in2[5];
    assign P[193] = in[5] ^ in2[5];
    assign G[194] = in[4] & in2[4];
    assign P[194] = in[4] ^ in2[4];
    assign G[195] = in[3] & in2[3];
    assign P[195] = in[3] ^ in2[3];
    assign G[196] = in[2] & in2[2];
    assign P[196] = in[2] ^ in2[2];
    assign G[197] = in[1] & in2[1];
    assign P[197] = in[1] ^ in2[1];
    assign G[198] = in[0] & in2[0];
    assign P[198] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign C[198] = G[197] | (P[197] & C[197]);
    assign cout = G[198] | (P[198] & C[198]);
    assign sum = P ^ C;
endmodule

module CLA198(output [197:0] sum, output cout, input [197:0] in1, input [197:0] in2;

    wire[197:0] G;
    wire[197:0] C;
    wire[197:0] P;

    assign G[0] = in[197] & in2[197];
    assign P[0] = in[197] ^ in2[197];
    assign G[1] = in[196] & in2[196];
    assign P[1] = in[196] ^ in2[196];
    assign G[2] = in[195] & in2[195];
    assign P[2] = in[195] ^ in2[195];
    assign G[3] = in[194] & in2[194];
    assign P[3] = in[194] ^ in2[194];
    assign G[4] = in[193] & in2[193];
    assign P[4] = in[193] ^ in2[193];
    assign G[5] = in[192] & in2[192];
    assign P[5] = in[192] ^ in2[192];
    assign G[6] = in[191] & in2[191];
    assign P[6] = in[191] ^ in2[191];
    assign G[7] = in[190] & in2[190];
    assign P[7] = in[190] ^ in2[190];
    assign G[8] = in[189] & in2[189];
    assign P[8] = in[189] ^ in2[189];
    assign G[9] = in[188] & in2[188];
    assign P[9] = in[188] ^ in2[188];
    assign G[10] = in[187] & in2[187];
    assign P[10] = in[187] ^ in2[187];
    assign G[11] = in[186] & in2[186];
    assign P[11] = in[186] ^ in2[186];
    assign G[12] = in[185] & in2[185];
    assign P[12] = in[185] ^ in2[185];
    assign G[13] = in[184] & in2[184];
    assign P[13] = in[184] ^ in2[184];
    assign G[14] = in[183] & in2[183];
    assign P[14] = in[183] ^ in2[183];
    assign G[15] = in[182] & in2[182];
    assign P[15] = in[182] ^ in2[182];
    assign G[16] = in[181] & in2[181];
    assign P[16] = in[181] ^ in2[181];
    assign G[17] = in[180] & in2[180];
    assign P[17] = in[180] ^ in2[180];
    assign G[18] = in[179] & in2[179];
    assign P[18] = in[179] ^ in2[179];
    assign G[19] = in[178] & in2[178];
    assign P[19] = in[178] ^ in2[178];
    assign G[20] = in[177] & in2[177];
    assign P[20] = in[177] ^ in2[177];
    assign G[21] = in[176] & in2[176];
    assign P[21] = in[176] ^ in2[176];
    assign G[22] = in[175] & in2[175];
    assign P[22] = in[175] ^ in2[175];
    assign G[23] = in[174] & in2[174];
    assign P[23] = in[174] ^ in2[174];
    assign G[24] = in[173] & in2[173];
    assign P[24] = in[173] ^ in2[173];
    assign G[25] = in[172] & in2[172];
    assign P[25] = in[172] ^ in2[172];
    assign G[26] = in[171] & in2[171];
    assign P[26] = in[171] ^ in2[171];
    assign G[27] = in[170] & in2[170];
    assign P[27] = in[170] ^ in2[170];
    assign G[28] = in[169] & in2[169];
    assign P[28] = in[169] ^ in2[169];
    assign G[29] = in[168] & in2[168];
    assign P[29] = in[168] ^ in2[168];
    assign G[30] = in[167] & in2[167];
    assign P[30] = in[167] ^ in2[167];
    assign G[31] = in[166] & in2[166];
    assign P[31] = in[166] ^ in2[166];
    assign G[32] = in[165] & in2[165];
    assign P[32] = in[165] ^ in2[165];
    assign G[33] = in[164] & in2[164];
    assign P[33] = in[164] ^ in2[164];
    assign G[34] = in[163] & in2[163];
    assign P[34] = in[163] ^ in2[163];
    assign G[35] = in[162] & in2[162];
    assign P[35] = in[162] ^ in2[162];
    assign G[36] = in[161] & in2[161];
    assign P[36] = in[161] ^ in2[161];
    assign G[37] = in[160] & in2[160];
    assign P[37] = in[160] ^ in2[160];
    assign G[38] = in[159] & in2[159];
    assign P[38] = in[159] ^ in2[159];
    assign G[39] = in[158] & in2[158];
    assign P[39] = in[158] ^ in2[158];
    assign G[40] = in[157] & in2[157];
    assign P[40] = in[157] ^ in2[157];
    assign G[41] = in[156] & in2[156];
    assign P[41] = in[156] ^ in2[156];
    assign G[42] = in[155] & in2[155];
    assign P[42] = in[155] ^ in2[155];
    assign G[43] = in[154] & in2[154];
    assign P[43] = in[154] ^ in2[154];
    assign G[44] = in[153] & in2[153];
    assign P[44] = in[153] ^ in2[153];
    assign G[45] = in[152] & in2[152];
    assign P[45] = in[152] ^ in2[152];
    assign G[46] = in[151] & in2[151];
    assign P[46] = in[151] ^ in2[151];
    assign G[47] = in[150] & in2[150];
    assign P[47] = in[150] ^ in2[150];
    assign G[48] = in[149] & in2[149];
    assign P[48] = in[149] ^ in2[149];
    assign G[49] = in[148] & in2[148];
    assign P[49] = in[148] ^ in2[148];
    assign G[50] = in[147] & in2[147];
    assign P[50] = in[147] ^ in2[147];
    assign G[51] = in[146] & in2[146];
    assign P[51] = in[146] ^ in2[146];
    assign G[52] = in[145] & in2[145];
    assign P[52] = in[145] ^ in2[145];
    assign G[53] = in[144] & in2[144];
    assign P[53] = in[144] ^ in2[144];
    assign G[54] = in[143] & in2[143];
    assign P[54] = in[143] ^ in2[143];
    assign G[55] = in[142] & in2[142];
    assign P[55] = in[142] ^ in2[142];
    assign G[56] = in[141] & in2[141];
    assign P[56] = in[141] ^ in2[141];
    assign G[57] = in[140] & in2[140];
    assign P[57] = in[140] ^ in2[140];
    assign G[58] = in[139] & in2[139];
    assign P[58] = in[139] ^ in2[139];
    assign G[59] = in[138] & in2[138];
    assign P[59] = in[138] ^ in2[138];
    assign G[60] = in[137] & in2[137];
    assign P[60] = in[137] ^ in2[137];
    assign G[61] = in[136] & in2[136];
    assign P[61] = in[136] ^ in2[136];
    assign G[62] = in[135] & in2[135];
    assign P[62] = in[135] ^ in2[135];
    assign G[63] = in[134] & in2[134];
    assign P[63] = in[134] ^ in2[134];
    assign G[64] = in[133] & in2[133];
    assign P[64] = in[133] ^ in2[133];
    assign G[65] = in[132] & in2[132];
    assign P[65] = in[132] ^ in2[132];
    assign G[66] = in[131] & in2[131];
    assign P[66] = in[131] ^ in2[131];
    assign G[67] = in[130] & in2[130];
    assign P[67] = in[130] ^ in2[130];
    assign G[68] = in[129] & in2[129];
    assign P[68] = in[129] ^ in2[129];
    assign G[69] = in[128] & in2[128];
    assign P[69] = in[128] ^ in2[128];
    assign G[70] = in[127] & in2[127];
    assign P[70] = in[127] ^ in2[127];
    assign G[71] = in[126] & in2[126];
    assign P[71] = in[126] ^ in2[126];
    assign G[72] = in[125] & in2[125];
    assign P[72] = in[125] ^ in2[125];
    assign G[73] = in[124] & in2[124];
    assign P[73] = in[124] ^ in2[124];
    assign G[74] = in[123] & in2[123];
    assign P[74] = in[123] ^ in2[123];
    assign G[75] = in[122] & in2[122];
    assign P[75] = in[122] ^ in2[122];
    assign G[76] = in[121] & in2[121];
    assign P[76] = in[121] ^ in2[121];
    assign G[77] = in[120] & in2[120];
    assign P[77] = in[120] ^ in2[120];
    assign G[78] = in[119] & in2[119];
    assign P[78] = in[119] ^ in2[119];
    assign G[79] = in[118] & in2[118];
    assign P[79] = in[118] ^ in2[118];
    assign G[80] = in[117] & in2[117];
    assign P[80] = in[117] ^ in2[117];
    assign G[81] = in[116] & in2[116];
    assign P[81] = in[116] ^ in2[116];
    assign G[82] = in[115] & in2[115];
    assign P[82] = in[115] ^ in2[115];
    assign G[83] = in[114] & in2[114];
    assign P[83] = in[114] ^ in2[114];
    assign G[84] = in[113] & in2[113];
    assign P[84] = in[113] ^ in2[113];
    assign G[85] = in[112] & in2[112];
    assign P[85] = in[112] ^ in2[112];
    assign G[86] = in[111] & in2[111];
    assign P[86] = in[111] ^ in2[111];
    assign G[87] = in[110] & in2[110];
    assign P[87] = in[110] ^ in2[110];
    assign G[88] = in[109] & in2[109];
    assign P[88] = in[109] ^ in2[109];
    assign G[89] = in[108] & in2[108];
    assign P[89] = in[108] ^ in2[108];
    assign G[90] = in[107] & in2[107];
    assign P[90] = in[107] ^ in2[107];
    assign G[91] = in[106] & in2[106];
    assign P[91] = in[106] ^ in2[106];
    assign G[92] = in[105] & in2[105];
    assign P[92] = in[105] ^ in2[105];
    assign G[93] = in[104] & in2[104];
    assign P[93] = in[104] ^ in2[104];
    assign G[94] = in[103] & in2[103];
    assign P[94] = in[103] ^ in2[103];
    assign G[95] = in[102] & in2[102];
    assign P[95] = in[102] ^ in2[102];
    assign G[96] = in[101] & in2[101];
    assign P[96] = in[101] ^ in2[101];
    assign G[97] = in[100] & in2[100];
    assign P[97] = in[100] ^ in2[100];
    assign G[98] = in[99] & in2[99];
    assign P[98] = in[99] ^ in2[99];
    assign G[99] = in[98] & in2[98];
    assign P[99] = in[98] ^ in2[98];
    assign G[100] = in[97] & in2[97];
    assign P[100] = in[97] ^ in2[97];
    assign G[101] = in[96] & in2[96];
    assign P[101] = in[96] ^ in2[96];
    assign G[102] = in[95] & in2[95];
    assign P[102] = in[95] ^ in2[95];
    assign G[103] = in[94] & in2[94];
    assign P[103] = in[94] ^ in2[94];
    assign G[104] = in[93] & in2[93];
    assign P[104] = in[93] ^ in2[93];
    assign G[105] = in[92] & in2[92];
    assign P[105] = in[92] ^ in2[92];
    assign G[106] = in[91] & in2[91];
    assign P[106] = in[91] ^ in2[91];
    assign G[107] = in[90] & in2[90];
    assign P[107] = in[90] ^ in2[90];
    assign G[108] = in[89] & in2[89];
    assign P[108] = in[89] ^ in2[89];
    assign G[109] = in[88] & in2[88];
    assign P[109] = in[88] ^ in2[88];
    assign G[110] = in[87] & in2[87];
    assign P[110] = in[87] ^ in2[87];
    assign G[111] = in[86] & in2[86];
    assign P[111] = in[86] ^ in2[86];
    assign G[112] = in[85] & in2[85];
    assign P[112] = in[85] ^ in2[85];
    assign G[113] = in[84] & in2[84];
    assign P[113] = in[84] ^ in2[84];
    assign G[114] = in[83] & in2[83];
    assign P[114] = in[83] ^ in2[83];
    assign G[115] = in[82] & in2[82];
    assign P[115] = in[82] ^ in2[82];
    assign G[116] = in[81] & in2[81];
    assign P[116] = in[81] ^ in2[81];
    assign G[117] = in[80] & in2[80];
    assign P[117] = in[80] ^ in2[80];
    assign G[118] = in[79] & in2[79];
    assign P[118] = in[79] ^ in2[79];
    assign G[119] = in[78] & in2[78];
    assign P[119] = in[78] ^ in2[78];
    assign G[120] = in[77] & in2[77];
    assign P[120] = in[77] ^ in2[77];
    assign G[121] = in[76] & in2[76];
    assign P[121] = in[76] ^ in2[76];
    assign G[122] = in[75] & in2[75];
    assign P[122] = in[75] ^ in2[75];
    assign G[123] = in[74] & in2[74];
    assign P[123] = in[74] ^ in2[74];
    assign G[124] = in[73] & in2[73];
    assign P[124] = in[73] ^ in2[73];
    assign G[125] = in[72] & in2[72];
    assign P[125] = in[72] ^ in2[72];
    assign G[126] = in[71] & in2[71];
    assign P[126] = in[71] ^ in2[71];
    assign G[127] = in[70] & in2[70];
    assign P[127] = in[70] ^ in2[70];
    assign G[128] = in[69] & in2[69];
    assign P[128] = in[69] ^ in2[69];
    assign G[129] = in[68] & in2[68];
    assign P[129] = in[68] ^ in2[68];
    assign G[130] = in[67] & in2[67];
    assign P[130] = in[67] ^ in2[67];
    assign G[131] = in[66] & in2[66];
    assign P[131] = in[66] ^ in2[66];
    assign G[132] = in[65] & in2[65];
    assign P[132] = in[65] ^ in2[65];
    assign G[133] = in[64] & in2[64];
    assign P[133] = in[64] ^ in2[64];
    assign G[134] = in[63] & in2[63];
    assign P[134] = in[63] ^ in2[63];
    assign G[135] = in[62] & in2[62];
    assign P[135] = in[62] ^ in2[62];
    assign G[136] = in[61] & in2[61];
    assign P[136] = in[61] ^ in2[61];
    assign G[137] = in[60] & in2[60];
    assign P[137] = in[60] ^ in2[60];
    assign G[138] = in[59] & in2[59];
    assign P[138] = in[59] ^ in2[59];
    assign G[139] = in[58] & in2[58];
    assign P[139] = in[58] ^ in2[58];
    assign G[140] = in[57] & in2[57];
    assign P[140] = in[57] ^ in2[57];
    assign G[141] = in[56] & in2[56];
    assign P[141] = in[56] ^ in2[56];
    assign G[142] = in[55] & in2[55];
    assign P[142] = in[55] ^ in2[55];
    assign G[143] = in[54] & in2[54];
    assign P[143] = in[54] ^ in2[54];
    assign G[144] = in[53] & in2[53];
    assign P[144] = in[53] ^ in2[53];
    assign G[145] = in[52] & in2[52];
    assign P[145] = in[52] ^ in2[52];
    assign G[146] = in[51] & in2[51];
    assign P[146] = in[51] ^ in2[51];
    assign G[147] = in[50] & in2[50];
    assign P[147] = in[50] ^ in2[50];
    assign G[148] = in[49] & in2[49];
    assign P[148] = in[49] ^ in2[49];
    assign G[149] = in[48] & in2[48];
    assign P[149] = in[48] ^ in2[48];
    assign G[150] = in[47] & in2[47];
    assign P[150] = in[47] ^ in2[47];
    assign G[151] = in[46] & in2[46];
    assign P[151] = in[46] ^ in2[46];
    assign G[152] = in[45] & in2[45];
    assign P[152] = in[45] ^ in2[45];
    assign G[153] = in[44] & in2[44];
    assign P[153] = in[44] ^ in2[44];
    assign G[154] = in[43] & in2[43];
    assign P[154] = in[43] ^ in2[43];
    assign G[155] = in[42] & in2[42];
    assign P[155] = in[42] ^ in2[42];
    assign G[156] = in[41] & in2[41];
    assign P[156] = in[41] ^ in2[41];
    assign G[157] = in[40] & in2[40];
    assign P[157] = in[40] ^ in2[40];
    assign G[158] = in[39] & in2[39];
    assign P[158] = in[39] ^ in2[39];
    assign G[159] = in[38] & in2[38];
    assign P[159] = in[38] ^ in2[38];
    assign G[160] = in[37] & in2[37];
    assign P[160] = in[37] ^ in2[37];
    assign G[161] = in[36] & in2[36];
    assign P[161] = in[36] ^ in2[36];
    assign G[162] = in[35] & in2[35];
    assign P[162] = in[35] ^ in2[35];
    assign G[163] = in[34] & in2[34];
    assign P[163] = in[34] ^ in2[34];
    assign G[164] = in[33] & in2[33];
    assign P[164] = in[33] ^ in2[33];
    assign G[165] = in[32] & in2[32];
    assign P[165] = in[32] ^ in2[32];
    assign G[166] = in[31] & in2[31];
    assign P[166] = in[31] ^ in2[31];
    assign G[167] = in[30] & in2[30];
    assign P[167] = in[30] ^ in2[30];
    assign G[168] = in[29] & in2[29];
    assign P[168] = in[29] ^ in2[29];
    assign G[169] = in[28] & in2[28];
    assign P[169] = in[28] ^ in2[28];
    assign G[170] = in[27] & in2[27];
    assign P[170] = in[27] ^ in2[27];
    assign G[171] = in[26] & in2[26];
    assign P[171] = in[26] ^ in2[26];
    assign G[172] = in[25] & in2[25];
    assign P[172] = in[25] ^ in2[25];
    assign G[173] = in[24] & in2[24];
    assign P[173] = in[24] ^ in2[24];
    assign G[174] = in[23] & in2[23];
    assign P[174] = in[23] ^ in2[23];
    assign G[175] = in[22] & in2[22];
    assign P[175] = in[22] ^ in2[22];
    assign G[176] = in[21] & in2[21];
    assign P[176] = in[21] ^ in2[21];
    assign G[177] = in[20] & in2[20];
    assign P[177] = in[20] ^ in2[20];
    assign G[178] = in[19] & in2[19];
    assign P[178] = in[19] ^ in2[19];
    assign G[179] = in[18] & in2[18];
    assign P[179] = in[18] ^ in2[18];
    assign G[180] = in[17] & in2[17];
    assign P[180] = in[17] ^ in2[17];
    assign G[181] = in[16] & in2[16];
    assign P[181] = in[16] ^ in2[16];
    assign G[182] = in[15] & in2[15];
    assign P[182] = in[15] ^ in2[15];
    assign G[183] = in[14] & in2[14];
    assign P[183] = in[14] ^ in2[14];
    assign G[184] = in[13] & in2[13];
    assign P[184] = in[13] ^ in2[13];
    assign G[185] = in[12] & in2[12];
    assign P[185] = in[12] ^ in2[12];
    assign G[186] = in[11] & in2[11];
    assign P[186] = in[11] ^ in2[11];
    assign G[187] = in[10] & in2[10];
    assign P[187] = in[10] ^ in2[10];
    assign G[188] = in[9] & in2[9];
    assign P[188] = in[9] ^ in2[9];
    assign G[189] = in[8] & in2[8];
    assign P[189] = in[8] ^ in2[8];
    assign G[190] = in[7] & in2[7];
    assign P[190] = in[7] ^ in2[7];
    assign G[191] = in[6] & in2[6];
    assign P[191] = in[6] ^ in2[6];
    assign G[192] = in[5] & in2[5];
    assign P[192] = in[5] ^ in2[5];
    assign G[193] = in[4] & in2[4];
    assign P[193] = in[4] ^ in2[4];
    assign G[194] = in[3] & in2[3];
    assign P[194] = in[3] ^ in2[3];
    assign G[195] = in[2] & in2[2];
    assign P[195] = in[2] ^ in2[2];
    assign G[196] = in[1] & in2[1];
    assign P[196] = in[1] ^ in2[1];
    assign G[197] = in[0] & in2[0];
    assign P[197] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign C[197] = G[196] | (P[196] & C[196]);
    assign cout = G[197] | (P[197] & C[197]);
    assign sum = P ^ C;
endmodule

module CLA197(output [196:0] sum, output cout, input [196:0] in1, input [196:0] in2;

    wire[196:0] G;
    wire[196:0] C;
    wire[196:0] P;

    assign G[0] = in[196] & in2[196];
    assign P[0] = in[196] ^ in2[196];
    assign G[1] = in[195] & in2[195];
    assign P[1] = in[195] ^ in2[195];
    assign G[2] = in[194] & in2[194];
    assign P[2] = in[194] ^ in2[194];
    assign G[3] = in[193] & in2[193];
    assign P[3] = in[193] ^ in2[193];
    assign G[4] = in[192] & in2[192];
    assign P[4] = in[192] ^ in2[192];
    assign G[5] = in[191] & in2[191];
    assign P[5] = in[191] ^ in2[191];
    assign G[6] = in[190] & in2[190];
    assign P[6] = in[190] ^ in2[190];
    assign G[7] = in[189] & in2[189];
    assign P[7] = in[189] ^ in2[189];
    assign G[8] = in[188] & in2[188];
    assign P[8] = in[188] ^ in2[188];
    assign G[9] = in[187] & in2[187];
    assign P[9] = in[187] ^ in2[187];
    assign G[10] = in[186] & in2[186];
    assign P[10] = in[186] ^ in2[186];
    assign G[11] = in[185] & in2[185];
    assign P[11] = in[185] ^ in2[185];
    assign G[12] = in[184] & in2[184];
    assign P[12] = in[184] ^ in2[184];
    assign G[13] = in[183] & in2[183];
    assign P[13] = in[183] ^ in2[183];
    assign G[14] = in[182] & in2[182];
    assign P[14] = in[182] ^ in2[182];
    assign G[15] = in[181] & in2[181];
    assign P[15] = in[181] ^ in2[181];
    assign G[16] = in[180] & in2[180];
    assign P[16] = in[180] ^ in2[180];
    assign G[17] = in[179] & in2[179];
    assign P[17] = in[179] ^ in2[179];
    assign G[18] = in[178] & in2[178];
    assign P[18] = in[178] ^ in2[178];
    assign G[19] = in[177] & in2[177];
    assign P[19] = in[177] ^ in2[177];
    assign G[20] = in[176] & in2[176];
    assign P[20] = in[176] ^ in2[176];
    assign G[21] = in[175] & in2[175];
    assign P[21] = in[175] ^ in2[175];
    assign G[22] = in[174] & in2[174];
    assign P[22] = in[174] ^ in2[174];
    assign G[23] = in[173] & in2[173];
    assign P[23] = in[173] ^ in2[173];
    assign G[24] = in[172] & in2[172];
    assign P[24] = in[172] ^ in2[172];
    assign G[25] = in[171] & in2[171];
    assign P[25] = in[171] ^ in2[171];
    assign G[26] = in[170] & in2[170];
    assign P[26] = in[170] ^ in2[170];
    assign G[27] = in[169] & in2[169];
    assign P[27] = in[169] ^ in2[169];
    assign G[28] = in[168] & in2[168];
    assign P[28] = in[168] ^ in2[168];
    assign G[29] = in[167] & in2[167];
    assign P[29] = in[167] ^ in2[167];
    assign G[30] = in[166] & in2[166];
    assign P[30] = in[166] ^ in2[166];
    assign G[31] = in[165] & in2[165];
    assign P[31] = in[165] ^ in2[165];
    assign G[32] = in[164] & in2[164];
    assign P[32] = in[164] ^ in2[164];
    assign G[33] = in[163] & in2[163];
    assign P[33] = in[163] ^ in2[163];
    assign G[34] = in[162] & in2[162];
    assign P[34] = in[162] ^ in2[162];
    assign G[35] = in[161] & in2[161];
    assign P[35] = in[161] ^ in2[161];
    assign G[36] = in[160] & in2[160];
    assign P[36] = in[160] ^ in2[160];
    assign G[37] = in[159] & in2[159];
    assign P[37] = in[159] ^ in2[159];
    assign G[38] = in[158] & in2[158];
    assign P[38] = in[158] ^ in2[158];
    assign G[39] = in[157] & in2[157];
    assign P[39] = in[157] ^ in2[157];
    assign G[40] = in[156] & in2[156];
    assign P[40] = in[156] ^ in2[156];
    assign G[41] = in[155] & in2[155];
    assign P[41] = in[155] ^ in2[155];
    assign G[42] = in[154] & in2[154];
    assign P[42] = in[154] ^ in2[154];
    assign G[43] = in[153] & in2[153];
    assign P[43] = in[153] ^ in2[153];
    assign G[44] = in[152] & in2[152];
    assign P[44] = in[152] ^ in2[152];
    assign G[45] = in[151] & in2[151];
    assign P[45] = in[151] ^ in2[151];
    assign G[46] = in[150] & in2[150];
    assign P[46] = in[150] ^ in2[150];
    assign G[47] = in[149] & in2[149];
    assign P[47] = in[149] ^ in2[149];
    assign G[48] = in[148] & in2[148];
    assign P[48] = in[148] ^ in2[148];
    assign G[49] = in[147] & in2[147];
    assign P[49] = in[147] ^ in2[147];
    assign G[50] = in[146] & in2[146];
    assign P[50] = in[146] ^ in2[146];
    assign G[51] = in[145] & in2[145];
    assign P[51] = in[145] ^ in2[145];
    assign G[52] = in[144] & in2[144];
    assign P[52] = in[144] ^ in2[144];
    assign G[53] = in[143] & in2[143];
    assign P[53] = in[143] ^ in2[143];
    assign G[54] = in[142] & in2[142];
    assign P[54] = in[142] ^ in2[142];
    assign G[55] = in[141] & in2[141];
    assign P[55] = in[141] ^ in2[141];
    assign G[56] = in[140] & in2[140];
    assign P[56] = in[140] ^ in2[140];
    assign G[57] = in[139] & in2[139];
    assign P[57] = in[139] ^ in2[139];
    assign G[58] = in[138] & in2[138];
    assign P[58] = in[138] ^ in2[138];
    assign G[59] = in[137] & in2[137];
    assign P[59] = in[137] ^ in2[137];
    assign G[60] = in[136] & in2[136];
    assign P[60] = in[136] ^ in2[136];
    assign G[61] = in[135] & in2[135];
    assign P[61] = in[135] ^ in2[135];
    assign G[62] = in[134] & in2[134];
    assign P[62] = in[134] ^ in2[134];
    assign G[63] = in[133] & in2[133];
    assign P[63] = in[133] ^ in2[133];
    assign G[64] = in[132] & in2[132];
    assign P[64] = in[132] ^ in2[132];
    assign G[65] = in[131] & in2[131];
    assign P[65] = in[131] ^ in2[131];
    assign G[66] = in[130] & in2[130];
    assign P[66] = in[130] ^ in2[130];
    assign G[67] = in[129] & in2[129];
    assign P[67] = in[129] ^ in2[129];
    assign G[68] = in[128] & in2[128];
    assign P[68] = in[128] ^ in2[128];
    assign G[69] = in[127] & in2[127];
    assign P[69] = in[127] ^ in2[127];
    assign G[70] = in[126] & in2[126];
    assign P[70] = in[126] ^ in2[126];
    assign G[71] = in[125] & in2[125];
    assign P[71] = in[125] ^ in2[125];
    assign G[72] = in[124] & in2[124];
    assign P[72] = in[124] ^ in2[124];
    assign G[73] = in[123] & in2[123];
    assign P[73] = in[123] ^ in2[123];
    assign G[74] = in[122] & in2[122];
    assign P[74] = in[122] ^ in2[122];
    assign G[75] = in[121] & in2[121];
    assign P[75] = in[121] ^ in2[121];
    assign G[76] = in[120] & in2[120];
    assign P[76] = in[120] ^ in2[120];
    assign G[77] = in[119] & in2[119];
    assign P[77] = in[119] ^ in2[119];
    assign G[78] = in[118] & in2[118];
    assign P[78] = in[118] ^ in2[118];
    assign G[79] = in[117] & in2[117];
    assign P[79] = in[117] ^ in2[117];
    assign G[80] = in[116] & in2[116];
    assign P[80] = in[116] ^ in2[116];
    assign G[81] = in[115] & in2[115];
    assign P[81] = in[115] ^ in2[115];
    assign G[82] = in[114] & in2[114];
    assign P[82] = in[114] ^ in2[114];
    assign G[83] = in[113] & in2[113];
    assign P[83] = in[113] ^ in2[113];
    assign G[84] = in[112] & in2[112];
    assign P[84] = in[112] ^ in2[112];
    assign G[85] = in[111] & in2[111];
    assign P[85] = in[111] ^ in2[111];
    assign G[86] = in[110] & in2[110];
    assign P[86] = in[110] ^ in2[110];
    assign G[87] = in[109] & in2[109];
    assign P[87] = in[109] ^ in2[109];
    assign G[88] = in[108] & in2[108];
    assign P[88] = in[108] ^ in2[108];
    assign G[89] = in[107] & in2[107];
    assign P[89] = in[107] ^ in2[107];
    assign G[90] = in[106] & in2[106];
    assign P[90] = in[106] ^ in2[106];
    assign G[91] = in[105] & in2[105];
    assign P[91] = in[105] ^ in2[105];
    assign G[92] = in[104] & in2[104];
    assign P[92] = in[104] ^ in2[104];
    assign G[93] = in[103] & in2[103];
    assign P[93] = in[103] ^ in2[103];
    assign G[94] = in[102] & in2[102];
    assign P[94] = in[102] ^ in2[102];
    assign G[95] = in[101] & in2[101];
    assign P[95] = in[101] ^ in2[101];
    assign G[96] = in[100] & in2[100];
    assign P[96] = in[100] ^ in2[100];
    assign G[97] = in[99] & in2[99];
    assign P[97] = in[99] ^ in2[99];
    assign G[98] = in[98] & in2[98];
    assign P[98] = in[98] ^ in2[98];
    assign G[99] = in[97] & in2[97];
    assign P[99] = in[97] ^ in2[97];
    assign G[100] = in[96] & in2[96];
    assign P[100] = in[96] ^ in2[96];
    assign G[101] = in[95] & in2[95];
    assign P[101] = in[95] ^ in2[95];
    assign G[102] = in[94] & in2[94];
    assign P[102] = in[94] ^ in2[94];
    assign G[103] = in[93] & in2[93];
    assign P[103] = in[93] ^ in2[93];
    assign G[104] = in[92] & in2[92];
    assign P[104] = in[92] ^ in2[92];
    assign G[105] = in[91] & in2[91];
    assign P[105] = in[91] ^ in2[91];
    assign G[106] = in[90] & in2[90];
    assign P[106] = in[90] ^ in2[90];
    assign G[107] = in[89] & in2[89];
    assign P[107] = in[89] ^ in2[89];
    assign G[108] = in[88] & in2[88];
    assign P[108] = in[88] ^ in2[88];
    assign G[109] = in[87] & in2[87];
    assign P[109] = in[87] ^ in2[87];
    assign G[110] = in[86] & in2[86];
    assign P[110] = in[86] ^ in2[86];
    assign G[111] = in[85] & in2[85];
    assign P[111] = in[85] ^ in2[85];
    assign G[112] = in[84] & in2[84];
    assign P[112] = in[84] ^ in2[84];
    assign G[113] = in[83] & in2[83];
    assign P[113] = in[83] ^ in2[83];
    assign G[114] = in[82] & in2[82];
    assign P[114] = in[82] ^ in2[82];
    assign G[115] = in[81] & in2[81];
    assign P[115] = in[81] ^ in2[81];
    assign G[116] = in[80] & in2[80];
    assign P[116] = in[80] ^ in2[80];
    assign G[117] = in[79] & in2[79];
    assign P[117] = in[79] ^ in2[79];
    assign G[118] = in[78] & in2[78];
    assign P[118] = in[78] ^ in2[78];
    assign G[119] = in[77] & in2[77];
    assign P[119] = in[77] ^ in2[77];
    assign G[120] = in[76] & in2[76];
    assign P[120] = in[76] ^ in2[76];
    assign G[121] = in[75] & in2[75];
    assign P[121] = in[75] ^ in2[75];
    assign G[122] = in[74] & in2[74];
    assign P[122] = in[74] ^ in2[74];
    assign G[123] = in[73] & in2[73];
    assign P[123] = in[73] ^ in2[73];
    assign G[124] = in[72] & in2[72];
    assign P[124] = in[72] ^ in2[72];
    assign G[125] = in[71] & in2[71];
    assign P[125] = in[71] ^ in2[71];
    assign G[126] = in[70] & in2[70];
    assign P[126] = in[70] ^ in2[70];
    assign G[127] = in[69] & in2[69];
    assign P[127] = in[69] ^ in2[69];
    assign G[128] = in[68] & in2[68];
    assign P[128] = in[68] ^ in2[68];
    assign G[129] = in[67] & in2[67];
    assign P[129] = in[67] ^ in2[67];
    assign G[130] = in[66] & in2[66];
    assign P[130] = in[66] ^ in2[66];
    assign G[131] = in[65] & in2[65];
    assign P[131] = in[65] ^ in2[65];
    assign G[132] = in[64] & in2[64];
    assign P[132] = in[64] ^ in2[64];
    assign G[133] = in[63] & in2[63];
    assign P[133] = in[63] ^ in2[63];
    assign G[134] = in[62] & in2[62];
    assign P[134] = in[62] ^ in2[62];
    assign G[135] = in[61] & in2[61];
    assign P[135] = in[61] ^ in2[61];
    assign G[136] = in[60] & in2[60];
    assign P[136] = in[60] ^ in2[60];
    assign G[137] = in[59] & in2[59];
    assign P[137] = in[59] ^ in2[59];
    assign G[138] = in[58] & in2[58];
    assign P[138] = in[58] ^ in2[58];
    assign G[139] = in[57] & in2[57];
    assign P[139] = in[57] ^ in2[57];
    assign G[140] = in[56] & in2[56];
    assign P[140] = in[56] ^ in2[56];
    assign G[141] = in[55] & in2[55];
    assign P[141] = in[55] ^ in2[55];
    assign G[142] = in[54] & in2[54];
    assign P[142] = in[54] ^ in2[54];
    assign G[143] = in[53] & in2[53];
    assign P[143] = in[53] ^ in2[53];
    assign G[144] = in[52] & in2[52];
    assign P[144] = in[52] ^ in2[52];
    assign G[145] = in[51] & in2[51];
    assign P[145] = in[51] ^ in2[51];
    assign G[146] = in[50] & in2[50];
    assign P[146] = in[50] ^ in2[50];
    assign G[147] = in[49] & in2[49];
    assign P[147] = in[49] ^ in2[49];
    assign G[148] = in[48] & in2[48];
    assign P[148] = in[48] ^ in2[48];
    assign G[149] = in[47] & in2[47];
    assign P[149] = in[47] ^ in2[47];
    assign G[150] = in[46] & in2[46];
    assign P[150] = in[46] ^ in2[46];
    assign G[151] = in[45] & in2[45];
    assign P[151] = in[45] ^ in2[45];
    assign G[152] = in[44] & in2[44];
    assign P[152] = in[44] ^ in2[44];
    assign G[153] = in[43] & in2[43];
    assign P[153] = in[43] ^ in2[43];
    assign G[154] = in[42] & in2[42];
    assign P[154] = in[42] ^ in2[42];
    assign G[155] = in[41] & in2[41];
    assign P[155] = in[41] ^ in2[41];
    assign G[156] = in[40] & in2[40];
    assign P[156] = in[40] ^ in2[40];
    assign G[157] = in[39] & in2[39];
    assign P[157] = in[39] ^ in2[39];
    assign G[158] = in[38] & in2[38];
    assign P[158] = in[38] ^ in2[38];
    assign G[159] = in[37] & in2[37];
    assign P[159] = in[37] ^ in2[37];
    assign G[160] = in[36] & in2[36];
    assign P[160] = in[36] ^ in2[36];
    assign G[161] = in[35] & in2[35];
    assign P[161] = in[35] ^ in2[35];
    assign G[162] = in[34] & in2[34];
    assign P[162] = in[34] ^ in2[34];
    assign G[163] = in[33] & in2[33];
    assign P[163] = in[33] ^ in2[33];
    assign G[164] = in[32] & in2[32];
    assign P[164] = in[32] ^ in2[32];
    assign G[165] = in[31] & in2[31];
    assign P[165] = in[31] ^ in2[31];
    assign G[166] = in[30] & in2[30];
    assign P[166] = in[30] ^ in2[30];
    assign G[167] = in[29] & in2[29];
    assign P[167] = in[29] ^ in2[29];
    assign G[168] = in[28] & in2[28];
    assign P[168] = in[28] ^ in2[28];
    assign G[169] = in[27] & in2[27];
    assign P[169] = in[27] ^ in2[27];
    assign G[170] = in[26] & in2[26];
    assign P[170] = in[26] ^ in2[26];
    assign G[171] = in[25] & in2[25];
    assign P[171] = in[25] ^ in2[25];
    assign G[172] = in[24] & in2[24];
    assign P[172] = in[24] ^ in2[24];
    assign G[173] = in[23] & in2[23];
    assign P[173] = in[23] ^ in2[23];
    assign G[174] = in[22] & in2[22];
    assign P[174] = in[22] ^ in2[22];
    assign G[175] = in[21] & in2[21];
    assign P[175] = in[21] ^ in2[21];
    assign G[176] = in[20] & in2[20];
    assign P[176] = in[20] ^ in2[20];
    assign G[177] = in[19] & in2[19];
    assign P[177] = in[19] ^ in2[19];
    assign G[178] = in[18] & in2[18];
    assign P[178] = in[18] ^ in2[18];
    assign G[179] = in[17] & in2[17];
    assign P[179] = in[17] ^ in2[17];
    assign G[180] = in[16] & in2[16];
    assign P[180] = in[16] ^ in2[16];
    assign G[181] = in[15] & in2[15];
    assign P[181] = in[15] ^ in2[15];
    assign G[182] = in[14] & in2[14];
    assign P[182] = in[14] ^ in2[14];
    assign G[183] = in[13] & in2[13];
    assign P[183] = in[13] ^ in2[13];
    assign G[184] = in[12] & in2[12];
    assign P[184] = in[12] ^ in2[12];
    assign G[185] = in[11] & in2[11];
    assign P[185] = in[11] ^ in2[11];
    assign G[186] = in[10] & in2[10];
    assign P[186] = in[10] ^ in2[10];
    assign G[187] = in[9] & in2[9];
    assign P[187] = in[9] ^ in2[9];
    assign G[188] = in[8] & in2[8];
    assign P[188] = in[8] ^ in2[8];
    assign G[189] = in[7] & in2[7];
    assign P[189] = in[7] ^ in2[7];
    assign G[190] = in[6] & in2[6];
    assign P[190] = in[6] ^ in2[6];
    assign G[191] = in[5] & in2[5];
    assign P[191] = in[5] ^ in2[5];
    assign G[192] = in[4] & in2[4];
    assign P[192] = in[4] ^ in2[4];
    assign G[193] = in[3] & in2[3];
    assign P[193] = in[3] ^ in2[3];
    assign G[194] = in[2] & in2[2];
    assign P[194] = in[2] ^ in2[2];
    assign G[195] = in[1] & in2[1];
    assign P[195] = in[1] ^ in2[1];
    assign G[196] = in[0] & in2[0];
    assign P[196] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign C[196] = G[195] | (P[195] & C[195]);
    assign cout = G[196] | (P[196] & C[196]);
    assign sum = P ^ C;
endmodule

module CLA196(output [195:0] sum, output cout, input [195:0] in1, input [195:0] in2;

    wire[195:0] G;
    wire[195:0] C;
    wire[195:0] P;

    assign G[0] = in[195] & in2[195];
    assign P[0] = in[195] ^ in2[195];
    assign G[1] = in[194] & in2[194];
    assign P[1] = in[194] ^ in2[194];
    assign G[2] = in[193] & in2[193];
    assign P[2] = in[193] ^ in2[193];
    assign G[3] = in[192] & in2[192];
    assign P[3] = in[192] ^ in2[192];
    assign G[4] = in[191] & in2[191];
    assign P[4] = in[191] ^ in2[191];
    assign G[5] = in[190] & in2[190];
    assign P[5] = in[190] ^ in2[190];
    assign G[6] = in[189] & in2[189];
    assign P[6] = in[189] ^ in2[189];
    assign G[7] = in[188] & in2[188];
    assign P[7] = in[188] ^ in2[188];
    assign G[8] = in[187] & in2[187];
    assign P[8] = in[187] ^ in2[187];
    assign G[9] = in[186] & in2[186];
    assign P[9] = in[186] ^ in2[186];
    assign G[10] = in[185] & in2[185];
    assign P[10] = in[185] ^ in2[185];
    assign G[11] = in[184] & in2[184];
    assign P[11] = in[184] ^ in2[184];
    assign G[12] = in[183] & in2[183];
    assign P[12] = in[183] ^ in2[183];
    assign G[13] = in[182] & in2[182];
    assign P[13] = in[182] ^ in2[182];
    assign G[14] = in[181] & in2[181];
    assign P[14] = in[181] ^ in2[181];
    assign G[15] = in[180] & in2[180];
    assign P[15] = in[180] ^ in2[180];
    assign G[16] = in[179] & in2[179];
    assign P[16] = in[179] ^ in2[179];
    assign G[17] = in[178] & in2[178];
    assign P[17] = in[178] ^ in2[178];
    assign G[18] = in[177] & in2[177];
    assign P[18] = in[177] ^ in2[177];
    assign G[19] = in[176] & in2[176];
    assign P[19] = in[176] ^ in2[176];
    assign G[20] = in[175] & in2[175];
    assign P[20] = in[175] ^ in2[175];
    assign G[21] = in[174] & in2[174];
    assign P[21] = in[174] ^ in2[174];
    assign G[22] = in[173] & in2[173];
    assign P[22] = in[173] ^ in2[173];
    assign G[23] = in[172] & in2[172];
    assign P[23] = in[172] ^ in2[172];
    assign G[24] = in[171] & in2[171];
    assign P[24] = in[171] ^ in2[171];
    assign G[25] = in[170] & in2[170];
    assign P[25] = in[170] ^ in2[170];
    assign G[26] = in[169] & in2[169];
    assign P[26] = in[169] ^ in2[169];
    assign G[27] = in[168] & in2[168];
    assign P[27] = in[168] ^ in2[168];
    assign G[28] = in[167] & in2[167];
    assign P[28] = in[167] ^ in2[167];
    assign G[29] = in[166] & in2[166];
    assign P[29] = in[166] ^ in2[166];
    assign G[30] = in[165] & in2[165];
    assign P[30] = in[165] ^ in2[165];
    assign G[31] = in[164] & in2[164];
    assign P[31] = in[164] ^ in2[164];
    assign G[32] = in[163] & in2[163];
    assign P[32] = in[163] ^ in2[163];
    assign G[33] = in[162] & in2[162];
    assign P[33] = in[162] ^ in2[162];
    assign G[34] = in[161] & in2[161];
    assign P[34] = in[161] ^ in2[161];
    assign G[35] = in[160] & in2[160];
    assign P[35] = in[160] ^ in2[160];
    assign G[36] = in[159] & in2[159];
    assign P[36] = in[159] ^ in2[159];
    assign G[37] = in[158] & in2[158];
    assign P[37] = in[158] ^ in2[158];
    assign G[38] = in[157] & in2[157];
    assign P[38] = in[157] ^ in2[157];
    assign G[39] = in[156] & in2[156];
    assign P[39] = in[156] ^ in2[156];
    assign G[40] = in[155] & in2[155];
    assign P[40] = in[155] ^ in2[155];
    assign G[41] = in[154] & in2[154];
    assign P[41] = in[154] ^ in2[154];
    assign G[42] = in[153] & in2[153];
    assign P[42] = in[153] ^ in2[153];
    assign G[43] = in[152] & in2[152];
    assign P[43] = in[152] ^ in2[152];
    assign G[44] = in[151] & in2[151];
    assign P[44] = in[151] ^ in2[151];
    assign G[45] = in[150] & in2[150];
    assign P[45] = in[150] ^ in2[150];
    assign G[46] = in[149] & in2[149];
    assign P[46] = in[149] ^ in2[149];
    assign G[47] = in[148] & in2[148];
    assign P[47] = in[148] ^ in2[148];
    assign G[48] = in[147] & in2[147];
    assign P[48] = in[147] ^ in2[147];
    assign G[49] = in[146] & in2[146];
    assign P[49] = in[146] ^ in2[146];
    assign G[50] = in[145] & in2[145];
    assign P[50] = in[145] ^ in2[145];
    assign G[51] = in[144] & in2[144];
    assign P[51] = in[144] ^ in2[144];
    assign G[52] = in[143] & in2[143];
    assign P[52] = in[143] ^ in2[143];
    assign G[53] = in[142] & in2[142];
    assign P[53] = in[142] ^ in2[142];
    assign G[54] = in[141] & in2[141];
    assign P[54] = in[141] ^ in2[141];
    assign G[55] = in[140] & in2[140];
    assign P[55] = in[140] ^ in2[140];
    assign G[56] = in[139] & in2[139];
    assign P[56] = in[139] ^ in2[139];
    assign G[57] = in[138] & in2[138];
    assign P[57] = in[138] ^ in2[138];
    assign G[58] = in[137] & in2[137];
    assign P[58] = in[137] ^ in2[137];
    assign G[59] = in[136] & in2[136];
    assign P[59] = in[136] ^ in2[136];
    assign G[60] = in[135] & in2[135];
    assign P[60] = in[135] ^ in2[135];
    assign G[61] = in[134] & in2[134];
    assign P[61] = in[134] ^ in2[134];
    assign G[62] = in[133] & in2[133];
    assign P[62] = in[133] ^ in2[133];
    assign G[63] = in[132] & in2[132];
    assign P[63] = in[132] ^ in2[132];
    assign G[64] = in[131] & in2[131];
    assign P[64] = in[131] ^ in2[131];
    assign G[65] = in[130] & in2[130];
    assign P[65] = in[130] ^ in2[130];
    assign G[66] = in[129] & in2[129];
    assign P[66] = in[129] ^ in2[129];
    assign G[67] = in[128] & in2[128];
    assign P[67] = in[128] ^ in2[128];
    assign G[68] = in[127] & in2[127];
    assign P[68] = in[127] ^ in2[127];
    assign G[69] = in[126] & in2[126];
    assign P[69] = in[126] ^ in2[126];
    assign G[70] = in[125] & in2[125];
    assign P[70] = in[125] ^ in2[125];
    assign G[71] = in[124] & in2[124];
    assign P[71] = in[124] ^ in2[124];
    assign G[72] = in[123] & in2[123];
    assign P[72] = in[123] ^ in2[123];
    assign G[73] = in[122] & in2[122];
    assign P[73] = in[122] ^ in2[122];
    assign G[74] = in[121] & in2[121];
    assign P[74] = in[121] ^ in2[121];
    assign G[75] = in[120] & in2[120];
    assign P[75] = in[120] ^ in2[120];
    assign G[76] = in[119] & in2[119];
    assign P[76] = in[119] ^ in2[119];
    assign G[77] = in[118] & in2[118];
    assign P[77] = in[118] ^ in2[118];
    assign G[78] = in[117] & in2[117];
    assign P[78] = in[117] ^ in2[117];
    assign G[79] = in[116] & in2[116];
    assign P[79] = in[116] ^ in2[116];
    assign G[80] = in[115] & in2[115];
    assign P[80] = in[115] ^ in2[115];
    assign G[81] = in[114] & in2[114];
    assign P[81] = in[114] ^ in2[114];
    assign G[82] = in[113] & in2[113];
    assign P[82] = in[113] ^ in2[113];
    assign G[83] = in[112] & in2[112];
    assign P[83] = in[112] ^ in2[112];
    assign G[84] = in[111] & in2[111];
    assign P[84] = in[111] ^ in2[111];
    assign G[85] = in[110] & in2[110];
    assign P[85] = in[110] ^ in2[110];
    assign G[86] = in[109] & in2[109];
    assign P[86] = in[109] ^ in2[109];
    assign G[87] = in[108] & in2[108];
    assign P[87] = in[108] ^ in2[108];
    assign G[88] = in[107] & in2[107];
    assign P[88] = in[107] ^ in2[107];
    assign G[89] = in[106] & in2[106];
    assign P[89] = in[106] ^ in2[106];
    assign G[90] = in[105] & in2[105];
    assign P[90] = in[105] ^ in2[105];
    assign G[91] = in[104] & in2[104];
    assign P[91] = in[104] ^ in2[104];
    assign G[92] = in[103] & in2[103];
    assign P[92] = in[103] ^ in2[103];
    assign G[93] = in[102] & in2[102];
    assign P[93] = in[102] ^ in2[102];
    assign G[94] = in[101] & in2[101];
    assign P[94] = in[101] ^ in2[101];
    assign G[95] = in[100] & in2[100];
    assign P[95] = in[100] ^ in2[100];
    assign G[96] = in[99] & in2[99];
    assign P[96] = in[99] ^ in2[99];
    assign G[97] = in[98] & in2[98];
    assign P[97] = in[98] ^ in2[98];
    assign G[98] = in[97] & in2[97];
    assign P[98] = in[97] ^ in2[97];
    assign G[99] = in[96] & in2[96];
    assign P[99] = in[96] ^ in2[96];
    assign G[100] = in[95] & in2[95];
    assign P[100] = in[95] ^ in2[95];
    assign G[101] = in[94] & in2[94];
    assign P[101] = in[94] ^ in2[94];
    assign G[102] = in[93] & in2[93];
    assign P[102] = in[93] ^ in2[93];
    assign G[103] = in[92] & in2[92];
    assign P[103] = in[92] ^ in2[92];
    assign G[104] = in[91] & in2[91];
    assign P[104] = in[91] ^ in2[91];
    assign G[105] = in[90] & in2[90];
    assign P[105] = in[90] ^ in2[90];
    assign G[106] = in[89] & in2[89];
    assign P[106] = in[89] ^ in2[89];
    assign G[107] = in[88] & in2[88];
    assign P[107] = in[88] ^ in2[88];
    assign G[108] = in[87] & in2[87];
    assign P[108] = in[87] ^ in2[87];
    assign G[109] = in[86] & in2[86];
    assign P[109] = in[86] ^ in2[86];
    assign G[110] = in[85] & in2[85];
    assign P[110] = in[85] ^ in2[85];
    assign G[111] = in[84] & in2[84];
    assign P[111] = in[84] ^ in2[84];
    assign G[112] = in[83] & in2[83];
    assign P[112] = in[83] ^ in2[83];
    assign G[113] = in[82] & in2[82];
    assign P[113] = in[82] ^ in2[82];
    assign G[114] = in[81] & in2[81];
    assign P[114] = in[81] ^ in2[81];
    assign G[115] = in[80] & in2[80];
    assign P[115] = in[80] ^ in2[80];
    assign G[116] = in[79] & in2[79];
    assign P[116] = in[79] ^ in2[79];
    assign G[117] = in[78] & in2[78];
    assign P[117] = in[78] ^ in2[78];
    assign G[118] = in[77] & in2[77];
    assign P[118] = in[77] ^ in2[77];
    assign G[119] = in[76] & in2[76];
    assign P[119] = in[76] ^ in2[76];
    assign G[120] = in[75] & in2[75];
    assign P[120] = in[75] ^ in2[75];
    assign G[121] = in[74] & in2[74];
    assign P[121] = in[74] ^ in2[74];
    assign G[122] = in[73] & in2[73];
    assign P[122] = in[73] ^ in2[73];
    assign G[123] = in[72] & in2[72];
    assign P[123] = in[72] ^ in2[72];
    assign G[124] = in[71] & in2[71];
    assign P[124] = in[71] ^ in2[71];
    assign G[125] = in[70] & in2[70];
    assign P[125] = in[70] ^ in2[70];
    assign G[126] = in[69] & in2[69];
    assign P[126] = in[69] ^ in2[69];
    assign G[127] = in[68] & in2[68];
    assign P[127] = in[68] ^ in2[68];
    assign G[128] = in[67] & in2[67];
    assign P[128] = in[67] ^ in2[67];
    assign G[129] = in[66] & in2[66];
    assign P[129] = in[66] ^ in2[66];
    assign G[130] = in[65] & in2[65];
    assign P[130] = in[65] ^ in2[65];
    assign G[131] = in[64] & in2[64];
    assign P[131] = in[64] ^ in2[64];
    assign G[132] = in[63] & in2[63];
    assign P[132] = in[63] ^ in2[63];
    assign G[133] = in[62] & in2[62];
    assign P[133] = in[62] ^ in2[62];
    assign G[134] = in[61] & in2[61];
    assign P[134] = in[61] ^ in2[61];
    assign G[135] = in[60] & in2[60];
    assign P[135] = in[60] ^ in2[60];
    assign G[136] = in[59] & in2[59];
    assign P[136] = in[59] ^ in2[59];
    assign G[137] = in[58] & in2[58];
    assign P[137] = in[58] ^ in2[58];
    assign G[138] = in[57] & in2[57];
    assign P[138] = in[57] ^ in2[57];
    assign G[139] = in[56] & in2[56];
    assign P[139] = in[56] ^ in2[56];
    assign G[140] = in[55] & in2[55];
    assign P[140] = in[55] ^ in2[55];
    assign G[141] = in[54] & in2[54];
    assign P[141] = in[54] ^ in2[54];
    assign G[142] = in[53] & in2[53];
    assign P[142] = in[53] ^ in2[53];
    assign G[143] = in[52] & in2[52];
    assign P[143] = in[52] ^ in2[52];
    assign G[144] = in[51] & in2[51];
    assign P[144] = in[51] ^ in2[51];
    assign G[145] = in[50] & in2[50];
    assign P[145] = in[50] ^ in2[50];
    assign G[146] = in[49] & in2[49];
    assign P[146] = in[49] ^ in2[49];
    assign G[147] = in[48] & in2[48];
    assign P[147] = in[48] ^ in2[48];
    assign G[148] = in[47] & in2[47];
    assign P[148] = in[47] ^ in2[47];
    assign G[149] = in[46] & in2[46];
    assign P[149] = in[46] ^ in2[46];
    assign G[150] = in[45] & in2[45];
    assign P[150] = in[45] ^ in2[45];
    assign G[151] = in[44] & in2[44];
    assign P[151] = in[44] ^ in2[44];
    assign G[152] = in[43] & in2[43];
    assign P[152] = in[43] ^ in2[43];
    assign G[153] = in[42] & in2[42];
    assign P[153] = in[42] ^ in2[42];
    assign G[154] = in[41] & in2[41];
    assign P[154] = in[41] ^ in2[41];
    assign G[155] = in[40] & in2[40];
    assign P[155] = in[40] ^ in2[40];
    assign G[156] = in[39] & in2[39];
    assign P[156] = in[39] ^ in2[39];
    assign G[157] = in[38] & in2[38];
    assign P[157] = in[38] ^ in2[38];
    assign G[158] = in[37] & in2[37];
    assign P[158] = in[37] ^ in2[37];
    assign G[159] = in[36] & in2[36];
    assign P[159] = in[36] ^ in2[36];
    assign G[160] = in[35] & in2[35];
    assign P[160] = in[35] ^ in2[35];
    assign G[161] = in[34] & in2[34];
    assign P[161] = in[34] ^ in2[34];
    assign G[162] = in[33] & in2[33];
    assign P[162] = in[33] ^ in2[33];
    assign G[163] = in[32] & in2[32];
    assign P[163] = in[32] ^ in2[32];
    assign G[164] = in[31] & in2[31];
    assign P[164] = in[31] ^ in2[31];
    assign G[165] = in[30] & in2[30];
    assign P[165] = in[30] ^ in2[30];
    assign G[166] = in[29] & in2[29];
    assign P[166] = in[29] ^ in2[29];
    assign G[167] = in[28] & in2[28];
    assign P[167] = in[28] ^ in2[28];
    assign G[168] = in[27] & in2[27];
    assign P[168] = in[27] ^ in2[27];
    assign G[169] = in[26] & in2[26];
    assign P[169] = in[26] ^ in2[26];
    assign G[170] = in[25] & in2[25];
    assign P[170] = in[25] ^ in2[25];
    assign G[171] = in[24] & in2[24];
    assign P[171] = in[24] ^ in2[24];
    assign G[172] = in[23] & in2[23];
    assign P[172] = in[23] ^ in2[23];
    assign G[173] = in[22] & in2[22];
    assign P[173] = in[22] ^ in2[22];
    assign G[174] = in[21] & in2[21];
    assign P[174] = in[21] ^ in2[21];
    assign G[175] = in[20] & in2[20];
    assign P[175] = in[20] ^ in2[20];
    assign G[176] = in[19] & in2[19];
    assign P[176] = in[19] ^ in2[19];
    assign G[177] = in[18] & in2[18];
    assign P[177] = in[18] ^ in2[18];
    assign G[178] = in[17] & in2[17];
    assign P[178] = in[17] ^ in2[17];
    assign G[179] = in[16] & in2[16];
    assign P[179] = in[16] ^ in2[16];
    assign G[180] = in[15] & in2[15];
    assign P[180] = in[15] ^ in2[15];
    assign G[181] = in[14] & in2[14];
    assign P[181] = in[14] ^ in2[14];
    assign G[182] = in[13] & in2[13];
    assign P[182] = in[13] ^ in2[13];
    assign G[183] = in[12] & in2[12];
    assign P[183] = in[12] ^ in2[12];
    assign G[184] = in[11] & in2[11];
    assign P[184] = in[11] ^ in2[11];
    assign G[185] = in[10] & in2[10];
    assign P[185] = in[10] ^ in2[10];
    assign G[186] = in[9] & in2[9];
    assign P[186] = in[9] ^ in2[9];
    assign G[187] = in[8] & in2[8];
    assign P[187] = in[8] ^ in2[8];
    assign G[188] = in[7] & in2[7];
    assign P[188] = in[7] ^ in2[7];
    assign G[189] = in[6] & in2[6];
    assign P[189] = in[6] ^ in2[6];
    assign G[190] = in[5] & in2[5];
    assign P[190] = in[5] ^ in2[5];
    assign G[191] = in[4] & in2[4];
    assign P[191] = in[4] ^ in2[4];
    assign G[192] = in[3] & in2[3];
    assign P[192] = in[3] ^ in2[3];
    assign G[193] = in[2] & in2[2];
    assign P[193] = in[2] ^ in2[2];
    assign G[194] = in[1] & in2[1];
    assign P[194] = in[1] ^ in2[1];
    assign G[195] = in[0] & in2[0];
    assign P[195] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign C[195] = G[194] | (P[194] & C[194]);
    assign cout = G[195] | (P[195] & C[195]);
    assign sum = P ^ C;
endmodule

module CLA195(output [194:0] sum, output cout, input [194:0] in1, input [194:0] in2;

    wire[194:0] G;
    wire[194:0] C;
    wire[194:0] P;

    assign G[0] = in[194] & in2[194];
    assign P[0] = in[194] ^ in2[194];
    assign G[1] = in[193] & in2[193];
    assign P[1] = in[193] ^ in2[193];
    assign G[2] = in[192] & in2[192];
    assign P[2] = in[192] ^ in2[192];
    assign G[3] = in[191] & in2[191];
    assign P[3] = in[191] ^ in2[191];
    assign G[4] = in[190] & in2[190];
    assign P[4] = in[190] ^ in2[190];
    assign G[5] = in[189] & in2[189];
    assign P[5] = in[189] ^ in2[189];
    assign G[6] = in[188] & in2[188];
    assign P[6] = in[188] ^ in2[188];
    assign G[7] = in[187] & in2[187];
    assign P[7] = in[187] ^ in2[187];
    assign G[8] = in[186] & in2[186];
    assign P[8] = in[186] ^ in2[186];
    assign G[9] = in[185] & in2[185];
    assign P[9] = in[185] ^ in2[185];
    assign G[10] = in[184] & in2[184];
    assign P[10] = in[184] ^ in2[184];
    assign G[11] = in[183] & in2[183];
    assign P[11] = in[183] ^ in2[183];
    assign G[12] = in[182] & in2[182];
    assign P[12] = in[182] ^ in2[182];
    assign G[13] = in[181] & in2[181];
    assign P[13] = in[181] ^ in2[181];
    assign G[14] = in[180] & in2[180];
    assign P[14] = in[180] ^ in2[180];
    assign G[15] = in[179] & in2[179];
    assign P[15] = in[179] ^ in2[179];
    assign G[16] = in[178] & in2[178];
    assign P[16] = in[178] ^ in2[178];
    assign G[17] = in[177] & in2[177];
    assign P[17] = in[177] ^ in2[177];
    assign G[18] = in[176] & in2[176];
    assign P[18] = in[176] ^ in2[176];
    assign G[19] = in[175] & in2[175];
    assign P[19] = in[175] ^ in2[175];
    assign G[20] = in[174] & in2[174];
    assign P[20] = in[174] ^ in2[174];
    assign G[21] = in[173] & in2[173];
    assign P[21] = in[173] ^ in2[173];
    assign G[22] = in[172] & in2[172];
    assign P[22] = in[172] ^ in2[172];
    assign G[23] = in[171] & in2[171];
    assign P[23] = in[171] ^ in2[171];
    assign G[24] = in[170] & in2[170];
    assign P[24] = in[170] ^ in2[170];
    assign G[25] = in[169] & in2[169];
    assign P[25] = in[169] ^ in2[169];
    assign G[26] = in[168] & in2[168];
    assign P[26] = in[168] ^ in2[168];
    assign G[27] = in[167] & in2[167];
    assign P[27] = in[167] ^ in2[167];
    assign G[28] = in[166] & in2[166];
    assign P[28] = in[166] ^ in2[166];
    assign G[29] = in[165] & in2[165];
    assign P[29] = in[165] ^ in2[165];
    assign G[30] = in[164] & in2[164];
    assign P[30] = in[164] ^ in2[164];
    assign G[31] = in[163] & in2[163];
    assign P[31] = in[163] ^ in2[163];
    assign G[32] = in[162] & in2[162];
    assign P[32] = in[162] ^ in2[162];
    assign G[33] = in[161] & in2[161];
    assign P[33] = in[161] ^ in2[161];
    assign G[34] = in[160] & in2[160];
    assign P[34] = in[160] ^ in2[160];
    assign G[35] = in[159] & in2[159];
    assign P[35] = in[159] ^ in2[159];
    assign G[36] = in[158] & in2[158];
    assign P[36] = in[158] ^ in2[158];
    assign G[37] = in[157] & in2[157];
    assign P[37] = in[157] ^ in2[157];
    assign G[38] = in[156] & in2[156];
    assign P[38] = in[156] ^ in2[156];
    assign G[39] = in[155] & in2[155];
    assign P[39] = in[155] ^ in2[155];
    assign G[40] = in[154] & in2[154];
    assign P[40] = in[154] ^ in2[154];
    assign G[41] = in[153] & in2[153];
    assign P[41] = in[153] ^ in2[153];
    assign G[42] = in[152] & in2[152];
    assign P[42] = in[152] ^ in2[152];
    assign G[43] = in[151] & in2[151];
    assign P[43] = in[151] ^ in2[151];
    assign G[44] = in[150] & in2[150];
    assign P[44] = in[150] ^ in2[150];
    assign G[45] = in[149] & in2[149];
    assign P[45] = in[149] ^ in2[149];
    assign G[46] = in[148] & in2[148];
    assign P[46] = in[148] ^ in2[148];
    assign G[47] = in[147] & in2[147];
    assign P[47] = in[147] ^ in2[147];
    assign G[48] = in[146] & in2[146];
    assign P[48] = in[146] ^ in2[146];
    assign G[49] = in[145] & in2[145];
    assign P[49] = in[145] ^ in2[145];
    assign G[50] = in[144] & in2[144];
    assign P[50] = in[144] ^ in2[144];
    assign G[51] = in[143] & in2[143];
    assign P[51] = in[143] ^ in2[143];
    assign G[52] = in[142] & in2[142];
    assign P[52] = in[142] ^ in2[142];
    assign G[53] = in[141] & in2[141];
    assign P[53] = in[141] ^ in2[141];
    assign G[54] = in[140] & in2[140];
    assign P[54] = in[140] ^ in2[140];
    assign G[55] = in[139] & in2[139];
    assign P[55] = in[139] ^ in2[139];
    assign G[56] = in[138] & in2[138];
    assign P[56] = in[138] ^ in2[138];
    assign G[57] = in[137] & in2[137];
    assign P[57] = in[137] ^ in2[137];
    assign G[58] = in[136] & in2[136];
    assign P[58] = in[136] ^ in2[136];
    assign G[59] = in[135] & in2[135];
    assign P[59] = in[135] ^ in2[135];
    assign G[60] = in[134] & in2[134];
    assign P[60] = in[134] ^ in2[134];
    assign G[61] = in[133] & in2[133];
    assign P[61] = in[133] ^ in2[133];
    assign G[62] = in[132] & in2[132];
    assign P[62] = in[132] ^ in2[132];
    assign G[63] = in[131] & in2[131];
    assign P[63] = in[131] ^ in2[131];
    assign G[64] = in[130] & in2[130];
    assign P[64] = in[130] ^ in2[130];
    assign G[65] = in[129] & in2[129];
    assign P[65] = in[129] ^ in2[129];
    assign G[66] = in[128] & in2[128];
    assign P[66] = in[128] ^ in2[128];
    assign G[67] = in[127] & in2[127];
    assign P[67] = in[127] ^ in2[127];
    assign G[68] = in[126] & in2[126];
    assign P[68] = in[126] ^ in2[126];
    assign G[69] = in[125] & in2[125];
    assign P[69] = in[125] ^ in2[125];
    assign G[70] = in[124] & in2[124];
    assign P[70] = in[124] ^ in2[124];
    assign G[71] = in[123] & in2[123];
    assign P[71] = in[123] ^ in2[123];
    assign G[72] = in[122] & in2[122];
    assign P[72] = in[122] ^ in2[122];
    assign G[73] = in[121] & in2[121];
    assign P[73] = in[121] ^ in2[121];
    assign G[74] = in[120] & in2[120];
    assign P[74] = in[120] ^ in2[120];
    assign G[75] = in[119] & in2[119];
    assign P[75] = in[119] ^ in2[119];
    assign G[76] = in[118] & in2[118];
    assign P[76] = in[118] ^ in2[118];
    assign G[77] = in[117] & in2[117];
    assign P[77] = in[117] ^ in2[117];
    assign G[78] = in[116] & in2[116];
    assign P[78] = in[116] ^ in2[116];
    assign G[79] = in[115] & in2[115];
    assign P[79] = in[115] ^ in2[115];
    assign G[80] = in[114] & in2[114];
    assign P[80] = in[114] ^ in2[114];
    assign G[81] = in[113] & in2[113];
    assign P[81] = in[113] ^ in2[113];
    assign G[82] = in[112] & in2[112];
    assign P[82] = in[112] ^ in2[112];
    assign G[83] = in[111] & in2[111];
    assign P[83] = in[111] ^ in2[111];
    assign G[84] = in[110] & in2[110];
    assign P[84] = in[110] ^ in2[110];
    assign G[85] = in[109] & in2[109];
    assign P[85] = in[109] ^ in2[109];
    assign G[86] = in[108] & in2[108];
    assign P[86] = in[108] ^ in2[108];
    assign G[87] = in[107] & in2[107];
    assign P[87] = in[107] ^ in2[107];
    assign G[88] = in[106] & in2[106];
    assign P[88] = in[106] ^ in2[106];
    assign G[89] = in[105] & in2[105];
    assign P[89] = in[105] ^ in2[105];
    assign G[90] = in[104] & in2[104];
    assign P[90] = in[104] ^ in2[104];
    assign G[91] = in[103] & in2[103];
    assign P[91] = in[103] ^ in2[103];
    assign G[92] = in[102] & in2[102];
    assign P[92] = in[102] ^ in2[102];
    assign G[93] = in[101] & in2[101];
    assign P[93] = in[101] ^ in2[101];
    assign G[94] = in[100] & in2[100];
    assign P[94] = in[100] ^ in2[100];
    assign G[95] = in[99] & in2[99];
    assign P[95] = in[99] ^ in2[99];
    assign G[96] = in[98] & in2[98];
    assign P[96] = in[98] ^ in2[98];
    assign G[97] = in[97] & in2[97];
    assign P[97] = in[97] ^ in2[97];
    assign G[98] = in[96] & in2[96];
    assign P[98] = in[96] ^ in2[96];
    assign G[99] = in[95] & in2[95];
    assign P[99] = in[95] ^ in2[95];
    assign G[100] = in[94] & in2[94];
    assign P[100] = in[94] ^ in2[94];
    assign G[101] = in[93] & in2[93];
    assign P[101] = in[93] ^ in2[93];
    assign G[102] = in[92] & in2[92];
    assign P[102] = in[92] ^ in2[92];
    assign G[103] = in[91] & in2[91];
    assign P[103] = in[91] ^ in2[91];
    assign G[104] = in[90] & in2[90];
    assign P[104] = in[90] ^ in2[90];
    assign G[105] = in[89] & in2[89];
    assign P[105] = in[89] ^ in2[89];
    assign G[106] = in[88] & in2[88];
    assign P[106] = in[88] ^ in2[88];
    assign G[107] = in[87] & in2[87];
    assign P[107] = in[87] ^ in2[87];
    assign G[108] = in[86] & in2[86];
    assign P[108] = in[86] ^ in2[86];
    assign G[109] = in[85] & in2[85];
    assign P[109] = in[85] ^ in2[85];
    assign G[110] = in[84] & in2[84];
    assign P[110] = in[84] ^ in2[84];
    assign G[111] = in[83] & in2[83];
    assign P[111] = in[83] ^ in2[83];
    assign G[112] = in[82] & in2[82];
    assign P[112] = in[82] ^ in2[82];
    assign G[113] = in[81] & in2[81];
    assign P[113] = in[81] ^ in2[81];
    assign G[114] = in[80] & in2[80];
    assign P[114] = in[80] ^ in2[80];
    assign G[115] = in[79] & in2[79];
    assign P[115] = in[79] ^ in2[79];
    assign G[116] = in[78] & in2[78];
    assign P[116] = in[78] ^ in2[78];
    assign G[117] = in[77] & in2[77];
    assign P[117] = in[77] ^ in2[77];
    assign G[118] = in[76] & in2[76];
    assign P[118] = in[76] ^ in2[76];
    assign G[119] = in[75] & in2[75];
    assign P[119] = in[75] ^ in2[75];
    assign G[120] = in[74] & in2[74];
    assign P[120] = in[74] ^ in2[74];
    assign G[121] = in[73] & in2[73];
    assign P[121] = in[73] ^ in2[73];
    assign G[122] = in[72] & in2[72];
    assign P[122] = in[72] ^ in2[72];
    assign G[123] = in[71] & in2[71];
    assign P[123] = in[71] ^ in2[71];
    assign G[124] = in[70] & in2[70];
    assign P[124] = in[70] ^ in2[70];
    assign G[125] = in[69] & in2[69];
    assign P[125] = in[69] ^ in2[69];
    assign G[126] = in[68] & in2[68];
    assign P[126] = in[68] ^ in2[68];
    assign G[127] = in[67] & in2[67];
    assign P[127] = in[67] ^ in2[67];
    assign G[128] = in[66] & in2[66];
    assign P[128] = in[66] ^ in2[66];
    assign G[129] = in[65] & in2[65];
    assign P[129] = in[65] ^ in2[65];
    assign G[130] = in[64] & in2[64];
    assign P[130] = in[64] ^ in2[64];
    assign G[131] = in[63] & in2[63];
    assign P[131] = in[63] ^ in2[63];
    assign G[132] = in[62] & in2[62];
    assign P[132] = in[62] ^ in2[62];
    assign G[133] = in[61] & in2[61];
    assign P[133] = in[61] ^ in2[61];
    assign G[134] = in[60] & in2[60];
    assign P[134] = in[60] ^ in2[60];
    assign G[135] = in[59] & in2[59];
    assign P[135] = in[59] ^ in2[59];
    assign G[136] = in[58] & in2[58];
    assign P[136] = in[58] ^ in2[58];
    assign G[137] = in[57] & in2[57];
    assign P[137] = in[57] ^ in2[57];
    assign G[138] = in[56] & in2[56];
    assign P[138] = in[56] ^ in2[56];
    assign G[139] = in[55] & in2[55];
    assign P[139] = in[55] ^ in2[55];
    assign G[140] = in[54] & in2[54];
    assign P[140] = in[54] ^ in2[54];
    assign G[141] = in[53] & in2[53];
    assign P[141] = in[53] ^ in2[53];
    assign G[142] = in[52] & in2[52];
    assign P[142] = in[52] ^ in2[52];
    assign G[143] = in[51] & in2[51];
    assign P[143] = in[51] ^ in2[51];
    assign G[144] = in[50] & in2[50];
    assign P[144] = in[50] ^ in2[50];
    assign G[145] = in[49] & in2[49];
    assign P[145] = in[49] ^ in2[49];
    assign G[146] = in[48] & in2[48];
    assign P[146] = in[48] ^ in2[48];
    assign G[147] = in[47] & in2[47];
    assign P[147] = in[47] ^ in2[47];
    assign G[148] = in[46] & in2[46];
    assign P[148] = in[46] ^ in2[46];
    assign G[149] = in[45] & in2[45];
    assign P[149] = in[45] ^ in2[45];
    assign G[150] = in[44] & in2[44];
    assign P[150] = in[44] ^ in2[44];
    assign G[151] = in[43] & in2[43];
    assign P[151] = in[43] ^ in2[43];
    assign G[152] = in[42] & in2[42];
    assign P[152] = in[42] ^ in2[42];
    assign G[153] = in[41] & in2[41];
    assign P[153] = in[41] ^ in2[41];
    assign G[154] = in[40] & in2[40];
    assign P[154] = in[40] ^ in2[40];
    assign G[155] = in[39] & in2[39];
    assign P[155] = in[39] ^ in2[39];
    assign G[156] = in[38] & in2[38];
    assign P[156] = in[38] ^ in2[38];
    assign G[157] = in[37] & in2[37];
    assign P[157] = in[37] ^ in2[37];
    assign G[158] = in[36] & in2[36];
    assign P[158] = in[36] ^ in2[36];
    assign G[159] = in[35] & in2[35];
    assign P[159] = in[35] ^ in2[35];
    assign G[160] = in[34] & in2[34];
    assign P[160] = in[34] ^ in2[34];
    assign G[161] = in[33] & in2[33];
    assign P[161] = in[33] ^ in2[33];
    assign G[162] = in[32] & in2[32];
    assign P[162] = in[32] ^ in2[32];
    assign G[163] = in[31] & in2[31];
    assign P[163] = in[31] ^ in2[31];
    assign G[164] = in[30] & in2[30];
    assign P[164] = in[30] ^ in2[30];
    assign G[165] = in[29] & in2[29];
    assign P[165] = in[29] ^ in2[29];
    assign G[166] = in[28] & in2[28];
    assign P[166] = in[28] ^ in2[28];
    assign G[167] = in[27] & in2[27];
    assign P[167] = in[27] ^ in2[27];
    assign G[168] = in[26] & in2[26];
    assign P[168] = in[26] ^ in2[26];
    assign G[169] = in[25] & in2[25];
    assign P[169] = in[25] ^ in2[25];
    assign G[170] = in[24] & in2[24];
    assign P[170] = in[24] ^ in2[24];
    assign G[171] = in[23] & in2[23];
    assign P[171] = in[23] ^ in2[23];
    assign G[172] = in[22] & in2[22];
    assign P[172] = in[22] ^ in2[22];
    assign G[173] = in[21] & in2[21];
    assign P[173] = in[21] ^ in2[21];
    assign G[174] = in[20] & in2[20];
    assign P[174] = in[20] ^ in2[20];
    assign G[175] = in[19] & in2[19];
    assign P[175] = in[19] ^ in2[19];
    assign G[176] = in[18] & in2[18];
    assign P[176] = in[18] ^ in2[18];
    assign G[177] = in[17] & in2[17];
    assign P[177] = in[17] ^ in2[17];
    assign G[178] = in[16] & in2[16];
    assign P[178] = in[16] ^ in2[16];
    assign G[179] = in[15] & in2[15];
    assign P[179] = in[15] ^ in2[15];
    assign G[180] = in[14] & in2[14];
    assign P[180] = in[14] ^ in2[14];
    assign G[181] = in[13] & in2[13];
    assign P[181] = in[13] ^ in2[13];
    assign G[182] = in[12] & in2[12];
    assign P[182] = in[12] ^ in2[12];
    assign G[183] = in[11] & in2[11];
    assign P[183] = in[11] ^ in2[11];
    assign G[184] = in[10] & in2[10];
    assign P[184] = in[10] ^ in2[10];
    assign G[185] = in[9] & in2[9];
    assign P[185] = in[9] ^ in2[9];
    assign G[186] = in[8] & in2[8];
    assign P[186] = in[8] ^ in2[8];
    assign G[187] = in[7] & in2[7];
    assign P[187] = in[7] ^ in2[7];
    assign G[188] = in[6] & in2[6];
    assign P[188] = in[6] ^ in2[6];
    assign G[189] = in[5] & in2[5];
    assign P[189] = in[5] ^ in2[5];
    assign G[190] = in[4] & in2[4];
    assign P[190] = in[4] ^ in2[4];
    assign G[191] = in[3] & in2[3];
    assign P[191] = in[3] ^ in2[3];
    assign G[192] = in[2] & in2[2];
    assign P[192] = in[2] ^ in2[2];
    assign G[193] = in[1] & in2[1];
    assign P[193] = in[1] ^ in2[1];
    assign G[194] = in[0] & in2[0];
    assign P[194] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign C[194] = G[193] | (P[193] & C[193]);
    assign cout = G[194] | (P[194] & C[194]);
    assign sum = P ^ C;
endmodule

module CLA194(output [193:0] sum, output cout, input [193:0] in1, input [193:0] in2;

    wire[193:0] G;
    wire[193:0] C;
    wire[193:0] P;

    assign G[0] = in[193] & in2[193];
    assign P[0] = in[193] ^ in2[193];
    assign G[1] = in[192] & in2[192];
    assign P[1] = in[192] ^ in2[192];
    assign G[2] = in[191] & in2[191];
    assign P[2] = in[191] ^ in2[191];
    assign G[3] = in[190] & in2[190];
    assign P[3] = in[190] ^ in2[190];
    assign G[4] = in[189] & in2[189];
    assign P[4] = in[189] ^ in2[189];
    assign G[5] = in[188] & in2[188];
    assign P[5] = in[188] ^ in2[188];
    assign G[6] = in[187] & in2[187];
    assign P[6] = in[187] ^ in2[187];
    assign G[7] = in[186] & in2[186];
    assign P[7] = in[186] ^ in2[186];
    assign G[8] = in[185] & in2[185];
    assign P[8] = in[185] ^ in2[185];
    assign G[9] = in[184] & in2[184];
    assign P[9] = in[184] ^ in2[184];
    assign G[10] = in[183] & in2[183];
    assign P[10] = in[183] ^ in2[183];
    assign G[11] = in[182] & in2[182];
    assign P[11] = in[182] ^ in2[182];
    assign G[12] = in[181] & in2[181];
    assign P[12] = in[181] ^ in2[181];
    assign G[13] = in[180] & in2[180];
    assign P[13] = in[180] ^ in2[180];
    assign G[14] = in[179] & in2[179];
    assign P[14] = in[179] ^ in2[179];
    assign G[15] = in[178] & in2[178];
    assign P[15] = in[178] ^ in2[178];
    assign G[16] = in[177] & in2[177];
    assign P[16] = in[177] ^ in2[177];
    assign G[17] = in[176] & in2[176];
    assign P[17] = in[176] ^ in2[176];
    assign G[18] = in[175] & in2[175];
    assign P[18] = in[175] ^ in2[175];
    assign G[19] = in[174] & in2[174];
    assign P[19] = in[174] ^ in2[174];
    assign G[20] = in[173] & in2[173];
    assign P[20] = in[173] ^ in2[173];
    assign G[21] = in[172] & in2[172];
    assign P[21] = in[172] ^ in2[172];
    assign G[22] = in[171] & in2[171];
    assign P[22] = in[171] ^ in2[171];
    assign G[23] = in[170] & in2[170];
    assign P[23] = in[170] ^ in2[170];
    assign G[24] = in[169] & in2[169];
    assign P[24] = in[169] ^ in2[169];
    assign G[25] = in[168] & in2[168];
    assign P[25] = in[168] ^ in2[168];
    assign G[26] = in[167] & in2[167];
    assign P[26] = in[167] ^ in2[167];
    assign G[27] = in[166] & in2[166];
    assign P[27] = in[166] ^ in2[166];
    assign G[28] = in[165] & in2[165];
    assign P[28] = in[165] ^ in2[165];
    assign G[29] = in[164] & in2[164];
    assign P[29] = in[164] ^ in2[164];
    assign G[30] = in[163] & in2[163];
    assign P[30] = in[163] ^ in2[163];
    assign G[31] = in[162] & in2[162];
    assign P[31] = in[162] ^ in2[162];
    assign G[32] = in[161] & in2[161];
    assign P[32] = in[161] ^ in2[161];
    assign G[33] = in[160] & in2[160];
    assign P[33] = in[160] ^ in2[160];
    assign G[34] = in[159] & in2[159];
    assign P[34] = in[159] ^ in2[159];
    assign G[35] = in[158] & in2[158];
    assign P[35] = in[158] ^ in2[158];
    assign G[36] = in[157] & in2[157];
    assign P[36] = in[157] ^ in2[157];
    assign G[37] = in[156] & in2[156];
    assign P[37] = in[156] ^ in2[156];
    assign G[38] = in[155] & in2[155];
    assign P[38] = in[155] ^ in2[155];
    assign G[39] = in[154] & in2[154];
    assign P[39] = in[154] ^ in2[154];
    assign G[40] = in[153] & in2[153];
    assign P[40] = in[153] ^ in2[153];
    assign G[41] = in[152] & in2[152];
    assign P[41] = in[152] ^ in2[152];
    assign G[42] = in[151] & in2[151];
    assign P[42] = in[151] ^ in2[151];
    assign G[43] = in[150] & in2[150];
    assign P[43] = in[150] ^ in2[150];
    assign G[44] = in[149] & in2[149];
    assign P[44] = in[149] ^ in2[149];
    assign G[45] = in[148] & in2[148];
    assign P[45] = in[148] ^ in2[148];
    assign G[46] = in[147] & in2[147];
    assign P[46] = in[147] ^ in2[147];
    assign G[47] = in[146] & in2[146];
    assign P[47] = in[146] ^ in2[146];
    assign G[48] = in[145] & in2[145];
    assign P[48] = in[145] ^ in2[145];
    assign G[49] = in[144] & in2[144];
    assign P[49] = in[144] ^ in2[144];
    assign G[50] = in[143] & in2[143];
    assign P[50] = in[143] ^ in2[143];
    assign G[51] = in[142] & in2[142];
    assign P[51] = in[142] ^ in2[142];
    assign G[52] = in[141] & in2[141];
    assign P[52] = in[141] ^ in2[141];
    assign G[53] = in[140] & in2[140];
    assign P[53] = in[140] ^ in2[140];
    assign G[54] = in[139] & in2[139];
    assign P[54] = in[139] ^ in2[139];
    assign G[55] = in[138] & in2[138];
    assign P[55] = in[138] ^ in2[138];
    assign G[56] = in[137] & in2[137];
    assign P[56] = in[137] ^ in2[137];
    assign G[57] = in[136] & in2[136];
    assign P[57] = in[136] ^ in2[136];
    assign G[58] = in[135] & in2[135];
    assign P[58] = in[135] ^ in2[135];
    assign G[59] = in[134] & in2[134];
    assign P[59] = in[134] ^ in2[134];
    assign G[60] = in[133] & in2[133];
    assign P[60] = in[133] ^ in2[133];
    assign G[61] = in[132] & in2[132];
    assign P[61] = in[132] ^ in2[132];
    assign G[62] = in[131] & in2[131];
    assign P[62] = in[131] ^ in2[131];
    assign G[63] = in[130] & in2[130];
    assign P[63] = in[130] ^ in2[130];
    assign G[64] = in[129] & in2[129];
    assign P[64] = in[129] ^ in2[129];
    assign G[65] = in[128] & in2[128];
    assign P[65] = in[128] ^ in2[128];
    assign G[66] = in[127] & in2[127];
    assign P[66] = in[127] ^ in2[127];
    assign G[67] = in[126] & in2[126];
    assign P[67] = in[126] ^ in2[126];
    assign G[68] = in[125] & in2[125];
    assign P[68] = in[125] ^ in2[125];
    assign G[69] = in[124] & in2[124];
    assign P[69] = in[124] ^ in2[124];
    assign G[70] = in[123] & in2[123];
    assign P[70] = in[123] ^ in2[123];
    assign G[71] = in[122] & in2[122];
    assign P[71] = in[122] ^ in2[122];
    assign G[72] = in[121] & in2[121];
    assign P[72] = in[121] ^ in2[121];
    assign G[73] = in[120] & in2[120];
    assign P[73] = in[120] ^ in2[120];
    assign G[74] = in[119] & in2[119];
    assign P[74] = in[119] ^ in2[119];
    assign G[75] = in[118] & in2[118];
    assign P[75] = in[118] ^ in2[118];
    assign G[76] = in[117] & in2[117];
    assign P[76] = in[117] ^ in2[117];
    assign G[77] = in[116] & in2[116];
    assign P[77] = in[116] ^ in2[116];
    assign G[78] = in[115] & in2[115];
    assign P[78] = in[115] ^ in2[115];
    assign G[79] = in[114] & in2[114];
    assign P[79] = in[114] ^ in2[114];
    assign G[80] = in[113] & in2[113];
    assign P[80] = in[113] ^ in2[113];
    assign G[81] = in[112] & in2[112];
    assign P[81] = in[112] ^ in2[112];
    assign G[82] = in[111] & in2[111];
    assign P[82] = in[111] ^ in2[111];
    assign G[83] = in[110] & in2[110];
    assign P[83] = in[110] ^ in2[110];
    assign G[84] = in[109] & in2[109];
    assign P[84] = in[109] ^ in2[109];
    assign G[85] = in[108] & in2[108];
    assign P[85] = in[108] ^ in2[108];
    assign G[86] = in[107] & in2[107];
    assign P[86] = in[107] ^ in2[107];
    assign G[87] = in[106] & in2[106];
    assign P[87] = in[106] ^ in2[106];
    assign G[88] = in[105] & in2[105];
    assign P[88] = in[105] ^ in2[105];
    assign G[89] = in[104] & in2[104];
    assign P[89] = in[104] ^ in2[104];
    assign G[90] = in[103] & in2[103];
    assign P[90] = in[103] ^ in2[103];
    assign G[91] = in[102] & in2[102];
    assign P[91] = in[102] ^ in2[102];
    assign G[92] = in[101] & in2[101];
    assign P[92] = in[101] ^ in2[101];
    assign G[93] = in[100] & in2[100];
    assign P[93] = in[100] ^ in2[100];
    assign G[94] = in[99] & in2[99];
    assign P[94] = in[99] ^ in2[99];
    assign G[95] = in[98] & in2[98];
    assign P[95] = in[98] ^ in2[98];
    assign G[96] = in[97] & in2[97];
    assign P[96] = in[97] ^ in2[97];
    assign G[97] = in[96] & in2[96];
    assign P[97] = in[96] ^ in2[96];
    assign G[98] = in[95] & in2[95];
    assign P[98] = in[95] ^ in2[95];
    assign G[99] = in[94] & in2[94];
    assign P[99] = in[94] ^ in2[94];
    assign G[100] = in[93] & in2[93];
    assign P[100] = in[93] ^ in2[93];
    assign G[101] = in[92] & in2[92];
    assign P[101] = in[92] ^ in2[92];
    assign G[102] = in[91] & in2[91];
    assign P[102] = in[91] ^ in2[91];
    assign G[103] = in[90] & in2[90];
    assign P[103] = in[90] ^ in2[90];
    assign G[104] = in[89] & in2[89];
    assign P[104] = in[89] ^ in2[89];
    assign G[105] = in[88] & in2[88];
    assign P[105] = in[88] ^ in2[88];
    assign G[106] = in[87] & in2[87];
    assign P[106] = in[87] ^ in2[87];
    assign G[107] = in[86] & in2[86];
    assign P[107] = in[86] ^ in2[86];
    assign G[108] = in[85] & in2[85];
    assign P[108] = in[85] ^ in2[85];
    assign G[109] = in[84] & in2[84];
    assign P[109] = in[84] ^ in2[84];
    assign G[110] = in[83] & in2[83];
    assign P[110] = in[83] ^ in2[83];
    assign G[111] = in[82] & in2[82];
    assign P[111] = in[82] ^ in2[82];
    assign G[112] = in[81] & in2[81];
    assign P[112] = in[81] ^ in2[81];
    assign G[113] = in[80] & in2[80];
    assign P[113] = in[80] ^ in2[80];
    assign G[114] = in[79] & in2[79];
    assign P[114] = in[79] ^ in2[79];
    assign G[115] = in[78] & in2[78];
    assign P[115] = in[78] ^ in2[78];
    assign G[116] = in[77] & in2[77];
    assign P[116] = in[77] ^ in2[77];
    assign G[117] = in[76] & in2[76];
    assign P[117] = in[76] ^ in2[76];
    assign G[118] = in[75] & in2[75];
    assign P[118] = in[75] ^ in2[75];
    assign G[119] = in[74] & in2[74];
    assign P[119] = in[74] ^ in2[74];
    assign G[120] = in[73] & in2[73];
    assign P[120] = in[73] ^ in2[73];
    assign G[121] = in[72] & in2[72];
    assign P[121] = in[72] ^ in2[72];
    assign G[122] = in[71] & in2[71];
    assign P[122] = in[71] ^ in2[71];
    assign G[123] = in[70] & in2[70];
    assign P[123] = in[70] ^ in2[70];
    assign G[124] = in[69] & in2[69];
    assign P[124] = in[69] ^ in2[69];
    assign G[125] = in[68] & in2[68];
    assign P[125] = in[68] ^ in2[68];
    assign G[126] = in[67] & in2[67];
    assign P[126] = in[67] ^ in2[67];
    assign G[127] = in[66] & in2[66];
    assign P[127] = in[66] ^ in2[66];
    assign G[128] = in[65] & in2[65];
    assign P[128] = in[65] ^ in2[65];
    assign G[129] = in[64] & in2[64];
    assign P[129] = in[64] ^ in2[64];
    assign G[130] = in[63] & in2[63];
    assign P[130] = in[63] ^ in2[63];
    assign G[131] = in[62] & in2[62];
    assign P[131] = in[62] ^ in2[62];
    assign G[132] = in[61] & in2[61];
    assign P[132] = in[61] ^ in2[61];
    assign G[133] = in[60] & in2[60];
    assign P[133] = in[60] ^ in2[60];
    assign G[134] = in[59] & in2[59];
    assign P[134] = in[59] ^ in2[59];
    assign G[135] = in[58] & in2[58];
    assign P[135] = in[58] ^ in2[58];
    assign G[136] = in[57] & in2[57];
    assign P[136] = in[57] ^ in2[57];
    assign G[137] = in[56] & in2[56];
    assign P[137] = in[56] ^ in2[56];
    assign G[138] = in[55] & in2[55];
    assign P[138] = in[55] ^ in2[55];
    assign G[139] = in[54] & in2[54];
    assign P[139] = in[54] ^ in2[54];
    assign G[140] = in[53] & in2[53];
    assign P[140] = in[53] ^ in2[53];
    assign G[141] = in[52] & in2[52];
    assign P[141] = in[52] ^ in2[52];
    assign G[142] = in[51] & in2[51];
    assign P[142] = in[51] ^ in2[51];
    assign G[143] = in[50] & in2[50];
    assign P[143] = in[50] ^ in2[50];
    assign G[144] = in[49] & in2[49];
    assign P[144] = in[49] ^ in2[49];
    assign G[145] = in[48] & in2[48];
    assign P[145] = in[48] ^ in2[48];
    assign G[146] = in[47] & in2[47];
    assign P[146] = in[47] ^ in2[47];
    assign G[147] = in[46] & in2[46];
    assign P[147] = in[46] ^ in2[46];
    assign G[148] = in[45] & in2[45];
    assign P[148] = in[45] ^ in2[45];
    assign G[149] = in[44] & in2[44];
    assign P[149] = in[44] ^ in2[44];
    assign G[150] = in[43] & in2[43];
    assign P[150] = in[43] ^ in2[43];
    assign G[151] = in[42] & in2[42];
    assign P[151] = in[42] ^ in2[42];
    assign G[152] = in[41] & in2[41];
    assign P[152] = in[41] ^ in2[41];
    assign G[153] = in[40] & in2[40];
    assign P[153] = in[40] ^ in2[40];
    assign G[154] = in[39] & in2[39];
    assign P[154] = in[39] ^ in2[39];
    assign G[155] = in[38] & in2[38];
    assign P[155] = in[38] ^ in2[38];
    assign G[156] = in[37] & in2[37];
    assign P[156] = in[37] ^ in2[37];
    assign G[157] = in[36] & in2[36];
    assign P[157] = in[36] ^ in2[36];
    assign G[158] = in[35] & in2[35];
    assign P[158] = in[35] ^ in2[35];
    assign G[159] = in[34] & in2[34];
    assign P[159] = in[34] ^ in2[34];
    assign G[160] = in[33] & in2[33];
    assign P[160] = in[33] ^ in2[33];
    assign G[161] = in[32] & in2[32];
    assign P[161] = in[32] ^ in2[32];
    assign G[162] = in[31] & in2[31];
    assign P[162] = in[31] ^ in2[31];
    assign G[163] = in[30] & in2[30];
    assign P[163] = in[30] ^ in2[30];
    assign G[164] = in[29] & in2[29];
    assign P[164] = in[29] ^ in2[29];
    assign G[165] = in[28] & in2[28];
    assign P[165] = in[28] ^ in2[28];
    assign G[166] = in[27] & in2[27];
    assign P[166] = in[27] ^ in2[27];
    assign G[167] = in[26] & in2[26];
    assign P[167] = in[26] ^ in2[26];
    assign G[168] = in[25] & in2[25];
    assign P[168] = in[25] ^ in2[25];
    assign G[169] = in[24] & in2[24];
    assign P[169] = in[24] ^ in2[24];
    assign G[170] = in[23] & in2[23];
    assign P[170] = in[23] ^ in2[23];
    assign G[171] = in[22] & in2[22];
    assign P[171] = in[22] ^ in2[22];
    assign G[172] = in[21] & in2[21];
    assign P[172] = in[21] ^ in2[21];
    assign G[173] = in[20] & in2[20];
    assign P[173] = in[20] ^ in2[20];
    assign G[174] = in[19] & in2[19];
    assign P[174] = in[19] ^ in2[19];
    assign G[175] = in[18] & in2[18];
    assign P[175] = in[18] ^ in2[18];
    assign G[176] = in[17] & in2[17];
    assign P[176] = in[17] ^ in2[17];
    assign G[177] = in[16] & in2[16];
    assign P[177] = in[16] ^ in2[16];
    assign G[178] = in[15] & in2[15];
    assign P[178] = in[15] ^ in2[15];
    assign G[179] = in[14] & in2[14];
    assign P[179] = in[14] ^ in2[14];
    assign G[180] = in[13] & in2[13];
    assign P[180] = in[13] ^ in2[13];
    assign G[181] = in[12] & in2[12];
    assign P[181] = in[12] ^ in2[12];
    assign G[182] = in[11] & in2[11];
    assign P[182] = in[11] ^ in2[11];
    assign G[183] = in[10] & in2[10];
    assign P[183] = in[10] ^ in2[10];
    assign G[184] = in[9] & in2[9];
    assign P[184] = in[9] ^ in2[9];
    assign G[185] = in[8] & in2[8];
    assign P[185] = in[8] ^ in2[8];
    assign G[186] = in[7] & in2[7];
    assign P[186] = in[7] ^ in2[7];
    assign G[187] = in[6] & in2[6];
    assign P[187] = in[6] ^ in2[6];
    assign G[188] = in[5] & in2[5];
    assign P[188] = in[5] ^ in2[5];
    assign G[189] = in[4] & in2[4];
    assign P[189] = in[4] ^ in2[4];
    assign G[190] = in[3] & in2[3];
    assign P[190] = in[3] ^ in2[3];
    assign G[191] = in[2] & in2[2];
    assign P[191] = in[2] ^ in2[2];
    assign G[192] = in[1] & in2[1];
    assign P[192] = in[1] ^ in2[1];
    assign G[193] = in[0] & in2[0];
    assign P[193] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign C[193] = G[192] | (P[192] & C[192]);
    assign cout = G[193] | (P[193] & C[193]);
    assign sum = P ^ C;
endmodule

module CLA193(output [192:0] sum, output cout, input [192:0] in1, input [192:0] in2;

    wire[192:0] G;
    wire[192:0] C;
    wire[192:0] P;

    assign G[0] = in[192] & in2[192];
    assign P[0] = in[192] ^ in2[192];
    assign G[1] = in[191] & in2[191];
    assign P[1] = in[191] ^ in2[191];
    assign G[2] = in[190] & in2[190];
    assign P[2] = in[190] ^ in2[190];
    assign G[3] = in[189] & in2[189];
    assign P[3] = in[189] ^ in2[189];
    assign G[4] = in[188] & in2[188];
    assign P[4] = in[188] ^ in2[188];
    assign G[5] = in[187] & in2[187];
    assign P[5] = in[187] ^ in2[187];
    assign G[6] = in[186] & in2[186];
    assign P[6] = in[186] ^ in2[186];
    assign G[7] = in[185] & in2[185];
    assign P[7] = in[185] ^ in2[185];
    assign G[8] = in[184] & in2[184];
    assign P[8] = in[184] ^ in2[184];
    assign G[9] = in[183] & in2[183];
    assign P[9] = in[183] ^ in2[183];
    assign G[10] = in[182] & in2[182];
    assign P[10] = in[182] ^ in2[182];
    assign G[11] = in[181] & in2[181];
    assign P[11] = in[181] ^ in2[181];
    assign G[12] = in[180] & in2[180];
    assign P[12] = in[180] ^ in2[180];
    assign G[13] = in[179] & in2[179];
    assign P[13] = in[179] ^ in2[179];
    assign G[14] = in[178] & in2[178];
    assign P[14] = in[178] ^ in2[178];
    assign G[15] = in[177] & in2[177];
    assign P[15] = in[177] ^ in2[177];
    assign G[16] = in[176] & in2[176];
    assign P[16] = in[176] ^ in2[176];
    assign G[17] = in[175] & in2[175];
    assign P[17] = in[175] ^ in2[175];
    assign G[18] = in[174] & in2[174];
    assign P[18] = in[174] ^ in2[174];
    assign G[19] = in[173] & in2[173];
    assign P[19] = in[173] ^ in2[173];
    assign G[20] = in[172] & in2[172];
    assign P[20] = in[172] ^ in2[172];
    assign G[21] = in[171] & in2[171];
    assign P[21] = in[171] ^ in2[171];
    assign G[22] = in[170] & in2[170];
    assign P[22] = in[170] ^ in2[170];
    assign G[23] = in[169] & in2[169];
    assign P[23] = in[169] ^ in2[169];
    assign G[24] = in[168] & in2[168];
    assign P[24] = in[168] ^ in2[168];
    assign G[25] = in[167] & in2[167];
    assign P[25] = in[167] ^ in2[167];
    assign G[26] = in[166] & in2[166];
    assign P[26] = in[166] ^ in2[166];
    assign G[27] = in[165] & in2[165];
    assign P[27] = in[165] ^ in2[165];
    assign G[28] = in[164] & in2[164];
    assign P[28] = in[164] ^ in2[164];
    assign G[29] = in[163] & in2[163];
    assign P[29] = in[163] ^ in2[163];
    assign G[30] = in[162] & in2[162];
    assign P[30] = in[162] ^ in2[162];
    assign G[31] = in[161] & in2[161];
    assign P[31] = in[161] ^ in2[161];
    assign G[32] = in[160] & in2[160];
    assign P[32] = in[160] ^ in2[160];
    assign G[33] = in[159] & in2[159];
    assign P[33] = in[159] ^ in2[159];
    assign G[34] = in[158] & in2[158];
    assign P[34] = in[158] ^ in2[158];
    assign G[35] = in[157] & in2[157];
    assign P[35] = in[157] ^ in2[157];
    assign G[36] = in[156] & in2[156];
    assign P[36] = in[156] ^ in2[156];
    assign G[37] = in[155] & in2[155];
    assign P[37] = in[155] ^ in2[155];
    assign G[38] = in[154] & in2[154];
    assign P[38] = in[154] ^ in2[154];
    assign G[39] = in[153] & in2[153];
    assign P[39] = in[153] ^ in2[153];
    assign G[40] = in[152] & in2[152];
    assign P[40] = in[152] ^ in2[152];
    assign G[41] = in[151] & in2[151];
    assign P[41] = in[151] ^ in2[151];
    assign G[42] = in[150] & in2[150];
    assign P[42] = in[150] ^ in2[150];
    assign G[43] = in[149] & in2[149];
    assign P[43] = in[149] ^ in2[149];
    assign G[44] = in[148] & in2[148];
    assign P[44] = in[148] ^ in2[148];
    assign G[45] = in[147] & in2[147];
    assign P[45] = in[147] ^ in2[147];
    assign G[46] = in[146] & in2[146];
    assign P[46] = in[146] ^ in2[146];
    assign G[47] = in[145] & in2[145];
    assign P[47] = in[145] ^ in2[145];
    assign G[48] = in[144] & in2[144];
    assign P[48] = in[144] ^ in2[144];
    assign G[49] = in[143] & in2[143];
    assign P[49] = in[143] ^ in2[143];
    assign G[50] = in[142] & in2[142];
    assign P[50] = in[142] ^ in2[142];
    assign G[51] = in[141] & in2[141];
    assign P[51] = in[141] ^ in2[141];
    assign G[52] = in[140] & in2[140];
    assign P[52] = in[140] ^ in2[140];
    assign G[53] = in[139] & in2[139];
    assign P[53] = in[139] ^ in2[139];
    assign G[54] = in[138] & in2[138];
    assign P[54] = in[138] ^ in2[138];
    assign G[55] = in[137] & in2[137];
    assign P[55] = in[137] ^ in2[137];
    assign G[56] = in[136] & in2[136];
    assign P[56] = in[136] ^ in2[136];
    assign G[57] = in[135] & in2[135];
    assign P[57] = in[135] ^ in2[135];
    assign G[58] = in[134] & in2[134];
    assign P[58] = in[134] ^ in2[134];
    assign G[59] = in[133] & in2[133];
    assign P[59] = in[133] ^ in2[133];
    assign G[60] = in[132] & in2[132];
    assign P[60] = in[132] ^ in2[132];
    assign G[61] = in[131] & in2[131];
    assign P[61] = in[131] ^ in2[131];
    assign G[62] = in[130] & in2[130];
    assign P[62] = in[130] ^ in2[130];
    assign G[63] = in[129] & in2[129];
    assign P[63] = in[129] ^ in2[129];
    assign G[64] = in[128] & in2[128];
    assign P[64] = in[128] ^ in2[128];
    assign G[65] = in[127] & in2[127];
    assign P[65] = in[127] ^ in2[127];
    assign G[66] = in[126] & in2[126];
    assign P[66] = in[126] ^ in2[126];
    assign G[67] = in[125] & in2[125];
    assign P[67] = in[125] ^ in2[125];
    assign G[68] = in[124] & in2[124];
    assign P[68] = in[124] ^ in2[124];
    assign G[69] = in[123] & in2[123];
    assign P[69] = in[123] ^ in2[123];
    assign G[70] = in[122] & in2[122];
    assign P[70] = in[122] ^ in2[122];
    assign G[71] = in[121] & in2[121];
    assign P[71] = in[121] ^ in2[121];
    assign G[72] = in[120] & in2[120];
    assign P[72] = in[120] ^ in2[120];
    assign G[73] = in[119] & in2[119];
    assign P[73] = in[119] ^ in2[119];
    assign G[74] = in[118] & in2[118];
    assign P[74] = in[118] ^ in2[118];
    assign G[75] = in[117] & in2[117];
    assign P[75] = in[117] ^ in2[117];
    assign G[76] = in[116] & in2[116];
    assign P[76] = in[116] ^ in2[116];
    assign G[77] = in[115] & in2[115];
    assign P[77] = in[115] ^ in2[115];
    assign G[78] = in[114] & in2[114];
    assign P[78] = in[114] ^ in2[114];
    assign G[79] = in[113] & in2[113];
    assign P[79] = in[113] ^ in2[113];
    assign G[80] = in[112] & in2[112];
    assign P[80] = in[112] ^ in2[112];
    assign G[81] = in[111] & in2[111];
    assign P[81] = in[111] ^ in2[111];
    assign G[82] = in[110] & in2[110];
    assign P[82] = in[110] ^ in2[110];
    assign G[83] = in[109] & in2[109];
    assign P[83] = in[109] ^ in2[109];
    assign G[84] = in[108] & in2[108];
    assign P[84] = in[108] ^ in2[108];
    assign G[85] = in[107] & in2[107];
    assign P[85] = in[107] ^ in2[107];
    assign G[86] = in[106] & in2[106];
    assign P[86] = in[106] ^ in2[106];
    assign G[87] = in[105] & in2[105];
    assign P[87] = in[105] ^ in2[105];
    assign G[88] = in[104] & in2[104];
    assign P[88] = in[104] ^ in2[104];
    assign G[89] = in[103] & in2[103];
    assign P[89] = in[103] ^ in2[103];
    assign G[90] = in[102] & in2[102];
    assign P[90] = in[102] ^ in2[102];
    assign G[91] = in[101] & in2[101];
    assign P[91] = in[101] ^ in2[101];
    assign G[92] = in[100] & in2[100];
    assign P[92] = in[100] ^ in2[100];
    assign G[93] = in[99] & in2[99];
    assign P[93] = in[99] ^ in2[99];
    assign G[94] = in[98] & in2[98];
    assign P[94] = in[98] ^ in2[98];
    assign G[95] = in[97] & in2[97];
    assign P[95] = in[97] ^ in2[97];
    assign G[96] = in[96] & in2[96];
    assign P[96] = in[96] ^ in2[96];
    assign G[97] = in[95] & in2[95];
    assign P[97] = in[95] ^ in2[95];
    assign G[98] = in[94] & in2[94];
    assign P[98] = in[94] ^ in2[94];
    assign G[99] = in[93] & in2[93];
    assign P[99] = in[93] ^ in2[93];
    assign G[100] = in[92] & in2[92];
    assign P[100] = in[92] ^ in2[92];
    assign G[101] = in[91] & in2[91];
    assign P[101] = in[91] ^ in2[91];
    assign G[102] = in[90] & in2[90];
    assign P[102] = in[90] ^ in2[90];
    assign G[103] = in[89] & in2[89];
    assign P[103] = in[89] ^ in2[89];
    assign G[104] = in[88] & in2[88];
    assign P[104] = in[88] ^ in2[88];
    assign G[105] = in[87] & in2[87];
    assign P[105] = in[87] ^ in2[87];
    assign G[106] = in[86] & in2[86];
    assign P[106] = in[86] ^ in2[86];
    assign G[107] = in[85] & in2[85];
    assign P[107] = in[85] ^ in2[85];
    assign G[108] = in[84] & in2[84];
    assign P[108] = in[84] ^ in2[84];
    assign G[109] = in[83] & in2[83];
    assign P[109] = in[83] ^ in2[83];
    assign G[110] = in[82] & in2[82];
    assign P[110] = in[82] ^ in2[82];
    assign G[111] = in[81] & in2[81];
    assign P[111] = in[81] ^ in2[81];
    assign G[112] = in[80] & in2[80];
    assign P[112] = in[80] ^ in2[80];
    assign G[113] = in[79] & in2[79];
    assign P[113] = in[79] ^ in2[79];
    assign G[114] = in[78] & in2[78];
    assign P[114] = in[78] ^ in2[78];
    assign G[115] = in[77] & in2[77];
    assign P[115] = in[77] ^ in2[77];
    assign G[116] = in[76] & in2[76];
    assign P[116] = in[76] ^ in2[76];
    assign G[117] = in[75] & in2[75];
    assign P[117] = in[75] ^ in2[75];
    assign G[118] = in[74] & in2[74];
    assign P[118] = in[74] ^ in2[74];
    assign G[119] = in[73] & in2[73];
    assign P[119] = in[73] ^ in2[73];
    assign G[120] = in[72] & in2[72];
    assign P[120] = in[72] ^ in2[72];
    assign G[121] = in[71] & in2[71];
    assign P[121] = in[71] ^ in2[71];
    assign G[122] = in[70] & in2[70];
    assign P[122] = in[70] ^ in2[70];
    assign G[123] = in[69] & in2[69];
    assign P[123] = in[69] ^ in2[69];
    assign G[124] = in[68] & in2[68];
    assign P[124] = in[68] ^ in2[68];
    assign G[125] = in[67] & in2[67];
    assign P[125] = in[67] ^ in2[67];
    assign G[126] = in[66] & in2[66];
    assign P[126] = in[66] ^ in2[66];
    assign G[127] = in[65] & in2[65];
    assign P[127] = in[65] ^ in2[65];
    assign G[128] = in[64] & in2[64];
    assign P[128] = in[64] ^ in2[64];
    assign G[129] = in[63] & in2[63];
    assign P[129] = in[63] ^ in2[63];
    assign G[130] = in[62] & in2[62];
    assign P[130] = in[62] ^ in2[62];
    assign G[131] = in[61] & in2[61];
    assign P[131] = in[61] ^ in2[61];
    assign G[132] = in[60] & in2[60];
    assign P[132] = in[60] ^ in2[60];
    assign G[133] = in[59] & in2[59];
    assign P[133] = in[59] ^ in2[59];
    assign G[134] = in[58] & in2[58];
    assign P[134] = in[58] ^ in2[58];
    assign G[135] = in[57] & in2[57];
    assign P[135] = in[57] ^ in2[57];
    assign G[136] = in[56] & in2[56];
    assign P[136] = in[56] ^ in2[56];
    assign G[137] = in[55] & in2[55];
    assign P[137] = in[55] ^ in2[55];
    assign G[138] = in[54] & in2[54];
    assign P[138] = in[54] ^ in2[54];
    assign G[139] = in[53] & in2[53];
    assign P[139] = in[53] ^ in2[53];
    assign G[140] = in[52] & in2[52];
    assign P[140] = in[52] ^ in2[52];
    assign G[141] = in[51] & in2[51];
    assign P[141] = in[51] ^ in2[51];
    assign G[142] = in[50] & in2[50];
    assign P[142] = in[50] ^ in2[50];
    assign G[143] = in[49] & in2[49];
    assign P[143] = in[49] ^ in2[49];
    assign G[144] = in[48] & in2[48];
    assign P[144] = in[48] ^ in2[48];
    assign G[145] = in[47] & in2[47];
    assign P[145] = in[47] ^ in2[47];
    assign G[146] = in[46] & in2[46];
    assign P[146] = in[46] ^ in2[46];
    assign G[147] = in[45] & in2[45];
    assign P[147] = in[45] ^ in2[45];
    assign G[148] = in[44] & in2[44];
    assign P[148] = in[44] ^ in2[44];
    assign G[149] = in[43] & in2[43];
    assign P[149] = in[43] ^ in2[43];
    assign G[150] = in[42] & in2[42];
    assign P[150] = in[42] ^ in2[42];
    assign G[151] = in[41] & in2[41];
    assign P[151] = in[41] ^ in2[41];
    assign G[152] = in[40] & in2[40];
    assign P[152] = in[40] ^ in2[40];
    assign G[153] = in[39] & in2[39];
    assign P[153] = in[39] ^ in2[39];
    assign G[154] = in[38] & in2[38];
    assign P[154] = in[38] ^ in2[38];
    assign G[155] = in[37] & in2[37];
    assign P[155] = in[37] ^ in2[37];
    assign G[156] = in[36] & in2[36];
    assign P[156] = in[36] ^ in2[36];
    assign G[157] = in[35] & in2[35];
    assign P[157] = in[35] ^ in2[35];
    assign G[158] = in[34] & in2[34];
    assign P[158] = in[34] ^ in2[34];
    assign G[159] = in[33] & in2[33];
    assign P[159] = in[33] ^ in2[33];
    assign G[160] = in[32] & in2[32];
    assign P[160] = in[32] ^ in2[32];
    assign G[161] = in[31] & in2[31];
    assign P[161] = in[31] ^ in2[31];
    assign G[162] = in[30] & in2[30];
    assign P[162] = in[30] ^ in2[30];
    assign G[163] = in[29] & in2[29];
    assign P[163] = in[29] ^ in2[29];
    assign G[164] = in[28] & in2[28];
    assign P[164] = in[28] ^ in2[28];
    assign G[165] = in[27] & in2[27];
    assign P[165] = in[27] ^ in2[27];
    assign G[166] = in[26] & in2[26];
    assign P[166] = in[26] ^ in2[26];
    assign G[167] = in[25] & in2[25];
    assign P[167] = in[25] ^ in2[25];
    assign G[168] = in[24] & in2[24];
    assign P[168] = in[24] ^ in2[24];
    assign G[169] = in[23] & in2[23];
    assign P[169] = in[23] ^ in2[23];
    assign G[170] = in[22] & in2[22];
    assign P[170] = in[22] ^ in2[22];
    assign G[171] = in[21] & in2[21];
    assign P[171] = in[21] ^ in2[21];
    assign G[172] = in[20] & in2[20];
    assign P[172] = in[20] ^ in2[20];
    assign G[173] = in[19] & in2[19];
    assign P[173] = in[19] ^ in2[19];
    assign G[174] = in[18] & in2[18];
    assign P[174] = in[18] ^ in2[18];
    assign G[175] = in[17] & in2[17];
    assign P[175] = in[17] ^ in2[17];
    assign G[176] = in[16] & in2[16];
    assign P[176] = in[16] ^ in2[16];
    assign G[177] = in[15] & in2[15];
    assign P[177] = in[15] ^ in2[15];
    assign G[178] = in[14] & in2[14];
    assign P[178] = in[14] ^ in2[14];
    assign G[179] = in[13] & in2[13];
    assign P[179] = in[13] ^ in2[13];
    assign G[180] = in[12] & in2[12];
    assign P[180] = in[12] ^ in2[12];
    assign G[181] = in[11] & in2[11];
    assign P[181] = in[11] ^ in2[11];
    assign G[182] = in[10] & in2[10];
    assign P[182] = in[10] ^ in2[10];
    assign G[183] = in[9] & in2[9];
    assign P[183] = in[9] ^ in2[9];
    assign G[184] = in[8] & in2[8];
    assign P[184] = in[8] ^ in2[8];
    assign G[185] = in[7] & in2[7];
    assign P[185] = in[7] ^ in2[7];
    assign G[186] = in[6] & in2[6];
    assign P[186] = in[6] ^ in2[6];
    assign G[187] = in[5] & in2[5];
    assign P[187] = in[5] ^ in2[5];
    assign G[188] = in[4] & in2[4];
    assign P[188] = in[4] ^ in2[4];
    assign G[189] = in[3] & in2[3];
    assign P[189] = in[3] ^ in2[3];
    assign G[190] = in[2] & in2[2];
    assign P[190] = in[2] ^ in2[2];
    assign G[191] = in[1] & in2[1];
    assign P[191] = in[1] ^ in2[1];
    assign G[192] = in[0] & in2[0];
    assign P[192] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign C[192] = G[191] | (P[191] & C[191]);
    assign cout = G[192] | (P[192] & C[192]);
    assign sum = P ^ C;
endmodule

module CLA192(output [191:0] sum, output cout, input [191:0] in1, input [191:0] in2;

    wire[191:0] G;
    wire[191:0] C;
    wire[191:0] P;

    assign G[0] = in[191] & in2[191];
    assign P[0] = in[191] ^ in2[191];
    assign G[1] = in[190] & in2[190];
    assign P[1] = in[190] ^ in2[190];
    assign G[2] = in[189] & in2[189];
    assign P[2] = in[189] ^ in2[189];
    assign G[3] = in[188] & in2[188];
    assign P[3] = in[188] ^ in2[188];
    assign G[4] = in[187] & in2[187];
    assign P[4] = in[187] ^ in2[187];
    assign G[5] = in[186] & in2[186];
    assign P[5] = in[186] ^ in2[186];
    assign G[6] = in[185] & in2[185];
    assign P[6] = in[185] ^ in2[185];
    assign G[7] = in[184] & in2[184];
    assign P[7] = in[184] ^ in2[184];
    assign G[8] = in[183] & in2[183];
    assign P[8] = in[183] ^ in2[183];
    assign G[9] = in[182] & in2[182];
    assign P[9] = in[182] ^ in2[182];
    assign G[10] = in[181] & in2[181];
    assign P[10] = in[181] ^ in2[181];
    assign G[11] = in[180] & in2[180];
    assign P[11] = in[180] ^ in2[180];
    assign G[12] = in[179] & in2[179];
    assign P[12] = in[179] ^ in2[179];
    assign G[13] = in[178] & in2[178];
    assign P[13] = in[178] ^ in2[178];
    assign G[14] = in[177] & in2[177];
    assign P[14] = in[177] ^ in2[177];
    assign G[15] = in[176] & in2[176];
    assign P[15] = in[176] ^ in2[176];
    assign G[16] = in[175] & in2[175];
    assign P[16] = in[175] ^ in2[175];
    assign G[17] = in[174] & in2[174];
    assign P[17] = in[174] ^ in2[174];
    assign G[18] = in[173] & in2[173];
    assign P[18] = in[173] ^ in2[173];
    assign G[19] = in[172] & in2[172];
    assign P[19] = in[172] ^ in2[172];
    assign G[20] = in[171] & in2[171];
    assign P[20] = in[171] ^ in2[171];
    assign G[21] = in[170] & in2[170];
    assign P[21] = in[170] ^ in2[170];
    assign G[22] = in[169] & in2[169];
    assign P[22] = in[169] ^ in2[169];
    assign G[23] = in[168] & in2[168];
    assign P[23] = in[168] ^ in2[168];
    assign G[24] = in[167] & in2[167];
    assign P[24] = in[167] ^ in2[167];
    assign G[25] = in[166] & in2[166];
    assign P[25] = in[166] ^ in2[166];
    assign G[26] = in[165] & in2[165];
    assign P[26] = in[165] ^ in2[165];
    assign G[27] = in[164] & in2[164];
    assign P[27] = in[164] ^ in2[164];
    assign G[28] = in[163] & in2[163];
    assign P[28] = in[163] ^ in2[163];
    assign G[29] = in[162] & in2[162];
    assign P[29] = in[162] ^ in2[162];
    assign G[30] = in[161] & in2[161];
    assign P[30] = in[161] ^ in2[161];
    assign G[31] = in[160] & in2[160];
    assign P[31] = in[160] ^ in2[160];
    assign G[32] = in[159] & in2[159];
    assign P[32] = in[159] ^ in2[159];
    assign G[33] = in[158] & in2[158];
    assign P[33] = in[158] ^ in2[158];
    assign G[34] = in[157] & in2[157];
    assign P[34] = in[157] ^ in2[157];
    assign G[35] = in[156] & in2[156];
    assign P[35] = in[156] ^ in2[156];
    assign G[36] = in[155] & in2[155];
    assign P[36] = in[155] ^ in2[155];
    assign G[37] = in[154] & in2[154];
    assign P[37] = in[154] ^ in2[154];
    assign G[38] = in[153] & in2[153];
    assign P[38] = in[153] ^ in2[153];
    assign G[39] = in[152] & in2[152];
    assign P[39] = in[152] ^ in2[152];
    assign G[40] = in[151] & in2[151];
    assign P[40] = in[151] ^ in2[151];
    assign G[41] = in[150] & in2[150];
    assign P[41] = in[150] ^ in2[150];
    assign G[42] = in[149] & in2[149];
    assign P[42] = in[149] ^ in2[149];
    assign G[43] = in[148] & in2[148];
    assign P[43] = in[148] ^ in2[148];
    assign G[44] = in[147] & in2[147];
    assign P[44] = in[147] ^ in2[147];
    assign G[45] = in[146] & in2[146];
    assign P[45] = in[146] ^ in2[146];
    assign G[46] = in[145] & in2[145];
    assign P[46] = in[145] ^ in2[145];
    assign G[47] = in[144] & in2[144];
    assign P[47] = in[144] ^ in2[144];
    assign G[48] = in[143] & in2[143];
    assign P[48] = in[143] ^ in2[143];
    assign G[49] = in[142] & in2[142];
    assign P[49] = in[142] ^ in2[142];
    assign G[50] = in[141] & in2[141];
    assign P[50] = in[141] ^ in2[141];
    assign G[51] = in[140] & in2[140];
    assign P[51] = in[140] ^ in2[140];
    assign G[52] = in[139] & in2[139];
    assign P[52] = in[139] ^ in2[139];
    assign G[53] = in[138] & in2[138];
    assign P[53] = in[138] ^ in2[138];
    assign G[54] = in[137] & in2[137];
    assign P[54] = in[137] ^ in2[137];
    assign G[55] = in[136] & in2[136];
    assign P[55] = in[136] ^ in2[136];
    assign G[56] = in[135] & in2[135];
    assign P[56] = in[135] ^ in2[135];
    assign G[57] = in[134] & in2[134];
    assign P[57] = in[134] ^ in2[134];
    assign G[58] = in[133] & in2[133];
    assign P[58] = in[133] ^ in2[133];
    assign G[59] = in[132] & in2[132];
    assign P[59] = in[132] ^ in2[132];
    assign G[60] = in[131] & in2[131];
    assign P[60] = in[131] ^ in2[131];
    assign G[61] = in[130] & in2[130];
    assign P[61] = in[130] ^ in2[130];
    assign G[62] = in[129] & in2[129];
    assign P[62] = in[129] ^ in2[129];
    assign G[63] = in[128] & in2[128];
    assign P[63] = in[128] ^ in2[128];
    assign G[64] = in[127] & in2[127];
    assign P[64] = in[127] ^ in2[127];
    assign G[65] = in[126] & in2[126];
    assign P[65] = in[126] ^ in2[126];
    assign G[66] = in[125] & in2[125];
    assign P[66] = in[125] ^ in2[125];
    assign G[67] = in[124] & in2[124];
    assign P[67] = in[124] ^ in2[124];
    assign G[68] = in[123] & in2[123];
    assign P[68] = in[123] ^ in2[123];
    assign G[69] = in[122] & in2[122];
    assign P[69] = in[122] ^ in2[122];
    assign G[70] = in[121] & in2[121];
    assign P[70] = in[121] ^ in2[121];
    assign G[71] = in[120] & in2[120];
    assign P[71] = in[120] ^ in2[120];
    assign G[72] = in[119] & in2[119];
    assign P[72] = in[119] ^ in2[119];
    assign G[73] = in[118] & in2[118];
    assign P[73] = in[118] ^ in2[118];
    assign G[74] = in[117] & in2[117];
    assign P[74] = in[117] ^ in2[117];
    assign G[75] = in[116] & in2[116];
    assign P[75] = in[116] ^ in2[116];
    assign G[76] = in[115] & in2[115];
    assign P[76] = in[115] ^ in2[115];
    assign G[77] = in[114] & in2[114];
    assign P[77] = in[114] ^ in2[114];
    assign G[78] = in[113] & in2[113];
    assign P[78] = in[113] ^ in2[113];
    assign G[79] = in[112] & in2[112];
    assign P[79] = in[112] ^ in2[112];
    assign G[80] = in[111] & in2[111];
    assign P[80] = in[111] ^ in2[111];
    assign G[81] = in[110] & in2[110];
    assign P[81] = in[110] ^ in2[110];
    assign G[82] = in[109] & in2[109];
    assign P[82] = in[109] ^ in2[109];
    assign G[83] = in[108] & in2[108];
    assign P[83] = in[108] ^ in2[108];
    assign G[84] = in[107] & in2[107];
    assign P[84] = in[107] ^ in2[107];
    assign G[85] = in[106] & in2[106];
    assign P[85] = in[106] ^ in2[106];
    assign G[86] = in[105] & in2[105];
    assign P[86] = in[105] ^ in2[105];
    assign G[87] = in[104] & in2[104];
    assign P[87] = in[104] ^ in2[104];
    assign G[88] = in[103] & in2[103];
    assign P[88] = in[103] ^ in2[103];
    assign G[89] = in[102] & in2[102];
    assign P[89] = in[102] ^ in2[102];
    assign G[90] = in[101] & in2[101];
    assign P[90] = in[101] ^ in2[101];
    assign G[91] = in[100] & in2[100];
    assign P[91] = in[100] ^ in2[100];
    assign G[92] = in[99] & in2[99];
    assign P[92] = in[99] ^ in2[99];
    assign G[93] = in[98] & in2[98];
    assign P[93] = in[98] ^ in2[98];
    assign G[94] = in[97] & in2[97];
    assign P[94] = in[97] ^ in2[97];
    assign G[95] = in[96] & in2[96];
    assign P[95] = in[96] ^ in2[96];
    assign G[96] = in[95] & in2[95];
    assign P[96] = in[95] ^ in2[95];
    assign G[97] = in[94] & in2[94];
    assign P[97] = in[94] ^ in2[94];
    assign G[98] = in[93] & in2[93];
    assign P[98] = in[93] ^ in2[93];
    assign G[99] = in[92] & in2[92];
    assign P[99] = in[92] ^ in2[92];
    assign G[100] = in[91] & in2[91];
    assign P[100] = in[91] ^ in2[91];
    assign G[101] = in[90] & in2[90];
    assign P[101] = in[90] ^ in2[90];
    assign G[102] = in[89] & in2[89];
    assign P[102] = in[89] ^ in2[89];
    assign G[103] = in[88] & in2[88];
    assign P[103] = in[88] ^ in2[88];
    assign G[104] = in[87] & in2[87];
    assign P[104] = in[87] ^ in2[87];
    assign G[105] = in[86] & in2[86];
    assign P[105] = in[86] ^ in2[86];
    assign G[106] = in[85] & in2[85];
    assign P[106] = in[85] ^ in2[85];
    assign G[107] = in[84] & in2[84];
    assign P[107] = in[84] ^ in2[84];
    assign G[108] = in[83] & in2[83];
    assign P[108] = in[83] ^ in2[83];
    assign G[109] = in[82] & in2[82];
    assign P[109] = in[82] ^ in2[82];
    assign G[110] = in[81] & in2[81];
    assign P[110] = in[81] ^ in2[81];
    assign G[111] = in[80] & in2[80];
    assign P[111] = in[80] ^ in2[80];
    assign G[112] = in[79] & in2[79];
    assign P[112] = in[79] ^ in2[79];
    assign G[113] = in[78] & in2[78];
    assign P[113] = in[78] ^ in2[78];
    assign G[114] = in[77] & in2[77];
    assign P[114] = in[77] ^ in2[77];
    assign G[115] = in[76] & in2[76];
    assign P[115] = in[76] ^ in2[76];
    assign G[116] = in[75] & in2[75];
    assign P[116] = in[75] ^ in2[75];
    assign G[117] = in[74] & in2[74];
    assign P[117] = in[74] ^ in2[74];
    assign G[118] = in[73] & in2[73];
    assign P[118] = in[73] ^ in2[73];
    assign G[119] = in[72] & in2[72];
    assign P[119] = in[72] ^ in2[72];
    assign G[120] = in[71] & in2[71];
    assign P[120] = in[71] ^ in2[71];
    assign G[121] = in[70] & in2[70];
    assign P[121] = in[70] ^ in2[70];
    assign G[122] = in[69] & in2[69];
    assign P[122] = in[69] ^ in2[69];
    assign G[123] = in[68] & in2[68];
    assign P[123] = in[68] ^ in2[68];
    assign G[124] = in[67] & in2[67];
    assign P[124] = in[67] ^ in2[67];
    assign G[125] = in[66] & in2[66];
    assign P[125] = in[66] ^ in2[66];
    assign G[126] = in[65] & in2[65];
    assign P[126] = in[65] ^ in2[65];
    assign G[127] = in[64] & in2[64];
    assign P[127] = in[64] ^ in2[64];
    assign G[128] = in[63] & in2[63];
    assign P[128] = in[63] ^ in2[63];
    assign G[129] = in[62] & in2[62];
    assign P[129] = in[62] ^ in2[62];
    assign G[130] = in[61] & in2[61];
    assign P[130] = in[61] ^ in2[61];
    assign G[131] = in[60] & in2[60];
    assign P[131] = in[60] ^ in2[60];
    assign G[132] = in[59] & in2[59];
    assign P[132] = in[59] ^ in2[59];
    assign G[133] = in[58] & in2[58];
    assign P[133] = in[58] ^ in2[58];
    assign G[134] = in[57] & in2[57];
    assign P[134] = in[57] ^ in2[57];
    assign G[135] = in[56] & in2[56];
    assign P[135] = in[56] ^ in2[56];
    assign G[136] = in[55] & in2[55];
    assign P[136] = in[55] ^ in2[55];
    assign G[137] = in[54] & in2[54];
    assign P[137] = in[54] ^ in2[54];
    assign G[138] = in[53] & in2[53];
    assign P[138] = in[53] ^ in2[53];
    assign G[139] = in[52] & in2[52];
    assign P[139] = in[52] ^ in2[52];
    assign G[140] = in[51] & in2[51];
    assign P[140] = in[51] ^ in2[51];
    assign G[141] = in[50] & in2[50];
    assign P[141] = in[50] ^ in2[50];
    assign G[142] = in[49] & in2[49];
    assign P[142] = in[49] ^ in2[49];
    assign G[143] = in[48] & in2[48];
    assign P[143] = in[48] ^ in2[48];
    assign G[144] = in[47] & in2[47];
    assign P[144] = in[47] ^ in2[47];
    assign G[145] = in[46] & in2[46];
    assign P[145] = in[46] ^ in2[46];
    assign G[146] = in[45] & in2[45];
    assign P[146] = in[45] ^ in2[45];
    assign G[147] = in[44] & in2[44];
    assign P[147] = in[44] ^ in2[44];
    assign G[148] = in[43] & in2[43];
    assign P[148] = in[43] ^ in2[43];
    assign G[149] = in[42] & in2[42];
    assign P[149] = in[42] ^ in2[42];
    assign G[150] = in[41] & in2[41];
    assign P[150] = in[41] ^ in2[41];
    assign G[151] = in[40] & in2[40];
    assign P[151] = in[40] ^ in2[40];
    assign G[152] = in[39] & in2[39];
    assign P[152] = in[39] ^ in2[39];
    assign G[153] = in[38] & in2[38];
    assign P[153] = in[38] ^ in2[38];
    assign G[154] = in[37] & in2[37];
    assign P[154] = in[37] ^ in2[37];
    assign G[155] = in[36] & in2[36];
    assign P[155] = in[36] ^ in2[36];
    assign G[156] = in[35] & in2[35];
    assign P[156] = in[35] ^ in2[35];
    assign G[157] = in[34] & in2[34];
    assign P[157] = in[34] ^ in2[34];
    assign G[158] = in[33] & in2[33];
    assign P[158] = in[33] ^ in2[33];
    assign G[159] = in[32] & in2[32];
    assign P[159] = in[32] ^ in2[32];
    assign G[160] = in[31] & in2[31];
    assign P[160] = in[31] ^ in2[31];
    assign G[161] = in[30] & in2[30];
    assign P[161] = in[30] ^ in2[30];
    assign G[162] = in[29] & in2[29];
    assign P[162] = in[29] ^ in2[29];
    assign G[163] = in[28] & in2[28];
    assign P[163] = in[28] ^ in2[28];
    assign G[164] = in[27] & in2[27];
    assign P[164] = in[27] ^ in2[27];
    assign G[165] = in[26] & in2[26];
    assign P[165] = in[26] ^ in2[26];
    assign G[166] = in[25] & in2[25];
    assign P[166] = in[25] ^ in2[25];
    assign G[167] = in[24] & in2[24];
    assign P[167] = in[24] ^ in2[24];
    assign G[168] = in[23] & in2[23];
    assign P[168] = in[23] ^ in2[23];
    assign G[169] = in[22] & in2[22];
    assign P[169] = in[22] ^ in2[22];
    assign G[170] = in[21] & in2[21];
    assign P[170] = in[21] ^ in2[21];
    assign G[171] = in[20] & in2[20];
    assign P[171] = in[20] ^ in2[20];
    assign G[172] = in[19] & in2[19];
    assign P[172] = in[19] ^ in2[19];
    assign G[173] = in[18] & in2[18];
    assign P[173] = in[18] ^ in2[18];
    assign G[174] = in[17] & in2[17];
    assign P[174] = in[17] ^ in2[17];
    assign G[175] = in[16] & in2[16];
    assign P[175] = in[16] ^ in2[16];
    assign G[176] = in[15] & in2[15];
    assign P[176] = in[15] ^ in2[15];
    assign G[177] = in[14] & in2[14];
    assign P[177] = in[14] ^ in2[14];
    assign G[178] = in[13] & in2[13];
    assign P[178] = in[13] ^ in2[13];
    assign G[179] = in[12] & in2[12];
    assign P[179] = in[12] ^ in2[12];
    assign G[180] = in[11] & in2[11];
    assign P[180] = in[11] ^ in2[11];
    assign G[181] = in[10] & in2[10];
    assign P[181] = in[10] ^ in2[10];
    assign G[182] = in[9] & in2[9];
    assign P[182] = in[9] ^ in2[9];
    assign G[183] = in[8] & in2[8];
    assign P[183] = in[8] ^ in2[8];
    assign G[184] = in[7] & in2[7];
    assign P[184] = in[7] ^ in2[7];
    assign G[185] = in[6] & in2[6];
    assign P[185] = in[6] ^ in2[6];
    assign G[186] = in[5] & in2[5];
    assign P[186] = in[5] ^ in2[5];
    assign G[187] = in[4] & in2[4];
    assign P[187] = in[4] ^ in2[4];
    assign G[188] = in[3] & in2[3];
    assign P[188] = in[3] ^ in2[3];
    assign G[189] = in[2] & in2[2];
    assign P[189] = in[2] ^ in2[2];
    assign G[190] = in[1] & in2[1];
    assign P[190] = in[1] ^ in2[1];
    assign G[191] = in[0] & in2[0];
    assign P[191] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign C[191] = G[190] | (P[190] & C[190]);
    assign cout = G[191] | (P[191] & C[191]);
    assign sum = P ^ C;
endmodule

module CLA191(output [190:0] sum, output cout, input [190:0] in1, input [190:0] in2;

    wire[190:0] G;
    wire[190:0] C;
    wire[190:0] P;

    assign G[0] = in[190] & in2[190];
    assign P[0] = in[190] ^ in2[190];
    assign G[1] = in[189] & in2[189];
    assign P[1] = in[189] ^ in2[189];
    assign G[2] = in[188] & in2[188];
    assign P[2] = in[188] ^ in2[188];
    assign G[3] = in[187] & in2[187];
    assign P[3] = in[187] ^ in2[187];
    assign G[4] = in[186] & in2[186];
    assign P[4] = in[186] ^ in2[186];
    assign G[5] = in[185] & in2[185];
    assign P[5] = in[185] ^ in2[185];
    assign G[6] = in[184] & in2[184];
    assign P[6] = in[184] ^ in2[184];
    assign G[7] = in[183] & in2[183];
    assign P[7] = in[183] ^ in2[183];
    assign G[8] = in[182] & in2[182];
    assign P[8] = in[182] ^ in2[182];
    assign G[9] = in[181] & in2[181];
    assign P[9] = in[181] ^ in2[181];
    assign G[10] = in[180] & in2[180];
    assign P[10] = in[180] ^ in2[180];
    assign G[11] = in[179] & in2[179];
    assign P[11] = in[179] ^ in2[179];
    assign G[12] = in[178] & in2[178];
    assign P[12] = in[178] ^ in2[178];
    assign G[13] = in[177] & in2[177];
    assign P[13] = in[177] ^ in2[177];
    assign G[14] = in[176] & in2[176];
    assign P[14] = in[176] ^ in2[176];
    assign G[15] = in[175] & in2[175];
    assign P[15] = in[175] ^ in2[175];
    assign G[16] = in[174] & in2[174];
    assign P[16] = in[174] ^ in2[174];
    assign G[17] = in[173] & in2[173];
    assign P[17] = in[173] ^ in2[173];
    assign G[18] = in[172] & in2[172];
    assign P[18] = in[172] ^ in2[172];
    assign G[19] = in[171] & in2[171];
    assign P[19] = in[171] ^ in2[171];
    assign G[20] = in[170] & in2[170];
    assign P[20] = in[170] ^ in2[170];
    assign G[21] = in[169] & in2[169];
    assign P[21] = in[169] ^ in2[169];
    assign G[22] = in[168] & in2[168];
    assign P[22] = in[168] ^ in2[168];
    assign G[23] = in[167] & in2[167];
    assign P[23] = in[167] ^ in2[167];
    assign G[24] = in[166] & in2[166];
    assign P[24] = in[166] ^ in2[166];
    assign G[25] = in[165] & in2[165];
    assign P[25] = in[165] ^ in2[165];
    assign G[26] = in[164] & in2[164];
    assign P[26] = in[164] ^ in2[164];
    assign G[27] = in[163] & in2[163];
    assign P[27] = in[163] ^ in2[163];
    assign G[28] = in[162] & in2[162];
    assign P[28] = in[162] ^ in2[162];
    assign G[29] = in[161] & in2[161];
    assign P[29] = in[161] ^ in2[161];
    assign G[30] = in[160] & in2[160];
    assign P[30] = in[160] ^ in2[160];
    assign G[31] = in[159] & in2[159];
    assign P[31] = in[159] ^ in2[159];
    assign G[32] = in[158] & in2[158];
    assign P[32] = in[158] ^ in2[158];
    assign G[33] = in[157] & in2[157];
    assign P[33] = in[157] ^ in2[157];
    assign G[34] = in[156] & in2[156];
    assign P[34] = in[156] ^ in2[156];
    assign G[35] = in[155] & in2[155];
    assign P[35] = in[155] ^ in2[155];
    assign G[36] = in[154] & in2[154];
    assign P[36] = in[154] ^ in2[154];
    assign G[37] = in[153] & in2[153];
    assign P[37] = in[153] ^ in2[153];
    assign G[38] = in[152] & in2[152];
    assign P[38] = in[152] ^ in2[152];
    assign G[39] = in[151] & in2[151];
    assign P[39] = in[151] ^ in2[151];
    assign G[40] = in[150] & in2[150];
    assign P[40] = in[150] ^ in2[150];
    assign G[41] = in[149] & in2[149];
    assign P[41] = in[149] ^ in2[149];
    assign G[42] = in[148] & in2[148];
    assign P[42] = in[148] ^ in2[148];
    assign G[43] = in[147] & in2[147];
    assign P[43] = in[147] ^ in2[147];
    assign G[44] = in[146] & in2[146];
    assign P[44] = in[146] ^ in2[146];
    assign G[45] = in[145] & in2[145];
    assign P[45] = in[145] ^ in2[145];
    assign G[46] = in[144] & in2[144];
    assign P[46] = in[144] ^ in2[144];
    assign G[47] = in[143] & in2[143];
    assign P[47] = in[143] ^ in2[143];
    assign G[48] = in[142] & in2[142];
    assign P[48] = in[142] ^ in2[142];
    assign G[49] = in[141] & in2[141];
    assign P[49] = in[141] ^ in2[141];
    assign G[50] = in[140] & in2[140];
    assign P[50] = in[140] ^ in2[140];
    assign G[51] = in[139] & in2[139];
    assign P[51] = in[139] ^ in2[139];
    assign G[52] = in[138] & in2[138];
    assign P[52] = in[138] ^ in2[138];
    assign G[53] = in[137] & in2[137];
    assign P[53] = in[137] ^ in2[137];
    assign G[54] = in[136] & in2[136];
    assign P[54] = in[136] ^ in2[136];
    assign G[55] = in[135] & in2[135];
    assign P[55] = in[135] ^ in2[135];
    assign G[56] = in[134] & in2[134];
    assign P[56] = in[134] ^ in2[134];
    assign G[57] = in[133] & in2[133];
    assign P[57] = in[133] ^ in2[133];
    assign G[58] = in[132] & in2[132];
    assign P[58] = in[132] ^ in2[132];
    assign G[59] = in[131] & in2[131];
    assign P[59] = in[131] ^ in2[131];
    assign G[60] = in[130] & in2[130];
    assign P[60] = in[130] ^ in2[130];
    assign G[61] = in[129] & in2[129];
    assign P[61] = in[129] ^ in2[129];
    assign G[62] = in[128] & in2[128];
    assign P[62] = in[128] ^ in2[128];
    assign G[63] = in[127] & in2[127];
    assign P[63] = in[127] ^ in2[127];
    assign G[64] = in[126] & in2[126];
    assign P[64] = in[126] ^ in2[126];
    assign G[65] = in[125] & in2[125];
    assign P[65] = in[125] ^ in2[125];
    assign G[66] = in[124] & in2[124];
    assign P[66] = in[124] ^ in2[124];
    assign G[67] = in[123] & in2[123];
    assign P[67] = in[123] ^ in2[123];
    assign G[68] = in[122] & in2[122];
    assign P[68] = in[122] ^ in2[122];
    assign G[69] = in[121] & in2[121];
    assign P[69] = in[121] ^ in2[121];
    assign G[70] = in[120] & in2[120];
    assign P[70] = in[120] ^ in2[120];
    assign G[71] = in[119] & in2[119];
    assign P[71] = in[119] ^ in2[119];
    assign G[72] = in[118] & in2[118];
    assign P[72] = in[118] ^ in2[118];
    assign G[73] = in[117] & in2[117];
    assign P[73] = in[117] ^ in2[117];
    assign G[74] = in[116] & in2[116];
    assign P[74] = in[116] ^ in2[116];
    assign G[75] = in[115] & in2[115];
    assign P[75] = in[115] ^ in2[115];
    assign G[76] = in[114] & in2[114];
    assign P[76] = in[114] ^ in2[114];
    assign G[77] = in[113] & in2[113];
    assign P[77] = in[113] ^ in2[113];
    assign G[78] = in[112] & in2[112];
    assign P[78] = in[112] ^ in2[112];
    assign G[79] = in[111] & in2[111];
    assign P[79] = in[111] ^ in2[111];
    assign G[80] = in[110] & in2[110];
    assign P[80] = in[110] ^ in2[110];
    assign G[81] = in[109] & in2[109];
    assign P[81] = in[109] ^ in2[109];
    assign G[82] = in[108] & in2[108];
    assign P[82] = in[108] ^ in2[108];
    assign G[83] = in[107] & in2[107];
    assign P[83] = in[107] ^ in2[107];
    assign G[84] = in[106] & in2[106];
    assign P[84] = in[106] ^ in2[106];
    assign G[85] = in[105] & in2[105];
    assign P[85] = in[105] ^ in2[105];
    assign G[86] = in[104] & in2[104];
    assign P[86] = in[104] ^ in2[104];
    assign G[87] = in[103] & in2[103];
    assign P[87] = in[103] ^ in2[103];
    assign G[88] = in[102] & in2[102];
    assign P[88] = in[102] ^ in2[102];
    assign G[89] = in[101] & in2[101];
    assign P[89] = in[101] ^ in2[101];
    assign G[90] = in[100] & in2[100];
    assign P[90] = in[100] ^ in2[100];
    assign G[91] = in[99] & in2[99];
    assign P[91] = in[99] ^ in2[99];
    assign G[92] = in[98] & in2[98];
    assign P[92] = in[98] ^ in2[98];
    assign G[93] = in[97] & in2[97];
    assign P[93] = in[97] ^ in2[97];
    assign G[94] = in[96] & in2[96];
    assign P[94] = in[96] ^ in2[96];
    assign G[95] = in[95] & in2[95];
    assign P[95] = in[95] ^ in2[95];
    assign G[96] = in[94] & in2[94];
    assign P[96] = in[94] ^ in2[94];
    assign G[97] = in[93] & in2[93];
    assign P[97] = in[93] ^ in2[93];
    assign G[98] = in[92] & in2[92];
    assign P[98] = in[92] ^ in2[92];
    assign G[99] = in[91] & in2[91];
    assign P[99] = in[91] ^ in2[91];
    assign G[100] = in[90] & in2[90];
    assign P[100] = in[90] ^ in2[90];
    assign G[101] = in[89] & in2[89];
    assign P[101] = in[89] ^ in2[89];
    assign G[102] = in[88] & in2[88];
    assign P[102] = in[88] ^ in2[88];
    assign G[103] = in[87] & in2[87];
    assign P[103] = in[87] ^ in2[87];
    assign G[104] = in[86] & in2[86];
    assign P[104] = in[86] ^ in2[86];
    assign G[105] = in[85] & in2[85];
    assign P[105] = in[85] ^ in2[85];
    assign G[106] = in[84] & in2[84];
    assign P[106] = in[84] ^ in2[84];
    assign G[107] = in[83] & in2[83];
    assign P[107] = in[83] ^ in2[83];
    assign G[108] = in[82] & in2[82];
    assign P[108] = in[82] ^ in2[82];
    assign G[109] = in[81] & in2[81];
    assign P[109] = in[81] ^ in2[81];
    assign G[110] = in[80] & in2[80];
    assign P[110] = in[80] ^ in2[80];
    assign G[111] = in[79] & in2[79];
    assign P[111] = in[79] ^ in2[79];
    assign G[112] = in[78] & in2[78];
    assign P[112] = in[78] ^ in2[78];
    assign G[113] = in[77] & in2[77];
    assign P[113] = in[77] ^ in2[77];
    assign G[114] = in[76] & in2[76];
    assign P[114] = in[76] ^ in2[76];
    assign G[115] = in[75] & in2[75];
    assign P[115] = in[75] ^ in2[75];
    assign G[116] = in[74] & in2[74];
    assign P[116] = in[74] ^ in2[74];
    assign G[117] = in[73] & in2[73];
    assign P[117] = in[73] ^ in2[73];
    assign G[118] = in[72] & in2[72];
    assign P[118] = in[72] ^ in2[72];
    assign G[119] = in[71] & in2[71];
    assign P[119] = in[71] ^ in2[71];
    assign G[120] = in[70] & in2[70];
    assign P[120] = in[70] ^ in2[70];
    assign G[121] = in[69] & in2[69];
    assign P[121] = in[69] ^ in2[69];
    assign G[122] = in[68] & in2[68];
    assign P[122] = in[68] ^ in2[68];
    assign G[123] = in[67] & in2[67];
    assign P[123] = in[67] ^ in2[67];
    assign G[124] = in[66] & in2[66];
    assign P[124] = in[66] ^ in2[66];
    assign G[125] = in[65] & in2[65];
    assign P[125] = in[65] ^ in2[65];
    assign G[126] = in[64] & in2[64];
    assign P[126] = in[64] ^ in2[64];
    assign G[127] = in[63] & in2[63];
    assign P[127] = in[63] ^ in2[63];
    assign G[128] = in[62] & in2[62];
    assign P[128] = in[62] ^ in2[62];
    assign G[129] = in[61] & in2[61];
    assign P[129] = in[61] ^ in2[61];
    assign G[130] = in[60] & in2[60];
    assign P[130] = in[60] ^ in2[60];
    assign G[131] = in[59] & in2[59];
    assign P[131] = in[59] ^ in2[59];
    assign G[132] = in[58] & in2[58];
    assign P[132] = in[58] ^ in2[58];
    assign G[133] = in[57] & in2[57];
    assign P[133] = in[57] ^ in2[57];
    assign G[134] = in[56] & in2[56];
    assign P[134] = in[56] ^ in2[56];
    assign G[135] = in[55] & in2[55];
    assign P[135] = in[55] ^ in2[55];
    assign G[136] = in[54] & in2[54];
    assign P[136] = in[54] ^ in2[54];
    assign G[137] = in[53] & in2[53];
    assign P[137] = in[53] ^ in2[53];
    assign G[138] = in[52] & in2[52];
    assign P[138] = in[52] ^ in2[52];
    assign G[139] = in[51] & in2[51];
    assign P[139] = in[51] ^ in2[51];
    assign G[140] = in[50] & in2[50];
    assign P[140] = in[50] ^ in2[50];
    assign G[141] = in[49] & in2[49];
    assign P[141] = in[49] ^ in2[49];
    assign G[142] = in[48] & in2[48];
    assign P[142] = in[48] ^ in2[48];
    assign G[143] = in[47] & in2[47];
    assign P[143] = in[47] ^ in2[47];
    assign G[144] = in[46] & in2[46];
    assign P[144] = in[46] ^ in2[46];
    assign G[145] = in[45] & in2[45];
    assign P[145] = in[45] ^ in2[45];
    assign G[146] = in[44] & in2[44];
    assign P[146] = in[44] ^ in2[44];
    assign G[147] = in[43] & in2[43];
    assign P[147] = in[43] ^ in2[43];
    assign G[148] = in[42] & in2[42];
    assign P[148] = in[42] ^ in2[42];
    assign G[149] = in[41] & in2[41];
    assign P[149] = in[41] ^ in2[41];
    assign G[150] = in[40] & in2[40];
    assign P[150] = in[40] ^ in2[40];
    assign G[151] = in[39] & in2[39];
    assign P[151] = in[39] ^ in2[39];
    assign G[152] = in[38] & in2[38];
    assign P[152] = in[38] ^ in2[38];
    assign G[153] = in[37] & in2[37];
    assign P[153] = in[37] ^ in2[37];
    assign G[154] = in[36] & in2[36];
    assign P[154] = in[36] ^ in2[36];
    assign G[155] = in[35] & in2[35];
    assign P[155] = in[35] ^ in2[35];
    assign G[156] = in[34] & in2[34];
    assign P[156] = in[34] ^ in2[34];
    assign G[157] = in[33] & in2[33];
    assign P[157] = in[33] ^ in2[33];
    assign G[158] = in[32] & in2[32];
    assign P[158] = in[32] ^ in2[32];
    assign G[159] = in[31] & in2[31];
    assign P[159] = in[31] ^ in2[31];
    assign G[160] = in[30] & in2[30];
    assign P[160] = in[30] ^ in2[30];
    assign G[161] = in[29] & in2[29];
    assign P[161] = in[29] ^ in2[29];
    assign G[162] = in[28] & in2[28];
    assign P[162] = in[28] ^ in2[28];
    assign G[163] = in[27] & in2[27];
    assign P[163] = in[27] ^ in2[27];
    assign G[164] = in[26] & in2[26];
    assign P[164] = in[26] ^ in2[26];
    assign G[165] = in[25] & in2[25];
    assign P[165] = in[25] ^ in2[25];
    assign G[166] = in[24] & in2[24];
    assign P[166] = in[24] ^ in2[24];
    assign G[167] = in[23] & in2[23];
    assign P[167] = in[23] ^ in2[23];
    assign G[168] = in[22] & in2[22];
    assign P[168] = in[22] ^ in2[22];
    assign G[169] = in[21] & in2[21];
    assign P[169] = in[21] ^ in2[21];
    assign G[170] = in[20] & in2[20];
    assign P[170] = in[20] ^ in2[20];
    assign G[171] = in[19] & in2[19];
    assign P[171] = in[19] ^ in2[19];
    assign G[172] = in[18] & in2[18];
    assign P[172] = in[18] ^ in2[18];
    assign G[173] = in[17] & in2[17];
    assign P[173] = in[17] ^ in2[17];
    assign G[174] = in[16] & in2[16];
    assign P[174] = in[16] ^ in2[16];
    assign G[175] = in[15] & in2[15];
    assign P[175] = in[15] ^ in2[15];
    assign G[176] = in[14] & in2[14];
    assign P[176] = in[14] ^ in2[14];
    assign G[177] = in[13] & in2[13];
    assign P[177] = in[13] ^ in2[13];
    assign G[178] = in[12] & in2[12];
    assign P[178] = in[12] ^ in2[12];
    assign G[179] = in[11] & in2[11];
    assign P[179] = in[11] ^ in2[11];
    assign G[180] = in[10] & in2[10];
    assign P[180] = in[10] ^ in2[10];
    assign G[181] = in[9] & in2[9];
    assign P[181] = in[9] ^ in2[9];
    assign G[182] = in[8] & in2[8];
    assign P[182] = in[8] ^ in2[8];
    assign G[183] = in[7] & in2[7];
    assign P[183] = in[7] ^ in2[7];
    assign G[184] = in[6] & in2[6];
    assign P[184] = in[6] ^ in2[6];
    assign G[185] = in[5] & in2[5];
    assign P[185] = in[5] ^ in2[5];
    assign G[186] = in[4] & in2[4];
    assign P[186] = in[4] ^ in2[4];
    assign G[187] = in[3] & in2[3];
    assign P[187] = in[3] ^ in2[3];
    assign G[188] = in[2] & in2[2];
    assign P[188] = in[2] ^ in2[2];
    assign G[189] = in[1] & in2[1];
    assign P[189] = in[1] ^ in2[1];
    assign G[190] = in[0] & in2[0];
    assign P[190] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign C[190] = G[189] | (P[189] & C[189]);
    assign cout = G[190] | (P[190] & C[190]);
    assign sum = P ^ C;
endmodule

module CLA190(output [189:0] sum, output cout, input [189:0] in1, input [189:0] in2;

    wire[189:0] G;
    wire[189:0] C;
    wire[189:0] P;

    assign G[0] = in[189] & in2[189];
    assign P[0] = in[189] ^ in2[189];
    assign G[1] = in[188] & in2[188];
    assign P[1] = in[188] ^ in2[188];
    assign G[2] = in[187] & in2[187];
    assign P[2] = in[187] ^ in2[187];
    assign G[3] = in[186] & in2[186];
    assign P[3] = in[186] ^ in2[186];
    assign G[4] = in[185] & in2[185];
    assign P[4] = in[185] ^ in2[185];
    assign G[5] = in[184] & in2[184];
    assign P[5] = in[184] ^ in2[184];
    assign G[6] = in[183] & in2[183];
    assign P[6] = in[183] ^ in2[183];
    assign G[7] = in[182] & in2[182];
    assign P[7] = in[182] ^ in2[182];
    assign G[8] = in[181] & in2[181];
    assign P[8] = in[181] ^ in2[181];
    assign G[9] = in[180] & in2[180];
    assign P[9] = in[180] ^ in2[180];
    assign G[10] = in[179] & in2[179];
    assign P[10] = in[179] ^ in2[179];
    assign G[11] = in[178] & in2[178];
    assign P[11] = in[178] ^ in2[178];
    assign G[12] = in[177] & in2[177];
    assign P[12] = in[177] ^ in2[177];
    assign G[13] = in[176] & in2[176];
    assign P[13] = in[176] ^ in2[176];
    assign G[14] = in[175] & in2[175];
    assign P[14] = in[175] ^ in2[175];
    assign G[15] = in[174] & in2[174];
    assign P[15] = in[174] ^ in2[174];
    assign G[16] = in[173] & in2[173];
    assign P[16] = in[173] ^ in2[173];
    assign G[17] = in[172] & in2[172];
    assign P[17] = in[172] ^ in2[172];
    assign G[18] = in[171] & in2[171];
    assign P[18] = in[171] ^ in2[171];
    assign G[19] = in[170] & in2[170];
    assign P[19] = in[170] ^ in2[170];
    assign G[20] = in[169] & in2[169];
    assign P[20] = in[169] ^ in2[169];
    assign G[21] = in[168] & in2[168];
    assign P[21] = in[168] ^ in2[168];
    assign G[22] = in[167] & in2[167];
    assign P[22] = in[167] ^ in2[167];
    assign G[23] = in[166] & in2[166];
    assign P[23] = in[166] ^ in2[166];
    assign G[24] = in[165] & in2[165];
    assign P[24] = in[165] ^ in2[165];
    assign G[25] = in[164] & in2[164];
    assign P[25] = in[164] ^ in2[164];
    assign G[26] = in[163] & in2[163];
    assign P[26] = in[163] ^ in2[163];
    assign G[27] = in[162] & in2[162];
    assign P[27] = in[162] ^ in2[162];
    assign G[28] = in[161] & in2[161];
    assign P[28] = in[161] ^ in2[161];
    assign G[29] = in[160] & in2[160];
    assign P[29] = in[160] ^ in2[160];
    assign G[30] = in[159] & in2[159];
    assign P[30] = in[159] ^ in2[159];
    assign G[31] = in[158] & in2[158];
    assign P[31] = in[158] ^ in2[158];
    assign G[32] = in[157] & in2[157];
    assign P[32] = in[157] ^ in2[157];
    assign G[33] = in[156] & in2[156];
    assign P[33] = in[156] ^ in2[156];
    assign G[34] = in[155] & in2[155];
    assign P[34] = in[155] ^ in2[155];
    assign G[35] = in[154] & in2[154];
    assign P[35] = in[154] ^ in2[154];
    assign G[36] = in[153] & in2[153];
    assign P[36] = in[153] ^ in2[153];
    assign G[37] = in[152] & in2[152];
    assign P[37] = in[152] ^ in2[152];
    assign G[38] = in[151] & in2[151];
    assign P[38] = in[151] ^ in2[151];
    assign G[39] = in[150] & in2[150];
    assign P[39] = in[150] ^ in2[150];
    assign G[40] = in[149] & in2[149];
    assign P[40] = in[149] ^ in2[149];
    assign G[41] = in[148] & in2[148];
    assign P[41] = in[148] ^ in2[148];
    assign G[42] = in[147] & in2[147];
    assign P[42] = in[147] ^ in2[147];
    assign G[43] = in[146] & in2[146];
    assign P[43] = in[146] ^ in2[146];
    assign G[44] = in[145] & in2[145];
    assign P[44] = in[145] ^ in2[145];
    assign G[45] = in[144] & in2[144];
    assign P[45] = in[144] ^ in2[144];
    assign G[46] = in[143] & in2[143];
    assign P[46] = in[143] ^ in2[143];
    assign G[47] = in[142] & in2[142];
    assign P[47] = in[142] ^ in2[142];
    assign G[48] = in[141] & in2[141];
    assign P[48] = in[141] ^ in2[141];
    assign G[49] = in[140] & in2[140];
    assign P[49] = in[140] ^ in2[140];
    assign G[50] = in[139] & in2[139];
    assign P[50] = in[139] ^ in2[139];
    assign G[51] = in[138] & in2[138];
    assign P[51] = in[138] ^ in2[138];
    assign G[52] = in[137] & in2[137];
    assign P[52] = in[137] ^ in2[137];
    assign G[53] = in[136] & in2[136];
    assign P[53] = in[136] ^ in2[136];
    assign G[54] = in[135] & in2[135];
    assign P[54] = in[135] ^ in2[135];
    assign G[55] = in[134] & in2[134];
    assign P[55] = in[134] ^ in2[134];
    assign G[56] = in[133] & in2[133];
    assign P[56] = in[133] ^ in2[133];
    assign G[57] = in[132] & in2[132];
    assign P[57] = in[132] ^ in2[132];
    assign G[58] = in[131] & in2[131];
    assign P[58] = in[131] ^ in2[131];
    assign G[59] = in[130] & in2[130];
    assign P[59] = in[130] ^ in2[130];
    assign G[60] = in[129] & in2[129];
    assign P[60] = in[129] ^ in2[129];
    assign G[61] = in[128] & in2[128];
    assign P[61] = in[128] ^ in2[128];
    assign G[62] = in[127] & in2[127];
    assign P[62] = in[127] ^ in2[127];
    assign G[63] = in[126] & in2[126];
    assign P[63] = in[126] ^ in2[126];
    assign G[64] = in[125] & in2[125];
    assign P[64] = in[125] ^ in2[125];
    assign G[65] = in[124] & in2[124];
    assign P[65] = in[124] ^ in2[124];
    assign G[66] = in[123] & in2[123];
    assign P[66] = in[123] ^ in2[123];
    assign G[67] = in[122] & in2[122];
    assign P[67] = in[122] ^ in2[122];
    assign G[68] = in[121] & in2[121];
    assign P[68] = in[121] ^ in2[121];
    assign G[69] = in[120] & in2[120];
    assign P[69] = in[120] ^ in2[120];
    assign G[70] = in[119] & in2[119];
    assign P[70] = in[119] ^ in2[119];
    assign G[71] = in[118] & in2[118];
    assign P[71] = in[118] ^ in2[118];
    assign G[72] = in[117] & in2[117];
    assign P[72] = in[117] ^ in2[117];
    assign G[73] = in[116] & in2[116];
    assign P[73] = in[116] ^ in2[116];
    assign G[74] = in[115] & in2[115];
    assign P[74] = in[115] ^ in2[115];
    assign G[75] = in[114] & in2[114];
    assign P[75] = in[114] ^ in2[114];
    assign G[76] = in[113] & in2[113];
    assign P[76] = in[113] ^ in2[113];
    assign G[77] = in[112] & in2[112];
    assign P[77] = in[112] ^ in2[112];
    assign G[78] = in[111] & in2[111];
    assign P[78] = in[111] ^ in2[111];
    assign G[79] = in[110] & in2[110];
    assign P[79] = in[110] ^ in2[110];
    assign G[80] = in[109] & in2[109];
    assign P[80] = in[109] ^ in2[109];
    assign G[81] = in[108] & in2[108];
    assign P[81] = in[108] ^ in2[108];
    assign G[82] = in[107] & in2[107];
    assign P[82] = in[107] ^ in2[107];
    assign G[83] = in[106] & in2[106];
    assign P[83] = in[106] ^ in2[106];
    assign G[84] = in[105] & in2[105];
    assign P[84] = in[105] ^ in2[105];
    assign G[85] = in[104] & in2[104];
    assign P[85] = in[104] ^ in2[104];
    assign G[86] = in[103] & in2[103];
    assign P[86] = in[103] ^ in2[103];
    assign G[87] = in[102] & in2[102];
    assign P[87] = in[102] ^ in2[102];
    assign G[88] = in[101] & in2[101];
    assign P[88] = in[101] ^ in2[101];
    assign G[89] = in[100] & in2[100];
    assign P[89] = in[100] ^ in2[100];
    assign G[90] = in[99] & in2[99];
    assign P[90] = in[99] ^ in2[99];
    assign G[91] = in[98] & in2[98];
    assign P[91] = in[98] ^ in2[98];
    assign G[92] = in[97] & in2[97];
    assign P[92] = in[97] ^ in2[97];
    assign G[93] = in[96] & in2[96];
    assign P[93] = in[96] ^ in2[96];
    assign G[94] = in[95] & in2[95];
    assign P[94] = in[95] ^ in2[95];
    assign G[95] = in[94] & in2[94];
    assign P[95] = in[94] ^ in2[94];
    assign G[96] = in[93] & in2[93];
    assign P[96] = in[93] ^ in2[93];
    assign G[97] = in[92] & in2[92];
    assign P[97] = in[92] ^ in2[92];
    assign G[98] = in[91] & in2[91];
    assign P[98] = in[91] ^ in2[91];
    assign G[99] = in[90] & in2[90];
    assign P[99] = in[90] ^ in2[90];
    assign G[100] = in[89] & in2[89];
    assign P[100] = in[89] ^ in2[89];
    assign G[101] = in[88] & in2[88];
    assign P[101] = in[88] ^ in2[88];
    assign G[102] = in[87] & in2[87];
    assign P[102] = in[87] ^ in2[87];
    assign G[103] = in[86] & in2[86];
    assign P[103] = in[86] ^ in2[86];
    assign G[104] = in[85] & in2[85];
    assign P[104] = in[85] ^ in2[85];
    assign G[105] = in[84] & in2[84];
    assign P[105] = in[84] ^ in2[84];
    assign G[106] = in[83] & in2[83];
    assign P[106] = in[83] ^ in2[83];
    assign G[107] = in[82] & in2[82];
    assign P[107] = in[82] ^ in2[82];
    assign G[108] = in[81] & in2[81];
    assign P[108] = in[81] ^ in2[81];
    assign G[109] = in[80] & in2[80];
    assign P[109] = in[80] ^ in2[80];
    assign G[110] = in[79] & in2[79];
    assign P[110] = in[79] ^ in2[79];
    assign G[111] = in[78] & in2[78];
    assign P[111] = in[78] ^ in2[78];
    assign G[112] = in[77] & in2[77];
    assign P[112] = in[77] ^ in2[77];
    assign G[113] = in[76] & in2[76];
    assign P[113] = in[76] ^ in2[76];
    assign G[114] = in[75] & in2[75];
    assign P[114] = in[75] ^ in2[75];
    assign G[115] = in[74] & in2[74];
    assign P[115] = in[74] ^ in2[74];
    assign G[116] = in[73] & in2[73];
    assign P[116] = in[73] ^ in2[73];
    assign G[117] = in[72] & in2[72];
    assign P[117] = in[72] ^ in2[72];
    assign G[118] = in[71] & in2[71];
    assign P[118] = in[71] ^ in2[71];
    assign G[119] = in[70] & in2[70];
    assign P[119] = in[70] ^ in2[70];
    assign G[120] = in[69] & in2[69];
    assign P[120] = in[69] ^ in2[69];
    assign G[121] = in[68] & in2[68];
    assign P[121] = in[68] ^ in2[68];
    assign G[122] = in[67] & in2[67];
    assign P[122] = in[67] ^ in2[67];
    assign G[123] = in[66] & in2[66];
    assign P[123] = in[66] ^ in2[66];
    assign G[124] = in[65] & in2[65];
    assign P[124] = in[65] ^ in2[65];
    assign G[125] = in[64] & in2[64];
    assign P[125] = in[64] ^ in2[64];
    assign G[126] = in[63] & in2[63];
    assign P[126] = in[63] ^ in2[63];
    assign G[127] = in[62] & in2[62];
    assign P[127] = in[62] ^ in2[62];
    assign G[128] = in[61] & in2[61];
    assign P[128] = in[61] ^ in2[61];
    assign G[129] = in[60] & in2[60];
    assign P[129] = in[60] ^ in2[60];
    assign G[130] = in[59] & in2[59];
    assign P[130] = in[59] ^ in2[59];
    assign G[131] = in[58] & in2[58];
    assign P[131] = in[58] ^ in2[58];
    assign G[132] = in[57] & in2[57];
    assign P[132] = in[57] ^ in2[57];
    assign G[133] = in[56] & in2[56];
    assign P[133] = in[56] ^ in2[56];
    assign G[134] = in[55] & in2[55];
    assign P[134] = in[55] ^ in2[55];
    assign G[135] = in[54] & in2[54];
    assign P[135] = in[54] ^ in2[54];
    assign G[136] = in[53] & in2[53];
    assign P[136] = in[53] ^ in2[53];
    assign G[137] = in[52] & in2[52];
    assign P[137] = in[52] ^ in2[52];
    assign G[138] = in[51] & in2[51];
    assign P[138] = in[51] ^ in2[51];
    assign G[139] = in[50] & in2[50];
    assign P[139] = in[50] ^ in2[50];
    assign G[140] = in[49] & in2[49];
    assign P[140] = in[49] ^ in2[49];
    assign G[141] = in[48] & in2[48];
    assign P[141] = in[48] ^ in2[48];
    assign G[142] = in[47] & in2[47];
    assign P[142] = in[47] ^ in2[47];
    assign G[143] = in[46] & in2[46];
    assign P[143] = in[46] ^ in2[46];
    assign G[144] = in[45] & in2[45];
    assign P[144] = in[45] ^ in2[45];
    assign G[145] = in[44] & in2[44];
    assign P[145] = in[44] ^ in2[44];
    assign G[146] = in[43] & in2[43];
    assign P[146] = in[43] ^ in2[43];
    assign G[147] = in[42] & in2[42];
    assign P[147] = in[42] ^ in2[42];
    assign G[148] = in[41] & in2[41];
    assign P[148] = in[41] ^ in2[41];
    assign G[149] = in[40] & in2[40];
    assign P[149] = in[40] ^ in2[40];
    assign G[150] = in[39] & in2[39];
    assign P[150] = in[39] ^ in2[39];
    assign G[151] = in[38] & in2[38];
    assign P[151] = in[38] ^ in2[38];
    assign G[152] = in[37] & in2[37];
    assign P[152] = in[37] ^ in2[37];
    assign G[153] = in[36] & in2[36];
    assign P[153] = in[36] ^ in2[36];
    assign G[154] = in[35] & in2[35];
    assign P[154] = in[35] ^ in2[35];
    assign G[155] = in[34] & in2[34];
    assign P[155] = in[34] ^ in2[34];
    assign G[156] = in[33] & in2[33];
    assign P[156] = in[33] ^ in2[33];
    assign G[157] = in[32] & in2[32];
    assign P[157] = in[32] ^ in2[32];
    assign G[158] = in[31] & in2[31];
    assign P[158] = in[31] ^ in2[31];
    assign G[159] = in[30] & in2[30];
    assign P[159] = in[30] ^ in2[30];
    assign G[160] = in[29] & in2[29];
    assign P[160] = in[29] ^ in2[29];
    assign G[161] = in[28] & in2[28];
    assign P[161] = in[28] ^ in2[28];
    assign G[162] = in[27] & in2[27];
    assign P[162] = in[27] ^ in2[27];
    assign G[163] = in[26] & in2[26];
    assign P[163] = in[26] ^ in2[26];
    assign G[164] = in[25] & in2[25];
    assign P[164] = in[25] ^ in2[25];
    assign G[165] = in[24] & in2[24];
    assign P[165] = in[24] ^ in2[24];
    assign G[166] = in[23] & in2[23];
    assign P[166] = in[23] ^ in2[23];
    assign G[167] = in[22] & in2[22];
    assign P[167] = in[22] ^ in2[22];
    assign G[168] = in[21] & in2[21];
    assign P[168] = in[21] ^ in2[21];
    assign G[169] = in[20] & in2[20];
    assign P[169] = in[20] ^ in2[20];
    assign G[170] = in[19] & in2[19];
    assign P[170] = in[19] ^ in2[19];
    assign G[171] = in[18] & in2[18];
    assign P[171] = in[18] ^ in2[18];
    assign G[172] = in[17] & in2[17];
    assign P[172] = in[17] ^ in2[17];
    assign G[173] = in[16] & in2[16];
    assign P[173] = in[16] ^ in2[16];
    assign G[174] = in[15] & in2[15];
    assign P[174] = in[15] ^ in2[15];
    assign G[175] = in[14] & in2[14];
    assign P[175] = in[14] ^ in2[14];
    assign G[176] = in[13] & in2[13];
    assign P[176] = in[13] ^ in2[13];
    assign G[177] = in[12] & in2[12];
    assign P[177] = in[12] ^ in2[12];
    assign G[178] = in[11] & in2[11];
    assign P[178] = in[11] ^ in2[11];
    assign G[179] = in[10] & in2[10];
    assign P[179] = in[10] ^ in2[10];
    assign G[180] = in[9] & in2[9];
    assign P[180] = in[9] ^ in2[9];
    assign G[181] = in[8] & in2[8];
    assign P[181] = in[8] ^ in2[8];
    assign G[182] = in[7] & in2[7];
    assign P[182] = in[7] ^ in2[7];
    assign G[183] = in[6] & in2[6];
    assign P[183] = in[6] ^ in2[6];
    assign G[184] = in[5] & in2[5];
    assign P[184] = in[5] ^ in2[5];
    assign G[185] = in[4] & in2[4];
    assign P[185] = in[4] ^ in2[4];
    assign G[186] = in[3] & in2[3];
    assign P[186] = in[3] ^ in2[3];
    assign G[187] = in[2] & in2[2];
    assign P[187] = in[2] ^ in2[2];
    assign G[188] = in[1] & in2[1];
    assign P[188] = in[1] ^ in2[1];
    assign G[189] = in[0] & in2[0];
    assign P[189] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign C[189] = G[188] | (P[188] & C[188]);
    assign cout = G[189] | (P[189] & C[189]);
    assign sum = P ^ C;
endmodule

module CLA189(output [188:0] sum, output cout, input [188:0] in1, input [188:0] in2;

    wire[188:0] G;
    wire[188:0] C;
    wire[188:0] P;

    assign G[0] = in[188] & in2[188];
    assign P[0] = in[188] ^ in2[188];
    assign G[1] = in[187] & in2[187];
    assign P[1] = in[187] ^ in2[187];
    assign G[2] = in[186] & in2[186];
    assign P[2] = in[186] ^ in2[186];
    assign G[3] = in[185] & in2[185];
    assign P[3] = in[185] ^ in2[185];
    assign G[4] = in[184] & in2[184];
    assign P[4] = in[184] ^ in2[184];
    assign G[5] = in[183] & in2[183];
    assign P[5] = in[183] ^ in2[183];
    assign G[6] = in[182] & in2[182];
    assign P[6] = in[182] ^ in2[182];
    assign G[7] = in[181] & in2[181];
    assign P[7] = in[181] ^ in2[181];
    assign G[8] = in[180] & in2[180];
    assign P[8] = in[180] ^ in2[180];
    assign G[9] = in[179] & in2[179];
    assign P[9] = in[179] ^ in2[179];
    assign G[10] = in[178] & in2[178];
    assign P[10] = in[178] ^ in2[178];
    assign G[11] = in[177] & in2[177];
    assign P[11] = in[177] ^ in2[177];
    assign G[12] = in[176] & in2[176];
    assign P[12] = in[176] ^ in2[176];
    assign G[13] = in[175] & in2[175];
    assign P[13] = in[175] ^ in2[175];
    assign G[14] = in[174] & in2[174];
    assign P[14] = in[174] ^ in2[174];
    assign G[15] = in[173] & in2[173];
    assign P[15] = in[173] ^ in2[173];
    assign G[16] = in[172] & in2[172];
    assign P[16] = in[172] ^ in2[172];
    assign G[17] = in[171] & in2[171];
    assign P[17] = in[171] ^ in2[171];
    assign G[18] = in[170] & in2[170];
    assign P[18] = in[170] ^ in2[170];
    assign G[19] = in[169] & in2[169];
    assign P[19] = in[169] ^ in2[169];
    assign G[20] = in[168] & in2[168];
    assign P[20] = in[168] ^ in2[168];
    assign G[21] = in[167] & in2[167];
    assign P[21] = in[167] ^ in2[167];
    assign G[22] = in[166] & in2[166];
    assign P[22] = in[166] ^ in2[166];
    assign G[23] = in[165] & in2[165];
    assign P[23] = in[165] ^ in2[165];
    assign G[24] = in[164] & in2[164];
    assign P[24] = in[164] ^ in2[164];
    assign G[25] = in[163] & in2[163];
    assign P[25] = in[163] ^ in2[163];
    assign G[26] = in[162] & in2[162];
    assign P[26] = in[162] ^ in2[162];
    assign G[27] = in[161] & in2[161];
    assign P[27] = in[161] ^ in2[161];
    assign G[28] = in[160] & in2[160];
    assign P[28] = in[160] ^ in2[160];
    assign G[29] = in[159] & in2[159];
    assign P[29] = in[159] ^ in2[159];
    assign G[30] = in[158] & in2[158];
    assign P[30] = in[158] ^ in2[158];
    assign G[31] = in[157] & in2[157];
    assign P[31] = in[157] ^ in2[157];
    assign G[32] = in[156] & in2[156];
    assign P[32] = in[156] ^ in2[156];
    assign G[33] = in[155] & in2[155];
    assign P[33] = in[155] ^ in2[155];
    assign G[34] = in[154] & in2[154];
    assign P[34] = in[154] ^ in2[154];
    assign G[35] = in[153] & in2[153];
    assign P[35] = in[153] ^ in2[153];
    assign G[36] = in[152] & in2[152];
    assign P[36] = in[152] ^ in2[152];
    assign G[37] = in[151] & in2[151];
    assign P[37] = in[151] ^ in2[151];
    assign G[38] = in[150] & in2[150];
    assign P[38] = in[150] ^ in2[150];
    assign G[39] = in[149] & in2[149];
    assign P[39] = in[149] ^ in2[149];
    assign G[40] = in[148] & in2[148];
    assign P[40] = in[148] ^ in2[148];
    assign G[41] = in[147] & in2[147];
    assign P[41] = in[147] ^ in2[147];
    assign G[42] = in[146] & in2[146];
    assign P[42] = in[146] ^ in2[146];
    assign G[43] = in[145] & in2[145];
    assign P[43] = in[145] ^ in2[145];
    assign G[44] = in[144] & in2[144];
    assign P[44] = in[144] ^ in2[144];
    assign G[45] = in[143] & in2[143];
    assign P[45] = in[143] ^ in2[143];
    assign G[46] = in[142] & in2[142];
    assign P[46] = in[142] ^ in2[142];
    assign G[47] = in[141] & in2[141];
    assign P[47] = in[141] ^ in2[141];
    assign G[48] = in[140] & in2[140];
    assign P[48] = in[140] ^ in2[140];
    assign G[49] = in[139] & in2[139];
    assign P[49] = in[139] ^ in2[139];
    assign G[50] = in[138] & in2[138];
    assign P[50] = in[138] ^ in2[138];
    assign G[51] = in[137] & in2[137];
    assign P[51] = in[137] ^ in2[137];
    assign G[52] = in[136] & in2[136];
    assign P[52] = in[136] ^ in2[136];
    assign G[53] = in[135] & in2[135];
    assign P[53] = in[135] ^ in2[135];
    assign G[54] = in[134] & in2[134];
    assign P[54] = in[134] ^ in2[134];
    assign G[55] = in[133] & in2[133];
    assign P[55] = in[133] ^ in2[133];
    assign G[56] = in[132] & in2[132];
    assign P[56] = in[132] ^ in2[132];
    assign G[57] = in[131] & in2[131];
    assign P[57] = in[131] ^ in2[131];
    assign G[58] = in[130] & in2[130];
    assign P[58] = in[130] ^ in2[130];
    assign G[59] = in[129] & in2[129];
    assign P[59] = in[129] ^ in2[129];
    assign G[60] = in[128] & in2[128];
    assign P[60] = in[128] ^ in2[128];
    assign G[61] = in[127] & in2[127];
    assign P[61] = in[127] ^ in2[127];
    assign G[62] = in[126] & in2[126];
    assign P[62] = in[126] ^ in2[126];
    assign G[63] = in[125] & in2[125];
    assign P[63] = in[125] ^ in2[125];
    assign G[64] = in[124] & in2[124];
    assign P[64] = in[124] ^ in2[124];
    assign G[65] = in[123] & in2[123];
    assign P[65] = in[123] ^ in2[123];
    assign G[66] = in[122] & in2[122];
    assign P[66] = in[122] ^ in2[122];
    assign G[67] = in[121] & in2[121];
    assign P[67] = in[121] ^ in2[121];
    assign G[68] = in[120] & in2[120];
    assign P[68] = in[120] ^ in2[120];
    assign G[69] = in[119] & in2[119];
    assign P[69] = in[119] ^ in2[119];
    assign G[70] = in[118] & in2[118];
    assign P[70] = in[118] ^ in2[118];
    assign G[71] = in[117] & in2[117];
    assign P[71] = in[117] ^ in2[117];
    assign G[72] = in[116] & in2[116];
    assign P[72] = in[116] ^ in2[116];
    assign G[73] = in[115] & in2[115];
    assign P[73] = in[115] ^ in2[115];
    assign G[74] = in[114] & in2[114];
    assign P[74] = in[114] ^ in2[114];
    assign G[75] = in[113] & in2[113];
    assign P[75] = in[113] ^ in2[113];
    assign G[76] = in[112] & in2[112];
    assign P[76] = in[112] ^ in2[112];
    assign G[77] = in[111] & in2[111];
    assign P[77] = in[111] ^ in2[111];
    assign G[78] = in[110] & in2[110];
    assign P[78] = in[110] ^ in2[110];
    assign G[79] = in[109] & in2[109];
    assign P[79] = in[109] ^ in2[109];
    assign G[80] = in[108] & in2[108];
    assign P[80] = in[108] ^ in2[108];
    assign G[81] = in[107] & in2[107];
    assign P[81] = in[107] ^ in2[107];
    assign G[82] = in[106] & in2[106];
    assign P[82] = in[106] ^ in2[106];
    assign G[83] = in[105] & in2[105];
    assign P[83] = in[105] ^ in2[105];
    assign G[84] = in[104] & in2[104];
    assign P[84] = in[104] ^ in2[104];
    assign G[85] = in[103] & in2[103];
    assign P[85] = in[103] ^ in2[103];
    assign G[86] = in[102] & in2[102];
    assign P[86] = in[102] ^ in2[102];
    assign G[87] = in[101] & in2[101];
    assign P[87] = in[101] ^ in2[101];
    assign G[88] = in[100] & in2[100];
    assign P[88] = in[100] ^ in2[100];
    assign G[89] = in[99] & in2[99];
    assign P[89] = in[99] ^ in2[99];
    assign G[90] = in[98] & in2[98];
    assign P[90] = in[98] ^ in2[98];
    assign G[91] = in[97] & in2[97];
    assign P[91] = in[97] ^ in2[97];
    assign G[92] = in[96] & in2[96];
    assign P[92] = in[96] ^ in2[96];
    assign G[93] = in[95] & in2[95];
    assign P[93] = in[95] ^ in2[95];
    assign G[94] = in[94] & in2[94];
    assign P[94] = in[94] ^ in2[94];
    assign G[95] = in[93] & in2[93];
    assign P[95] = in[93] ^ in2[93];
    assign G[96] = in[92] & in2[92];
    assign P[96] = in[92] ^ in2[92];
    assign G[97] = in[91] & in2[91];
    assign P[97] = in[91] ^ in2[91];
    assign G[98] = in[90] & in2[90];
    assign P[98] = in[90] ^ in2[90];
    assign G[99] = in[89] & in2[89];
    assign P[99] = in[89] ^ in2[89];
    assign G[100] = in[88] & in2[88];
    assign P[100] = in[88] ^ in2[88];
    assign G[101] = in[87] & in2[87];
    assign P[101] = in[87] ^ in2[87];
    assign G[102] = in[86] & in2[86];
    assign P[102] = in[86] ^ in2[86];
    assign G[103] = in[85] & in2[85];
    assign P[103] = in[85] ^ in2[85];
    assign G[104] = in[84] & in2[84];
    assign P[104] = in[84] ^ in2[84];
    assign G[105] = in[83] & in2[83];
    assign P[105] = in[83] ^ in2[83];
    assign G[106] = in[82] & in2[82];
    assign P[106] = in[82] ^ in2[82];
    assign G[107] = in[81] & in2[81];
    assign P[107] = in[81] ^ in2[81];
    assign G[108] = in[80] & in2[80];
    assign P[108] = in[80] ^ in2[80];
    assign G[109] = in[79] & in2[79];
    assign P[109] = in[79] ^ in2[79];
    assign G[110] = in[78] & in2[78];
    assign P[110] = in[78] ^ in2[78];
    assign G[111] = in[77] & in2[77];
    assign P[111] = in[77] ^ in2[77];
    assign G[112] = in[76] & in2[76];
    assign P[112] = in[76] ^ in2[76];
    assign G[113] = in[75] & in2[75];
    assign P[113] = in[75] ^ in2[75];
    assign G[114] = in[74] & in2[74];
    assign P[114] = in[74] ^ in2[74];
    assign G[115] = in[73] & in2[73];
    assign P[115] = in[73] ^ in2[73];
    assign G[116] = in[72] & in2[72];
    assign P[116] = in[72] ^ in2[72];
    assign G[117] = in[71] & in2[71];
    assign P[117] = in[71] ^ in2[71];
    assign G[118] = in[70] & in2[70];
    assign P[118] = in[70] ^ in2[70];
    assign G[119] = in[69] & in2[69];
    assign P[119] = in[69] ^ in2[69];
    assign G[120] = in[68] & in2[68];
    assign P[120] = in[68] ^ in2[68];
    assign G[121] = in[67] & in2[67];
    assign P[121] = in[67] ^ in2[67];
    assign G[122] = in[66] & in2[66];
    assign P[122] = in[66] ^ in2[66];
    assign G[123] = in[65] & in2[65];
    assign P[123] = in[65] ^ in2[65];
    assign G[124] = in[64] & in2[64];
    assign P[124] = in[64] ^ in2[64];
    assign G[125] = in[63] & in2[63];
    assign P[125] = in[63] ^ in2[63];
    assign G[126] = in[62] & in2[62];
    assign P[126] = in[62] ^ in2[62];
    assign G[127] = in[61] & in2[61];
    assign P[127] = in[61] ^ in2[61];
    assign G[128] = in[60] & in2[60];
    assign P[128] = in[60] ^ in2[60];
    assign G[129] = in[59] & in2[59];
    assign P[129] = in[59] ^ in2[59];
    assign G[130] = in[58] & in2[58];
    assign P[130] = in[58] ^ in2[58];
    assign G[131] = in[57] & in2[57];
    assign P[131] = in[57] ^ in2[57];
    assign G[132] = in[56] & in2[56];
    assign P[132] = in[56] ^ in2[56];
    assign G[133] = in[55] & in2[55];
    assign P[133] = in[55] ^ in2[55];
    assign G[134] = in[54] & in2[54];
    assign P[134] = in[54] ^ in2[54];
    assign G[135] = in[53] & in2[53];
    assign P[135] = in[53] ^ in2[53];
    assign G[136] = in[52] & in2[52];
    assign P[136] = in[52] ^ in2[52];
    assign G[137] = in[51] & in2[51];
    assign P[137] = in[51] ^ in2[51];
    assign G[138] = in[50] & in2[50];
    assign P[138] = in[50] ^ in2[50];
    assign G[139] = in[49] & in2[49];
    assign P[139] = in[49] ^ in2[49];
    assign G[140] = in[48] & in2[48];
    assign P[140] = in[48] ^ in2[48];
    assign G[141] = in[47] & in2[47];
    assign P[141] = in[47] ^ in2[47];
    assign G[142] = in[46] & in2[46];
    assign P[142] = in[46] ^ in2[46];
    assign G[143] = in[45] & in2[45];
    assign P[143] = in[45] ^ in2[45];
    assign G[144] = in[44] & in2[44];
    assign P[144] = in[44] ^ in2[44];
    assign G[145] = in[43] & in2[43];
    assign P[145] = in[43] ^ in2[43];
    assign G[146] = in[42] & in2[42];
    assign P[146] = in[42] ^ in2[42];
    assign G[147] = in[41] & in2[41];
    assign P[147] = in[41] ^ in2[41];
    assign G[148] = in[40] & in2[40];
    assign P[148] = in[40] ^ in2[40];
    assign G[149] = in[39] & in2[39];
    assign P[149] = in[39] ^ in2[39];
    assign G[150] = in[38] & in2[38];
    assign P[150] = in[38] ^ in2[38];
    assign G[151] = in[37] & in2[37];
    assign P[151] = in[37] ^ in2[37];
    assign G[152] = in[36] & in2[36];
    assign P[152] = in[36] ^ in2[36];
    assign G[153] = in[35] & in2[35];
    assign P[153] = in[35] ^ in2[35];
    assign G[154] = in[34] & in2[34];
    assign P[154] = in[34] ^ in2[34];
    assign G[155] = in[33] & in2[33];
    assign P[155] = in[33] ^ in2[33];
    assign G[156] = in[32] & in2[32];
    assign P[156] = in[32] ^ in2[32];
    assign G[157] = in[31] & in2[31];
    assign P[157] = in[31] ^ in2[31];
    assign G[158] = in[30] & in2[30];
    assign P[158] = in[30] ^ in2[30];
    assign G[159] = in[29] & in2[29];
    assign P[159] = in[29] ^ in2[29];
    assign G[160] = in[28] & in2[28];
    assign P[160] = in[28] ^ in2[28];
    assign G[161] = in[27] & in2[27];
    assign P[161] = in[27] ^ in2[27];
    assign G[162] = in[26] & in2[26];
    assign P[162] = in[26] ^ in2[26];
    assign G[163] = in[25] & in2[25];
    assign P[163] = in[25] ^ in2[25];
    assign G[164] = in[24] & in2[24];
    assign P[164] = in[24] ^ in2[24];
    assign G[165] = in[23] & in2[23];
    assign P[165] = in[23] ^ in2[23];
    assign G[166] = in[22] & in2[22];
    assign P[166] = in[22] ^ in2[22];
    assign G[167] = in[21] & in2[21];
    assign P[167] = in[21] ^ in2[21];
    assign G[168] = in[20] & in2[20];
    assign P[168] = in[20] ^ in2[20];
    assign G[169] = in[19] & in2[19];
    assign P[169] = in[19] ^ in2[19];
    assign G[170] = in[18] & in2[18];
    assign P[170] = in[18] ^ in2[18];
    assign G[171] = in[17] & in2[17];
    assign P[171] = in[17] ^ in2[17];
    assign G[172] = in[16] & in2[16];
    assign P[172] = in[16] ^ in2[16];
    assign G[173] = in[15] & in2[15];
    assign P[173] = in[15] ^ in2[15];
    assign G[174] = in[14] & in2[14];
    assign P[174] = in[14] ^ in2[14];
    assign G[175] = in[13] & in2[13];
    assign P[175] = in[13] ^ in2[13];
    assign G[176] = in[12] & in2[12];
    assign P[176] = in[12] ^ in2[12];
    assign G[177] = in[11] & in2[11];
    assign P[177] = in[11] ^ in2[11];
    assign G[178] = in[10] & in2[10];
    assign P[178] = in[10] ^ in2[10];
    assign G[179] = in[9] & in2[9];
    assign P[179] = in[9] ^ in2[9];
    assign G[180] = in[8] & in2[8];
    assign P[180] = in[8] ^ in2[8];
    assign G[181] = in[7] & in2[7];
    assign P[181] = in[7] ^ in2[7];
    assign G[182] = in[6] & in2[6];
    assign P[182] = in[6] ^ in2[6];
    assign G[183] = in[5] & in2[5];
    assign P[183] = in[5] ^ in2[5];
    assign G[184] = in[4] & in2[4];
    assign P[184] = in[4] ^ in2[4];
    assign G[185] = in[3] & in2[3];
    assign P[185] = in[3] ^ in2[3];
    assign G[186] = in[2] & in2[2];
    assign P[186] = in[2] ^ in2[2];
    assign G[187] = in[1] & in2[1];
    assign P[187] = in[1] ^ in2[1];
    assign G[188] = in[0] & in2[0];
    assign P[188] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign C[188] = G[187] | (P[187] & C[187]);
    assign cout = G[188] | (P[188] & C[188]);
    assign sum = P ^ C;
endmodule

module CLA188(output [187:0] sum, output cout, input [187:0] in1, input [187:0] in2;

    wire[187:0] G;
    wire[187:0] C;
    wire[187:0] P;

    assign G[0] = in[187] & in2[187];
    assign P[0] = in[187] ^ in2[187];
    assign G[1] = in[186] & in2[186];
    assign P[1] = in[186] ^ in2[186];
    assign G[2] = in[185] & in2[185];
    assign P[2] = in[185] ^ in2[185];
    assign G[3] = in[184] & in2[184];
    assign P[3] = in[184] ^ in2[184];
    assign G[4] = in[183] & in2[183];
    assign P[4] = in[183] ^ in2[183];
    assign G[5] = in[182] & in2[182];
    assign P[5] = in[182] ^ in2[182];
    assign G[6] = in[181] & in2[181];
    assign P[6] = in[181] ^ in2[181];
    assign G[7] = in[180] & in2[180];
    assign P[7] = in[180] ^ in2[180];
    assign G[8] = in[179] & in2[179];
    assign P[8] = in[179] ^ in2[179];
    assign G[9] = in[178] & in2[178];
    assign P[9] = in[178] ^ in2[178];
    assign G[10] = in[177] & in2[177];
    assign P[10] = in[177] ^ in2[177];
    assign G[11] = in[176] & in2[176];
    assign P[11] = in[176] ^ in2[176];
    assign G[12] = in[175] & in2[175];
    assign P[12] = in[175] ^ in2[175];
    assign G[13] = in[174] & in2[174];
    assign P[13] = in[174] ^ in2[174];
    assign G[14] = in[173] & in2[173];
    assign P[14] = in[173] ^ in2[173];
    assign G[15] = in[172] & in2[172];
    assign P[15] = in[172] ^ in2[172];
    assign G[16] = in[171] & in2[171];
    assign P[16] = in[171] ^ in2[171];
    assign G[17] = in[170] & in2[170];
    assign P[17] = in[170] ^ in2[170];
    assign G[18] = in[169] & in2[169];
    assign P[18] = in[169] ^ in2[169];
    assign G[19] = in[168] & in2[168];
    assign P[19] = in[168] ^ in2[168];
    assign G[20] = in[167] & in2[167];
    assign P[20] = in[167] ^ in2[167];
    assign G[21] = in[166] & in2[166];
    assign P[21] = in[166] ^ in2[166];
    assign G[22] = in[165] & in2[165];
    assign P[22] = in[165] ^ in2[165];
    assign G[23] = in[164] & in2[164];
    assign P[23] = in[164] ^ in2[164];
    assign G[24] = in[163] & in2[163];
    assign P[24] = in[163] ^ in2[163];
    assign G[25] = in[162] & in2[162];
    assign P[25] = in[162] ^ in2[162];
    assign G[26] = in[161] & in2[161];
    assign P[26] = in[161] ^ in2[161];
    assign G[27] = in[160] & in2[160];
    assign P[27] = in[160] ^ in2[160];
    assign G[28] = in[159] & in2[159];
    assign P[28] = in[159] ^ in2[159];
    assign G[29] = in[158] & in2[158];
    assign P[29] = in[158] ^ in2[158];
    assign G[30] = in[157] & in2[157];
    assign P[30] = in[157] ^ in2[157];
    assign G[31] = in[156] & in2[156];
    assign P[31] = in[156] ^ in2[156];
    assign G[32] = in[155] & in2[155];
    assign P[32] = in[155] ^ in2[155];
    assign G[33] = in[154] & in2[154];
    assign P[33] = in[154] ^ in2[154];
    assign G[34] = in[153] & in2[153];
    assign P[34] = in[153] ^ in2[153];
    assign G[35] = in[152] & in2[152];
    assign P[35] = in[152] ^ in2[152];
    assign G[36] = in[151] & in2[151];
    assign P[36] = in[151] ^ in2[151];
    assign G[37] = in[150] & in2[150];
    assign P[37] = in[150] ^ in2[150];
    assign G[38] = in[149] & in2[149];
    assign P[38] = in[149] ^ in2[149];
    assign G[39] = in[148] & in2[148];
    assign P[39] = in[148] ^ in2[148];
    assign G[40] = in[147] & in2[147];
    assign P[40] = in[147] ^ in2[147];
    assign G[41] = in[146] & in2[146];
    assign P[41] = in[146] ^ in2[146];
    assign G[42] = in[145] & in2[145];
    assign P[42] = in[145] ^ in2[145];
    assign G[43] = in[144] & in2[144];
    assign P[43] = in[144] ^ in2[144];
    assign G[44] = in[143] & in2[143];
    assign P[44] = in[143] ^ in2[143];
    assign G[45] = in[142] & in2[142];
    assign P[45] = in[142] ^ in2[142];
    assign G[46] = in[141] & in2[141];
    assign P[46] = in[141] ^ in2[141];
    assign G[47] = in[140] & in2[140];
    assign P[47] = in[140] ^ in2[140];
    assign G[48] = in[139] & in2[139];
    assign P[48] = in[139] ^ in2[139];
    assign G[49] = in[138] & in2[138];
    assign P[49] = in[138] ^ in2[138];
    assign G[50] = in[137] & in2[137];
    assign P[50] = in[137] ^ in2[137];
    assign G[51] = in[136] & in2[136];
    assign P[51] = in[136] ^ in2[136];
    assign G[52] = in[135] & in2[135];
    assign P[52] = in[135] ^ in2[135];
    assign G[53] = in[134] & in2[134];
    assign P[53] = in[134] ^ in2[134];
    assign G[54] = in[133] & in2[133];
    assign P[54] = in[133] ^ in2[133];
    assign G[55] = in[132] & in2[132];
    assign P[55] = in[132] ^ in2[132];
    assign G[56] = in[131] & in2[131];
    assign P[56] = in[131] ^ in2[131];
    assign G[57] = in[130] & in2[130];
    assign P[57] = in[130] ^ in2[130];
    assign G[58] = in[129] & in2[129];
    assign P[58] = in[129] ^ in2[129];
    assign G[59] = in[128] & in2[128];
    assign P[59] = in[128] ^ in2[128];
    assign G[60] = in[127] & in2[127];
    assign P[60] = in[127] ^ in2[127];
    assign G[61] = in[126] & in2[126];
    assign P[61] = in[126] ^ in2[126];
    assign G[62] = in[125] & in2[125];
    assign P[62] = in[125] ^ in2[125];
    assign G[63] = in[124] & in2[124];
    assign P[63] = in[124] ^ in2[124];
    assign G[64] = in[123] & in2[123];
    assign P[64] = in[123] ^ in2[123];
    assign G[65] = in[122] & in2[122];
    assign P[65] = in[122] ^ in2[122];
    assign G[66] = in[121] & in2[121];
    assign P[66] = in[121] ^ in2[121];
    assign G[67] = in[120] & in2[120];
    assign P[67] = in[120] ^ in2[120];
    assign G[68] = in[119] & in2[119];
    assign P[68] = in[119] ^ in2[119];
    assign G[69] = in[118] & in2[118];
    assign P[69] = in[118] ^ in2[118];
    assign G[70] = in[117] & in2[117];
    assign P[70] = in[117] ^ in2[117];
    assign G[71] = in[116] & in2[116];
    assign P[71] = in[116] ^ in2[116];
    assign G[72] = in[115] & in2[115];
    assign P[72] = in[115] ^ in2[115];
    assign G[73] = in[114] & in2[114];
    assign P[73] = in[114] ^ in2[114];
    assign G[74] = in[113] & in2[113];
    assign P[74] = in[113] ^ in2[113];
    assign G[75] = in[112] & in2[112];
    assign P[75] = in[112] ^ in2[112];
    assign G[76] = in[111] & in2[111];
    assign P[76] = in[111] ^ in2[111];
    assign G[77] = in[110] & in2[110];
    assign P[77] = in[110] ^ in2[110];
    assign G[78] = in[109] & in2[109];
    assign P[78] = in[109] ^ in2[109];
    assign G[79] = in[108] & in2[108];
    assign P[79] = in[108] ^ in2[108];
    assign G[80] = in[107] & in2[107];
    assign P[80] = in[107] ^ in2[107];
    assign G[81] = in[106] & in2[106];
    assign P[81] = in[106] ^ in2[106];
    assign G[82] = in[105] & in2[105];
    assign P[82] = in[105] ^ in2[105];
    assign G[83] = in[104] & in2[104];
    assign P[83] = in[104] ^ in2[104];
    assign G[84] = in[103] & in2[103];
    assign P[84] = in[103] ^ in2[103];
    assign G[85] = in[102] & in2[102];
    assign P[85] = in[102] ^ in2[102];
    assign G[86] = in[101] & in2[101];
    assign P[86] = in[101] ^ in2[101];
    assign G[87] = in[100] & in2[100];
    assign P[87] = in[100] ^ in2[100];
    assign G[88] = in[99] & in2[99];
    assign P[88] = in[99] ^ in2[99];
    assign G[89] = in[98] & in2[98];
    assign P[89] = in[98] ^ in2[98];
    assign G[90] = in[97] & in2[97];
    assign P[90] = in[97] ^ in2[97];
    assign G[91] = in[96] & in2[96];
    assign P[91] = in[96] ^ in2[96];
    assign G[92] = in[95] & in2[95];
    assign P[92] = in[95] ^ in2[95];
    assign G[93] = in[94] & in2[94];
    assign P[93] = in[94] ^ in2[94];
    assign G[94] = in[93] & in2[93];
    assign P[94] = in[93] ^ in2[93];
    assign G[95] = in[92] & in2[92];
    assign P[95] = in[92] ^ in2[92];
    assign G[96] = in[91] & in2[91];
    assign P[96] = in[91] ^ in2[91];
    assign G[97] = in[90] & in2[90];
    assign P[97] = in[90] ^ in2[90];
    assign G[98] = in[89] & in2[89];
    assign P[98] = in[89] ^ in2[89];
    assign G[99] = in[88] & in2[88];
    assign P[99] = in[88] ^ in2[88];
    assign G[100] = in[87] & in2[87];
    assign P[100] = in[87] ^ in2[87];
    assign G[101] = in[86] & in2[86];
    assign P[101] = in[86] ^ in2[86];
    assign G[102] = in[85] & in2[85];
    assign P[102] = in[85] ^ in2[85];
    assign G[103] = in[84] & in2[84];
    assign P[103] = in[84] ^ in2[84];
    assign G[104] = in[83] & in2[83];
    assign P[104] = in[83] ^ in2[83];
    assign G[105] = in[82] & in2[82];
    assign P[105] = in[82] ^ in2[82];
    assign G[106] = in[81] & in2[81];
    assign P[106] = in[81] ^ in2[81];
    assign G[107] = in[80] & in2[80];
    assign P[107] = in[80] ^ in2[80];
    assign G[108] = in[79] & in2[79];
    assign P[108] = in[79] ^ in2[79];
    assign G[109] = in[78] & in2[78];
    assign P[109] = in[78] ^ in2[78];
    assign G[110] = in[77] & in2[77];
    assign P[110] = in[77] ^ in2[77];
    assign G[111] = in[76] & in2[76];
    assign P[111] = in[76] ^ in2[76];
    assign G[112] = in[75] & in2[75];
    assign P[112] = in[75] ^ in2[75];
    assign G[113] = in[74] & in2[74];
    assign P[113] = in[74] ^ in2[74];
    assign G[114] = in[73] & in2[73];
    assign P[114] = in[73] ^ in2[73];
    assign G[115] = in[72] & in2[72];
    assign P[115] = in[72] ^ in2[72];
    assign G[116] = in[71] & in2[71];
    assign P[116] = in[71] ^ in2[71];
    assign G[117] = in[70] & in2[70];
    assign P[117] = in[70] ^ in2[70];
    assign G[118] = in[69] & in2[69];
    assign P[118] = in[69] ^ in2[69];
    assign G[119] = in[68] & in2[68];
    assign P[119] = in[68] ^ in2[68];
    assign G[120] = in[67] & in2[67];
    assign P[120] = in[67] ^ in2[67];
    assign G[121] = in[66] & in2[66];
    assign P[121] = in[66] ^ in2[66];
    assign G[122] = in[65] & in2[65];
    assign P[122] = in[65] ^ in2[65];
    assign G[123] = in[64] & in2[64];
    assign P[123] = in[64] ^ in2[64];
    assign G[124] = in[63] & in2[63];
    assign P[124] = in[63] ^ in2[63];
    assign G[125] = in[62] & in2[62];
    assign P[125] = in[62] ^ in2[62];
    assign G[126] = in[61] & in2[61];
    assign P[126] = in[61] ^ in2[61];
    assign G[127] = in[60] & in2[60];
    assign P[127] = in[60] ^ in2[60];
    assign G[128] = in[59] & in2[59];
    assign P[128] = in[59] ^ in2[59];
    assign G[129] = in[58] & in2[58];
    assign P[129] = in[58] ^ in2[58];
    assign G[130] = in[57] & in2[57];
    assign P[130] = in[57] ^ in2[57];
    assign G[131] = in[56] & in2[56];
    assign P[131] = in[56] ^ in2[56];
    assign G[132] = in[55] & in2[55];
    assign P[132] = in[55] ^ in2[55];
    assign G[133] = in[54] & in2[54];
    assign P[133] = in[54] ^ in2[54];
    assign G[134] = in[53] & in2[53];
    assign P[134] = in[53] ^ in2[53];
    assign G[135] = in[52] & in2[52];
    assign P[135] = in[52] ^ in2[52];
    assign G[136] = in[51] & in2[51];
    assign P[136] = in[51] ^ in2[51];
    assign G[137] = in[50] & in2[50];
    assign P[137] = in[50] ^ in2[50];
    assign G[138] = in[49] & in2[49];
    assign P[138] = in[49] ^ in2[49];
    assign G[139] = in[48] & in2[48];
    assign P[139] = in[48] ^ in2[48];
    assign G[140] = in[47] & in2[47];
    assign P[140] = in[47] ^ in2[47];
    assign G[141] = in[46] & in2[46];
    assign P[141] = in[46] ^ in2[46];
    assign G[142] = in[45] & in2[45];
    assign P[142] = in[45] ^ in2[45];
    assign G[143] = in[44] & in2[44];
    assign P[143] = in[44] ^ in2[44];
    assign G[144] = in[43] & in2[43];
    assign P[144] = in[43] ^ in2[43];
    assign G[145] = in[42] & in2[42];
    assign P[145] = in[42] ^ in2[42];
    assign G[146] = in[41] & in2[41];
    assign P[146] = in[41] ^ in2[41];
    assign G[147] = in[40] & in2[40];
    assign P[147] = in[40] ^ in2[40];
    assign G[148] = in[39] & in2[39];
    assign P[148] = in[39] ^ in2[39];
    assign G[149] = in[38] & in2[38];
    assign P[149] = in[38] ^ in2[38];
    assign G[150] = in[37] & in2[37];
    assign P[150] = in[37] ^ in2[37];
    assign G[151] = in[36] & in2[36];
    assign P[151] = in[36] ^ in2[36];
    assign G[152] = in[35] & in2[35];
    assign P[152] = in[35] ^ in2[35];
    assign G[153] = in[34] & in2[34];
    assign P[153] = in[34] ^ in2[34];
    assign G[154] = in[33] & in2[33];
    assign P[154] = in[33] ^ in2[33];
    assign G[155] = in[32] & in2[32];
    assign P[155] = in[32] ^ in2[32];
    assign G[156] = in[31] & in2[31];
    assign P[156] = in[31] ^ in2[31];
    assign G[157] = in[30] & in2[30];
    assign P[157] = in[30] ^ in2[30];
    assign G[158] = in[29] & in2[29];
    assign P[158] = in[29] ^ in2[29];
    assign G[159] = in[28] & in2[28];
    assign P[159] = in[28] ^ in2[28];
    assign G[160] = in[27] & in2[27];
    assign P[160] = in[27] ^ in2[27];
    assign G[161] = in[26] & in2[26];
    assign P[161] = in[26] ^ in2[26];
    assign G[162] = in[25] & in2[25];
    assign P[162] = in[25] ^ in2[25];
    assign G[163] = in[24] & in2[24];
    assign P[163] = in[24] ^ in2[24];
    assign G[164] = in[23] & in2[23];
    assign P[164] = in[23] ^ in2[23];
    assign G[165] = in[22] & in2[22];
    assign P[165] = in[22] ^ in2[22];
    assign G[166] = in[21] & in2[21];
    assign P[166] = in[21] ^ in2[21];
    assign G[167] = in[20] & in2[20];
    assign P[167] = in[20] ^ in2[20];
    assign G[168] = in[19] & in2[19];
    assign P[168] = in[19] ^ in2[19];
    assign G[169] = in[18] & in2[18];
    assign P[169] = in[18] ^ in2[18];
    assign G[170] = in[17] & in2[17];
    assign P[170] = in[17] ^ in2[17];
    assign G[171] = in[16] & in2[16];
    assign P[171] = in[16] ^ in2[16];
    assign G[172] = in[15] & in2[15];
    assign P[172] = in[15] ^ in2[15];
    assign G[173] = in[14] & in2[14];
    assign P[173] = in[14] ^ in2[14];
    assign G[174] = in[13] & in2[13];
    assign P[174] = in[13] ^ in2[13];
    assign G[175] = in[12] & in2[12];
    assign P[175] = in[12] ^ in2[12];
    assign G[176] = in[11] & in2[11];
    assign P[176] = in[11] ^ in2[11];
    assign G[177] = in[10] & in2[10];
    assign P[177] = in[10] ^ in2[10];
    assign G[178] = in[9] & in2[9];
    assign P[178] = in[9] ^ in2[9];
    assign G[179] = in[8] & in2[8];
    assign P[179] = in[8] ^ in2[8];
    assign G[180] = in[7] & in2[7];
    assign P[180] = in[7] ^ in2[7];
    assign G[181] = in[6] & in2[6];
    assign P[181] = in[6] ^ in2[6];
    assign G[182] = in[5] & in2[5];
    assign P[182] = in[5] ^ in2[5];
    assign G[183] = in[4] & in2[4];
    assign P[183] = in[4] ^ in2[4];
    assign G[184] = in[3] & in2[3];
    assign P[184] = in[3] ^ in2[3];
    assign G[185] = in[2] & in2[2];
    assign P[185] = in[2] ^ in2[2];
    assign G[186] = in[1] & in2[1];
    assign P[186] = in[1] ^ in2[1];
    assign G[187] = in[0] & in2[0];
    assign P[187] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign C[187] = G[186] | (P[186] & C[186]);
    assign cout = G[187] | (P[187] & C[187]);
    assign sum = P ^ C;
endmodule

module CLA187(output [186:0] sum, output cout, input [186:0] in1, input [186:0] in2;

    wire[186:0] G;
    wire[186:0] C;
    wire[186:0] P;

    assign G[0] = in[186] & in2[186];
    assign P[0] = in[186] ^ in2[186];
    assign G[1] = in[185] & in2[185];
    assign P[1] = in[185] ^ in2[185];
    assign G[2] = in[184] & in2[184];
    assign P[2] = in[184] ^ in2[184];
    assign G[3] = in[183] & in2[183];
    assign P[3] = in[183] ^ in2[183];
    assign G[4] = in[182] & in2[182];
    assign P[4] = in[182] ^ in2[182];
    assign G[5] = in[181] & in2[181];
    assign P[5] = in[181] ^ in2[181];
    assign G[6] = in[180] & in2[180];
    assign P[6] = in[180] ^ in2[180];
    assign G[7] = in[179] & in2[179];
    assign P[7] = in[179] ^ in2[179];
    assign G[8] = in[178] & in2[178];
    assign P[8] = in[178] ^ in2[178];
    assign G[9] = in[177] & in2[177];
    assign P[9] = in[177] ^ in2[177];
    assign G[10] = in[176] & in2[176];
    assign P[10] = in[176] ^ in2[176];
    assign G[11] = in[175] & in2[175];
    assign P[11] = in[175] ^ in2[175];
    assign G[12] = in[174] & in2[174];
    assign P[12] = in[174] ^ in2[174];
    assign G[13] = in[173] & in2[173];
    assign P[13] = in[173] ^ in2[173];
    assign G[14] = in[172] & in2[172];
    assign P[14] = in[172] ^ in2[172];
    assign G[15] = in[171] & in2[171];
    assign P[15] = in[171] ^ in2[171];
    assign G[16] = in[170] & in2[170];
    assign P[16] = in[170] ^ in2[170];
    assign G[17] = in[169] & in2[169];
    assign P[17] = in[169] ^ in2[169];
    assign G[18] = in[168] & in2[168];
    assign P[18] = in[168] ^ in2[168];
    assign G[19] = in[167] & in2[167];
    assign P[19] = in[167] ^ in2[167];
    assign G[20] = in[166] & in2[166];
    assign P[20] = in[166] ^ in2[166];
    assign G[21] = in[165] & in2[165];
    assign P[21] = in[165] ^ in2[165];
    assign G[22] = in[164] & in2[164];
    assign P[22] = in[164] ^ in2[164];
    assign G[23] = in[163] & in2[163];
    assign P[23] = in[163] ^ in2[163];
    assign G[24] = in[162] & in2[162];
    assign P[24] = in[162] ^ in2[162];
    assign G[25] = in[161] & in2[161];
    assign P[25] = in[161] ^ in2[161];
    assign G[26] = in[160] & in2[160];
    assign P[26] = in[160] ^ in2[160];
    assign G[27] = in[159] & in2[159];
    assign P[27] = in[159] ^ in2[159];
    assign G[28] = in[158] & in2[158];
    assign P[28] = in[158] ^ in2[158];
    assign G[29] = in[157] & in2[157];
    assign P[29] = in[157] ^ in2[157];
    assign G[30] = in[156] & in2[156];
    assign P[30] = in[156] ^ in2[156];
    assign G[31] = in[155] & in2[155];
    assign P[31] = in[155] ^ in2[155];
    assign G[32] = in[154] & in2[154];
    assign P[32] = in[154] ^ in2[154];
    assign G[33] = in[153] & in2[153];
    assign P[33] = in[153] ^ in2[153];
    assign G[34] = in[152] & in2[152];
    assign P[34] = in[152] ^ in2[152];
    assign G[35] = in[151] & in2[151];
    assign P[35] = in[151] ^ in2[151];
    assign G[36] = in[150] & in2[150];
    assign P[36] = in[150] ^ in2[150];
    assign G[37] = in[149] & in2[149];
    assign P[37] = in[149] ^ in2[149];
    assign G[38] = in[148] & in2[148];
    assign P[38] = in[148] ^ in2[148];
    assign G[39] = in[147] & in2[147];
    assign P[39] = in[147] ^ in2[147];
    assign G[40] = in[146] & in2[146];
    assign P[40] = in[146] ^ in2[146];
    assign G[41] = in[145] & in2[145];
    assign P[41] = in[145] ^ in2[145];
    assign G[42] = in[144] & in2[144];
    assign P[42] = in[144] ^ in2[144];
    assign G[43] = in[143] & in2[143];
    assign P[43] = in[143] ^ in2[143];
    assign G[44] = in[142] & in2[142];
    assign P[44] = in[142] ^ in2[142];
    assign G[45] = in[141] & in2[141];
    assign P[45] = in[141] ^ in2[141];
    assign G[46] = in[140] & in2[140];
    assign P[46] = in[140] ^ in2[140];
    assign G[47] = in[139] & in2[139];
    assign P[47] = in[139] ^ in2[139];
    assign G[48] = in[138] & in2[138];
    assign P[48] = in[138] ^ in2[138];
    assign G[49] = in[137] & in2[137];
    assign P[49] = in[137] ^ in2[137];
    assign G[50] = in[136] & in2[136];
    assign P[50] = in[136] ^ in2[136];
    assign G[51] = in[135] & in2[135];
    assign P[51] = in[135] ^ in2[135];
    assign G[52] = in[134] & in2[134];
    assign P[52] = in[134] ^ in2[134];
    assign G[53] = in[133] & in2[133];
    assign P[53] = in[133] ^ in2[133];
    assign G[54] = in[132] & in2[132];
    assign P[54] = in[132] ^ in2[132];
    assign G[55] = in[131] & in2[131];
    assign P[55] = in[131] ^ in2[131];
    assign G[56] = in[130] & in2[130];
    assign P[56] = in[130] ^ in2[130];
    assign G[57] = in[129] & in2[129];
    assign P[57] = in[129] ^ in2[129];
    assign G[58] = in[128] & in2[128];
    assign P[58] = in[128] ^ in2[128];
    assign G[59] = in[127] & in2[127];
    assign P[59] = in[127] ^ in2[127];
    assign G[60] = in[126] & in2[126];
    assign P[60] = in[126] ^ in2[126];
    assign G[61] = in[125] & in2[125];
    assign P[61] = in[125] ^ in2[125];
    assign G[62] = in[124] & in2[124];
    assign P[62] = in[124] ^ in2[124];
    assign G[63] = in[123] & in2[123];
    assign P[63] = in[123] ^ in2[123];
    assign G[64] = in[122] & in2[122];
    assign P[64] = in[122] ^ in2[122];
    assign G[65] = in[121] & in2[121];
    assign P[65] = in[121] ^ in2[121];
    assign G[66] = in[120] & in2[120];
    assign P[66] = in[120] ^ in2[120];
    assign G[67] = in[119] & in2[119];
    assign P[67] = in[119] ^ in2[119];
    assign G[68] = in[118] & in2[118];
    assign P[68] = in[118] ^ in2[118];
    assign G[69] = in[117] & in2[117];
    assign P[69] = in[117] ^ in2[117];
    assign G[70] = in[116] & in2[116];
    assign P[70] = in[116] ^ in2[116];
    assign G[71] = in[115] & in2[115];
    assign P[71] = in[115] ^ in2[115];
    assign G[72] = in[114] & in2[114];
    assign P[72] = in[114] ^ in2[114];
    assign G[73] = in[113] & in2[113];
    assign P[73] = in[113] ^ in2[113];
    assign G[74] = in[112] & in2[112];
    assign P[74] = in[112] ^ in2[112];
    assign G[75] = in[111] & in2[111];
    assign P[75] = in[111] ^ in2[111];
    assign G[76] = in[110] & in2[110];
    assign P[76] = in[110] ^ in2[110];
    assign G[77] = in[109] & in2[109];
    assign P[77] = in[109] ^ in2[109];
    assign G[78] = in[108] & in2[108];
    assign P[78] = in[108] ^ in2[108];
    assign G[79] = in[107] & in2[107];
    assign P[79] = in[107] ^ in2[107];
    assign G[80] = in[106] & in2[106];
    assign P[80] = in[106] ^ in2[106];
    assign G[81] = in[105] & in2[105];
    assign P[81] = in[105] ^ in2[105];
    assign G[82] = in[104] & in2[104];
    assign P[82] = in[104] ^ in2[104];
    assign G[83] = in[103] & in2[103];
    assign P[83] = in[103] ^ in2[103];
    assign G[84] = in[102] & in2[102];
    assign P[84] = in[102] ^ in2[102];
    assign G[85] = in[101] & in2[101];
    assign P[85] = in[101] ^ in2[101];
    assign G[86] = in[100] & in2[100];
    assign P[86] = in[100] ^ in2[100];
    assign G[87] = in[99] & in2[99];
    assign P[87] = in[99] ^ in2[99];
    assign G[88] = in[98] & in2[98];
    assign P[88] = in[98] ^ in2[98];
    assign G[89] = in[97] & in2[97];
    assign P[89] = in[97] ^ in2[97];
    assign G[90] = in[96] & in2[96];
    assign P[90] = in[96] ^ in2[96];
    assign G[91] = in[95] & in2[95];
    assign P[91] = in[95] ^ in2[95];
    assign G[92] = in[94] & in2[94];
    assign P[92] = in[94] ^ in2[94];
    assign G[93] = in[93] & in2[93];
    assign P[93] = in[93] ^ in2[93];
    assign G[94] = in[92] & in2[92];
    assign P[94] = in[92] ^ in2[92];
    assign G[95] = in[91] & in2[91];
    assign P[95] = in[91] ^ in2[91];
    assign G[96] = in[90] & in2[90];
    assign P[96] = in[90] ^ in2[90];
    assign G[97] = in[89] & in2[89];
    assign P[97] = in[89] ^ in2[89];
    assign G[98] = in[88] & in2[88];
    assign P[98] = in[88] ^ in2[88];
    assign G[99] = in[87] & in2[87];
    assign P[99] = in[87] ^ in2[87];
    assign G[100] = in[86] & in2[86];
    assign P[100] = in[86] ^ in2[86];
    assign G[101] = in[85] & in2[85];
    assign P[101] = in[85] ^ in2[85];
    assign G[102] = in[84] & in2[84];
    assign P[102] = in[84] ^ in2[84];
    assign G[103] = in[83] & in2[83];
    assign P[103] = in[83] ^ in2[83];
    assign G[104] = in[82] & in2[82];
    assign P[104] = in[82] ^ in2[82];
    assign G[105] = in[81] & in2[81];
    assign P[105] = in[81] ^ in2[81];
    assign G[106] = in[80] & in2[80];
    assign P[106] = in[80] ^ in2[80];
    assign G[107] = in[79] & in2[79];
    assign P[107] = in[79] ^ in2[79];
    assign G[108] = in[78] & in2[78];
    assign P[108] = in[78] ^ in2[78];
    assign G[109] = in[77] & in2[77];
    assign P[109] = in[77] ^ in2[77];
    assign G[110] = in[76] & in2[76];
    assign P[110] = in[76] ^ in2[76];
    assign G[111] = in[75] & in2[75];
    assign P[111] = in[75] ^ in2[75];
    assign G[112] = in[74] & in2[74];
    assign P[112] = in[74] ^ in2[74];
    assign G[113] = in[73] & in2[73];
    assign P[113] = in[73] ^ in2[73];
    assign G[114] = in[72] & in2[72];
    assign P[114] = in[72] ^ in2[72];
    assign G[115] = in[71] & in2[71];
    assign P[115] = in[71] ^ in2[71];
    assign G[116] = in[70] & in2[70];
    assign P[116] = in[70] ^ in2[70];
    assign G[117] = in[69] & in2[69];
    assign P[117] = in[69] ^ in2[69];
    assign G[118] = in[68] & in2[68];
    assign P[118] = in[68] ^ in2[68];
    assign G[119] = in[67] & in2[67];
    assign P[119] = in[67] ^ in2[67];
    assign G[120] = in[66] & in2[66];
    assign P[120] = in[66] ^ in2[66];
    assign G[121] = in[65] & in2[65];
    assign P[121] = in[65] ^ in2[65];
    assign G[122] = in[64] & in2[64];
    assign P[122] = in[64] ^ in2[64];
    assign G[123] = in[63] & in2[63];
    assign P[123] = in[63] ^ in2[63];
    assign G[124] = in[62] & in2[62];
    assign P[124] = in[62] ^ in2[62];
    assign G[125] = in[61] & in2[61];
    assign P[125] = in[61] ^ in2[61];
    assign G[126] = in[60] & in2[60];
    assign P[126] = in[60] ^ in2[60];
    assign G[127] = in[59] & in2[59];
    assign P[127] = in[59] ^ in2[59];
    assign G[128] = in[58] & in2[58];
    assign P[128] = in[58] ^ in2[58];
    assign G[129] = in[57] & in2[57];
    assign P[129] = in[57] ^ in2[57];
    assign G[130] = in[56] & in2[56];
    assign P[130] = in[56] ^ in2[56];
    assign G[131] = in[55] & in2[55];
    assign P[131] = in[55] ^ in2[55];
    assign G[132] = in[54] & in2[54];
    assign P[132] = in[54] ^ in2[54];
    assign G[133] = in[53] & in2[53];
    assign P[133] = in[53] ^ in2[53];
    assign G[134] = in[52] & in2[52];
    assign P[134] = in[52] ^ in2[52];
    assign G[135] = in[51] & in2[51];
    assign P[135] = in[51] ^ in2[51];
    assign G[136] = in[50] & in2[50];
    assign P[136] = in[50] ^ in2[50];
    assign G[137] = in[49] & in2[49];
    assign P[137] = in[49] ^ in2[49];
    assign G[138] = in[48] & in2[48];
    assign P[138] = in[48] ^ in2[48];
    assign G[139] = in[47] & in2[47];
    assign P[139] = in[47] ^ in2[47];
    assign G[140] = in[46] & in2[46];
    assign P[140] = in[46] ^ in2[46];
    assign G[141] = in[45] & in2[45];
    assign P[141] = in[45] ^ in2[45];
    assign G[142] = in[44] & in2[44];
    assign P[142] = in[44] ^ in2[44];
    assign G[143] = in[43] & in2[43];
    assign P[143] = in[43] ^ in2[43];
    assign G[144] = in[42] & in2[42];
    assign P[144] = in[42] ^ in2[42];
    assign G[145] = in[41] & in2[41];
    assign P[145] = in[41] ^ in2[41];
    assign G[146] = in[40] & in2[40];
    assign P[146] = in[40] ^ in2[40];
    assign G[147] = in[39] & in2[39];
    assign P[147] = in[39] ^ in2[39];
    assign G[148] = in[38] & in2[38];
    assign P[148] = in[38] ^ in2[38];
    assign G[149] = in[37] & in2[37];
    assign P[149] = in[37] ^ in2[37];
    assign G[150] = in[36] & in2[36];
    assign P[150] = in[36] ^ in2[36];
    assign G[151] = in[35] & in2[35];
    assign P[151] = in[35] ^ in2[35];
    assign G[152] = in[34] & in2[34];
    assign P[152] = in[34] ^ in2[34];
    assign G[153] = in[33] & in2[33];
    assign P[153] = in[33] ^ in2[33];
    assign G[154] = in[32] & in2[32];
    assign P[154] = in[32] ^ in2[32];
    assign G[155] = in[31] & in2[31];
    assign P[155] = in[31] ^ in2[31];
    assign G[156] = in[30] & in2[30];
    assign P[156] = in[30] ^ in2[30];
    assign G[157] = in[29] & in2[29];
    assign P[157] = in[29] ^ in2[29];
    assign G[158] = in[28] & in2[28];
    assign P[158] = in[28] ^ in2[28];
    assign G[159] = in[27] & in2[27];
    assign P[159] = in[27] ^ in2[27];
    assign G[160] = in[26] & in2[26];
    assign P[160] = in[26] ^ in2[26];
    assign G[161] = in[25] & in2[25];
    assign P[161] = in[25] ^ in2[25];
    assign G[162] = in[24] & in2[24];
    assign P[162] = in[24] ^ in2[24];
    assign G[163] = in[23] & in2[23];
    assign P[163] = in[23] ^ in2[23];
    assign G[164] = in[22] & in2[22];
    assign P[164] = in[22] ^ in2[22];
    assign G[165] = in[21] & in2[21];
    assign P[165] = in[21] ^ in2[21];
    assign G[166] = in[20] & in2[20];
    assign P[166] = in[20] ^ in2[20];
    assign G[167] = in[19] & in2[19];
    assign P[167] = in[19] ^ in2[19];
    assign G[168] = in[18] & in2[18];
    assign P[168] = in[18] ^ in2[18];
    assign G[169] = in[17] & in2[17];
    assign P[169] = in[17] ^ in2[17];
    assign G[170] = in[16] & in2[16];
    assign P[170] = in[16] ^ in2[16];
    assign G[171] = in[15] & in2[15];
    assign P[171] = in[15] ^ in2[15];
    assign G[172] = in[14] & in2[14];
    assign P[172] = in[14] ^ in2[14];
    assign G[173] = in[13] & in2[13];
    assign P[173] = in[13] ^ in2[13];
    assign G[174] = in[12] & in2[12];
    assign P[174] = in[12] ^ in2[12];
    assign G[175] = in[11] & in2[11];
    assign P[175] = in[11] ^ in2[11];
    assign G[176] = in[10] & in2[10];
    assign P[176] = in[10] ^ in2[10];
    assign G[177] = in[9] & in2[9];
    assign P[177] = in[9] ^ in2[9];
    assign G[178] = in[8] & in2[8];
    assign P[178] = in[8] ^ in2[8];
    assign G[179] = in[7] & in2[7];
    assign P[179] = in[7] ^ in2[7];
    assign G[180] = in[6] & in2[6];
    assign P[180] = in[6] ^ in2[6];
    assign G[181] = in[5] & in2[5];
    assign P[181] = in[5] ^ in2[5];
    assign G[182] = in[4] & in2[4];
    assign P[182] = in[4] ^ in2[4];
    assign G[183] = in[3] & in2[3];
    assign P[183] = in[3] ^ in2[3];
    assign G[184] = in[2] & in2[2];
    assign P[184] = in[2] ^ in2[2];
    assign G[185] = in[1] & in2[1];
    assign P[185] = in[1] ^ in2[1];
    assign G[186] = in[0] & in2[0];
    assign P[186] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign C[186] = G[185] | (P[185] & C[185]);
    assign cout = G[186] | (P[186] & C[186]);
    assign sum = P ^ C;
endmodule

module CLA186(output [185:0] sum, output cout, input [185:0] in1, input [185:0] in2;

    wire[185:0] G;
    wire[185:0] C;
    wire[185:0] P;

    assign G[0] = in[185] & in2[185];
    assign P[0] = in[185] ^ in2[185];
    assign G[1] = in[184] & in2[184];
    assign P[1] = in[184] ^ in2[184];
    assign G[2] = in[183] & in2[183];
    assign P[2] = in[183] ^ in2[183];
    assign G[3] = in[182] & in2[182];
    assign P[3] = in[182] ^ in2[182];
    assign G[4] = in[181] & in2[181];
    assign P[4] = in[181] ^ in2[181];
    assign G[5] = in[180] & in2[180];
    assign P[5] = in[180] ^ in2[180];
    assign G[6] = in[179] & in2[179];
    assign P[6] = in[179] ^ in2[179];
    assign G[7] = in[178] & in2[178];
    assign P[7] = in[178] ^ in2[178];
    assign G[8] = in[177] & in2[177];
    assign P[8] = in[177] ^ in2[177];
    assign G[9] = in[176] & in2[176];
    assign P[9] = in[176] ^ in2[176];
    assign G[10] = in[175] & in2[175];
    assign P[10] = in[175] ^ in2[175];
    assign G[11] = in[174] & in2[174];
    assign P[11] = in[174] ^ in2[174];
    assign G[12] = in[173] & in2[173];
    assign P[12] = in[173] ^ in2[173];
    assign G[13] = in[172] & in2[172];
    assign P[13] = in[172] ^ in2[172];
    assign G[14] = in[171] & in2[171];
    assign P[14] = in[171] ^ in2[171];
    assign G[15] = in[170] & in2[170];
    assign P[15] = in[170] ^ in2[170];
    assign G[16] = in[169] & in2[169];
    assign P[16] = in[169] ^ in2[169];
    assign G[17] = in[168] & in2[168];
    assign P[17] = in[168] ^ in2[168];
    assign G[18] = in[167] & in2[167];
    assign P[18] = in[167] ^ in2[167];
    assign G[19] = in[166] & in2[166];
    assign P[19] = in[166] ^ in2[166];
    assign G[20] = in[165] & in2[165];
    assign P[20] = in[165] ^ in2[165];
    assign G[21] = in[164] & in2[164];
    assign P[21] = in[164] ^ in2[164];
    assign G[22] = in[163] & in2[163];
    assign P[22] = in[163] ^ in2[163];
    assign G[23] = in[162] & in2[162];
    assign P[23] = in[162] ^ in2[162];
    assign G[24] = in[161] & in2[161];
    assign P[24] = in[161] ^ in2[161];
    assign G[25] = in[160] & in2[160];
    assign P[25] = in[160] ^ in2[160];
    assign G[26] = in[159] & in2[159];
    assign P[26] = in[159] ^ in2[159];
    assign G[27] = in[158] & in2[158];
    assign P[27] = in[158] ^ in2[158];
    assign G[28] = in[157] & in2[157];
    assign P[28] = in[157] ^ in2[157];
    assign G[29] = in[156] & in2[156];
    assign P[29] = in[156] ^ in2[156];
    assign G[30] = in[155] & in2[155];
    assign P[30] = in[155] ^ in2[155];
    assign G[31] = in[154] & in2[154];
    assign P[31] = in[154] ^ in2[154];
    assign G[32] = in[153] & in2[153];
    assign P[32] = in[153] ^ in2[153];
    assign G[33] = in[152] & in2[152];
    assign P[33] = in[152] ^ in2[152];
    assign G[34] = in[151] & in2[151];
    assign P[34] = in[151] ^ in2[151];
    assign G[35] = in[150] & in2[150];
    assign P[35] = in[150] ^ in2[150];
    assign G[36] = in[149] & in2[149];
    assign P[36] = in[149] ^ in2[149];
    assign G[37] = in[148] & in2[148];
    assign P[37] = in[148] ^ in2[148];
    assign G[38] = in[147] & in2[147];
    assign P[38] = in[147] ^ in2[147];
    assign G[39] = in[146] & in2[146];
    assign P[39] = in[146] ^ in2[146];
    assign G[40] = in[145] & in2[145];
    assign P[40] = in[145] ^ in2[145];
    assign G[41] = in[144] & in2[144];
    assign P[41] = in[144] ^ in2[144];
    assign G[42] = in[143] & in2[143];
    assign P[42] = in[143] ^ in2[143];
    assign G[43] = in[142] & in2[142];
    assign P[43] = in[142] ^ in2[142];
    assign G[44] = in[141] & in2[141];
    assign P[44] = in[141] ^ in2[141];
    assign G[45] = in[140] & in2[140];
    assign P[45] = in[140] ^ in2[140];
    assign G[46] = in[139] & in2[139];
    assign P[46] = in[139] ^ in2[139];
    assign G[47] = in[138] & in2[138];
    assign P[47] = in[138] ^ in2[138];
    assign G[48] = in[137] & in2[137];
    assign P[48] = in[137] ^ in2[137];
    assign G[49] = in[136] & in2[136];
    assign P[49] = in[136] ^ in2[136];
    assign G[50] = in[135] & in2[135];
    assign P[50] = in[135] ^ in2[135];
    assign G[51] = in[134] & in2[134];
    assign P[51] = in[134] ^ in2[134];
    assign G[52] = in[133] & in2[133];
    assign P[52] = in[133] ^ in2[133];
    assign G[53] = in[132] & in2[132];
    assign P[53] = in[132] ^ in2[132];
    assign G[54] = in[131] & in2[131];
    assign P[54] = in[131] ^ in2[131];
    assign G[55] = in[130] & in2[130];
    assign P[55] = in[130] ^ in2[130];
    assign G[56] = in[129] & in2[129];
    assign P[56] = in[129] ^ in2[129];
    assign G[57] = in[128] & in2[128];
    assign P[57] = in[128] ^ in2[128];
    assign G[58] = in[127] & in2[127];
    assign P[58] = in[127] ^ in2[127];
    assign G[59] = in[126] & in2[126];
    assign P[59] = in[126] ^ in2[126];
    assign G[60] = in[125] & in2[125];
    assign P[60] = in[125] ^ in2[125];
    assign G[61] = in[124] & in2[124];
    assign P[61] = in[124] ^ in2[124];
    assign G[62] = in[123] & in2[123];
    assign P[62] = in[123] ^ in2[123];
    assign G[63] = in[122] & in2[122];
    assign P[63] = in[122] ^ in2[122];
    assign G[64] = in[121] & in2[121];
    assign P[64] = in[121] ^ in2[121];
    assign G[65] = in[120] & in2[120];
    assign P[65] = in[120] ^ in2[120];
    assign G[66] = in[119] & in2[119];
    assign P[66] = in[119] ^ in2[119];
    assign G[67] = in[118] & in2[118];
    assign P[67] = in[118] ^ in2[118];
    assign G[68] = in[117] & in2[117];
    assign P[68] = in[117] ^ in2[117];
    assign G[69] = in[116] & in2[116];
    assign P[69] = in[116] ^ in2[116];
    assign G[70] = in[115] & in2[115];
    assign P[70] = in[115] ^ in2[115];
    assign G[71] = in[114] & in2[114];
    assign P[71] = in[114] ^ in2[114];
    assign G[72] = in[113] & in2[113];
    assign P[72] = in[113] ^ in2[113];
    assign G[73] = in[112] & in2[112];
    assign P[73] = in[112] ^ in2[112];
    assign G[74] = in[111] & in2[111];
    assign P[74] = in[111] ^ in2[111];
    assign G[75] = in[110] & in2[110];
    assign P[75] = in[110] ^ in2[110];
    assign G[76] = in[109] & in2[109];
    assign P[76] = in[109] ^ in2[109];
    assign G[77] = in[108] & in2[108];
    assign P[77] = in[108] ^ in2[108];
    assign G[78] = in[107] & in2[107];
    assign P[78] = in[107] ^ in2[107];
    assign G[79] = in[106] & in2[106];
    assign P[79] = in[106] ^ in2[106];
    assign G[80] = in[105] & in2[105];
    assign P[80] = in[105] ^ in2[105];
    assign G[81] = in[104] & in2[104];
    assign P[81] = in[104] ^ in2[104];
    assign G[82] = in[103] & in2[103];
    assign P[82] = in[103] ^ in2[103];
    assign G[83] = in[102] & in2[102];
    assign P[83] = in[102] ^ in2[102];
    assign G[84] = in[101] & in2[101];
    assign P[84] = in[101] ^ in2[101];
    assign G[85] = in[100] & in2[100];
    assign P[85] = in[100] ^ in2[100];
    assign G[86] = in[99] & in2[99];
    assign P[86] = in[99] ^ in2[99];
    assign G[87] = in[98] & in2[98];
    assign P[87] = in[98] ^ in2[98];
    assign G[88] = in[97] & in2[97];
    assign P[88] = in[97] ^ in2[97];
    assign G[89] = in[96] & in2[96];
    assign P[89] = in[96] ^ in2[96];
    assign G[90] = in[95] & in2[95];
    assign P[90] = in[95] ^ in2[95];
    assign G[91] = in[94] & in2[94];
    assign P[91] = in[94] ^ in2[94];
    assign G[92] = in[93] & in2[93];
    assign P[92] = in[93] ^ in2[93];
    assign G[93] = in[92] & in2[92];
    assign P[93] = in[92] ^ in2[92];
    assign G[94] = in[91] & in2[91];
    assign P[94] = in[91] ^ in2[91];
    assign G[95] = in[90] & in2[90];
    assign P[95] = in[90] ^ in2[90];
    assign G[96] = in[89] & in2[89];
    assign P[96] = in[89] ^ in2[89];
    assign G[97] = in[88] & in2[88];
    assign P[97] = in[88] ^ in2[88];
    assign G[98] = in[87] & in2[87];
    assign P[98] = in[87] ^ in2[87];
    assign G[99] = in[86] & in2[86];
    assign P[99] = in[86] ^ in2[86];
    assign G[100] = in[85] & in2[85];
    assign P[100] = in[85] ^ in2[85];
    assign G[101] = in[84] & in2[84];
    assign P[101] = in[84] ^ in2[84];
    assign G[102] = in[83] & in2[83];
    assign P[102] = in[83] ^ in2[83];
    assign G[103] = in[82] & in2[82];
    assign P[103] = in[82] ^ in2[82];
    assign G[104] = in[81] & in2[81];
    assign P[104] = in[81] ^ in2[81];
    assign G[105] = in[80] & in2[80];
    assign P[105] = in[80] ^ in2[80];
    assign G[106] = in[79] & in2[79];
    assign P[106] = in[79] ^ in2[79];
    assign G[107] = in[78] & in2[78];
    assign P[107] = in[78] ^ in2[78];
    assign G[108] = in[77] & in2[77];
    assign P[108] = in[77] ^ in2[77];
    assign G[109] = in[76] & in2[76];
    assign P[109] = in[76] ^ in2[76];
    assign G[110] = in[75] & in2[75];
    assign P[110] = in[75] ^ in2[75];
    assign G[111] = in[74] & in2[74];
    assign P[111] = in[74] ^ in2[74];
    assign G[112] = in[73] & in2[73];
    assign P[112] = in[73] ^ in2[73];
    assign G[113] = in[72] & in2[72];
    assign P[113] = in[72] ^ in2[72];
    assign G[114] = in[71] & in2[71];
    assign P[114] = in[71] ^ in2[71];
    assign G[115] = in[70] & in2[70];
    assign P[115] = in[70] ^ in2[70];
    assign G[116] = in[69] & in2[69];
    assign P[116] = in[69] ^ in2[69];
    assign G[117] = in[68] & in2[68];
    assign P[117] = in[68] ^ in2[68];
    assign G[118] = in[67] & in2[67];
    assign P[118] = in[67] ^ in2[67];
    assign G[119] = in[66] & in2[66];
    assign P[119] = in[66] ^ in2[66];
    assign G[120] = in[65] & in2[65];
    assign P[120] = in[65] ^ in2[65];
    assign G[121] = in[64] & in2[64];
    assign P[121] = in[64] ^ in2[64];
    assign G[122] = in[63] & in2[63];
    assign P[122] = in[63] ^ in2[63];
    assign G[123] = in[62] & in2[62];
    assign P[123] = in[62] ^ in2[62];
    assign G[124] = in[61] & in2[61];
    assign P[124] = in[61] ^ in2[61];
    assign G[125] = in[60] & in2[60];
    assign P[125] = in[60] ^ in2[60];
    assign G[126] = in[59] & in2[59];
    assign P[126] = in[59] ^ in2[59];
    assign G[127] = in[58] & in2[58];
    assign P[127] = in[58] ^ in2[58];
    assign G[128] = in[57] & in2[57];
    assign P[128] = in[57] ^ in2[57];
    assign G[129] = in[56] & in2[56];
    assign P[129] = in[56] ^ in2[56];
    assign G[130] = in[55] & in2[55];
    assign P[130] = in[55] ^ in2[55];
    assign G[131] = in[54] & in2[54];
    assign P[131] = in[54] ^ in2[54];
    assign G[132] = in[53] & in2[53];
    assign P[132] = in[53] ^ in2[53];
    assign G[133] = in[52] & in2[52];
    assign P[133] = in[52] ^ in2[52];
    assign G[134] = in[51] & in2[51];
    assign P[134] = in[51] ^ in2[51];
    assign G[135] = in[50] & in2[50];
    assign P[135] = in[50] ^ in2[50];
    assign G[136] = in[49] & in2[49];
    assign P[136] = in[49] ^ in2[49];
    assign G[137] = in[48] & in2[48];
    assign P[137] = in[48] ^ in2[48];
    assign G[138] = in[47] & in2[47];
    assign P[138] = in[47] ^ in2[47];
    assign G[139] = in[46] & in2[46];
    assign P[139] = in[46] ^ in2[46];
    assign G[140] = in[45] & in2[45];
    assign P[140] = in[45] ^ in2[45];
    assign G[141] = in[44] & in2[44];
    assign P[141] = in[44] ^ in2[44];
    assign G[142] = in[43] & in2[43];
    assign P[142] = in[43] ^ in2[43];
    assign G[143] = in[42] & in2[42];
    assign P[143] = in[42] ^ in2[42];
    assign G[144] = in[41] & in2[41];
    assign P[144] = in[41] ^ in2[41];
    assign G[145] = in[40] & in2[40];
    assign P[145] = in[40] ^ in2[40];
    assign G[146] = in[39] & in2[39];
    assign P[146] = in[39] ^ in2[39];
    assign G[147] = in[38] & in2[38];
    assign P[147] = in[38] ^ in2[38];
    assign G[148] = in[37] & in2[37];
    assign P[148] = in[37] ^ in2[37];
    assign G[149] = in[36] & in2[36];
    assign P[149] = in[36] ^ in2[36];
    assign G[150] = in[35] & in2[35];
    assign P[150] = in[35] ^ in2[35];
    assign G[151] = in[34] & in2[34];
    assign P[151] = in[34] ^ in2[34];
    assign G[152] = in[33] & in2[33];
    assign P[152] = in[33] ^ in2[33];
    assign G[153] = in[32] & in2[32];
    assign P[153] = in[32] ^ in2[32];
    assign G[154] = in[31] & in2[31];
    assign P[154] = in[31] ^ in2[31];
    assign G[155] = in[30] & in2[30];
    assign P[155] = in[30] ^ in2[30];
    assign G[156] = in[29] & in2[29];
    assign P[156] = in[29] ^ in2[29];
    assign G[157] = in[28] & in2[28];
    assign P[157] = in[28] ^ in2[28];
    assign G[158] = in[27] & in2[27];
    assign P[158] = in[27] ^ in2[27];
    assign G[159] = in[26] & in2[26];
    assign P[159] = in[26] ^ in2[26];
    assign G[160] = in[25] & in2[25];
    assign P[160] = in[25] ^ in2[25];
    assign G[161] = in[24] & in2[24];
    assign P[161] = in[24] ^ in2[24];
    assign G[162] = in[23] & in2[23];
    assign P[162] = in[23] ^ in2[23];
    assign G[163] = in[22] & in2[22];
    assign P[163] = in[22] ^ in2[22];
    assign G[164] = in[21] & in2[21];
    assign P[164] = in[21] ^ in2[21];
    assign G[165] = in[20] & in2[20];
    assign P[165] = in[20] ^ in2[20];
    assign G[166] = in[19] & in2[19];
    assign P[166] = in[19] ^ in2[19];
    assign G[167] = in[18] & in2[18];
    assign P[167] = in[18] ^ in2[18];
    assign G[168] = in[17] & in2[17];
    assign P[168] = in[17] ^ in2[17];
    assign G[169] = in[16] & in2[16];
    assign P[169] = in[16] ^ in2[16];
    assign G[170] = in[15] & in2[15];
    assign P[170] = in[15] ^ in2[15];
    assign G[171] = in[14] & in2[14];
    assign P[171] = in[14] ^ in2[14];
    assign G[172] = in[13] & in2[13];
    assign P[172] = in[13] ^ in2[13];
    assign G[173] = in[12] & in2[12];
    assign P[173] = in[12] ^ in2[12];
    assign G[174] = in[11] & in2[11];
    assign P[174] = in[11] ^ in2[11];
    assign G[175] = in[10] & in2[10];
    assign P[175] = in[10] ^ in2[10];
    assign G[176] = in[9] & in2[9];
    assign P[176] = in[9] ^ in2[9];
    assign G[177] = in[8] & in2[8];
    assign P[177] = in[8] ^ in2[8];
    assign G[178] = in[7] & in2[7];
    assign P[178] = in[7] ^ in2[7];
    assign G[179] = in[6] & in2[6];
    assign P[179] = in[6] ^ in2[6];
    assign G[180] = in[5] & in2[5];
    assign P[180] = in[5] ^ in2[5];
    assign G[181] = in[4] & in2[4];
    assign P[181] = in[4] ^ in2[4];
    assign G[182] = in[3] & in2[3];
    assign P[182] = in[3] ^ in2[3];
    assign G[183] = in[2] & in2[2];
    assign P[183] = in[2] ^ in2[2];
    assign G[184] = in[1] & in2[1];
    assign P[184] = in[1] ^ in2[1];
    assign G[185] = in[0] & in2[0];
    assign P[185] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign C[185] = G[184] | (P[184] & C[184]);
    assign cout = G[185] | (P[185] & C[185]);
    assign sum = P ^ C;
endmodule

module CLA185(output [184:0] sum, output cout, input [184:0] in1, input [184:0] in2;

    wire[184:0] G;
    wire[184:0] C;
    wire[184:0] P;

    assign G[0] = in[184] & in2[184];
    assign P[0] = in[184] ^ in2[184];
    assign G[1] = in[183] & in2[183];
    assign P[1] = in[183] ^ in2[183];
    assign G[2] = in[182] & in2[182];
    assign P[2] = in[182] ^ in2[182];
    assign G[3] = in[181] & in2[181];
    assign P[3] = in[181] ^ in2[181];
    assign G[4] = in[180] & in2[180];
    assign P[4] = in[180] ^ in2[180];
    assign G[5] = in[179] & in2[179];
    assign P[5] = in[179] ^ in2[179];
    assign G[6] = in[178] & in2[178];
    assign P[6] = in[178] ^ in2[178];
    assign G[7] = in[177] & in2[177];
    assign P[7] = in[177] ^ in2[177];
    assign G[8] = in[176] & in2[176];
    assign P[8] = in[176] ^ in2[176];
    assign G[9] = in[175] & in2[175];
    assign P[9] = in[175] ^ in2[175];
    assign G[10] = in[174] & in2[174];
    assign P[10] = in[174] ^ in2[174];
    assign G[11] = in[173] & in2[173];
    assign P[11] = in[173] ^ in2[173];
    assign G[12] = in[172] & in2[172];
    assign P[12] = in[172] ^ in2[172];
    assign G[13] = in[171] & in2[171];
    assign P[13] = in[171] ^ in2[171];
    assign G[14] = in[170] & in2[170];
    assign P[14] = in[170] ^ in2[170];
    assign G[15] = in[169] & in2[169];
    assign P[15] = in[169] ^ in2[169];
    assign G[16] = in[168] & in2[168];
    assign P[16] = in[168] ^ in2[168];
    assign G[17] = in[167] & in2[167];
    assign P[17] = in[167] ^ in2[167];
    assign G[18] = in[166] & in2[166];
    assign P[18] = in[166] ^ in2[166];
    assign G[19] = in[165] & in2[165];
    assign P[19] = in[165] ^ in2[165];
    assign G[20] = in[164] & in2[164];
    assign P[20] = in[164] ^ in2[164];
    assign G[21] = in[163] & in2[163];
    assign P[21] = in[163] ^ in2[163];
    assign G[22] = in[162] & in2[162];
    assign P[22] = in[162] ^ in2[162];
    assign G[23] = in[161] & in2[161];
    assign P[23] = in[161] ^ in2[161];
    assign G[24] = in[160] & in2[160];
    assign P[24] = in[160] ^ in2[160];
    assign G[25] = in[159] & in2[159];
    assign P[25] = in[159] ^ in2[159];
    assign G[26] = in[158] & in2[158];
    assign P[26] = in[158] ^ in2[158];
    assign G[27] = in[157] & in2[157];
    assign P[27] = in[157] ^ in2[157];
    assign G[28] = in[156] & in2[156];
    assign P[28] = in[156] ^ in2[156];
    assign G[29] = in[155] & in2[155];
    assign P[29] = in[155] ^ in2[155];
    assign G[30] = in[154] & in2[154];
    assign P[30] = in[154] ^ in2[154];
    assign G[31] = in[153] & in2[153];
    assign P[31] = in[153] ^ in2[153];
    assign G[32] = in[152] & in2[152];
    assign P[32] = in[152] ^ in2[152];
    assign G[33] = in[151] & in2[151];
    assign P[33] = in[151] ^ in2[151];
    assign G[34] = in[150] & in2[150];
    assign P[34] = in[150] ^ in2[150];
    assign G[35] = in[149] & in2[149];
    assign P[35] = in[149] ^ in2[149];
    assign G[36] = in[148] & in2[148];
    assign P[36] = in[148] ^ in2[148];
    assign G[37] = in[147] & in2[147];
    assign P[37] = in[147] ^ in2[147];
    assign G[38] = in[146] & in2[146];
    assign P[38] = in[146] ^ in2[146];
    assign G[39] = in[145] & in2[145];
    assign P[39] = in[145] ^ in2[145];
    assign G[40] = in[144] & in2[144];
    assign P[40] = in[144] ^ in2[144];
    assign G[41] = in[143] & in2[143];
    assign P[41] = in[143] ^ in2[143];
    assign G[42] = in[142] & in2[142];
    assign P[42] = in[142] ^ in2[142];
    assign G[43] = in[141] & in2[141];
    assign P[43] = in[141] ^ in2[141];
    assign G[44] = in[140] & in2[140];
    assign P[44] = in[140] ^ in2[140];
    assign G[45] = in[139] & in2[139];
    assign P[45] = in[139] ^ in2[139];
    assign G[46] = in[138] & in2[138];
    assign P[46] = in[138] ^ in2[138];
    assign G[47] = in[137] & in2[137];
    assign P[47] = in[137] ^ in2[137];
    assign G[48] = in[136] & in2[136];
    assign P[48] = in[136] ^ in2[136];
    assign G[49] = in[135] & in2[135];
    assign P[49] = in[135] ^ in2[135];
    assign G[50] = in[134] & in2[134];
    assign P[50] = in[134] ^ in2[134];
    assign G[51] = in[133] & in2[133];
    assign P[51] = in[133] ^ in2[133];
    assign G[52] = in[132] & in2[132];
    assign P[52] = in[132] ^ in2[132];
    assign G[53] = in[131] & in2[131];
    assign P[53] = in[131] ^ in2[131];
    assign G[54] = in[130] & in2[130];
    assign P[54] = in[130] ^ in2[130];
    assign G[55] = in[129] & in2[129];
    assign P[55] = in[129] ^ in2[129];
    assign G[56] = in[128] & in2[128];
    assign P[56] = in[128] ^ in2[128];
    assign G[57] = in[127] & in2[127];
    assign P[57] = in[127] ^ in2[127];
    assign G[58] = in[126] & in2[126];
    assign P[58] = in[126] ^ in2[126];
    assign G[59] = in[125] & in2[125];
    assign P[59] = in[125] ^ in2[125];
    assign G[60] = in[124] & in2[124];
    assign P[60] = in[124] ^ in2[124];
    assign G[61] = in[123] & in2[123];
    assign P[61] = in[123] ^ in2[123];
    assign G[62] = in[122] & in2[122];
    assign P[62] = in[122] ^ in2[122];
    assign G[63] = in[121] & in2[121];
    assign P[63] = in[121] ^ in2[121];
    assign G[64] = in[120] & in2[120];
    assign P[64] = in[120] ^ in2[120];
    assign G[65] = in[119] & in2[119];
    assign P[65] = in[119] ^ in2[119];
    assign G[66] = in[118] & in2[118];
    assign P[66] = in[118] ^ in2[118];
    assign G[67] = in[117] & in2[117];
    assign P[67] = in[117] ^ in2[117];
    assign G[68] = in[116] & in2[116];
    assign P[68] = in[116] ^ in2[116];
    assign G[69] = in[115] & in2[115];
    assign P[69] = in[115] ^ in2[115];
    assign G[70] = in[114] & in2[114];
    assign P[70] = in[114] ^ in2[114];
    assign G[71] = in[113] & in2[113];
    assign P[71] = in[113] ^ in2[113];
    assign G[72] = in[112] & in2[112];
    assign P[72] = in[112] ^ in2[112];
    assign G[73] = in[111] & in2[111];
    assign P[73] = in[111] ^ in2[111];
    assign G[74] = in[110] & in2[110];
    assign P[74] = in[110] ^ in2[110];
    assign G[75] = in[109] & in2[109];
    assign P[75] = in[109] ^ in2[109];
    assign G[76] = in[108] & in2[108];
    assign P[76] = in[108] ^ in2[108];
    assign G[77] = in[107] & in2[107];
    assign P[77] = in[107] ^ in2[107];
    assign G[78] = in[106] & in2[106];
    assign P[78] = in[106] ^ in2[106];
    assign G[79] = in[105] & in2[105];
    assign P[79] = in[105] ^ in2[105];
    assign G[80] = in[104] & in2[104];
    assign P[80] = in[104] ^ in2[104];
    assign G[81] = in[103] & in2[103];
    assign P[81] = in[103] ^ in2[103];
    assign G[82] = in[102] & in2[102];
    assign P[82] = in[102] ^ in2[102];
    assign G[83] = in[101] & in2[101];
    assign P[83] = in[101] ^ in2[101];
    assign G[84] = in[100] & in2[100];
    assign P[84] = in[100] ^ in2[100];
    assign G[85] = in[99] & in2[99];
    assign P[85] = in[99] ^ in2[99];
    assign G[86] = in[98] & in2[98];
    assign P[86] = in[98] ^ in2[98];
    assign G[87] = in[97] & in2[97];
    assign P[87] = in[97] ^ in2[97];
    assign G[88] = in[96] & in2[96];
    assign P[88] = in[96] ^ in2[96];
    assign G[89] = in[95] & in2[95];
    assign P[89] = in[95] ^ in2[95];
    assign G[90] = in[94] & in2[94];
    assign P[90] = in[94] ^ in2[94];
    assign G[91] = in[93] & in2[93];
    assign P[91] = in[93] ^ in2[93];
    assign G[92] = in[92] & in2[92];
    assign P[92] = in[92] ^ in2[92];
    assign G[93] = in[91] & in2[91];
    assign P[93] = in[91] ^ in2[91];
    assign G[94] = in[90] & in2[90];
    assign P[94] = in[90] ^ in2[90];
    assign G[95] = in[89] & in2[89];
    assign P[95] = in[89] ^ in2[89];
    assign G[96] = in[88] & in2[88];
    assign P[96] = in[88] ^ in2[88];
    assign G[97] = in[87] & in2[87];
    assign P[97] = in[87] ^ in2[87];
    assign G[98] = in[86] & in2[86];
    assign P[98] = in[86] ^ in2[86];
    assign G[99] = in[85] & in2[85];
    assign P[99] = in[85] ^ in2[85];
    assign G[100] = in[84] & in2[84];
    assign P[100] = in[84] ^ in2[84];
    assign G[101] = in[83] & in2[83];
    assign P[101] = in[83] ^ in2[83];
    assign G[102] = in[82] & in2[82];
    assign P[102] = in[82] ^ in2[82];
    assign G[103] = in[81] & in2[81];
    assign P[103] = in[81] ^ in2[81];
    assign G[104] = in[80] & in2[80];
    assign P[104] = in[80] ^ in2[80];
    assign G[105] = in[79] & in2[79];
    assign P[105] = in[79] ^ in2[79];
    assign G[106] = in[78] & in2[78];
    assign P[106] = in[78] ^ in2[78];
    assign G[107] = in[77] & in2[77];
    assign P[107] = in[77] ^ in2[77];
    assign G[108] = in[76] & in2[76];
    assign P[108] = in[76] ^ in2[76];
    assign G[109] = in[75] & in2[75];
    assign P[109] = in[75] ^ in2[75];
    assign G[110] = in[74] & in2[74];
    assign P[110] = in[74] ^ in2[74];
    assign G[111] = in[73] & in2[73];
    assign P[111] = in[73] ^ in2[73];
    assign G[112] = in[72] & in2[72];
    assign P[112] = in[72] ^ in2[72];
    assign G[113] = in[71] & in2[71];
    assign P[113] = in[71] ^ in2[71];
    assign G[114] = in[70] & in2[70];
    assign P[114] = in[70] ^ in2[70];
    assign G[115] = in[69] & in2[69];
    assign P[115] = in[69] ^ in2[69];
    assign G[116] = in[68] & in2[68];
    assign P[116] = in[68] ^ in2[68];
    assign G[117] = in[67] & in2[67];
    assign P[117] = in[67] ^ in2[67];
    assign G[118] = in[66] & in2[66];
    assign P[118] = in[66] ^ in2[66];
    assign G[119] = in[65] & in2[65];
    assign P[119] = in[65] ^ in2[65];
    assign G[120] = in[64] & in2[64];
    assign P[120] = in[64] ^ in2[64];
    assign G[121] = in[63] & in2[63];
    assign P[121] = in[63] ^ in2[63];
    assign G[122] = in[62] & in2[62];
    assign P[122] = in[62] ^ in2[62];
    assign G[123] = in[61] & in2[61];
    assign P[123] = in[61] ^ in2[61];
    assign G[124] = in[60] & in2[60];
    assign P[124] = in[60] ^ in2[60];
    assign G[125] = in[59] & in2[59];
    assign P[125] = in[59] ^ in2[59];
    assign G[126] = in[58] & in2[58];
    assign P[126] = in[58] ^ in2[58];
    assign G[127] = in[57] & in2[57];
    assign P[127] = in[57] ^ in2[57];
    assign G[128] = in[56] & in2[56];
    assign P[128] = in[56] ^ in2[56];
    assign G[129] = in[55] & in2[55];
    assign P[129] = in[55] ^ in2[55];
    assign G[130] = in[54] & in2[54];
    assign P[130] = in[54] ^ in2[54];
    assign G[131] = in[53] & in2[53];
    assign P[131] = in[53] ^ in2[53];
    assign G[132] = in[52] & in2[52];
    assign P[132] = in[52] ^ in2[52];
    assign G[133] = in[51] & in2[51];
    assign P[133] = in[51] ^ in2[51];
    assign G[134] = in[50] & in2[50];
    assign P[134] = in[50] ^ in2[50];
    assign G[135] = in[49] & in2[49];
    assign P[135] = in[49] ^ in2[49];
    assign G[136] = in[48] & in2[48];
    assign P[136] = in[48] ^ in2[48];
    assign G[137] = in[47] & in2[47];
    assign P[137] = in[47] ^ in2[47];
    assign G[138] = in[46] & in2[46];
    assign P[138] = in[46] ^ in2[46];
    assign G[139] = in[45] & in2[45];
    assign P[139] = in[45] ^ in2[45];
    assign G[140] = in[44] & in2[44];
    assign P[140] = in[44] ^ in2[44];
    assign G[141] = in[43] & in2[43];
    assign P[141] = in[43] ^ in2[43];
    assign G[142] = in[42] & in2[42];
    assign P[142] = in[42] ^ in2[42];
    assign G[143] = in[41] & in2[41];
    assign P[143] = in[41] ^ in2[41];
    assign G[144] = in[40] & in2[40];
    assign P[144] = in[40] ^ in2[40];
    assign G[145] = in[39] & in2[39];
    assign P[145] = in[39] ^ in2[39];
    assign G[146] = in[38] & in2[38];
    assign P[146] = in[38] ^ in2[38];
    assign G[147] = in[37] & in2[37];
    assign P[147] = in[37] ^ in2[37];
    assign G[148] = in[36] & in2[36];
    assign P[148] = in[36] ^ in2[36];
    assign G[149] = in[35] & in2[35];
    assign P[149] = in[35] ^ in2[35];
    assign G[150] = in[34] & in2[34];
    assign P[150] = in[34] ^ in2[34];
    assign G[151] = in[33] & in2[33];
    assign P[151] = in[33] ^ in2[33];
    assign G[152] = in[32] & in2[32];
    assign P[152] = in[32] ^ in2[32];
    assign G[153] = in[31] & in2[31];
    assign P[153] = in[31] ^ in2[31];
    assign G[154] = in[30] & in2[30];
    assign P[154] = in[30] ^ in2[30];
    assign G[155] = in[29] & in2[29];
    assign P[155] = in[29] ^ in2[29];
    assign G[156] = in[28] & in2[28];
    assign P[156] = in[28] ^ in2[28];
    assign G[157] = in[27] & in2[27];
    assign P[157] = in[27] ^ in2[27];
    assign G[158] = in[26] & in2[26];
    assign P[158] = in[26] ^ in2[26];
    assign G[159] = in[25] & in2[25];
    assign P[159] = in[25] ^ in2[25];
    assign G[160] = in[24] & in2[24];
    assign P[160] = in[24] ^ in2[24];
    assign G[161] = in[23] & in2[23];
    assign P[161] = in[23] ^ in2[23];
    assign G[162] = in[22] & in2[22];
    assign P[162] = in[22] ^ in2[22];
    assign G[163] = in[21] & in2[21];
    assign P[163] = in[21] ^ in2[21];
    assign G[164] = in[20] & in2[20];
    assign P[164] = in[20] ^ in2[20];
    assign G[165] = in[19] & in2[19];
    assign P[165] = in[19] ^ in2[19];
    assign G[166] = in[18] & in2[18];
    assign P[166] = in[18] ^ in2[18];
    assign G[167] = in[17] & in2[17];
    assign P[167] = in[17] ^ in2[17];
    assign G[168] = in[16] & in2[16];
    assign P[168] = in[16] ^ in2[16];
    assign G[169] = in[15] & in2[15];
    assign P[169] = in[15] ^ in2[15];
    assign G[170] = in[14] & in2[14];
    assign P[170] = in[14] ^ in2[14];
    assign G[171] = in[13] & in2[13];
    assign P[171] = in[13] ^ in2[13];
    assign G[172] = in[12] & in2[12];
    assign P[172] = in[12] ^ in2[12];
    assign G[173] = in[11] & in2[11];
    assign P[173] = in[11] ^ in2[11];
    assign G[174] = in[10] & in2[10];
    assign P[174] = in[10] ^ in2[10];
    assign G[175] = in[9] & in2[9];
    assign P[175] = in[9] ^ in2[9];
    assign G[176] = in[8] & in2[8];
    assign P[176] = in[8] ^ in2[8];
    assign G[177] = in[7] & in2[7];
    assign P[177] = in[7] ^ in2[7];
    assign G[178] = in[6] & in2[6];
    assign P[178] = in[6] ^ in2[6];
    assign G[179] = in[5] & in2[5];
    assign P[179] = in[5] ^ in2[5];
    assign G[180] = in[4] & in2[4];
    assign P[180] = in[4] ^ in2[4];
    assign G[181] = in[3] & in2[3];
    assign P[181] = in[3] ^ in2[3];
    assign G[182] = in[2] & in2[2];
    assign P[182] = in[2] ^ in2[2];
    assign G[183] = in[1] & in2[1];
    assign P[183] = in[1] ^ in2[1];
    assign G[184] = in[0] & in2[0];
    assign P[184] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign C[184] = G[183] | (P[183] & C[183]);
    assign cout = G[184] | (P[184] & C[184]);
    assign sum = P ^ C;
endmodule

module CLA184(output [183:0] sum, output cout, input [183:0] in1, input [183:0] in2;

    wire[183:0] G;
    wire[183:0] C;
    wire[183:0] P;

    assign G[0] = in[183] & in2[183];
    assign P[0] = in[183] ^ in2[183];
    assign G[1] = in[182] & in2[182];
    assign P[1] = in[182] ^ in2[182];
    assign G[2] = in[181] & in2[181];
    assign P[2] = in[181] ^ in2[181];
    assign G[3] = in[180] & in2[180];
    assign P[3] = in[180] ^ in2[180];
    assign G[4] = in[179] & in2[179];
    assign P[4] = in[179] ^ in2[179];
    assign G[5] = in[178] & in2[178];
    assign P[5] = in[178] ^ in2[178];
    assign G[6] = in[177] & in2[177];
    assign P[6] = in[177] ^ in2[177];
    assign G[7] = in[176] & in2[176];
    assign P[7] = in[176] ^ in2[176];
    assign G[8] = in[175] & in2[175];
    assign P[8] = in[175] ^ in2[175];
    assign G[9] = in[174] & in2[174];
    assign P[9] = in[174] ^ in2[174];
    assign G[10] = in[173] & in2[173];
    assign P[10] = in[173] ^ in2[173];
    assign G[11] = in[172] & in2[172];
    assign P[11] = in[172] ^ in2[172];
    assign G[12] = in[171] & in2[171];
    assign P[12] = in[171] ^ in2[171];
    assign G[13] = in[170] & in2[170];
    assign P[13] = in[170] ^ in2[170];
    assign G[14] = in[169] & in2[169];
    assign P[14] = in[169] ^ in2[169];
    assign G[15] = in[168] & in2[168];
    assign P[15] = in[168] ^ in2[168];
    assign G[16] = in[167] & in2[167];
    assign P[16] = in[167] ^ in2[167];
    assign G[17] = in[166] & in2[166];
    assign P[17] = in[166] ^ in2[166];
    assign G[18] = in[165] & in2[165];
    assign P[18] = in[165] ^ in2[165];
    assign G[19] = in[164] & in2[164];
    assign P[19] = in[164] ^ in2[164];
    assign G[20] = in[163] & in2[163];
    assign P[20] = in[163] ^ in2[163];
    assign G[21] = in[162] & in2[162];
    assign P[21] = in[162] ^ in2[162];
    assign G[22] = in[161] & in2[161];
    assign P[22] = in[161] ^ in2[161];
    assign G[23] = in[160] & in2[160];
    assign P[23] = in[160] ^ in2[160];
    assign G[24] = in[159] & in2[159];
    assign P[24] = in[159] ^ in2[159];
    assign G[25] = in[158] & in2[158];
    assign P[25] = in[158] ^ in2[158];
    assign G[26] = in[157] & in2[157];
    assign P[26] = in[157] ^ in2[157];
    assign G[27] = in[156] & in2[156];
    assign P[27] = in[156] ^ in2[156];
    assign G[28] = in[155] & in2[155];
    assign P[28] = in[155] ^ in2[155];
    assign G[29] = in[154] & in2[154];
    assign P[29] = in[154] ^ in2[154];
    assign G[30] = in[153] & in2[153];
    assign P[30] = in[153] ^ in2[153];
    assign G[31] = in[152] & in2[152];
    assign P[31] = in[152] ^ in2[152];
    assign G[32] = in[151] & in2[151];
    assign P[32] = in[151] ^ in2[151];
    assign G[33] = in[150] & in2[150];
    assign P[33] = in[150] ^ in2[150];
    assign G[34] = in[149] & in2[149];
    assign P[34] = in[149] ^ in2[149];
    assign G[35] = in[148] & in2[148];
    assign P[35] = in[148] ^ in2[148];
    assign G[36] = in[147] & in2[147];
    assign P[36] = in[147] ^ in2[147];
    assign G[37] = in[146] & in2[146];
    assign P[37] = in[146] ^ in2[146];
    assign G[38] = in[145] & in2[145];
    assign P[38] = in[145] ^ in2[145];
    assign G[39] = in[144] & in2[144];
    assign P[39] = in[144] ^ in2[144];
    assign G[40] = in[143] & in2[143];
    assign P[40] = in[143] ^ in2[143];
    assign G[41] = in[142] & in2[142];
    assign P[41] = in[142] ^ in2[142];
    assign G[42] = in[141] & in2[141];
    assign P[42] = in[141] ^ in2[141];
    assign G[43] = in[140] & in2[140];
    assign P[43] = in[140] ^ in2[140];
    assign G[44] = in[139] & in2[139];
    assign P[44] = in[139] ^ in2[139];
    assign G[45] = in[138] & in2[138];
    assign P[45] = in[138] ^ in2[138];
    assign G[46] = in[137] & in2[137];
    assign P[46] = in[137] ^ in2[137];
    assign G[47] = in[136] & in2[136];
    assign P[47] = in[136] ^ in2[136];
    assign G[48] = in[135] & in2[135];
    assign P[48] = in[135] ^ in2[135];
    assign G[49] = in[134] & in2[134];
    assign P[49] = in[134] ^ in2[134];
    assign G[50] = in[133] & in2[133];
    assign P[50] = in[133] ^ in2[133];
    assign G[51] = in[132] & in2[132];
    assign P[51] = in[132] ^ in2[132];
    assign G[52] = in[131] & in2[131];
    assign P[52] = in[131] ^ in2[131];
    assign G[53] = in[130] & in2[130];
    assign P[53] = in[130] ^ in2[130];
    assign G[54] = in[129] & in2[129];
    assign P[54] = in[129] ^ in2[129];
    assign G[55] = in[128] & in2[128];
    assign P[55] = in[128] ^ in2[128];
    assign G[56] = in[127] & in2[127];
    assign P[56] = in[127] ^ in2[127];
    assign G[57] = in[126] & in2[126];
    assign P[57] = in[126] ^ in2[126];
    assign G[58] = in[125] & in2[125];
    assign P[58] = in[125] ^ in2[125];
    assign G[59] = in[124] & in2[124];
    assign P[59] = in[124] ^ in2[124];
    assign G[60] = in[123] & in2[123];
    assign P[60] = in[123] ^ in2[123];
    assign G[61] = in[122] & in2[122];
    assign P[61] = in[122] ^ in2[122];
    assign G[62] = in[121] & in2[121];
    assign P[62] = in[121] ^ in2[121];
    assign G[63] = in[120] & in2[120];
    assign P[63] = in[120] ^ in2[120];
    assign G[64] = in[119] & in2[119];
    assign P[64] = in[119] ^ in2[119];
    assign G[65] = in[118] & in2[118];
    assign P[65] = in[118] ^ in2[118];
    assign G[66] = in[117] & in2[117];
    assign P[66] = in[117] ^ in2[117];
    assign G[67] = in[116] & in2[116];
    assign P[67] = in[116] ^ in2[116];
    assign G[68] = in[115] & in2[115];
    assign P[68] = in[115] ^ in2[115];
    assign G[69] = in[114] & in2[114];
    assign P[69] = in[114] ^ in2[114];
    assign G[70] = in[113] & in2[113];
    assign P[70] = in[113] ^ in2[113];
    assign G[71] = in[112] & in2[112];
    assign P[71] = in[112] ^ in2[112];
    assign G[72] = in[111] & in2[111];
    assign P[72] = in[111] ^ in2[111];
    assign G[73] = in[110] & in2[110];
    assign P[73] = in[110] ^ in2[110];
    assign G[74] = in[109] & in2[109];
    assign P[74] = in[109] ^ in2[109];
    assign G[75] = in[108] & in2[108];
    assign P[75] = in[108] ^ in2[108];
    assign G[76] = in[107] & in2[107];
    assign P[76] = in[107] ^ in2[107];
    assign G[77] = in[106] & in2[106];
    assign P[77] = in[106] ^ in2[106];
    assign G[78] = in[105] & in2[105];
    assign P[78] = in[105] ^ in2[105];
    assign G[79] = in[104] & in2[104];
    assign P[79] = in[104] ^ in2[104];
    assign G[80] = in[103] & in2[103];
    assign P[80] = in[103] ^ in2[103];
    assign G[81] = in[102] & in2[102];
    assign P[81] = in[102] ^ in2[102];
    assign G[82] = in[101] & in2[101];
    assign P[82] = in[101] ^ in2[101];
    assign G[83] = in[100] & in2[100];
    assign P[83] = in[100] ^ in2[100];
    assign G[84] = in[99] & in2[99];
    assign P[84] = in[99] ^ in2[99];
    assign G[85] = in[98] & in2[98];
    assign P[85] = in[98] ^ in2[98];
    assign G[86] = in[97] & in2[97];
    assign P[86] = in[97] ^ in2[97];
    assign G[87] = in[96] & in2[96];
    assign P[87] = in[96] ^ in2[96];
    assign G[88] = in[95] & in2[95];
    assign P[88] = in[95] ^ in2[95];
    assign G[89] = in[94] & in2[94];
    assign P[89] = in[94] ^ in2[94];
    assign G[90] = in[93] & in2[93];
    assign P[90] = in[93] ^ in2[93];
    assign G[91] = in[92] & in2[92];
    assign P[91] = in[92] ^ in2[92];
    assign G[92] = in[91] & in2[91];
    assign P[92] = in[91] ^ in2[91];
    assign G[93] = in[90] & in2[90];
    assign P[93] = in[90] ^ in2[90];
    assign G[94] = in[89] & in2[89];
    assign P[94] = in[89] ^ in2[89];
    assign G[95] = in[88] & in2[88];
    assign P[95] = in[88] ^ in2[88];
    assign G[96] = in[87] & in2[87];
    assign P[96] = in[87] ^ in2[87];
    assign G[97] = in[86] & in2[86];
    assign P[97] = in[86] ^ in2[86];
    assign G[98] = in[85] & in2[85];
    assign P[98] = in[85] ^ in2[85];
    assign G[99] = in[84] & in2[84];
    assign P[99] = in[84] ^ in2[84];
    assign G[100] = in[83] & in2[83];
    assign P[100] = in[83] ^ in2[83];
    assign G[101] = in[82] & in2[82];
    assign P[101] = in[82] ^ in2[82];
    assign G[102] = in[81] & in2[81];
    assign P[102] = in[81] ^ in2[81];
    assign G[103] = in[80] & in2[80];
    assign P[103] = in[80] ^ in2[80];
    assign G[104] = in[79] & in2[79];
    assign P[104] = in[79] ^ in2[79];
    assign G[105] = in[78] & in2[78];
    assign P[105] = in[78] ^ in2[78];
    assign G[106] = in[77] & in2[77];
    assign P[106] = in[77] ^ in2[77];
    assign G[107] = in[76] & in2[76];
    assign P[107] = in[76] ^ in2[76];
    assign G[108] = in[75] & in2[75];
    assign P[108] = in[75] ^ in2[75];
    assign G[109] = in[74] & in2[74];
    assign P[109] = in[74] ^ in2[74];
    assign G[110] = in[73] & in2[73];
    assign P[110] = in[73] ^ in2[73];
    assign G[111] = in[72] & in2[72];
    assign P[111] = in[72] ^ in2[72];
    assign G[112] = in[71] & in2[71];
    assign P[112] = in[71] ^ in2[71];
    assign G[113] = in[70] & in2[70];
    assign P[113] = in[70] ^ in2[70];
    assign G[114] = in[69] & in2[69];
    assign P[114] = in[69] ^ in2[69];
    assign G[115] = in[68] & in2[68];
    assign P[115] = in[68] ^ in2[68];
    assign G[116] = in[67] & in2[67];
    assign P[116] = in[67] ^ in2[67];
    assign G[117] = in[66] & in2[66];
    assign P[117] = in[66] ^ in2[66];
    assign G[118] = in[65] & in2[65];
    assign P[118] = in[65] ^ in2[65];
    assign G[119] = in[64] & in2[64];
    assign P[119] = in[64] ^ in2[64];
    assign G[120] = in[63] & in2[63];
    assign P[120] = in[63] ^ in2[63];
    assign G[121] = in[62] & in2[62];
    assign P[121] = in[62] ^ in2[62];
    assign G[122] = in[61] & in2[61];
    assign P[122] = in[61] ^ in2[61];
    assign G[123] = in[60] & in2[60];
    assign P[123] = in[60] ^ in2[60];
    assign G[124] = in[59] & in2[59];
    assign P[124] = in[59] ^ in2[59];
    assign G[125] = in[58] & in2[58];
    assign P[125] = in[58] ^ in2[58];
    assign G[126] = in[57] & in2[57];
    assign P[126] = in[57] ^ in2[57];
    assign G[127] = in[56] & in2[56];
    assign P[127] = in[56] ^ in2[56];
    assign G[128] = in[55] & in2[55];
    assign P[128] = in[55] ^ in2[55];
    assign G[129] = in[54] & in2[54];
    assign P[129] = in[54] ^ in2[54];
    assign G[130] = in[53] & in2[53];
    assign P[130] = in[53] ^ in2[53];
    assign G[131] = in[52] & in2[52];
    assign P[131] = in[52] ^ in2[52];
    assign G[132] = in[51] & in2[51];
    assign P[132] = in[51] ^ in2[51];
    assign G[133] = in[50] & in2[50];
    assign P[133] = in[50] ^ in2[50];
    assign G[134] = in[49] & in2[49];
    assign P[134] = in[49] ^ in2[49];
    assign G[135] = in[48] & in2[48];
    assign P[135] = in[48] ^ in2[48];
    assign G[136] = in[47] & in2[47];
    assign P[136] = in[47] ^ in2[47];
    assign G[137] = in[46] & in2[46];
    assign P[137] = in[46] ^ in2[46];
    assign G[138] = in[45] & in2[45];
    assign P[138] = in[45] ^ in2[45];
    assign G[139] = in[44] & in2[44];
    assign P[139] = in[44] ^ in2[44];
    assign G[140] = in[43] & in2[43];
    assign P[140] = in[43] ^ in2[43];
    assign G[141] = in[42] & in2[42];
    assign P[141] = in[42] ^ in2[42];
    assign G[142] = in[41] & in2[41];
    assign P[142] = in[41] ^ in2[41];
    assign G[143] = in[40] & in2[40];
    assign P[143] = in[40] ^ in2[40];
    assign G[144] = in[39] & in2[39];
    assign P[144] = in[39] ^ in2[39];
    assign G[145] = in[38] & in2[38];
    assign P[145] = in[38] ^ in2[38];
    assign G[146] = in[37] & in2[37];
    assign P[146] = in[37] ^ in2[37];
    assign G[147] = in[36] & in2[36];
    assign P[147] = in[36] ^ in2[36];
    assign G[148] = in[35] & in2[35];
    assign P[148] = in[35] ^ in2[35];
    assign G[149] = in[34] & in2[34];
    assign P[149] = in[34] ^ in2[34];
    assign G[150] = in[33] & in2[33];
    assign P[150] = in[33] ^ in2[33];
    assign G[151] = in[32] & in2[32];
    assign P[151] = in[32] ^ in2[32];
    assign G[152] = in[31] & in2[31];
    assign P[152] = in[31] ^ in2[31];
    assign G[153] = in[30] & in2[30];
    assign P[153] = in[30] ^ in2[30];
    assign G[154] = in[29] & in2[29];
    assign P[154] = in[29] ^ in2[29];
    assign G[155] = in[28] & in2[28];
    assign P[155] = in[28] ^ in2[28];
    assign G[156] = in[27] & in2[27];
    assign P[156] = in[27] ^ in2[27];
    assign G[157] = in[26] & in2[26];
    assign P[157] = in[26] ^ in2[26];
    assign G[158] = in[25] & in2[25];
    assign P[158] = in[25] ^ in2[25];
    assign G[159] = in[24] & in2[24];
    assign P[159] = in[24] ^ in2[24];
    assign G[160] = in[23] & in2[23];
    assign P[160] = in[23] ^ in2[23];
    assign G[161] = in[22] & in2[22];
    assign P[161] = in[22] ^ in2[22];
    assign G[162] = in[21] & in2[21];
    assign P[162] = in[21] ^ in2[21];
    assign G[163] = in[20] & in2[20];
    assign P[163] = in[20] ^ in2[20];
    assign G[164] = in[19] & in2[19];
    assign P[164] = in[19] ^ in2[19];
    assign G[165] = in[18] & in2[18];
    assign P[165] = in[18] ^ in2[18];
    assign G[166] = in[17] & in2[17];
    assign P[166] = in[17] ^ in2[17];
    assign G[167] = in[16] & in2[16];
    assign P[167] = in[16] ^ in2[16];
    assign G[168] = in[15] & in2[15];
    assign P[168] = in[15] ^ in2[15];
    assign G[169] = in[14] & in2[14];
    assign P[169] = in[14] ^ in2[14];
    assign G[170] = in[13] & in2[13];
    assign P[170] = in[13] ^ in2[13];
    assign G[171] = in[12] & in2[12];
    assign P[171] = in[12] ^ in2[12];
    assign G[172] = in[11] & in2[11];
    assign P[172] = in[11] ^ in2[11];
    assign G[173] = in[10] & in2[10];
    assign P[173] = in[10] ^ in2[10];
    assign G[174] = in[9] & in2[9];
    assign P[174] = in[9] ^ in2[9];
    assign G[175] = in[8] & in2[8];
    assign P[175] = in[8] ^ in2[8];
    assign G[176] = in[7] & in2[7];
    assign P[176] = in[7] ^ in2[7];
    assign G[177] = in[6] & in2[6];
    assign P[177] = in[6] ^ in2[6];
    assign G[178] = in[5] & in2[5];
    assign P[178] = in[5] ^ in2[5];
    assign G[179] = in[4] & in2[4];
    assign P[179] = in[4] ^ in2[4];
    assign G[180] = in[3] & in2[3];
    assign P[180] = in[3] ^ in2[3];
    assign G[181] = in[2] & in2[2];
    assign P[181] = in[2] ^ in2[2];
    assign G[182] = in[1] & in2[1];
    assign P[182] = in[1] ^ in2[1];
    assign G[183] = in[0] & in2[0];
    assign P[183] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign C[183] = G[182] | (P[182] & C[182]);
    assign cout = G[183] | (P[183] & C[183]);
    assign sum = P ^ C;
endmodule

module CLA183(output [182:0] sum, output cout, input [182:0] in1, input [182:0] in2;

    wire[182:0] G;
    wire[182:0] C;
    wire[182:0] P;

    assign G[0] = in[182] & in2[182];
    assign P[0] = in[182] ^ in2[182];
    assign G[1] = in[181] & in2[181];
    assign P[1] = in[181] ^ in2[181];
    assign G[2] = in[180] & in2[180];
    assign P[2] = in[180] ^ in2[180];
    assign G[3] = in[179] & in2[179];
    assign P[3] = in[179] ^ in2[179];
    assign G[4] = in[178] & in2[178];
    assign P[4] = in[178] ^ in2[178];
    assign G[5] = in[177] & in2[177];
    assign P[5] = in[177] ^ in2[177];
    assign G[6] = in[176] & in2[176];
    assign P[6] = in[176] ^ in2[176];
    assign G[7] = in[175] & in2[175];
    assign P[7] = in[175] ^ in2[175];
    assign G[8] = in[174] & in2[174];
    assign P[8] = in[174] ^ in2[174];
    assign G[9] = in[173] & in2[173];
    assign P[9] = in[173] ^ in2[173];
    assign G[10] = in[172] & in2[172];
    assign P[10] = in[172] ^ in2[172];
    assign G[11] = in[171] & in2[171];
    assign P[11] = in[171] ^ in2[171];
    assign G[12] = in[170] & in2[170];
    assign P[12] = in[170] ^ in2[170];
    assign G[13] = in[169] & in2[169];
    assign P[13] = in[169] ^ in2[169];
    assign G[14] = in[168] & in2[168];
    assign P[14] = in[168] ^ in2[168];
    assign G[15] = in[167] & in2[167];
    assign P[15] = in[167] ^ in2[167];
    assign G[16] = in[166] & in2[166];
    assign P[16] = in[166] ^ in2[166];
    assign G[17] = in[165] & in2[165];
    assign P[17] = in[165] ^ in2[165];
    assign G[18] = in[164] & in2[164];
    assign P[18] = in[164] ^ in2[164];
    assign G[19] = in[163] & in2[163];
    assign P[19] = in[163] ^ in2[163];
    assign G[20] = in[162] & in2[162];
    assign P[20] = in[162] ^ in2[162];
    assign G[21] = in[161] & in2[161];
    assign P[21] = in[161] ^ in2[161];
    assign G[22] = in[160] & in2[160];
    assign P[22] = in[160] ^ in2[160];
    assign G[23] = in[159] & in2[159];
    assign P[23] = in[159] ^ in2[159];
    assign G[24] = in[158] & in2[158];
    assign P[24] = in[158] ^ in2[158];
    assign G[25] = in[157] & in2[157];
    assign P[25] = in[157] ^ in2[157];
    assign G[26] = in[156] & in2[156];
    assign P[26] = in[156] ^ in2[156];
    assign G[27] = in[155] & in2[155];
    assign P[27] = in[155] ^ in2[155];
    assign G[28] = in[154] & in2[154];
    assign P[28] = in[154] ^ in2[154];
    assign G[29] = in[153] & in2[153];
    assign P[29] = in[153] ^ in2[153];
    assign G[30] = in[152] & in2[152];
    assign P[30] = in[152] ^ in2[152];
    assign G[31] = in[151] & in2[151];
    assign P[31] = in[151] ^ in2[151];
    assign G[32] = in[150] & in2[150];
    assign P[32] = in[150] ^ in2[150];
    assign G[33] = in[149] & in2[149];
    assign P[33] = in[149] ^ in2[149];
    assign G[34] = in[148] & in2[148];
    assign P[34] = in[148] ^ in2[148];
    assign G[35] = in[147] & in2[147];
    assign P[35] = in[147] ^ in2[147];
    assign G[36] = in[146] & in2[146];
    assign P[36] = in[146] ^ in2[146];
    assign G[37] = in[145] & in2[145];
    assign P[37] = in[145] ^ in2[145];
    assign G[38] = in[144] & in2[144];
    assign P[38] = in[144] ^ in2[144];
    assign G[39] = in[143] & in2[143];
    assign P[39] = in[143] ^ in2[143];
    assign G[40] = in[142] & in2[142];
    assign P[40] = in[142] ^ in2[142];
    assign G[41] = in[141] & in2[141];
    assign P[41] = in[141] ^ in2[141];
    assign G[42] = in[140] & in2[140];
    assign P[42] = in[140] ^ in2[140];
    assign G[43] = in[139] & in2[139];
    assign P[43] = in[139] ^ in2[139];
    assign G[44] = in[138] & in2[138];
    assign P[44] = in[138] ^ in2[138];
    assign G[45] = in[137] & in2[137];
    assign P[45] = in[137] ^ in2[137];
    assign G[46] = in[136] & in2[136];
    assign P[46] = in[136] ^ in2[136];
    assign G[47] = in[135] & in2[135];
    assign P[47] = in[135] ^ in2[135];
    assign G[48] = in[134] & in2[134];
    assign P[48] = in[134] ^ in2[134];
    assign G[49] = in[133] & in2[133];
    assign P[49] = in[133] ^ in2[133];
    assign G[50] = in[132] & in2[132];
    assign P[50] = in[132] ^ in2[132];
    assign G[51] = in[131] & in2[131];
    assign P[51] = in[131] ^ in2[131];
    assign G[52] = in[130] & in2[130];
    assign P[52] = in[130] ^ in2[130];
    assign G[53] = in[129] & in2[129];
    assign P[53] = in[129] ^ in2[129];
    assign G[54] = in[128] & in2[128];
    assign P[54] = in[128] ^ in2[128];
    assign G[55] = in[127] & in2[127];
    assign P[55] = in[127] ^ in2[127];
    assign G[56] = in[126] & in2[126];
    assign P[56] = in[126] ^ in2[126];
    assign G[57] = in[125] & in2[125];
    assign P[57] = in[125] ^ in2[125];
    assign G[58] = in[124] & in2[124];
    assign P[58] = in[124] ^ in2[124];
    assign G[59] = in[123] & in2[123];
    assign P[59] = in[123] ^ in2[123];
    assign G[60] = in[122] & in2[122];
    assign P[60] = in[122] ^ in2[122];
    assign G[61] = in[121] & in2[121];
    assign P[61] = in[121] ^ in2[121];
    assign G[62] = in[120] & in2[120];
    assign P[62] = in[120] ^ in2[120];
    assign G[63] = in[119] & in2[119];
    assign P[63] = in[119] ^ in2[119];
    assign G[64] = in[118] & in2[118];
    assign P[64] = in[118] ^ in2[118];
    assign G[65] = in[117] & in2[117];
    assign P[65] = in[117] ^ in2[117];
    assign G[66] = in[116] & in2[116];
    assign P[66] = in[116] ^ in2[116];
    assign G[67] = in[115] & in2[115];
    assign P[67] = in[115] ^ in2[115];
    assign G[68] = in[114] & in2[114];
    assign P[68] = in[114] ^ in2[114];
    assign G[69] = in[113] & in2[113];
    assign P[69] = in[113] ^ in2[113];
    assign G[70] = in[112] & in2[112];
    assign P[70] = in[112] ^ in2[112];
    assign G[71] = in[111] & in2[111];
    assign P[71] = in[111] ^ in2[111];
    assign G[72] = in[110] & in2[110];
    assign P[72] = in[110] ^ in2[110];
    assign G[73] = in[109] & in2[109];
    assign P[73] = in[109] ^ in2[109];
    assign G[74] = in[108] & in2[108];
    assign P[74] = in[108] ^ in2[108];
    assign G[75] = in[107] & in2[107];
    assign P[75] = in[107] ^ in2[107];
    assign G[76] = in[106] & in2[106];
    assign P[76] = in[106] ^ in2[106];
    assign G[77] = in[105] & in2[105];
    assign P[77] = in[105] ^ in2[105];
    assign G[78] = in[104] & in2[104];
    assign P[78] = in[104] ^ in2[104];
    assign G[79] = in[103] & in2[103];
    assign P[79] = in[103] ^ in2[103];
    assign G[80] = in[102] & in2[102];
    assign P[80] = in[102] ^ in2[102];
    assign G[81] = in[101] & in2[101];
    assign P[81] = in[101] ^ in2[101];
    assign G[82] = in[100] & in2[100];
    assign P[82] = in[100] ^ in2[100];
    assign G[83] = in[99] & in2[99];
    assign P[83] = in[99] ^ in2[99];
    assign G[84] = in[98] & in2[98];
    assign P[84] = in[98] ^ in2[98];
    assign G[85] = in[97] & in2[97];
    assign P[85] = in[97] ^ in2[97];
    assign G[86] = in[96] & in2[96];
    assign P[86] = in[96] ^ in2[96];
    assign G[87] = in[95] & in2[95];
    assign P[87] = in[95] ^ in2[95];
    assign G[88] = in[94] & in2[94];
    assign P[88] = in[94] ^ in2[94];
    assign G[89] = in[93] & in2[93];
    assign P[89] = in[93] ^ in2[93];
    assign G[90] = in[92] & in2[92];
    assign P[90] = in[92] ^ in2[92];
    assign G[91] = in[91] & in2[91];
    assign P[91] = in[91] ^ in2[91];
    assign G[92] = in[90] & in2[90];
    assign P[92] = in[90] ^ in2[90];
    assign G[93] = in[89] & in2[89];
    assign P[93] = in[89] ^ in2[89];
    assign G[94] = in[88] & in2[88];
    assign P[94] = in[88] ^ in2[88];
    assign G[95] = in[87] & in2[87];
    assign P[95] = in[87] ^ in2[87];
    assign G[96] = in[86] & in2[86];
    assign P[96] = in[86] ^ in2[86];
    assign G[97] = in[85] & in2[85];
    assign P[97] = in[85] ^ in2[85];
    assign G[98] = in[84] & in2[84];
    assign P[98] = in[84] ^ in2[84];
    assign G[99] = in[83] & in2[83];
    assign P[99] = in[83] ^ in2[83];
    assign G[100] = in[82] & in2[82];
    assign P[100] = in[82] ^ in2[82];
    assign G[101] = in[81] & in2[81];
    assign P[101] = in[81] ^ in2[81];
    assign G[102] = in[80] & in2[80];
    assign P[102] = in[80] ^ in2[80];
    assign G[103] = in[79] & in2[79];
    assign P[103] = in[79] ^ in2[79];
    assign G[104] = in[78] & in2[78];
    assign P[104] = in[78] ^ in2[78];
    assign G[105] = in[77] & in2[77];
    assign P[105] = in[77] ^ in2[77];
    assign G[106] = in[76] & in2[76];
    assign P[106] = in[76] ^ in2[76];
    assign G[107] = in[75] & in2[75];
    assign P[107] = in[75] ^ in2[75];
    assign G[108] = in[74] & in2[74];
    assign P[108] = in[74] ^ in2[74];
    assign G[109] = in[73] & in2[73];
    assign P[109] = in[73] ^ in2[73];
    assign G[110] = in[72] & in2[72];
    assign P[110] = in[72] ^ in2[72];
    assign G[111] = in[71] & in2[71];
    assign P[111] = in[71] ^ in2[71];
    assign G[112] = in[70] & in2[70];
    assign P[112] = in[70] ^ in2[70];
    assign G[113] = in[69] & in2[69];
    assign P[113] = in[69] ^ in2[69];
    assign G[114] = in[68] & in2[68];
    assign P[114] = in[68] ^ in2[68];
    assign G[115] = in[67] & in2[67];
    assign P[115] = in[67] ^ in2[67];
    assign G[116] = in[66] & in2[66];
    assign P[116] = in[66] ^ in2[66];
    assign G[117] = in[65] & in2[65];
    assign P[117] = in[65] ^ in2[65];
    assign G[118] = in[64] & in2[64];
    assign P[118] = in[64] ^ in2[64];
    assign G[119] = in[63] & in2[63];
    assign P[119] = in[63] ^ in2[63];
    assign G[120] = in[62] & in2[62];
    assign P[120] = in[62] ^ in2[62];
    assign G[121] = in[61] & in2[61];
    assign P[121] = in[61] ^ in2[61];
    assign G[122] = in[60] & in2[60];
    assign P[122] = in[60] ^ in2[60];
    assign G[123] = in[59] & in2[59];
    assign P[123] = in[59] ^ in2[59];
    assign G[124] = in[58] & in2[58];
    assign P[124] = in[58] ^ in2[58];
    assign G[125] = in[57] & in2[57];
    assign P[125] = in[57] ^ in2[57];
    assign G[126] = in[56] & in2[56];
    assign P[126] = in[56] ^ in2[56];
    assign G[127] = in[55] & in2[55];
    assign P[127] = in[55] ^ in2[55];
    assign G[128] = in[54] & in2[54];
    assign P[128] = in[54] ^ in2[54];
    assign G[129] = in[53] & in2[53];
    assign P[129] = in[53] ^ in2[53];
    assign G[130] = in[52] & in2[52];
    assign P[130] = in[52] ^ in2[52];
    assign G[131] = in[51] & in2[51];
    assign P[131] = in[51] ^ in2[51];
    assign G[132] = in[50] & in2[50];
    assign P[132] = in[50] ^ in2[50];
    assign G[133] = in[49] & in2[49];
    assign P[133] = in[49] ^ in2[49];
    assign G[134] = in[48] & in2[48];
    assign P[134] = in[48] ^ in2[48];
    assign G[135] = in[47] & in2[47];
    assign P[135] = in[47] ^ in2[47];
    assign G[136] = in[46] & in2[46];
    assign P[136] = in[46] ^ in2[46];
    assign G[137] = in[45] & in2[45];
    assign P[137] = in[45] ^ in2[45];
    assign G[138] = in[44] & in2[44];
    assign P[138] = in[44] ^ in2[44];
    assign G[139] = in[43] & in2[43];
    assign P[139] = in[43] ^ in2[43];
    assign G[140] = in[42] & in2[42];
    assign P[140] = in[42] ^ in2[42];
    assign G[141] = in[41] & in2[41];
    assign P[141] = in[41] ^ in2[41];
    assign G[142] = in[40] & in2[40];
    assign P[142] = in[40] ^ in2[40];
    assign G[143] = in[39] & in2[39];
    assign P[143] = in[39] ^ in2[39];
    assign G[144] = in[38] & in2[38];
    assign P[144] = in[38] ^ in2[38];
    assign G[145] = in[37] & in2[37];
    assign P[145] = in[37] ^ in2[37];
    assign G[146] = in[36] & in2[36];
    assign P[146] = in[36] ^ in2[36];
    assign G[147] = in[35] & in2[35];
    assign P[147] = in[35] ^ in2[35];
    assign G[148] = in[34] & in2[34];
    assign P[148] = in[34] ^ in2[34];
    assign G[149] = in[33] & in2[33];
    assign P[149] = in[33] ^ in2[33];
    assign G[150] = in[32] & in2[32];
    assign P[150] = in[32] ^ in2[32];
    assign G[151] = in[31] & in2[31];
    assign P[151] = in[31] ^ in2[31];
    assign G[152] = in[30] & in2[30];
    assign P[152] = in[30] ^ in2[30];
    assign G[153] = in[29] & in2[29];
    assign P[153] = in[29] ^ in2[29];
    assign G[154] = in[28] & in2[28];
    assign P[154] = in[28] ^ in2[28];
    assign G[155] = in[27] & in2[27];
    assign P[155] = in[27] ^ in2[27];
    assign G[156] = in[26] & in2[26];
    assign P[156] = in[26] ^ in2[26];
    assign G[157] = in[25] & in2[25];
    assign P[157] = in[25] ^ in2[25];
    assign G[158] = in[24] & in2[24];
    assign P[158] = in[24] ^ in2[24];
    assign G[159] = in[23] & in2[23];
    assign P[159] = in[23] ^ in2[23];
    assign G[160] = in[22] & in2[22];
    assign P[160] = in[22] ^ in2[22];
    assign G[161] = in[21] & in2[21];
    assign P[161] = in[21] ^ in2[21];
    assign G[162] = in[20] & in2[20];
    assign P[162] = in[20] ^ in2[20];
    assign G[163] = in[19] & in2[19];
    assign P[163] = in[19] ^ in2[19];
    assign G[164] = in[18] & in2[18];
    assign P[164] = in[18] ^ in2[18];
    assign G[165] = in[17] & in2[17];
    assign P[165] = in[17] ^ in2[17];
    assign G[166] = in[16] & in2[16];
    assign P[166] = in[16] ^ in2[16];
    assign G[167] = in[15] & in2[15];
    assign P[167] = in[15] ^ in2[15];
    assign G[168] = in[14] & in2[14];
    assign P[168] = in[14] ^ in2[14];
    assign G[169] = in[13] & in2[13];
    assign P[169] = in[13] ^ in2[13];
    assign G[170] = in[12] & in2[12];
    assign P[170] = in[12] ^ in2[12];
    assign G[171] = in[11] & in2[11];
    assign P[171] = in[11] ^ in2[11];
    assign G[172] = in[10] & in2[10];
    assign P[172] = in[10] ^ in2[10];
    assign G[173] = in[9] & in2[9];
    assign P[173] = in[9] ^ in2[9];
    assign G[174] = in[8] & in2[8];
    assign P[174] = in[8] ^ in2[8];
    assign G[175] = in[7] & in2[7];
    assign P[175] = in[7] ^ in2[7];
    assign G[176] = in[6] & in2[6];
    assign P[176] = in[6] ^ in2[6];
    assign G[177] = in[5] & in2[5];
    assign P[177] = in[5] ^ in2[5];
    assign G[178] = in[4] & in2[4];
    assign P[178] = in[4] ^ in2[4];
    assign G[179] = in[3] & in2[3];
    assign P[179] = in[3] ^ in2[3];
    assign G[180] = in[2] & in2[2];
    assign P[180] = in[2] ^ in2[2];
    assign G[181] = in[1] & in2[1];
    assign P[181] = in[1] ^ in2[1];
    assign G[182] = in[0] & in2[0];
    assign P[182] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign C[182] = G[181] | (P[181] & C[181]);
    assign cout = G[182] | (P[182] & C[182]);
    assign sum = P ^ C;
endmodule

module CLA182(output [181:0] sum, output cout, input [181:0] in1, input [181:0] in2;

    wire[181:0] G;
    wire[181:0] C;
    wire[181:0] P;

    assign G[0] = in[181] & in2[181];
    assign P[0] = in[181] ^ in2[181];
    assign G[1] = in[180] & in2[180];
    assign P[1] = in[180] ^ in2[180];
    assign G[2] = in[179] & in2[179];
    assign P[2] = in[179] ^ in2[179];
    assign G[3] = in[178] & in2[178];
    assign P[3] = in[178] ^ in2[178];
    assign G[4] = in[177] & in2[177];
    assign P[4] = in[177] ^ in2[177];
    assign G[5] = in[176] & in2[176];
    assign P[5] = in[176] ^ in2[176];
    assign G[6] = in[175] & in2[175];
    assign P[6] = in[175] ^ in2[175];
    assign G[7] = in[174] & in2[174];
    assign P[7] = in[174] ^ in2[174];
    assign G[8] = in[173] & in2[173];
    assign P[8] = in[173] ^ in2[173];
    assign G[9] = in[172] & in2[172];
    assign P[9] = in[172] ^ in2[172];
    assign G[10] = in[171] & in2[171];
    assign P[10] = in[171] ^ in2[171];
    assign G[11] = in[170] & in2[170];
    assign P[11] = in[170] ^ in2[170];
    assign G[12] = in[169] & in2[169];
    assign P[12] = in[169] ^ in2[169];
    assign G[13] = in[168] & in2[168];
    assign P[13] = in[168] ^ in2[168];
    assign G[14] = in[167] & in2[167];
    assign P[14] = in[167] ^ in2[167];
    assign G[15] = in[166] & in2[166];
    assign P[15] = in[166] ^ in2[166];
    assign G[16] = in[165] & in2[165];
    assign P[16] = in[165] ^ in2[165];
    assign G[17] = in[164] & in2[164];
    assign P[17] = in[164] ^ in2[164];
    assign G[18] = in[163] & in2[163];
    assign P[18] = in[163] ^ in2[163];
    assign G[19] = in[162] & in2[162];
    assign P[19] = in[162] ^ in2[162];
    assign G[20] = in[161] & in2[161];
    assign P[20] = in[161] ^ in2[161];
    assign G[21] = in[160] & in2[160];
    assign P[21] = in[160] ^ in2[160];
    assign G[22] = in[159] & in2[159];
    assign P[22] = in[159] ^ in2[159];
    assign G[23] = in[158] & in2[158];
    assign P[23] = in[158] ^ in2[158];
    assign G[24] = in[157] & in2[157];
    assign P[24] = in[157] ^ in2[157];
    assign G[25] = in[156] & in2[156];
    assign P[25] = in[156] ^ in2[156];
    assign G[26] = in[155] & in2[155];
    assign P[26] = in[155] ^ in2[155];
    assign G[27] = in[154] & in2[154];
    assign P[27] = in[154] ^ in2[154];
    assign G[28] = in[153] & in2[153];
    assign P[28] = in[153] ^ in2[153];
    assign G[29] = in[152] & in2[152];
    assign P[29] = in[152] ^ in2[152];
    assign G[30] = in[151] & in2[151];
    assign P[30] = in[151] ^ in2[151];
    assign G[31] = in[150] & in2[150];
    assign P[31] = in[150] ^ in2[150];
    assign G[32] = in[149] & in2[149];
    assign P[32] = in[149] ^ in2[149];
    assign G[33] = in[148] & in2[148];
    assign P[33] = in[148] ^ in2[148];
    assign G[34] = in[147] & in2[147];
    assign P[34] = in[147] ^ in2[147];
    assign G[35] = in[146] & in2[146];
    assign P[35] = in[146] ^ in2[146];
    assign G[36] = in[145] & in2[145];
    assign P[36] = in[145] ^ in2[145];
    assign G[37] = in[144] & in2[144];
    assign P[37] = in[144] ^ in2[144];
    assign G[38] = in[143] & in2[143];
    assign P[38] = in[143] ^ in2[143];
    assign G[39] = in[142] & in2[142];
    assign P[39] = in[142] ^ in2[142];
    assign G[40] = in[141] & in2[141];
    assign P[40] = in[141] ^ in2[141];
    assign G[41] = in[140] & in2[140];
    assign P[41] = in[140] ^ in2[140];
    assign G[42] = in[139] & in2[139];
    assign P[42] = in[139] ^ in2[139];
    assign G[43] = in[138] & in2[138];
    assign P[43] = in[138] ^ in2[138];
    assign G[44] = in[137] & in2[137];
    assign P[44] = in[137] ^ in2[137];
    assign G[45] = in[136] & in2[136];
    assign P[45] = in[136] ^ in2[136];
    assign G[46] = in[135] & in2[135];
    assign P[46] = in[135] ^ in2[135];
    assign G[47] = in[134] & in2[134];
    assign P[47] = in[134] ^ in2[134];
    assign G[48] = in[133] & in2[133];
    assign P[48] = in[133] ^ in2[133];
    assign G[49] = in[132] & in2[132];
    assign P[49] = in[132] ^ in2[132];
    assign G[50] = in[131] & in2[131];
    assign P[50] = in[131] ^ in2[131];
    assign G[51] = in[130] & in2[130];
    assign P[51] = in[130] ^ in2[130];
    assign G[52] = in[129] & in2[129];
    assign P[52] = in[129] ^ in2[129];
    assign G[53] = in[128] & in2[128];
    assign P[53] = in[128] ^ in2[128];
    assign G[54] = in[127] & in2[127];
    assign P[54] = in[127] ^ in2[127];
    assign G[55] = in[126] & in2[126];
    assign P[55] = in[126] ^ in2[126];
    assign G[56] = in[125] & in2[125];
    assign P[56] = in[125] ^ in2[125];
    assign G[57] = in[124] & in2[124];
    assign P[57] = in[124] ^ in2[124];
    assign G[58] = in[123] & in2[123];
    assign P[58] = in[123] ^ in2[123];
    assign G[59] = in[122] & in2[122];
    assign P[59] = in[122] ^ in2[122];
    assign G[60] = in[121] & in2[121];
    assign P[60] = in[121] ^ in2[121];
    assign G[61] = in[120] & in2[120];
    assign P[61] = in[120] ^ in2[120];
    assign G[62] = in[119] & in2[119];
    assign P[62] = in[119] ^ in2[119];
    assign G[63] = in[118] & in2[118];
    assign P[63] = in[118] ^ in2[118];
    assign G[64] = in[117] & in2[117];
    assign P[64] = in[117] ^ in2[117];
    assign G[65] = in[116] & in2[116];
    assign P[65] = in[116] ^ in2[116];
    assign G[66] = in[115] & in2[115];
    assign P[66] = in[115] ^ in2[115];
    assign G[67] = in[114] & in2[114];
    assign P[67] = in[114] ^ in2[114];
    assign G[68] = in[113] & in2[113];
    assign P[68] = in[113] ^ in2[113];
    assign G[69] = in[112] & in2[112];
    assign P[69] = in[112] ^ in2[112];
    assign G[70] = in[111] & in2[111];
    assign P[70] = in[111] ^ in2[111];
    assign G[71] = in[110] & in2[110];
    assign P[71] = in[110] ^ in2[110];
    assign G[72] = in[109] & in2[109];
    assign P[72] = in[109] ^ in2[109];
    assign G[73] = in[108] & in2[108];
    assign P[73] = in[108] ^ in2[108];
    assign G[74] = in[107] & in2[107];
    assign P[74] = in[107] ^ in2[107];
    assign G[75] = in[106] & in2[106];
    assign P[75] = in[106] ^ in2[106];
    assign G[76] = in[105] & in2[105];
    assign P[76] = in[105] ^ in2[105];
    assign G[77] = in[104] & in2[104];
    assign P[77] = in[104] ^ in2[104];
    assign G[78] = in[103] & in2[103];
    assign P[78] = in[103] ^ in2[103];
    assign G[79] = in[102] & in2[102];
    assign P[79] = in[102] ^ in2[102];
    assign G[80] = in[101] & in2[101];
    assign P[80] = in[101] ^ in2[101];
    assign G[81] = in[100] & in2[100];
    assign P[81] = in[100] ^ in2[100];
    assign G[82] = in[99] & in2[99];
    assign P[82] = in[99] ^ in2[99];
    assign G[83] = in[98] & in2[98];
    assign P[83] = in[98] ^ in2[98];
    assign G[84] = in[97] & in2[97];
    assign P[84] = in[97] ^ in2[97];
    assign G[85] = in[96] & in2[96];
    assign P[85] = in[96] ^ in2[96];
    assign G[86] = in[95] & in2[95];
    assign P[86] = in[95] ^ in2[95];
    assign G[87] = in[94] & in2[94];
    assign P[87] = in[94] ^ in2[94];
    assign G[88] = in[93] & in2[93];
    assign P[88] = in[93] ^ in2[93];
    assign G[89] = in[92] & in2[92];
    assign P[89] = in[92] ^ in2[92];
    assign G[90] = in[91] & in2[91];
    assign P[90] = in[91] ^ in2[91];
    assign G[91] = in[90] & in2[90];
    assign P[91] = in[90] ^ in2[90];
    assign G[92] = in[89] & in2[89];
    assign P[92] = in[89] ^ in2[89];
    assign G[93] = in[88] & in2[88];
    assign P[93] = in[88] ^ in2[88];
    assign G[94] = in[87] & in2[87];
    assign P[94] = in[87] ^ in2[87];
    assign G[95] = in[86] & in2[86];
    assign P[95] = in[86] ^ in2[86];
    assign G[96] = in[85] & in2[85];
    assign P[96] = in[85] ^ in2[85];
    assign G[97] = in[84] & in2[84];
    assign P[97] = in[84] ^ in2[84];
    assign G[98] = in[83] & in2[83];
    assign P[98] = in[83] ^ in2[83];
    assign G[99] = in[82] & in2[82];
    assign P[99] = in[82] ^ in2[82];
    assign G[100] = in[81] & in2[81];
    assign P[100] = in[81] ^ in2[81];
    assign G[101] = in[80] & in2[80];
    assign P[101] = in[80] ^ in2[80];
    assign G[102] = in[79] & in2[79];
    assign P[102] = in[79] ^ in2[79];
    assign G[103] = in[78] & in2[78];
    assign P[103] = in[78] ^ in2[78];
    assign G[104] = in[77] & in2[77];
    assign P[104] = in[77] ^ in2[77];
    assign G[105] = in[76] & in2[76];
    assign P[105] = in[76] ^ in2[76];
    assign G[106] = in[75] & in2[75];
    assign P[106] = in[75] ^ in2[75];
    assign G[107] = in[74] & in2[74];
    assign P[107] = in[74] ^ in2[74];
    assign G[108] = in[73] & in2[73];
    assign P[108] = in[73] ^ in2[73];
    assign G[109] = in[72] & in2[72];
    assign P[109] = in[72] ^ in2[72];
    assign G[110] = in[71] & in2[71];
    assign P[110] = in[71] ^ in2[71];
    assign G[111] = in[70] & in2[70];
    assign P[111] = in[70] ^ in2[70];
    assign G[112] = in[69] & in2[69];
    assign P[112] = in[69] ^ in2[69];
    assign G[113] = in[68] & in2[68];
    assign P[113] = in[68] ^ in2[68];
    assign G[114] = in[67] & in2[67];
    assign P[114] = in[67] ^ in2[67];
    assign G[115] = in[66] & in2[66];
    assign P[115] = in[66] ^ in2[66];
    assign G[116] = in[65] & in2[65];
    assign P[116] = in[65] ^ in2[65];
    assign G[117] = in[64] & in2[64];
    assign P[117] = in[64] ^ in2[64];
    assign G[118] = in[63] & in2[63];
    assign P[118] = in[63] ^ in2[63];
    assign G[119] = in[62] & in2[62];
    assign P[119] = in[62] ^ in2[62];
    assign G[120] = in[61] & in2[61];
    assign P[120] = in[61] ^ in2[61];
    assign G[121] = in[60] & in2[60];
    assign P[121] = in[60] ^ in2[60];
    assign G[122] = in[59] & in2[59];
    assign P[122] = in[59] ^ in2[59];
    assign G[123] = in[58] & in2[58];
    assign P[123] = in[58] ^ in2[58];
    assign G[124] = in[57] & in2[57];
    assign P[124] = in[57] ^ in2[57];
    assign G[125] = in[56] & in2[56];
    assign P[125] = in[56] ^ in2[56];
    assign G[126] = in[55] & in2[55];
    assign P[126] = in[55] ^ in2[55];
    assign G[127] = in[54] & in2[54];
    assign P[127] = in[54] ^ in2[54];
    assign G[128] = in[53] & in2[53];
    assign P[128] = in[53] ^ in2[53];
    assign G[129] = in[52] & in2[52];
    assign P[129] = in[52] ^ in2[52];
    assign G[130] = in[51] & in2[51];
    assign P[130] = in[51] ^ in2[51];
    assign G[131] = in[50] & in2[50];
    assign P[131] = in[50] ^ in2[50];
    assign G[132] = in[49] & in2[49];
    assign P[132] = in[49] ^ in2[49];
    assign G[133] = in[48] & in2[48];
    assign P[133] = in[48] ^ in2[48];
    assign G[134] = in[47] & in2[47];
    assign P[134] = in[47] ^ in2[47];
    assign G[135] = in[46] & in2[46];
    assign P[135] = in[46] ^ in2[46];
    assign G[136] = in[45] & in2[45];
    assign P[136] = in[45] ^ in2[45];
    assign G[137] = in[44] & in2[44];
    assign P[137] = in[44] ^ in2[44];
    assign G[138] = in[43] & in2[43];
    assign P[138] = in[43] ^ in2[43];
    assign G[139] = in[42] & in2[42];
    assign P[139] = in[42] ^ in2[42];
    assign G[140] = in[41] & in2[41];
    assign P[140] = in[41] ^ in2[41];
    assign G[141] = in[40] & in2[40];
    assign P[141] = in[40] ^ in2[40];
    assign G[142] = in[39] & in2[39];
    assign P[142] = in[39] ^ in2[39];
    assign G[143] = in[38] & in2[38];
    assign P[143] = in[38] ^ in2[38];
    assign G[144] = in[37] & in2[37];
    assign P[144] = in[37] ^ in2[37];
    assign G[145] = in[36] & in2[36];
    assign P[145] = in[36] ^ in2[36];
    assign G[146] = in[35] & in2[35];
    assign P[146] = in[35] ^ in2[35];
    assign G[147] = in[34] & in2[34];
    assign P[147] = in[34] ^ in2[34];
    assign G[148] = in[33] & in2[33];
    assign P[148] = in[33] ^ in2[33];
    assign G[149] = in[32] & in2[32];
    assign P[149] = in[32] ^ in2[32];
    assign G[150] = in[31] & in2[31];
    assign P[150] = in[31] ^ in2[31];
    assign G[151] = in[30] & in2[30];
    assign P[151] = in[30] ^ in2[30];
    assign G[152] = in[29] & in2[29];
    assign P[152] = in[29] ^ in2[29];
    assign G[153] = in[28] & in2[28];
    assign P[153] = in[28] ^ in2[28];
    assign G[154] = in[27] & in2[27];
    assign P[154] = in[27] ^ in2[27];
    assign G[155] = in[26] & in2[26];
    assign P[155] = in[26] ^ in2[26];
    assign G[156] = in[25] & in2[25];
    assign P[156] = in[25] ^ in2[25];
    assign G[157] = in[24] & in2[24];
    assign P[157] = in[24] ^ in2[24];
    assign G[158] = in[23] & in2[23];
    assign P[158] = in[23] ^ in2[23];
    assign G[159] = in[22] & in2[22];
    assign P[159] = in[22] ^ in2[22];
    assign G[160] = in[21] & in2[21];
    assign P[160] = in[21] ^ in2[21];
    assign G[161] = in[20] & in2[20];
    assign P[161] = in[20] ^ in2[20];
    assign G[162] = in[19] & in2[19];
    assign P[162] = in[19] ^ in2[19];
    assign G[163] = in[18] & in2[18];
    assign P[163] = in[18] ^ in2[18];
    assign G[164] = in[17] & in2[17];
    assign P[164] = in[17] ^ in2[17];
    assign G[165] = in[16] & in2[16];
    assign P[165] = in[16] ^ in2[16];
    assign G[166] = in[15] & in2[15];
    assign P[166] = in[15] ^ in2[15];
    assign G[167] = in[14] & in2[14];
    assign P[167] = in[14] ^ in2[14];
    assign G[168] = in[13] & in2[13];
    assign P[168] = in[13] ^ in2[13];
    assign G[169] = in[12] & in2[12];
    assign P[169] = in[12] ^ in2[12];
    assign G[170] = in[11] & in2[11];
    assign P[170] = in[11] ^ in2[11];
    assign G[171] = in[10] & in2[10];
    assign P[171] = in[10] ^ in2[10];
    assign G[172] = in[9] & in2[9];
    assign P[172] = in[9] ^ in2[9];
    assign G[173] = in[8] & in2[8];
    assign P[173] = in[8] ^ in2[8];
    assign G[174] = in[7] & in2[7];
    assign P[174] = in[7] ^ in2[7];
    assign G[175] = in[6] & in2[6];
    assign P[175] = in[6] ^ in2[6];
    assign G[176] = in[5] & in2[5];
    assign P[176] = in[5] ^ in2[5];
    assign G[177] = in[4] & in2[4];
    assign P[177] = in[4] ^ in2[4];
    assign G[178] = in[3] & in2[3];
    assign P[178] = in[3] ^ in2[3];
    assign G[179] = in[2] & in2[2];
    assign P[179] = in[2] ^ in2[2];
    assign G[180] = in[1] & in2[1];
    assign P[180] = in[1] ^ in2[1];
    assign G[181] = in[0] & in2[0];
    assign P[181] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign C[181] = G[180] | (P[180] & C[180]);
    assign cout = G[181] | (P[181] & C[181]);
    assign sum = P ^ C;
endmodule

module CLA181(output [180:0] sum, output cout, input [180:0] in1, input [180:0] in2;

    wire[180:0] G;
    wire[180:0] C;
    wire[180:0] P;

    assign G[0] = in[180] & in2[180];
    assign P[0] = in[180] ^ in2[180];
    assign G[1] = in[179] & in2[179];
    assign P[1] = in[179] ^ in2[179];
    assign G[2] = in[178] & in2[178];
    assign P[2] = in[178] ^ in2[178];
    assign G[3] = in[177] & in2[177];
    assign P[3] = in[177] ^ in2[177];
    assign G[4] = in[176] & in2[176];
    assign P[4] = in[176] ^ in2[176];
    assign G[5] = in[175] & in2[175];
    assign P[5] = in[175] ^ in2[175];
    assign G[6] = in[174] & in2[174];
    assign P[6] = in[174] ^ in2[174];
    assign G[7] = in[173] & in2[173];
    assign P[7] = in[173] ^ in2[173];
    assign G[8] = in[172] & in2[172];
    assign P[8] = in[172] ^ in2[172];
    assign G[9] = in[171] & in2[171];
    assign P[9] = in[171] ^ in2[171];
    assign G[10] = in[170] & in2[170];
    assign P[10] = in[170] ^ in2[170];
    assign G[11] = in[169] & in2[169];
    assign P[11] = in[169] ^ in2[169];
    assign G[12] = in[168] & in2[168];
    assign P[12] = in[168] ^ in2[168];
    assign G[13] = in[167] & in2[167];
    assign P[13] = in[167] ^ in2[167];
    assign G[14] = in[166] & in2[166];
    assign P[14] = in[166] ^ in2[166];
    assign G[15] = in[165] & in2[165];
    assign P[15] = in[165] ^ in2[165];
    assign G[16] = in[164] & in2[164];
    assign P[16] = in[164] ^ in2[164];
    assign G[17] = in[163] & in2[163];
    assign P[17] = in[163] ^ in2[163];
    assign G[18] = in[162] & in2[162];
    assign P[18] = in[162] ^ in2[162];
    assign G[19] = in[161] & in2[161];
    assign P[19] = in[161] ^ in2[161];
    assign G[20] = in[160] & in2[160];
    assign P[20] = in[160] ^ in2[160];
    assign G[21] = in[159] & in2[159];
    assign P[21] = in[159] ^ in2[159];
    assign G[22] = in[158] & in2[158];
    assign P[22] = in[158] ^ in2[158];
    assign G[23] = in[157] & in2[157];
    assign P[23] = in[157] ^ in2[157];
    assign G[24] = in[156] & in2[156];
    assign P[24] = in[156] ^ in2[156];
    assign G[25] = in[155] & in2[155];
    assign P[25] = in[155] ^ in2[155];
    assign G[26] = in[154] & in2[154];
    assign P[26] = in[154] ^ in2[154];
    assign G[27] = in[153] & in2[153];
    assign P[27] = in[153] ^ in2[153];
    assign G[28] = in[152] & in2[152];
    assign P[28] = in[152] ^ in2[152];
    assign G[29] = in[151] & in2[151];
    assign P[29] = in[151] ^ in2[151];
    assign G[30] = in[150] & in2[150];
    assign P[30] = in[150] ^ in2[150];
    assign G[31] = in[149] & in2[149];
    assign P[31] = in[149] ^ in2[149];
    assign G[32] = in[148] & in2[148];
    assign P[32] = in[148] ^ in2[148];
    assign G[33] = in[147] & in2[147];
    assign P[33] = in[147] ^ in2[147];
    assign G[34] = in[146] & in2[146];
    assign P[34] = in[146] ^ in2[146];
    assign G[35] = in[145] & in2[145];
    assign P[35] = in[145] ^ in2[145];
    assign G[36] = in[144] & in2[144];
    assign P[36] = in[144] ^ in2[144];
    assign G[37] = in[143] & in2[143];
    assign P[37] = in[143] ^ in2[143];
    assign G[38] = in[142] & in2[142];
    assign P[38] = in[142] ^ in2[142];
    assign G[39] = in[141] & in2[141];
    assign P[39] = in[141] ^ in2[141];
    assign G[40] = in[140] & in2[140];
    assign P[40] = in[140] ^ in2[140];
    assign G[41] = in[139] & in2[139];
    assign P[41] = in[139] ^ in2[139];
    assign G[42] = in[138] & in2[138];
    assign P[42] = in[138] ^ in2[138];
    assign G[43] = in[137] & in2[137];
    assign P[43] = in[137] ^ in2[137];
    assign G[44] = in[136] & in2[136];
    assign P[44] = in[136] ^ in2[136];
    assign G[45] = in[135] & in2[135];
    assign P[45] = in[135] ^ in2[135];
    assign G[46] = in[134] & in2[134];
    assign P[46] = in[134] ^ in2[134];
    assign G[47] = in[133] & in2[133];
    assign P[47] = in[133] ^ in2[133];
    assign G[48] = in[132] & in2[132];
    assign P[48] = in[132] ^ in2[132];
    assign G[49] = in[131] & in2[131];
    assign P[49] = in[131] ^ in2[131];
    assign G[50] = in[130] & in2[130];
    assign P[50] = in[130] ^ in2[130];
    assign G[51] = in[129] & in2[129];
    assign P[51] = in[129] ^ in2[129];
    assign G[52] = in[128] & in2[128];
    assign P[52] = in[128] ^ in2[128];
    assign G[53] = in[127] & in2[127];
    assign P[53] = in[127] ^ in2[127];
    assign G[54] = in[126] & in2[126];
    assign P[54] = in[126] ^ in2[126];
    assign G[55] = in[125] & in2[125];
    assign P[55] = in[125] ^ in2[125];
    assign G[56] = in[124] & in2[124];
    assign P[56] = in[124] ^ in2[124];
    assign G[57] = in[123] & in2[123];
    assign P[57] = in[123] ^ in2[123];
    assign G[58] = in[122] & in2[122];
    assign P[58] = in[122] ^ in2[122];
    assign G[59] = in[121] & in2[121];
    assign P[59] = in[121] ^ in2[121];
    assign G[60] = in[120] & in2[120];
    assign P[60] = in[120] ^ in2[120];
    assign G[61] = in[119] & in2[119];
    assign P[61] = in[119] ^ in2[119];
    assign G[62] = in[118] & in2[118];
    assign P[62] = in[118] ^ in2[118];
    assign G[63] = in[117] & in2[117];
    assign P[63] = in[117] ^ in2[117];
    assign G[64] = in[116] & in2[116];
    assign P[64] = in[116] ^ in2[116];
    assign G[65] = in[115] & in2[115];
    assign P[65] = in[115] ^ in2[115];
    assign G[66] = in[114] & in2[114];
    assign P[66] = in[114] ^ in2[114];
    assign G[67] = in[113] & in2[113];
    assign P[67] = in[113] ^ in2[113];
    assign G[68] = in[112] & in2[112];
    assign P[68] = in[112] ^ in2[112];
    assign G[69] = in[111] & in2[111];
    assign P[69] = in[111] ^ in2[111];
    assign G[70] = in[110] & in2[110];
    assign P[70] = in[110] ^ in2[110];
    assign G[71] = in[109] & in2[109];
    assign P[71] = in[109] ^ in2[109];
    assign G[72] = in[108] & in2[108];
    assign P[72] = in[108] ^ in2[108];
    assign G[73] = in[107] & in2[107];
    assign P[73] = in[107] ^ in2[107];
    assign G[74] = in[106] & in2[106];
    assign P[74] = in[106] ^ in2[106];
    assign G[75] = in[105] & in2[105];
    assign P[75] = in[105] ^ in2[105];
    assign G[76] = in[104] & in2[104];
    assign P[76] = in[104] ^ in2[104];
    assign G[77] = in[103] & in2[103];
    assign P[77] = in[103] ^ in2[103];
    assign G[78] = in[102] & in2[102];
    assign P[78] = in[102] ^ in2[102];
    assign G[79] = in[101] & in2[101];
    assign P[79] = in[101] ^ in2[101];
    assign G[80] = in[100] & in2[100];
    assign P[80] = in[100] ^ in2[100];
    assign G[81] = in[99] & in2[99];
    assign P[81] = in[99] ^ in2[99];
    assign G[82] = in[98] & in2[98];
    assign P[82] = in[98] ^ in2[98];
    assign G[83] = in[97] & in2[97];
    assign P[83] = in[97] ^ in2[97];
    assign G[84] = in[96] & in2[96];
    assign P[84] = in[96] ^ in2[96];
    assign G[85] = in[95] & in2[95];
    assign P[85] = in[95] ^ in2[95];
    assign G[86] = in[94] & in2[94];
    assign P[86] = in[94] ^ in2[94];
    assign G[87] = in[93] & in2[93];
    assign P[87] = in[93] ^ in2[93];
    assign G[88] = in[92] & in2[92];
    assign P[88] = in[92] ^ in2[92];
    assign G[89] = in[91] & in2[91];
    assign P[89] = in[91] ^ in2[91];
    assign G[90] = in[90] & in2[90];
    assign P[90] = in[90] ^ in2[90];
    assign G[91] = in[89] & in2[89];
    assign P[91] = in[89] ^ in2[89];
    assign G[92] = in[88] & in2[88];
    assign P[92] = in[88] ^ in2[88];
    assign G[93] = in[87] & in2[87];
    assign P[93] = in[87] ^ in2[87];
    assign G[94] = in[86] & in2[86];
    assign P[94] = in[86] ^ in2[86];
    assign G[95] = in[85] & in2[85];
    assign P[95] = in[85] ^ in2[85];
    assign G[96] = in[84] & in2[84];
    assign P[96] = in[84] ^ in2[84];
    assign G[97] = in[83] & in2[83];
    assign P[97] = in[83] ^ in2[83];
    assign G[98] = in[82] & in2[82];
    assign P[98] = in[82] ^ in2[82];
    assign G[99] = in[81] & in2[81];
    assign P[99] = in[81] ^ in2[81];
    assign G[100] = in[80] & in2[80];
    assign P[100] = in[80] ^ in2[80];
    assign G[101] = in[79] & in2[79];
    assign P[101] = in[79] ^ in2[79];
    assign G[102] = in[78] & in2[78];
    assign P[102] = in[78] ^ in2[78];
    assign G[103] = in[77] & in2[77];
    assign P[103] = in[77] ^ in2[77];
    assign G[104] = in[76] & in2[76];
    assign P[104] = in[76] ^ in2[76];
    assign G[105] = in[75] & in2[75];
    assign P[105] = in[75] ^ in2[75];
    assign G[106] = in[74] & in2[74];
    assign P[106] = in[74] ^ in2[74];
    assign G[107] = in[73] & in2[73];
    assign P[107] = in[73] ^ in2[73];
    assign G[108] = in[72] & in2[72];
    assign P[108] = in[72] ^ in2[72];
    assign G[109] = in[71] & in2[71];
    assign P[109] = in[71] ^ in2[71];
    assign G[110] = in[70] & in2[70];
    assign P[110] = in[70] ^ in2[70];
    assign G[111] = in[69] & in2[69];
    assign P[111] = in[69] ^ in2[69];
    assign G[112] = in[68] & in2[68];
    assign P[112] = in[68] ^ in2[68];
    assign G[113] = in[67] & in2[67];
    assign P[113] = in[67] ^ in2[67];
    assign G[114] = in[66] & in2[66];
    assign P[114] = in[66] ^ in2[66];
    assign G[115] = in[65] & in2[65];
    assign P[115] = in[65] ^ in2[65];
    assign G[116] = in[64] & in2[64];
    assign P[116] = in[64] ^ in2[64];
    assign G[117] = in[63] & in2[63];
    assign P[117] = in[63] ^ in2[63];
    assign G[118] = in[62] & in2[62];
    assign P[118] = in[62] ^ in2[62];
    assign G[119] = in[61] & in2[61];
    assign P[119] = in[61] ^ in2[61];
    assign G[120] = in[60] & in2[60];
    assign P[120] = in[60] ^ in2[60];
    assign G[121] = in[59] & in2[59];
    assign P[121] = in[59] ^ in2[59];
    assign G[122] = in[58] & in2[58];
    assign P[122] = in[58] ^ in2[58];
    assign G[123] = in[57] & in2[57];
    assign P[123] = in[57] ^ in2[57];
    assign G[124] = in[56] & in2[56];
    assign P[124] = in[56] ^ in2[56];
    assign G[125] = in[55] & in2[55];
    assign P[125] = in[55] ^ in2[55];
    assign G[126] = in[54] & in2[54];
    assign P[126] = in[54] ^ in2[54];
    assign G[127] = in[53] & in2[53];
    assign P[127] = in[53] ^ in2[53];
    assign G[128] = in[52] & in2[52];
    assign P[128] = in[52] ^ in2[52];
    assign G[129] = in[51] & in2[51];
    assign P[129] = in[51] ^ in2[51];
    assign G[130] = in[50] & in2[50];
    assign P[130] = in[50] ^ in2[50];
    assign G[131] = in[49] & in2[49];
    assign P[131] = in[49] ^ in2[49];
    assign G[132] = in[48] & in2[48];
    assign P[132] = in[48] ^ in2[48];
    assign G[133] = in[47] & in2[47];
    assign P[133] = in[47] ^ in2[47];
    assign G[134] = in[46] & in2[46];
    assign P[134] = in[46] ^ in2[46];
    assign G[135] = in[45] & in2[45];
    assign P[135] = in[45] ^ in2[45];
    assign G[136] = in[44] & in2[44];
    assign P[136] = in[44] ^ in2[44];
    assign G[137] = in[43] & in2[43];
    assign P[137] = in[43] ^ in2[43];
    assign G[138] = in[42] & in2[42];
    assign P[138] = in[42] ^ in2[42];
    assign G[139] = in[41] & in2[41];
    assign P[139] = in[41] ^ in2[41];
    assign G[140] = in[40] & in2[40];
    assign P[140] = in[40] ^ in2[40];
    assign G[141] = in[39] & in2[39];
    assign P[141] = in[39] ^ in2[39];
    assign G[142] = in[38] & in2[38];
    assign P[142] = in[38] ^ in2[38];
    assign G[143] = in[37] & in2[37];
    assign P[143] = in[37] ^ in2[37];
    assign G[144] = in[36] & in2[36];
    assign P[144] = in[36] ^ in2[36];
    assign G[145] = in[35] & in2[35];
    assign P[145] = in[35] ^ in2[35];
    assign G[146] = in[34] & in2[34];
    assign P[146] = in[34] ^ in2[34];
    assign G[147] = in[33] & in2[33];
    assign P[147] = in[33] ^ in2[33];
    assign G[148] = in[32] & in2[32];
    assign P[148] = in[32] ^ in2[32];
    assign G[149] = in[31] & in2[31];
    assign P[149] = in[31] ^ in2[31];
    assign G[150] = in[30] & in2[30];
    assign P[150] = in[30] ^ in2[30];
    assign G[151] = in[29] & in2[29];
    assign P[151] = in[29] ^ in2[29];
    assign G[152] = in[28] & in2[28];
    assign P[152] = in[28] ^ in2[28];
    assign G[153] = in[27] & in2[27];
    assign P[153] = in[27] ^ in2[27];
    assign G[154] = in[26] & in2[26];
    assign P[154] = in[26] ^ in2[26];
    assign G[155] = in[25] & in2[25];
    assign P[155] = in[25] ^ in2[25];
    assign G[156] = in[24] & in2[24];
    assign P[156] = in[24] ^ in2[24];
    assign G[157] = in[23] & in2[23];
    assign P[157] = in[23] ^ in2[23];
    assign G[158] = in[22] & in2[22];
    assign P[158] = in[22] ^ in2[22];
    assign G[159] = in[21] & in2[21];
    assign P[159] = in[21] ^ in2[21];
    assign G[160] = in[20] & in2[20];
    assign P[160] = in[20] ^ in2[20];
    assign G[161] = in[19] & in2[19];
    assign P[161] = in[19] ^ in2[19];
    assign G[162] = in[18] & in2[18];
    assign P[162] = in[18] ^ in2[18];
    assign G[163] = in[17] & in2[17];
    assign P[163] = in[17] ^ in2[17];
    assign G[164] = in[16] & in2[16];
    assign P[164] = in[16] ^ in2[16];
    assign G[165] = in[15] & in2[15];
    assign P[165] = in[15] ^ in2[15];
    assign G[166] = in[14] & in2[14];
    assign P[166] = in[14] ^ in2[14];
    assign G[167] = in[13] & in2[13];
    assign P[167] = in[13] ^ in2[13];
    assign G[168] = in[12] & in2[12];
    assign P[168] = in[12] ^ in2[12];
    assign G[169] = in[11] & in2[11];
    assign P[169] = in[11] ^ in2[11];
    assign G[170] = in[10] & in2[10];
    assign P[170] = in[10] ^ in2[10];
    assign G[171] = in[9] & in2[9];
    assign P[171] = in[9] ^ in2[9];
    assign G[172] = in[8] & in2[8];
    assign P[172] = in[8] ^ in2[8];
    assign G[173] = in[7] & in2[7];
    assign P[173] = in[7] ^ in2[7];
    assign G[174] = in[6] & in2[6];
    assign P[174] = in[6] ^ in2[6];
    assign G[175] = in[5] & in2[5];
    assign P[175] = in[5] ^ in2[5];
    assign G[176] = in[4] & in2[4];
    assign P[176] = in[4] ^ in2[4];
    assign G[177] = in[3] & in2[3];
    assign P[177] = in[3] ^ in2[3];
    assign G[178] = in[2] & in2[2];
    assign P[178] = in[2] ^ in2[2];
    assign G[179] = in[1] & in2[1];
    assign P[179] = in[1] ^ in2[1];
    assign G[180] = in[0] & in2[0];
    assign P[180] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign C[180] = G[179] | (P[179] & C[179]);
    assign cout = G[180] | (P[180] & C[180]);
    assign sum = P ^ C;
endmodule

module CLA180(output [179:0] sum, output cout, input [179:0] in1, input [179:0] in2;

    wire[179:0] G;
    wire[179:0] C;
    wire[179:0] P;

    assign G[0] = in[179] & in2[179];
    assign P[0] = in[179] ^ in2[179];
    assign G[1] = in[178] & in2[178];
    assign P[1] = in[178] ^ in2[178];
    assign G[2] = in[177] & in2[177];
    assign P[2] = in[177] ^ in2[177];
    assign G[3] = in[176] & in2[176];
    assign P[3] = in[176] ^ in2[176];
    assign G[4] = in[175] & in2[175];
    assign P[4] = in[175] ^ in2[175];
    assign G[5] = in[174] & in2[174];
    assign P[5] = in[174] ^ in2[174];
    assign G[6] = in[173] & in2[173];
    assign P[6] = in[173] ^ in2[173];
    assign G[7] = in[172] & in2[172];
    assign P[7] = in[172] ^ in2[172];
    assign G[8] = in[171] & in2[171];
    assign P[8] = in[171] ^ in2[171];
    assign G[9] = in[170] & in2[170];
    assign P[9] = in[170] ^ in2[170];
    assign G[10] = in[169] & in2[169];
    assign P[10] = in[169] ^ in2[169];
    assign G[11] = in[168] & in2[168];
    assign P[11] = in[168] ^ in2[168];
    assign G[12] = in[167] & in2[167];
    assign P[12] = in[167] ^ in2[167];
    assign G[13] = in[166] & in2[166];
    assign P[13] = in[166] ^ in2[166];
    assign G[14] = in[165] & in2[165];
    assign P[14] = in[165] ^ in2[165];
    assign G[15] = in[164] & in2[164];
    assign P[15] = in[164] ^ in2[164];
    assign G[16] = in[163] & in2[163];
    assign P[16] = in[163] ^ in2[163];
    assign G[17] = in[162] & in2[162];
    assign P[17] = in[162] ^ in2[162];
    assign G[18] = in[161] & in2[161];
    assign P[18] = in[161] ^ in2[161];
    assign G[19] = in[160] & in2[160];
    assign P[19] = in[160] ^ in2[160];
    assign G[20] = in[159] & in2[159];
    assign P[20] = in[159] ^ in2[159];
    assign G[21] = in[158] & in2[158];
    assign P[21] = in[158] ^ in2[158];
    assign G[22] = in[157] & in2[157];
    assign P[22] = in[157] ^ in2[157];
    assign G[23] = in[156] & in2[156];
    assign P[23] = in[156] ^ in2[156];
    assign G[24] = in[155] & in2[155];
    assign P[24] = in[155] ^ in2[155];
    assign G[25] = in[154] & in2[154];
    assign P[25] = in[154] ^ in2[154];
    assign G[26] = in[153] & in2[153];
    assign P[26] = in[153] ^ in2[153];
    assign G[27] = in[152] & in2[152];
    assign P[27] = in[152] ^ in2[152];
    assign G[28] = in[151] & in2[151];
    assign P[28] = in[151] ^ in2[151];
    assign G[29] = in[150] & in2[150];
    assign P[29] = in[150] ^ in2[150];
    assign G[30] = in[149] & in2[149];
    assign P[30] = in[149] ^ in2[149];
    assign G[31] = in[148] & in2[148];
    assign P[31] = in[148] ^ in2[148];
    assign G[32] = in[147] & in2[147];
    assign P[32] = in[147] ^ in2[147];
    assign G[33] = in[146] & in2[146];
    assign P[33] = in[146] ^ in2[146];
    assign G[34] = in[145] & in2[145];
    assign P[34] = in[145] ^ in2[145];
    assign G[35] = in[144] & in2[144];
    assign P[35] = in[144] ^ in2[144];
    assign G[36] = in[143] & in2[143];
    assign P[36] = in[143] ^ in2[143];
    assign G[37] = in[142] & in2[142];
    assign P[37] = in[142] ^ in2[142];
    assign G[38] = in[141] & in2[141];
    assign P[38] = in[141] ^ in2[141];
    assign G[39] = in[140] & in2[140];
    assign P[39] = in[140] ^ in2[140];
    assign G[40] = in[139] & in2[139];
    assign P[40] = in[139] ^ in2[139];
    assign G[41] = in[138] & in2[138];
    assign P[41] = in[138] ^ in2[138];
    assign G[42] = in[137] & in2[137];
    assign P[42] = in[137] ^ in2[137];
    assign G[43] = in[136] & in2[136];
    assign P[43] = in[136] ^ in2[136];
    assign G[44] = in[135] & in2[135];
    assign P[44] = in[135] ^ in2[135];
    assign G[45] = in[134] & in2[134];
    assign P[45] = in[134] ^ in2[134];
    assign G[46] = in[133] & in2[133];
    assign P[46] = in[133] ^ in2[133];
    assign G[47] = in[132] & in2[132];
    assign P[47] = in[132] ^ in2[132];
    assign G[48] = in[131] & in2[131];
    assign P[48] = in[131] ^ in2[131];
    assign G[49] = in[130] & in2[130];
    assign P[49] = in[130] ^ in2[130];
    assign G[50] = in[129] & in2[129];
    assign P[50] = in[129] ^ in2[129];
    assign G[51] = in[128] & in2[128];
    assign P[51] = in[128] ^ in2[128];
    assign G[52] = in[127] & in2[127];
    assign P[52] = in[127] ^ in2[127];
    assign G[53] = in[126] & in2[126];
    assign P[53] = in[126] ^ in2[126];
    assign G[54] = in[125] & in2[125];
    assign P[54] = in[125] ^ in2[125];
    assign G[55] = in[124] & in2[124];
    assign P[55] = in[124] ^ in2[124];
    assign G[56] = in[123] & in2[123];
    assign P[56] = in[123] ^ in2[123];
    assign G[57] = in[122] & in2[122];
    assign P[57] = in[122] ^ in2[122];
    assign G[58] = in[121] & in2[121];
    assign P[58] = in[121] ^ in2[121];
    assign G[59] = in[120] & in2[120];
    assign P[59] = in[120] ^ in2[120];
    assign G[60] = in[119] & in2[119];
    assign P[60] = in[119] ^ in2[119];
    assign G[61] = in[118] & in2[118];
    assign P[61] = in[118] ^ in2[118];
    assign G[62] = in[117] & in2[117];
    assign P[62] = in[117] ^ in2[117];
    assign G[63] = in[116] & in2[116];
    assign P[63] = in[116] ^ in2[116];
    assign G[64] = in[115] & in2[115];
    assign P[64] = in[115] ^ in2[115];
    assign G[65] = in[114] & in2[114];
    assign P[65] = in[114] ^ in2[114];
    assign G[66] = in[113] & in2[113];
    assign P[66] = in[113] ^ in2[113];
    assign G[67] = in[112] & in2[112];
    assign P[67] = in[112] ^ in2[112];
    assign G[68] = in[111] & in2[111];
    assign P[68] = in[111] ^ in2[111];
    assign G[69] = in[110] & in2[110];
    assign P[69] = in[110] ^ in2[110];
    assign G[70] = in[109] & in2[109];
    assign P[70] = in[109] ^ in2[109];
    assign G[71] = in[108] & in2[108];
    assign P[71] = in[108] ^ in2[108];
    assign G[72] = in[107] & in2[107];
    assign P[72] = in[107] ^ in2[107];
    assign G[73] = in[106] & in2[106];
    assign P[73] = in[106] ^ in2[106];
    assign G[74] = in[105] & in2[105];
    assign P[74] = in[105] ^ in2[105];
    assign G[75] = in[104] & in2[104];
    assign P[75] = in[104] ^ in2[104];
    assign G[76] = in[103] & in2[103];
    assign P[76] = in[103] ^ in2[103];
    assign G[77] = in[102] & in2[102];
    assign P[77] = in[102] ^ in2[102];
    assign G[78] = in[101] & in2[101];
    assign P[78] = in[101] ^ in2[101];
    assign G[79] = in[100] & in2[100];
    assign P[79] = in[100] ^ in2[100];
    assign G[80] = in[99] & in2[99];
    assign P[80] = in[99] ^ in2[99];
    assign G[81] = in[98] & in2[98];
    assign P[81] = in[98] ^ in2[98];
    assign G[82] = in[97] & in2[97];
    assign P[82] = in[97] ^ in2[97];
    assign G[83] = in[96] & in2[96];
    assign P[83] = in[96] ^ in2[96];
    assign G[84] = in[95] & in2[95];
    assign P[84] = in[95] ^ in2[95];
    assign G[85] = in[94] & in2[94];
    assign P[85] = in[94] ^ in2[94];
    assign G[86] = in[93] & in2[93];
    assign P[86] = in[93] ^ in2[93];
    assign G[87] = in[92] & in2[92];
    assign P[87] = in[92] ^ in2[92];
    assign G[88] = in[91] & in2[91];
    assign P[88] = in[91] ^ in2[91];
    assign G[89] = in[90] & in2[90];
    assign P[89] = in[90] ^ in2[90];
    assign G[90] = in[89] & in2[89];
    assign P[90] = in[89] ^ in2[89];
    assign G[91] = in[88] & in2[88];
    assign P[91] = in[88] ^ in2[88];
    assign G[92] = in[87] & in2[87];
    assign P[92] = in[87] ^ in2[87];
    assign G[93] = in[86] & in2[86];
    assign P[93] = in[86] ^ in2[86];
    assign G[94] = in[85] & in2[85];
    assign P[94] = in[85] ^ in2[85];
    assign G[95] = in[84] & in2[84];
    assign P[95] = in[84] ^ in2[84];
    assign G[96] = in[83] & in2[83];
    assign P[96] = in[83] ^ in2[83];
    assign G[97] = in[82] & in2[82];
    assign P[97] = in[82] ^ in2[82];
    assign G[98] = in[81] & in2[81];
    assign P[98] = in[81] ^ in2[81];
    assign G[99] = in[80] & in2[80];
    assign P[99] = in[80] ^ in2[80];
    assign G[100] = in[79] & in2[79];
    assign P[100] = in[79] ^ in2[79];
    assign G[101] = in[78] & in2[78];
    assign P[101] = in[78] ^ in2[78];
    assign G[102] = in[77] & in2[77];
    assign P[102] = in[77] ^ in2[77];
    assign G[103] = in[76] & in2[76];
    assign P[103] = in[76] ^ in2[76];
    assign G[104] = in[75] & in2[75];
    assign P[104] = in[75] ^ in2[75];
    assign G[105] = in[74] & in2[74];
    assign P[105] = in[74] ^ in2[74];
    assign G[106] = in[73] & in2[73];
    assign P[106] = in[73] ^ in2[73];
    assign G[107] = in[72] & in2[72];
    assign P[107] = in[72] ^ in2[72];
    assign G[108] = in[71] & in2[71];
    assign P[108] = in[71] ^ in2[71];
    assign G[109] = in[70] & in2[70];
    assign P[109] = in[70] ^ in2[70];
    assign G[110] = in[69] & in2[69];
    assign P[110] = in[69] ^ in2[69];
    assign G[111] = in[68] & in2[68];
    assign P[111] = in[68] ^ in2[68];
    assign G[112] = in[67] & in2[67];
    assign P[112] = in[67] ^ in2[67];
    assign G[113] = in[66] & in2[66];
    assign P[113] = in[66] ^ in2[66];
    assign G[114] = in[65] & in2[65];
    assign P[114] = in[65] ^ in2[65];
    assign G[115] = in[64] & in2[64];
    assign P[115] = in[64] ^ in2[64];
    assign G[116] = in[63] & in2[63];
    assign P[116] = in[63] ^ in2[63];
    assign G[117] = in[62] & in2[62];
    assign P[117] = in[62] ^ in2[62];
    assign G[118] = in[61] & in2[61];
    assign P[118] = in[61] ^ in2[61];
    assign G[119] = in[60] & in2[60];
    assign P[119] = in[60] ^ in2[60];
    assign G[120] = in[59] & in2[59];
    assign P[120] = in[59] ^ in2[59];
    assign G[121] = in[58] & in2[58];
    assign P[121] = in[58] ^ in2[58];
    assign G[122] = in[57] & in2[57];
    assign P[122] = in[57] ^ in2[57];
    assign G[123] = in[56] & in2[56];
    assign P[123] = in[56] ^ in2[56];
    assign G[124] = in[55] & in2[55];
    assign P[124] = in[55] ^ in2[55];
    assign G[125] = in[54] & in2[54];
    assign P[125] = in[54] ^ in2[54];
    assign G[126] = in[53] & in2[53];
    assign P[126] = in[53] ^ in2[53];
    assign G[127] = in[52] & in2[52];
    assign P[127] = in[52] ^ in2[52];
    assign G[128] = in[51] & in2[51];
    assign P[128] = in[51] ^ in2[51];
    assign G[129] = in[50] & in2[50];
    assign P[129] = in[50] ^ in2[50];
    assign G[130] = in[49] & in2[49];
    assign P[130] = in[49] ^ in2[49];
    assign G[131] = in[48] & in2[48];
    assign P[131] = in[48] ^ in2[48];
    assign G[132] = in[47] & in2[47];
    assign P[132] = in[47] ^ in2[47];
    assign G[133] = in[46] & in2[46];
    assign P[133] = in[46] ^ in2[46];
    assign G[134] = in[45] & in2[45];
    assign P[134] = in[45] ^ in2[45];
    assign G[135] = in[44] & in2[44];
    assign P[135] = in[44] ^ in2[44];
    assign G[136] = in[43] & in2[43];
    assign P[136] = in[43] ^ in2[43];
    assign G[137] = in[42] & in2[42];
    assign P[137] = in[42] ^ in2[42];
    assign G[138] = in[41] & in2[41];
    assign P[138] = in[41] ^ in2[41];
    assign G[139] = in[40] & in2[40];
    assign P[139] = in[40] ^ in2[40];
    assign G[140] = in[39] & in2[39];
    assign P[140] = in[39] ^ in2[39];
    assign G[141] = in[38] & in2[38];
    assign P[141] = in[38] ^ in2[38];
    assign G[142] = in[37] & in2[37];
    assign P[142] = in[37] ^ in2[37];
    assign G[143] = in[36] & in2[36];
    assign P[143] = in[36] ^ in2[36];
    assign G[144] = in[35] & in2[35];
    assign P[144] = in[35] ^ in2[35];
    assign G[145] = in[34] & in2[34];
    assign P[145] = in[34] ^ in2[34];
    assign G[146] = in[33] & in2[33];
    assign P[146] = in[33] ^ in2[33];
    assign G[147] = in[32] & in2[32];
    assign P[147] = in[32] ^ in2[32];
    assign G[148] = in[31] & in2[31];
    assign P[148] = in[31] ^ in2[31];
    assign G[149] = in[30] & in2[30];
    assign P[149] = in[30] ^ in2[30];
    assign G[150] = in[29] & in2[29];
    assign P[150] = in[29] ^ in2[29];
    assign G[151] = in[28] & in2[28];
    assign P[151] = in[28] ^ in2[28];
    assign G[152] = in[27] & in2[27];
    assign P[152] = in[27] ^ in2[27];
    assign G[153] = in[26] & in2[26];
    assign P[153] = in[26] ^ in2[26];
    assign G[154] = in[25] & in2[25];
    assign P[154] = in[25] ^ in2[25];
    assign G[155] = in[24] & in2[24];
    assign P[155] = in[24] ^ in2[24];
    assign G[156] = in[23] & in2[23];
    assign P[156] = in[23] ^ in2[23];
    assign G[157] = in[22] & in2[22];
    assign P[157] = in[22] ^ in2[22];
    assign G[158] = in[21] & in2[21];
    assign P[158] = in[21] ^ in2[21];
    assign G[159] = in[20] & in2[20];
    assign P[159] = in[20] ^ in2[20];
    assign G[160] = in[19] & in2[19];
    assign P[160] = in[19] ^ in2[19];
    assign G[161] = in[18] & in2[18];
    assign P[161] = in[18] ^ in2[18];
    assign G[162] = in[17] & in2[17];
    assign P[162] = in[17] ^ in2[17];
    assign G[163] = in[16] & in2[16];
    assign P[163] = in[16] ^ in2[16];
    assign G[164] = in[15] & in2[15];
    assign P[164] = in[15] ^ in2[15];
    assign G[165] = in[14] & in2[14];
    assign P[165] = in[14] ^ in2[14];
    assign G[166] = in[13] & in2[13];
    assign P[166] = in[13] ^ in2[13];
    assign G[167] = in[12] & in2[12];
    assign P[167] = in[12] ^ in2[12];
    assign G[168] = in[11] & in2[11];
    assign P[168] = in[11] ^ in2[11];
    assign G[169] = in[10] & in2[10];
    assign P[169] = in[10] ^ in2[10];
    assign G[170] = in[9] & in2[9];
    assign P[170] = in[9] ^ in2[9];
    assign G[171] = in[8] & in2[8];
    assign P[171] = in[8] ^ in2[8];
    assign G[172] = in[7] & in2[7];
    assign P[172] = in[7] ^ in2[7];
    assign G[173] = in[6] & in2[6];
    assign P[173] = in[6] ^ in2[6];
    assign G[174] = in[5] & in2[5];
    assign P[174] = in[5] ^ in2[5];
    assign G[175] = in[4] & in2[4];
    assign P[175] = in[4] ^ in2[4];
    assign G[176] = in[3] & in2[3];
    assign P[176] = in[3] ^ in2[3];
    assign G[177] = in[2] & in2[2];
    assign P[177] = in[2] ^ in2[2];
    assign G[178] = in[1] & in2[1];
    assign P[178] = in[1] ^ in2[1];
    assign G[179] = in[0] & in2[0];
    assign P[179] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign C[179] = G[178] | (P[178] & C[178]);
    assign cout = G[179] | (P[179] & C[179]);
    assign sum = P ^ C;
endmodule

module CLA179(output [178:0] sum, output cout, input [178:0] in1, input [178:0] in2;

    wire[178:0] G;
    wire[178:0] C;
    wire[178:0] P;

    assign G[0] = in[178] & in2[178];
    assign P[0] = in[178] ^ in2[178];
    assign G[1] = in[177] & in2[177];
    assign P[1] = in[177] ^ in2[177];
    assign G[2] = in[176] & in2[176];
    assign P[2] = in[176] ^ in2[176];
    assign G[3] = in[175] & in2[175];
    assign P[3] = in[175] ^ in2[175];
    assign G[4] = in[174] & in2[174];
    assign P[4] = in[174] ^ in2[174];
    assign G[5] = in[173] & in2[173];
    assign P[5] = in[173] ^ in2[173];
    assign G[6] = in[172] & in2[172];
    assign P[6] = in[172] ^ in2[172];
    assign G[7] = in[171] & in2[171];
    assign P[7] = in[171] ^ in2[171];
    assign G[8] = in[170] & in2[170];
    assign P[8] = in[170] ^ in2[170];
    assign G[9] = in[169] & in2[169];
    assign P[9] = in[169] ^ in2[169];
    assign G[10] = in[168] & in2[168];
    assign P[10] = in[168] ^ in2[168];
    assign G[11] = in[167] & in2[167];
    assign P[11] = in[167] ^ in2[167];
    assign G[12] = in[166] & in2[166];
    assign P[12] = in[166] ^ in2[166];
    assign G[13] = in[165] & in2[165];
    assign P[13] = in[165] ^ in2[165];
    assign G[14] = in[164] & in2[164];
    assign P[14] = in[164] ^ in2[164];
    assign G[15] = in[163] & in2[163];
    assign P[15] = in[163] ^ in2[163];
    assign G[16] = in[162] & in2[162];
    assign P[16] = in[162] ^ in2[162];
    assign G[17] = in[161] & in2[161];
    assign P[17] = in[161] ^ in2[161];
    assign G[18] = in[160] & in2[160];
    assign P[18] = in[160] ^ in2[160];
    assign G[19] = in[159] & in2[159];
    assign P[19] = in[159] ^ in2[159];
    assign G[20] = in[158] & in2[158];
    assign P[20] = in[158] ^ in2[158];
    assign G[21] = in[157] & in2[157];
    assign P[21] = in[157] ^ in2[157];
    assign G[22] = in[156] & in2[156];
    assign P[22] = in[156] ^ in2[156];
    assign G[23] = in[155] & in2[155];
    assign P[23] = in[155] ^ in2[155];
    assign G[24] = in[154] & in2[154];
    assign P[24] = in[154] ^ in2[154];
    assign G[25] = in[153] & in2[153];
    assign P[25] = in[153] ^ in2[153];
    assign G[26] = in[152] & in2[152];
    assign P[26] = in[152] ^ in2[152];
    assign G[27] = in[151] & in2[151];
    assign P[27] = in[151] ^ in2[151];
    assign G[28] = in[150] & in2[150];
    assign P[28] = in[150] ^ in2[150];
    assign G[29] = in[149] & in2[149];
    assign P[29] = in[149] ^ in2[149];
    assign G[30] = in[148] & in2[148];
    assign P[30] = in[148] ^ in2[148];
    assign G[31] = in[147] & in2[147];
    assign P[31] = in[147] ^ in2[147];
    assign G[32] = in[146] & in2[146];
    assign P[32] = in[146] ^ in2[146];
    assign G[33] = in[145] & in2[145];
    assign P[33] = in[145] ^ in2[145];
    assign G[34] = in[144] & in2[144];
    assign P[34] = in[144] ^ in2[144];
    assign G[35] = in[143] & in2[143];
    assign P[35] = in[143] ^ in2[143];
    assign G[36] = in[142] & in2[142];
    assign P[36] = in[142] ^ in2[142];
    assign G[37] = in[141] & in2[141];
    assign P[37] = in[141] ^ in2[141];
    assign G[38] = in[140] & in2[140];
    assign P[38] = in[140] ^ in2[140];
    assign G[39] = in[139] & in2[139];
    assign P[39] = in[139] ^ in2[139];
    assign G[40] = in[138] & in2[138];
    assign P[40] = in[138] ^ in2[138];
    assign G[41] = in[137] & in2[137];
    assign P[41] = in[137] ^ in2[137];
    assign G[42] = in[136] & in2[136];
    assign P[42] = in[136] ^ in2[136];
    assign G[43] = in[135] & in2[135];
    assign P[43] = in[135] ^ in2[135];
    assign G[44] = in[134] & in2[134];
    assign P[44] = in[134] ^ in2[134];
    assign G[45] = in[133] & in2[133];
    assign P[45] = in[133] ^ in2[133];
    assign G[46] = in[132] & in2[132];
    assign P[46] = in[132] ^ in2[132];
    assign G[47] = in[131] & in2[131];
    assign P[47] = in[131] ^ in2[131];
    assign G[48] = in[130] & in2[130];
    assign P[48] = in[130] ^ in2[130];
    assign G[49] = in[129] & in2[129];
    assign P[49] = in[129] ^ in2[129];
    assign G[50] = in[128] & in2[128];
    assign P[50] = in[128] ^ in2[128];
    assign G[51] = in[127] & in2[127];
    assign P[51] = in[127] ^ in2[127];
    assign G[52] = in[126] & in2[126];
    assign P[52] = in[126] ^ in2[126];
    assign G[53] = in[125] & in2[125];
    assign P[53] = in[125] ^ in2[125];
    assign G[54] = in[124] & in2[124];
    assign P[54] = in[124] ^ in2[124];
    assign G[55] = in[123] & in2[123];
    assign P[55] = in[123] ^ in2[123];
    assign G[56] = in[122] & in2[122];
    assign P[56] = in[122] ^ in2[122];
    assign G[57] = in[121] & in2[121];
    assign P[57] = in[121] ^ in2[121];
    assign G[58] = in[120] & in2[120];
    assign P[58] = in[120] ^ in2[120];
    assign G[59] = in[119] & in2[119];
    assign P[59] = in[119] ^ in2[119];
    assign G[60] = in[118] & in2[118];
    assign P[60] = in[118] ^ in2[118];
    assign G[61] = in[117] & in2[117];
    assign P[61] = in[117] ^ in2[117];
    assign G[62] = in[116] & in2[116];
    assign P[62] = in[116] ^ in2[116];
    assign G[63] = in[115] & in2[115];
    assign P[63] = in[115] ^ in2[115];
    assign G[64] = in[114] & in2[114];
    assign P[64] = in[114] ^ in2[114];
    assign G[65] = in[113] & in2[113];
    assign P[65] = in[113] ^ in2[113];
    assign G[66] = in[112] & in2[112];
    assign P[66] = in[112] ^ in2[112];
    assign G[67] = in[111] & in2[111];
    assign P[67] = in[111] ^ in2[111];
    assign G[68] = in[110] & in2[110];
    assign P[68] = in[110] ^ in2[110];
    assign G[69] = in[109] & in2[109];
    assign P[69] = in[109] ^ in2[109];
    assign G[70] = in[108] & in2[108];
    assign P[70] = in[108] ^ in2[108];
    assign G[71] = in[107] & in2[107];
    assign P[71] = in[107] ^ in2[107];
    assign G[72] = in[106] & in2[106];
    assign P[72] = in[106] ^ in2[106];
    assign G[73] = in[105] & in2[105];
    assign P[73] = in[105] ^ in2[105];
    assign G[74] = in[104] & in2[104];
    assign P[74] = in[104] ^ in2[104];
    assign G[75] = in[103] & in2[103];
    assign P[75] = in[103] ^ in2[103];
    assign G[76] = in[102] & in2[102];
    assign P[76] = in[102] ^ in2[102];
    assign G[77] = in[101] & in2[101];
    assign P[77] = in[101] ^ in2[101];
    assign G[78] = in[100] & in2[100];
    assign P[78] = in[100] ^ in2[100];
    assign G[79] = in[99] & in2[99];
    assign P[79] = in[99] ^ in2[99];
    assign G[80] = in[98] & in2[98];
    assign P[80] = in[98] ^ in2[98];
    assign G[81] = in[97] & in2[97];
    assign P[81] = in[97] ^ in2[97];
    assign G[82] = in[96] & in2[96];
    assign P[82] = in[96] ^ in2[96];
    assign G[83] = in[95] & in2[95];
    assign P[83] = in[95] ^ in2[95];
    assign G[84] = in[94] & in2[94];
    assign P[84] = in[94] ^ in2[94];
    assign G[85] = in[93] & in2[93];
    assign P[85] = in[93] ^ in2[93];
    assign G[86] = in[92] & in2[92];
    assign P[86] = in[92] ^ in2[92];
    assign G[87] = in[91] & in2[91];
    assign P[87] = in[91] ^ in2[91];
    assign G[88] = in[90] & in2[90];
    assign P[88] = in[90] ^ in2[90];
    assign G[89] = in[89] & in2[89];
    assign P[89] = in[89] ^ in2[89];
    assign G[90] = in[88] & in2[88];
    assign P[90] = in[88] ^ in2[88];
    assign G[91] = in[87] & in2[87];
    assign P[91] = in[87] ^ in2[87];
    assign G[92] = in[86] & in2[86];
    assign P[92] = in[86] ^ in2[86];
    assign G[93] = in[85] & in2[85];
    assign P[93] = in[85] ^ in2[85];
    assign G[94] = in[84] & in2[84];
    assign P[94] = in[84] ^ in2[84];
    assign G[95] = in[83] & in2[83];
    assign P[95] = in[83] ^ in2[83];
    assign G[96] = in[82] & in2[82];
    assign P[96] = in[82] ^ in2[82];
    assign G[97] = in[81] & in2[81];
    assign P[97] = in[81] ^ in2[81];
    assign G[98] = in[80] & in2[80];
    assign P[98] = in[80] ^ in2[80];
    assign G[99] = in[79] & in2[79];
    assign P[99] = in[79] ^ in2[79];
    assign G[100] = in[78] & in2[78];
    assign P[100] = in[78] ^ in2[78];
    assign G[101] = in[77] & in2[77];
    assign P[101] = in[77] ^ in2[77];
    assign G[102] = in[76] & in2[76];
    assign P[102] = in[76] ^ in2[76];
    assign G[103] = in[75] & in2[75];
    assign P[103] = in[75] ^ in2[75];
    assign G[104] = in[74] & in2[74];
    assign P[104] = in[74] ^ in2[74];
    assign G[105] = in[73] & in2[73];
    assign P[105] = in[73] ^ in2[73];
    assign G[106] = in[72] & in2[72];
    assign P[106] = in[72] ^ in2[72];
    assign G[107] = in[71] & in2[71];
    assign P[107] = in[71] ^ in2[71];
    assign G[108] = in[70] & in2[70];
    assign P[108] = in[70] ^ in2[70];
    assign G[109] = in[69] & in2[69];
    assign P[109] = in[69] ^ in2[69];
    assign G[110] = in[68] & in2[68];
    assign P[110] = in[68] ^ in2[68];
    assign G[111] = in[67] & in2[67];
    assign P[111] = in[67] ^ in2[67];
    assign G[112] = in[66] & in2[66];
    assign P[112] = in[66] ^ in2[66];
    assign G[113] = in[65] & in2[65];
    assign P[113] = in[65] ^ in2[65];
    assign G[114] = in[64] & in2[64];
    assign P[114] = in[64] ^ in2[64];
    assign G[115] = in[63] & in2[63];
    assign P[115] = in[63] ^ in2[63];
    assign G[116] = in[62] & in2[62];
    assign P[116] = in[62] ^ in2[62];
    assign G[117] = in[61] & in2[61];
    assign P[117] = in[61] ^ in2[61];
    assign G[118] = in[60] & in2[60];
    assign P[118] = in[60] ^ in2[60];
    assign G[119] = in[59] & in2[59];
    assign P[119] = in[59] ^ in2[59];
    assign G[120] = in[58] & in2[58];
    assign P[120] = in[58] ^ in2[58];
    assign G[121] = in[57] & in2[57];
    assign P[121] = in[57] ^ in2[57];
    assign G[122] = in[56] & in2[56];
    assign P[122] = in[56] ^ in2[56];
    assign G[123] = in[55] & in2[55];
    assign P[123] = in[55] ^ in2[55];
    assign G[124] = in[54] & in2[54];
    assign P[124] = in[54] ^ in2[54];
    assign G[125] = in[53] & in2[53];
    assign P[125] = in[53] ^ in2[53];
    assign G[126] = in[52] & in2[52];
    assign P[126] = in[52] ^ in2[52];
    assign G[127] = in[51] & in2[51];
    assign P[127] = in[51] ^ in2[51];
    assign G[128] = in[50] & in2[50];
    assign P[128] = in[50] ^ in2[50];
    assign G[129] = in[49] & in2[49];
    assign P[129] = in[49] ^ in2[49];
    assign G[130] = in[48] & in2[48];
    assign P[130] = in[48] ^ in2[48];
    assign G[131] = in[47] & in2[47];
    assign P[131] = in[47] ^ in2[47];
    assign G[132] = in[46] & in2[46];
    assign P[132] = in[46] ^ in2[46];
    assign G[133] = in[45] & in2[45];
    assign P[133] = in[45] ^ in2[45];
    assign G[134] = in[44] & in2[44];
    assign P[134] = in[44] ^ in2[44];
    assign G[135] = in[43] & in2[43];
    assign P[135] = in[43] ^ in2[43];
    assign G[136] = in[42] & in2[42];
    assign P[136] = in[42] ^ in2[42];
    assign G[137] = in[41] & in2[41];
    assign P[137] = in[41] ^ in2[41];
    assign G[138] = in[40] & in2[40];
    assign P[138] = in[40] ^ in2[40];
    assign G[139] = in[39] & in2[39];
    assign P[139] = in[39] ^ in2[39];
    assign G[140] = in[38] & in2[38];
    assign P[140] = in[38] ^ in2[38];
    assign G[141] = in[37] & in2[37];
    assign P[141] = in[37] ^ in2[37];
    assign G[142] = in[36] & in2[36];
    assign P[142] = in[36] ^ in2[36];
    assign G[143] = in[35] & in2[35];
    assign P[143] = in[35] ^ in2[35];
    assign G[144] = in[34] & in2[34];
    assign P[144] = in[34] ^ in2[34];
    assign G[145] = in[33] & in2[33];
    assign P[145] = in[33] ^ in2[33];
    assign G[146] = in[32] & in2[32];
    assign P[146] = in[32] ^ in2[32];
    assign G[147] = in[31] & in2[31];
    assign P[147] = in[31] ^ in2[31];
    assign G[148] = in[30] & in2[30];
    assign P[148] = in[30] ^ in2[30];
    assign G[149] = in[29] & in2[29];
    assign P[149] = in[29] ^ in2[29];
    assign G[150] = in[28] & in2[28];
    assign P[150] = in[28] ^ in2[28];
    assign G[151] = in[27] & in2[27];
    assign P[151] = in[27] ^ in2[27];
    assign G[152] = in[26] & in2[26];
    assign P[152] = in[26] ^ in2[26];
    assign G[153] = in[25] & in2[25];
    assign P[153] = in[25] ^ in2[25];
    assign G[154] = in[24] & in2[24];
    assign P[154] = in[24] ^ in2[24];
    assign G[155] = in[23] & in2[23];
    assign P[155] = in[23] ^ in2[23];
    assign G[156] = in[22] & in2[22];
    assign P[156] = in[22] ^ in2[22];
    assign G[157] = in[21] & in2[21];
    assign P[157] = in[21] ^ in2[21];
    assign G[158] = in[20] & in2[20];
    assign P[158] = in[20] ^ in2[20];
    assign G[159] = in[19] & in2[19];
    assign P[159] = in[19] ^ in2[19];
    assign G[160] = in[18] & in2[18];
    assign P[160] = in[18] ^ in2[18];
    assign G[161] = in[17] & in2[17];
    assign P[161] = in[17] ^ in2[17];
    assign G[162] = in[16] & in2[16];
    assign P[162] = in[16] ^ in2[16];
    assign G[163] = in[15] & in2[15];
    assign P[163] = in[15] ^ in2[15];
    assign G[164] = in[14] & in2[14];
    assign P[164] = in[14] ^ in2[14];
    assign G[165] = in[13] & in2[13];
    assign P[165] = in[13] ^ in2[13];
    assign G[166] = in[12] & in2[12];
    assign P[166] = in[12] ^ in2[12];
    assign G[167] = in[11] & in2[11];
    assign P[167] = in[11] ^ in2[11];
    assign G[168] = in[10] & in2[10];
    assign P[168] = in[10] ^ in2[10];
    assign G[169] = in[9] & in2[9];
    assign P[169] = in[9] ^ in2[9];
    assign G[170] = in[8] & in2[8];
    assign P[170] = in[8] ^ in2[8];
    assign G[171] = in[7] & in2[7];
    assign P[171] = in[7] ^ in2[7];
    assign G[172] = in[6] & in2[6];
    assign P[172] = in[6] ^ in2[6];
    assign G[173] = in[5] & in2[5];
    assign P[173] = in[5] ^ in2[5];
    assign G[174] = in[4] & in2[4];
    assign P[174] = in[4] ^ in2[4];
    assign G[175] = in[3] & in2[3];
    assign P[175] = in[3] ^ in2[3];
    assign G[176] = in[2] & in2[2];
    assign P[176] = in[2] ^ in2[2];
    assign G[177] = in[1] & in2[1];
    assign P[177] = in[1] ^ in2[1];
    assign G[178] = in[0] & in2[0];
    assign P[178] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign C[178] = G[177] | (P[177] & C[177]);
    assign cout = G[178] | (P[178] & C[178]);
    assign sum = P ^ C;
endmodule

module CLA178(output [177:0] sum, output cout, input [177:0] in1, input [177:0] in2;

    wire[177:0] G;
    wire[177:0] C;
    wire[177:0] P;

    assign G[0] = in[177] & in2[177];
    assign P[0] = in[177] ^ in2[177];
    assign G[1] = in[176] & in2[176];
    assign P[1] = in[176] ^ in2[176];
    assign G[2] = in[175] & in2[175];
    assign P[2] = in[175] ^ in2[175];
    assign G[3] = in[174] & in2[174];
    assign P[3] = in[174] ^ in2[174];
    assign G[4] = in[173] & in2[173];
    assign P[4] = in[173] ^ in2[173];
    assign G[5] = in[172] & in2[172];
    assign P[5] = in[172] ^ in2[172];
    assign G[6] = in[171] & in2[171];
    assign P[6] = in[171] ^ in2[171];
    assign G[7] = in[170] & in2[170];
    assign P[7] = in[170] ^ in2[170];
    assign G[8] = in[169] & in2[169];
    assign P[8] = in[169] ^ in2[169];
    assign G[9] = in[168] & in2[168];
    assign P[9] = in[168] ^ in2[168];
    assign G[10] = in[167] & in2[167];
    assign P[10] = in[167] ^ in2[167];
    assign G[11] = in[166] & in2[166];
    assign P[11] = in[166] ^ in2[166];
    assign G[12] = in[165] & in2[165];
    assign P[12] = in[165] ^ in2[165];
    assign G[13] = in[164] & in2[164];
    assign P[13] = in[164] ^ in2[164];
    assign G[14] = in[163] & in2[163];
    assign P[14] = in[163] ^ in2[163];
    assign G[15] = in[162] & in2[162];
    assign P[15] = in[162] ^ in2[162];
    assign G[16] = in[161] & in2[161];
    assign P[16] = in[161] ^ in2[161];
    assign G[17] = in[160] & in2[160];
    assign P[17] = in[160] ^ in2[160];
    assign G[18] = in[159] & in2[159];
    assign P[18] = in[159] ^ in2[159];
    assign G[19] = in[158] & in2[158];
    assign P[19] = in[158] ^ in2[158];
    assign G[20] = in[157] & in2[157];
    assign P[20] = in[157] ^ in2[157];
    assign G[21] = in[156] & in2[156];
    assign P[21] = in[156] ^ in2[156];
    assign G[22] = in[155] & in2[155];
    assign P[22] = in[155] ^ in2[155];
    assign G[23] = in[154] & in2[154];
    assign P[23] = in[154] ^ in2[154];
    assign G[24] = in[153] & in2[153];
    assign P[24] = in[153] ^ in2[153];
    assign G[25] = in[152] & in2[152];
    assign P[25] = in[152] ^ in2[152];
    assign G[26] = in[151] & in2[151];
    assign P[26] = in[151] ^ in2[151];
    assign G[27] = in[150] & in2[150];
    assign P[27] = in[150] ^ in2[150];
    assign G[28] = in[149] & in2[149];
    assign P[28] = in[149] ^ in2[149];
    assign G[29] = in[148] & in2[148];
    assign P[29] = in[148] ^ in2[148];
    assign G[30] = in[147] & in2[147];
    assign P[30] = in[147] ^ in2[147];
    assign G[31] = in[146] & in2[146];
    assign P[31] = in[146] ^ in2[146];
    assign G[32] = in[145] & in2[145];
    assign P[32] = in[145] ^ in2[145];
    assign G[33] = in[144] & in2[144];
    assign P[33] = in[144] ^ in2[144];
    assign G[34] = in[143] & in2[143];
    assign P[34] = in[143] ^ in2[143];
    assign G[35] = in[142] & in2[142];
    assign P[35] = in[142] ^ in2[142];
    assign G[36] = in[141] & in2[141];
    assign P[36] = in[141] ^ in2[141];
    assign G[37] = in[140] & in2[140];
    assign P[37] = in[140] ^ in2[140];
    assign G[38] = in[139] & in2[139];
    assign P[38] = in[139] ^ in2[139];
    assign G[39] = in[138] & in2[138];
    assign P[39] = in[138] ^ in2[138];
    assign G[40] = in[137] & in2[137];
    assign P[40] = in[137] ^ in2[137];
    assign G[41] = in[136] & in2[136];
    assign P[41] = in[136] ^ in2[136];
    assign G[42] = in[135] & in2[135];
    assign P[42] = in[135] ^ in2[135];
    assign G[43] = in[134] & in2[134];
    assign P[43] = in[134] ^ in2[134];
    assign G[44] = in[133] & in2[133];
    assign P[44] = in[133] ^ in2[133];
    assign G[45] = in[132] & in2[132];
    assign P[45] = in[132] ^ in2[132];
    assign G[46] = in[131] & in2[131];
    assign P[46] = in[131] ^ in2[131];
    assign G[47] = in[130] & in2[130];
    assign P[47] = in[130] ^ in2[130];
    assign G[48] = in[129] & in2[129];
    assign P[48] = in[129] ^ in2[129];
    assign G[49] = in[128] & in2[128];
    assign P[49] = in[128] ^ in2[128];
    assign G[50] = in[127] & in2[127];
    assign P[50] = in[127] ^ in2[127];
    assign G[51] = in[126] & in2[126];
    assign P[51] = in[126] ^ in2[126];
    assign G[52] = in[125] & in2[125];
    assign P[52] = in[125] ^ in2[125];
    assign G[53] = in[124] & in2[124];
    assign P[53] = in[124] ^ in2[124];
    assign G[54] = in[123] & in2[123];
    assign P[54] = in[123] ^ in2[123];
    assign G[55] = in[122] & in2[122];
    assign P[55] = in[122] ^ in2[122];
    assign G[56] = in[121] & in2[121];
    assign P[56] = in[121] ^ in2[121];
    assign G[57] = in[120] & in2[120];
    assign P[57] = in[120] ^ in2[120];
    assign G[58] = in[119] & in2[119];
    assign P[58] = in[119] ^ in2[119];
    assign G[59] = in[118] & in2[118];
    assign P[59] = in[118] ^ in2[118];
    assign G[60] = in[117] & in2[117];
    assign P[60] = in[117] ^ in2[117];
    assign G[61] = in[116] & in2[116];
    assign P[61] = in[116] ^ in2[116];
    assign G[62] = in[115] & in2[115];
    assign P[62] = in[115] ^ in2[115];
    assign G[63] = in[114] & in2[114];
    assign P[63] = in[114] ^ in2[114];
    assign G[64] = in[113] & in2[113];
    assign P[64] = in[113] ^ in2[113];
    assign G[65] = in[112] & in2[112];
    assign P[65] = in[112] ^ in2[112];
    assign G[66] = in[111] & in2[111];
    assign P[66] = in[111] ^ in2[111];
    assign G[67] = in[110] & in2[110];
    assign P[67] = in[110] ^ in2[110];
    assign G[68] = in[109] & in2[109];
    assign P[68] = in[109] ^ in2[109];
    assign G[69] = in[108] & in2[108];
    assign P[69] = in[108] ^ in2[108];
    assign G[70] = in[107] & in2[107];
    assign P[70] = in[107] ^ in2[107];
    assign G[71] = in[106] & in2[106];
    assign P[71] = in[106] ^ in2[106];
    assign G[72] = in[105] & in2[105];
    assign P[72] = in[105] ^ in2[105];
    assign G[73] = in[104] & in2[104];
    assign P[73] = in[104] ^ in2[104];
    assign G[74] = in[103] & in2[103];
    assign P[74] = in[103] ^ in2[103];
    assign G[75] = in[102] & in2[102];
    assign P[75] = in[102] ^ in2[102];
    assign G[76] = in[101] & in2[101];
    assign P[76] = in[101] ^ in2[101];
    assign G[77] = in[100] & in2[100];
    assign P[77] = in[100] ^ in2[100];
    assign G[78] = in[99] & in2[99];
    assign P[78] = in[99] ^ in2[99];
    assign G[79] = in[98] & in2[98];
    assign P[79] = in[98] ^ in2[98];
    assign G[80] = in[97] & in2[97];
    assign P[80] = in[97] ^ in2[97];
    assign G[81] = in[96] & in2[96];
    assign P[81] = in[96] ^ in2[96];
    assign G[82] = in[95] & in2[95];
    assign P[82] = in[95] ^ in2[95];
    assign G[83] = in[94] & in2[94];
    assign P[83] = in[94] ^ in2[94];
    assign G[84] = in[93] & in2[93];
    assign P[84] = in[93] ^ in2[93];
    assign G[85] = in[92] & in2[92];
    assign P[85] = in[92] ^ in2[92];
    assign G[86] = in[91] & in2[91];
    assign P[86] = in[91] ^ in2[91];
    assign G[87] = in[90] & in2[90];
    assign P[87] = in[90] ^ in2[90];
    assign G[88] = in[89] & in2[89];
    assign P[88] = in[89] ^ in2[89];
    assign G[89] = in[88] & in2[88];
    assign P[89] = in[88] ^ in2[88];
    assign G[90] = in[87] & in2[87];
    assign P[90] = in[87] ^ in2[87];
    assign G[91] = in[86] & in2[86];
    assign P[91] = in[86] ^ in2[86];
    assign G[92] = in[85] & in2[85];
    assign P[92] = in[85] ^ in2[85];
    assign G[93] = in[84] & in2[84];
    assign P[93] = in[84] ^ in2[84];
    assign G[94] = in[83] & in2[83];
    assign P[94] = in[83] ^ in2[83];
    assign G[95] = in[82] & in2[82];
    assign P[95] = in[82] ^ in2[82];
    assign G[96] = in[81] & in2[81];
    assign P[96] = in[81] ^ in2[81];
    assign G[97] = in[80] & in2[80];
    assign P[97] = in[80] ^ in2[80];
    assign G[98] = in[79] & in2[79];
    assign P[98] = in[79] ^ in2[79];
    assign G[99] = in[78] & in2[78];
    assign P[99] = in[78] ^ in2[78];
    assign G[100] = in[77] & in2[77];
    assign P[100] = in[77] ^ in2[77];
    assign G[101] = in[76] & in2[76];
    assign P[101] = in[76] ^ in2[76];
    assign G[102] = in[75] & in2[75];
    assign P[102] = in[75] ^ in2[75];
    assign G[103] = in[74] & in2[74];
    assign P[103] = in[74] ^ in2[74];
    assign G[104] = in[73] & in2[73];
    assign P[104] = in[73] ^ in2[73];
    assign G[105] = in[72] & in2[72];
    assign P[105] = in[72] ^ in2[72];
    assign G[106] = in[71] & in2[71];
    assign P[106] = in[71] ^ in2[71];
    assign G[107] = in[70] & in2[70];
    assign P[107] = in[70] ^ in2[70];
    assign G[108] = in[69] & in2[69];
    assign P[108] = in[69] ^ in2[69];
    assign G[109] = in[68] & in2[68];
    assign P[109] = in[68] ^ in2[68];
    assign G[110] = in[67] & in2[67];
    assign P[110] = in[67] ^ in2[67];
    assign G[111] = in[66] & in2[66];
    assign P[111] = in[66] ^ in2[66];
    assign G[112] = in[65] & in2[65];
    assign P[112] = in[65] ^ in2[65];
    assign G[113] = in[64] & in2[64];
    assign P[113] = in[64] ^ in2[64];
    assign G[114] = in[63] & in2[63];
    assign P[114] = in[63] ^ in2[63];
    assign G[115] = in[62] & in2[62];
    assign P[115] = in[62] ^ in2[62];
    assign G[116] = in[61] & in2[61];
    assign P[116] = in[61] ^ in2[61];
    assign G[117] = in[60] & in2[60];
    assign P[117] = in[60] ^ in2[60];
    assign G[118] = in[59] & in2[59];
    assign P[118] = in[59] ^ in2[59];
    assign G[119] = in[58] & in2[58];
    assign P[119] = in[58] ^ in2[58];
    assign G[120] = in[57] & in2[57];
    assign P[120] = in[57] ^ in2[57];
    assign G[121] = in[56] & in2[56];
    assign P[121] = in[56] ^ in2[56];
    assign G[122] = in[55] & in2[55];
    assign P[122] = in[55] ^ in2[55];
    assign G[123] = in[54] & in2[54];
    assign P[123] = in[54] ^ in2[54];
    assign G[124] = in[53] & in2[53];
    assign P[124] = in[53] ^ in2[53];
    assign G[125] = in[52] & in2[52];
    assign P[125] = in[52] ^ in2[52];
    assign G[126] = in[51] & in2[51];
    assign P[126] = in[51] ^ in2[51];
    assign G[127] = in[50] & in2[50];
    assign P[127] = in[50] ^ in2[50];
    assign G[128] = in[49] & in2[49];
    assign P[128] = in[49] ^ in2[49];
    assign G[129] = in[48] & in2[48];
    assign P[129] = in[48] ^ in2[48];
    assign G[130] = in[47] & in2[47];
    assign P[130] = in[47] ^ in2[47];
    assign G[131] = in[46] & in2[46];
    assign P[131] = in[46] ^ in2[46];
    assign G[132] = in[45] & in2[45];
    assign P[132] = in[45] ^ in2[45];
    assign G[133] = in[44] & in2[44];
    assign P[133] = in[44] ^ in2[44];
    assign G[134] = in[43] & in2[43];
    assign P[134] = in[43] ^ in2[43];
    assign G[135] = in[42] & in2[42];
    assign P[135] = in[42] ^ in2[42];
    assign G[136] = in[41] & in2[41];
    assign P[136] = in[41] ^ in2[41];
    assign G[137] = in[40] & in2[40];
    assign P[137] = in[40] ^ in2[40];
    assign G[138] = in[39] & in2[39];
    assign P[138] = in[39] ^ in2[39];
    assign G[139] = in[38] & in2[38];
    assign P[139] = in[38] ^ in2[38];
    assign G[140] = in[37] & in2[37];
    assign P[140] = in[37] ^ in2[37];
    assign G[141] = in[36] & in2[36];
    assign P[141] = in[36] ^ in2[36];
    assign G[142] = in[35] & in2[35];
    assign P[142] = in[35] ^ in2[35];
    assign G[143] = in[34] & in2[34];
    assign P[143] = in[34] ^ in2[34];
    assign G[144] = in[33] & in2[33];
    assign P[144] = in[33] ^ in2[33];
    assign G[145] = in[32] & in2[32];
    assign P[145] = in[32] ^ in2[32];
    assign G[146] = in[31] & in2[31];
    assign P[146] = in[31] ^ in2[31];
    assign G[147] = in[30] & in2[30];
    assign P[147] = in[30] ^ in2[30];
    assign G[148] = in[29] & in2[29];
    assign P[148] = in[29] ^ in2[29];
    assign G[149] = in[28] & in2[28];
    assign P[149] = in[28] ^ in2[28];
    assign G[150] = in[27] & in2[27];
    assign P[150] = in[27] ^ in2[27];
    assign G[151] = in[26] & in2[26];
    assign P[151] = in[26] ^ in2[26];
    assign G[152] = in[25] & in2[25];
    assign P[152] = in[25] ^ in2[25];
    assign G[153] = in[24] & in2[24];
    assign P[153] = in[24] ^ in2[24];
    assign G[154] = in[23] & in2[23];
    assign P[154] = in[23] ^ in2[23];
    assign G[155] = in[22] & in2[22];
    assign P[155] = in[22] ^ in2[22];
    assign G[156] = in[21] & in2[21];
    assign P[156] = in[21] ^ in2[21];
    assign G[157] = in[20] & in2[20];
    assign P[157] = in[20] ^ in2[20];
    assign G[158] = in[19] & in2[19];
    assign P[158] = in[19] ^ in2[19];
    assign G[159] = in[18] & in2[18];
    assign P[159] = in[18] ^ in2[18];
    assign G[160] = in[17] & in2[17];
    assign P[160] = in[17] ^ in2[17];
    assign G[161] = in[16] & in2[16];
    assign P[161] = in[16] ^ in2[16];
    assign G[162] = in[15] & in2[15];
    assign P[162] = in[15] ^ in2[15];
    assign G[163] = in[14] & in2[14];
    assign P[163] = in[14] ^ in2[14];
    assign G[164] = in[13] & in2[13];
    assign P[164] = in[13] ^ in2[13];
    assign G[165] = in[12] & in2[12];
    assign P[165] = in[12] ^ in2[12];
    assign G[166] = in[11] & in2[11];
    assign P[166] = in[11] ^ in2[11];
    assign G[167] = in[10] & in2[10];
    assign P[167] = in[10] ^ in2[10];
    assign G[168] = in[9] & in2[9];
    assign P[168] = in[9] ^ in2[9];
    assign G[169] = in[8] & in2[8];
    assign P[169] = in[8] ^ in2[8];
    assign G[170] = in[7] & in2[7];
    assign P[170] = in[7] ^ in2[7];
    assign G[171] = in[6] & in2[6];
    assign P[171] = in[6] ^ in2[6];
    assign G[172] = in[5] & in2[5];
    assign P[172] = in[5] ^ in2[5];
    assign G[173] = in[4] & in2[4];
    assign P[173] = in[4] ^ in2[4];
    assign G[174] = in[3] & in2[3];
    assign P[174] = in[3] ^ in2[3];
    assign G[175] = in[2] & in2[2];
    assign P[175] = in[2] ^ in2[2];
    assign G[176] = in[1] & in2[1];
    assign P[176] = in[1] ^ in2[1];
    assign G[177] = in[0] & in2[0];
    assign P[177] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign C[177] = G[176] | (P[176] & C[176]);
    assign cout = G[177] | (P[177] & C[177]);
    assign sum = P ^ C;
endmodule

module CLA177(output [176:0] sum, output cout, input [176:0] in1, input [176:0] in2;

    wire[176:0] G;
    wire[176:0] C;
    wire[176:0] P;

    assign G[0] = in[176] & in2[176];
    assign P[0] = in[176] ^ in2[176];
    assign G[1] = in[175] & in2[175];
    assign P[1] = in[175] ^ in2[175];
    assign G[2] = in[174] & in2[174];
    assign P[2] = in[174] ^ in2[174];
    assign G[3] = in[173] & in2[173];
    assign P[3] = in[173] ^ in2[173];
    assign G[4] = in[172] & in2[172];
    assign P[4] = in[172] ^ in2[172];
    assign G[5] = in[171] & in2[171];
    assign P[5] = in[171] ^ in2[171];
    assign G[6] = in[170] & in2[170];
    assign P[6] = in[170] ^ in2[170];
    assign G[7] = in[169] & in2[169];
    assign P[7] = in[169] ^ in2[169];
    assign G[8] = in[168] & in2[168];
    assign P[8] = in[168] ^ in2[168];
    assign G[9] = in[167] & in2[167];
    assign P[9] = in[167] ^ in2[167];
    assign G[10] = in[166] & in2[166];
    assign P[10] = in[166] ^ in2[166];
    assign G[11] = in[165] & in2[165];
    assign P[11] = in[165] ^ in2[165];
    assign G[12] = in[164] & in2[164];
    assign P[12] = in[164] ^ in2[164];
    assign G[13] = in[163] & in2[163];
    assign P[13] = in[163] ^ in2[163];
    assign G[14] = in[162] & in2[162];
    assign P[14] = in[162] ^ in2[162];
    assign G[15] = in[161] & in2[161];
    assign P[15] = in[161] ^ in2[161];
    assign G[16] = in[160] & in2[160];
    assign P[16] = in[160] ^ in2[160];
    assign G[17] = in[159] & in2[159];
    assign P[17] = in[159] ^ in2[159];
    assign G[18] = in[158] & in2[158];
    assign P[18] = in[158] ^ in2[158];
    assign G[19] = in[157] & in2[157];
    assign P[19] = in[157] ^ in2[157];
    assign G[20] = in[156] & in2[156];
    assign P[20] = in[156] ^ in2[156];
    assign G[21] = in[155] & in2[155];
    assign P[21] = in[155] ^ in2[155];
    assign G[22] = in[154] & in2[154];
    assign P[22] = in[154] ^ in2[154];
    assign G[23] = in[153] & in2[153];
    assign P[23] = in[153] ^ in2[153];
    assign G[24] = in[152] & in2[152];
    assign P[24] = in[152] ^ in2[152];
    assign G[25] = in[151] & in2[151];
    assign P[25] = in[151] ^ in2[151];
    assign G[26] = in[150] & in2[150];
    assign P[26] = in[150] ^ in2[150];
    assign G[27] = in[149] & in2[149];
    assign P[27] = in[149] ^ in2[149];
    assign G[28] = in[148] & in2[148];
    assign P[28] = in[148] ^ in2[148];
    assign G[29] = in[147] & in2[147];
    assign P[29] = in[147] ^ in2[147];
    assign G[30] = in[146] & in2[146];
    assign P[30] = in[146] ^ in2[146];
    assign G[31] = in[145] & in2[145];
    assign P[31] = in[145] ^ in2[145];
    assign G[32] = in[144] & in2[144];
    assign P[32] = in[144] ^ in2[144];
    assign G[33] = in[143] & in2[143];
    assign P[33] = in[143] ^ in2[143];
    assign G[34] = in[142] & in2[142];
    assign P[34] = in[142] ^ in2[142];
    assign G[35] = in[141] & in2[141];
    assign P[35] = in[141] ^ in2[141];
    assign G[36] = in[140] & in2[140];
    assign P[36] = in[140] ^ in2[140];
    assign G[37] = in[139] & in2[139];
    assign P[37] = in[139] ^ in2[139];
    assign G[38] = in[138] & in2[138];
    assign P[38] = in[138] ^ in2[138];
    assign G[39] = in[137] & in2[137];
    assign P[39] = in[137] ^ in2[137];
    assign G[40] = in[136] & in2[136];
    assign P[40] = in[136] ^ in2[136];
    assign G[41] = in[135] & in2[135];
    assign P[41] = in[135] ^ in2[135];
    assign G[42] = in[134] & in2[134];
    assign P[42] = in[134] ^ in2[134];
    assign G[43] = in[133] & in2[133];
    assign P[43] = in[133] ^ in2[133];
    assign G[44] = in[132] & in2[132];
    assign P[44] = in[132] ^ in2[132];
    assign G[45] = in[131] & in2[131];
    assign P[45] = in[131] ^ in2[131];
    assign G[46] = in[130] & in2[130];
    assign P[46] = in[130] ^ in2[130];
    assign G[47] = in[129] & in2[129];
    assign P[47] = in[129] ^ in2[129];
    assign G[48] = in[128] & in2[128];
    assign P[48] = in[128] ^ in2[128];
    assign G[49] = in[127] & in2[127];
    assign P[49] = in[127] ^ in2[127];
    assign G[50] = in[126] & in2[126];
    assign P[50] = in[126] ^ in2[126];
    assign G[51] = in[125] & in2[125];
    assign P[51] = in[125] ^ in2[125];
    assign G[52] = in[124] & in2[124];
    assign P[52] = in[124] ^ in2[124];
    assign G[53] = in[123] & in2[123];
    assign P[53] = in[123] ^ in2[123];
    assign G[54] = in[122] & in2[122];
    assign P[54] = in[122] ^ in2[122];
    assign G[55] = in[121] & in2[121];
    assign P[55] = in[121] ^ in2[121];
    assign G[56] = in[120] & in2[120];
    assign P[56] = in[120] ^ in2[120];
    assign G[57] = in[119] & in2[119];
    assign P[57] = in[119] ^ in2[119];
    assign G[58] = in[118] & in2[118];
    assign P[58] = in[118] ^ in2[118];
    assign G[59] = in[117] & in2[117];
    assign P[59] = in[117] ^ in2[117];
    assign G[60] = in[116] & in2[116];
    assign P[60] = in[116] ^ in2[116];
    assign G[61] = in[115] & in2[115];
    assign P[61] = in[115] ^ in2[115];
    assign G[62] = in[114] & in2[114];
    assign P[62] = in[114] ^ in2[114];
    assign G[63] = in[113] & in2[113];
    assign P[63] = in[113] ^ in2[113];
    assign G[64] = in[112] & in2[112];
    assign P[64] = in[112] ^ in2[112];
    assign G[65] = in[111] & in2[111];
    assign P[65] = in[111] ^ in2[111];
    assign G[66] = in[110] & in2[110];
    assign P[66] = in[110] ^ in2[110];
    assign G[67] = in[109] & in2[109];
    assign P[67] = in[109] ^ in2[109];
    assign G[68] = in[108] & in2[108];
    assign P[68] = in[108] ^ in2[108];
    assign G[69] = in[107] & in2[107];
    assign P[69] = in[107] ^ in2[107];
    assign G[70] = in[106] & in2[106];
    assign P[70] = in[106] ^ in2[106];
    assign G[71] = in[105] & in2[105];
    assign P[71] = in[105] ^ in2[105];
    assign G[72] = in[104] & in2[104];
    assign P[72] = in[104] ^ in2[104];
    assign G[73] = in[103] & in2[103];
    assign P[73] = in[103] ^ in2[103];
    assign G[74] = in[102] & in2[102];
    assign P[74] = in[102] ^ in2[102];
    assign G[75] = in[101] & in2[101];
    assign P[75] = in[101] ^ in2[101];
    assign G[76] = in[100] & in2[100];
    assign P[76] = in[100] ^ in2[100];
    assign G[77] = in[99] & in2[99];
    assign P[77] = in[99] ^ in2[99];
    assign G[78] = in[98] & in2[98];
    assign P[78] = in[98] ^ in2[98];
    assign G[79] = in[97] & in2[97];
    assign P[79] = in[97] ^ in2[97];
    assign G[80] = in[96] & in2[96];
    assign P[80] = in[96] ^ in2[96];
    assign G[81] = in[95] & in2[95];
    assign P[81] = in[95] ^ in2[95];
    assign G[82] = in[94] & in2[94];
    assign P[82] = in[94] ^ in2[94];
    assign G[83] = in[93] & in2[93];
    assign P[83] = in[93] ^ in2[93];
    assign G[84] = in[92] & in2[92];
    assign P[84] = in[92] ^ in2[92];
    assign G[85] = in[91] & in2[91];
    assign P[85] = in[91] ^ in2[91];
    assign G[86] = in[90] & in2[90];
    assign P[86] = in[90] ^ in2[90];
    assign G[87] = in[89] & in2[89];
    assign P[87] = in[89] ^ in2[89];
    assign G[88] = in[88] & in2[88];
    assign P[88] = in[88] ^ in2[88];
    assign G[89] = in[87] & in2[87];
    assign P[89] = in[87] ^ in2[87];
    assign G[90] = in[86] & in2[86];
    assign P[90] = in[86] ^ in2[86];
    assign G[91] = in[85] & in2[85];
    assign P[91] = in[85] ^ in2[85];
    assign G[92] = in[84] & in2[84];
    assign P[92] = in[84] ^ in2[84];
    assign G[93] = in[83] & in2[83];
    assign P[93] = in[83] ^ in2[83];
    assign G[94] = in[82] & in2[82];
    assign P[94] = in[82] ^ in2[82];
    assign G[95] = in[81] & in2[81];
    assign P[95] = in[81] ^ in2[81];
    assign G[96] = in[80] & in2[80];
    assign P[96] = in[80] ^ in2[80];
    assign G[97] = in[79] & in2[79];
    assign P[97] = in[79] ^ in2[79];
    assign G[98] = in[78] & in2[78];
    assign P[98] = in[78] ^ in2[78];
    assign G[99] = in[77] & in2[77];
    assign P[99] = in[77] ^ in2[77];
    assign G[100] = in[76] & in2[76];
    assign P[100] = in[76] ^ in2[76];
    assign G[101] = in[75] & in2[75];
    assign P[101] = in[75] ^ in2[75];
    assign G[102] = in[74] & in2[74];
    assign P[102] = in[74] ^ in2[74];
    assign G[103] = in[73] & in2[73];
    assign P[103] = in[73] ^ in2[73];
    assign G[104] = in[72] & in2[72];
    assign P[104] = in[72] ^ in2[72];
    assign G[105] = in[71] & in2[71];
    assign P[105] = in[71] ^ in2[71];
    assign G[106] = in[70] & in2[70];
    assign P[106] = in[70] ^ in2[70];
    assign G[107] = in[69] & in2[69];
    assign P[107] = in[69] ^ in2[69];
    assign G[108] = in[68] & in2[68];
    assign P[108] = in[68] ^ in2[68];
    assign G[109] = in[67] & in2[67];
    assign P[109] = in[67] ^ in2[67];
    assign G[110] = in[66] & in2[66];
    assign P[110] = in[66] ^ in2[66];
    assign G[111] = in[65] & in2[65];
    assign P[111] = in[65] ^ in2[65];
    assign G[112] = in[64] & in2[64];
    assign P[112] = in[64] ^ in2[64];
    assign G[113] = in[63] & in2[63];
    assign P[113] = in[63] ^ in2[63];
    assign G[114] = in[62] & in2[62];
    assign P[114] = in[62] ^ in2[62];
    assign G[115] = in[61] & in2[61];
    assign P[115] = in[61] ^ in2[61];
    assign G[116] = in[60] & in2[60];
    assign P[116] = in[60] ^ in2[60];
    assign G[117] = in[59] & in2[59];
    assign P[117] = in[59] ^ in2[59];
    assign G[118] = in[58] & in2[58];
    assign P[118] = in[58] ^ in2[58];
    assign G[119] = in[57] & in2[57];
    assign P[119] = in[57] ^ in2[57];
    assign G[120] = in[56] & in2[56];
    assign P[120] = in[56] ^ in2[56];
    assign G[121] = in[55] & in2[55];
    assign P[121] = in[55] ^ in2[55];
    assign G[122] = in[54] & in2[54];
    assign P[122] = in[54] ^ in2[54];
    assign G[123] = in[53] & in2[53];
    assign P[123] = in[53] ^ in2[53];
    assign G[124] = in[52] & in2[52];
    assign P[124] = in[52] ^ in2[52];
    assign G[125] = in[51] & in2[51];
    assign P[125] = in[51] ^ in2[51];
    assign G[126] = in[50] & in2[50];
    assign P[126] = in[50] ^ in2[50];
    assign G[127] = in[49] & in2[49];
    assign P[127] = in[49] ^ in2[49];
    assign G[128] = in[48] & in2[48];
    assign P[128] = in[48] ^ in2[48];
    assign G[129] = in[47] & in2[47];
    assign P[129] = in[47] ^ in2[47];
    assign G[130] = in[46] & in2[46];
    assign P[130] = in[46] ^ in2[46];
    assign G[131] = in[45] & in2[45];
    assign P[131] = in[45] ^ in2[45];
    assign G[132] = in[44] & in2[44];
    assign P[132] = in[44] ^ in2[44];
    assign G[133] = in[43] & in2[43];
    assign P[133] = in[43] ^ in2[43];
    assign G[134] = in[42] & in2[42];
    assign P[134] = in[42] ^ in2[42];
    assign G[135] = in[41] & in2[41];
    assign P[135] = in[41] ^ in2[41];
    assign G[136] = in[40] & in2[40];
    assign P[136] = in[40] ^ in2[40];
    assign G[137] = in[39] & in2[39];
    assign P[137] = in[39] ^ in2[39];
    assign G[138] = in[38] & in2[38];
    assign P[138] = in[38] ^ in2[38];
    assign G[139] = in[37] & in2[37];
    assign P[139] = in[37] ^ in2[37];
    assign G[140] = in[36] & in2[36];
    assign P[140] = in[36] ^ in2[36];
    assign G[141] = in[35] & in2[35];
    assign P[141] = in[35] ^ in2[35];
    assign G[142] = in[34] & in2[34];
    assign P[142] = in[34] ^ in2[34];
    assign G[143] = in[33] & in2[33];
    assign P[143] = in[33] ^ in2[33];
    assign G[144] = in[32] & in2[32];
    assign P[144] = in[32] ^ in2[32];
    assign G[145] = in[31] & in2[31];
    assign P[145] = in[31] ^ in2[31];
    assign G[146] = in[30] & in2[30];
    assign P[146] = in[30] ^ in2[30];
    assign G[147] = in[29] & in2[29];
    assign P[147] = in[29] ^ in2[29];
    assign G[148] = in[28] & in2[28];
    assign P[148] = in[28] ^ in2[28];
    assign G[149] = in[27] & in2[27];
    assign P[149] = in[27] ^ in2[27];
    assign G[150] = in[26] & in2[26];
    assign P[150] = in[26] ^ in2[26];
    assign G[151] = in[25] & in2[25];
    assign P[151] = in[25] ^ in2[25];
    assign G[152] = in[24] & in2[24];
    assign P[152] = in[24] ^ in2[24];
    assign G[153] = in[23] & in2[23];
    assign P[153] = in[23] ^ in2[23];
    assign G[154] = in[22] & in2[22];
    assign P[154] = in[22] ^ in2[22];
    assign G[155] = in[21] & in2[21];
    assign P[155] = in[21] ^ in2[21];
    assign G[156] = in[20] & in2[20];
    assign P[156] = in[20] ^ in2[20];
    assign G[157] = in[19] & in2[19];
    assign P[157] = in[19] ^ in2[19];
    assign G[158] = in[18] & in2[18];
    assign P[158] = in[18] ^ in2[18];
    assign G[159] = in[17] & in2[17];
    assign P[159] = in[17] ^ in2[17];
    assign G[160] = in[16] & in2[16];
    assign P[160] = in[16] ^ in2[16];
    assign G[161] = in[15] & in2[15];
    assign P[161] = in[15] ^ in2[15];
    assign G[162] = in[14] & in2[14];
    assign P[162] = in[14] ^ in2[14];
    assign G[163] = in[13] & in2[13];
    assign P[163] = in[13] ^ in2[13];
    assign G[164] = in[12] & in2[12];
    assign P[164] = in[12] ^ in2[12];
    assign G[165] = in[11] & in2[11];
    assign P[165] = in[11] ^ in2[11];
    assign G[166] = in[10] & in2[10];
    assign P[166] = in[10] ^ in2[10];
    assign G[167] = in[9] & in2[9];
    assign P[167] = in[9] ^ in2[9];
    assign G[168] = in[8] & in2[8];
    assign P[168] = in[8] ^ in2[8];
    assign G[169] = in[7] & in2[7];
    assign P[169] = in[7] ^ in2[7];
    assign G[170] = in[6] & in2[6];
    assign P[170] = in[6] ^ in2[6];
    assign G[171] = in[5] & in2[5];
    assign P[171] = in[5] ^ in2[5];
    assign G[172] = in[4] & in2[4];
    assign P[172] = in[4] ^ in2[4];
    assign G[173] = in[3] & in2[3];
    assign P[173] = in[3] ^ in2[3];
    assign G[174] = in[2] & in2[2];
    assign P[174] = in[2] ^ in2[2];
    assign G[175] = in[1] & in2[1];
    assign P[175] = in[1] ^ in2[1];
    assign G[176] = in[0] & in2[0];
    assign P[176] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign C[176] = G[175] | (P[175] & C[175]);
    assign cout = G[176] | (P[176] & C[176]);
    assign sum = P ^ C;
endmodule

module CLA176(output [175:0] sum, output cout, input [175:0] in1, input [175:0] in2;

    wire[175:0] G;
    wire[175:0] C;
    wire[175:0] P;

    assign G[0] = in[175] & in2[175];
    assign P[0] = in[175] ^ in2[175];
    assign G[1] = in[174] & in2[174];
    assign P[1] = in[174] ^ in2[174];
    assign G[2] = in[173] & in2[173];
    assign P[2] = in[173] ^ in2[173];
    assign G[3] = in[172] & in2[172];
    assign P[3] = in[172] ^ in2[172];
    assign G[4] = in[171] & in2[171];
    assign P[4] = in[171] ^ in2[171];
    assign G[5] = in[170] & in2[170];
    assign P[5] = in[170] ^ in2[170];
    assign G[6] = in[169] & in2[169];
    assign P[6] = in[169] ^ in2[169];
    assign G[7] = in[168] & in2[168];
    assign P[7] = in[168] ^ in2[168];
    assign G[8] = in[167] & in2[167];
    assign P[8] = in[167] ^ in2[167];
    assign G[9] = in[166] & in2[166];
    assign P[9] = in[166] ^ in2[166];
    assign G[10] = in[165] & in2[165];
    assign P[10] = in[165] ^ in2[165];
    assign G[11] = in[164] & in2[164];
    assign P[11] = in[164] ^ in2[164];
    assign G[12] = in[163] & in2[163];
    assign P[12] = in[163] ^ in2[163];
    assign G[13] = in[162] & in2[162];
    assign P[13] = in[162] ^ in2[162];
    assign G[14] = in[161] & in2[161];
    assign P[14] = in[161] ^ in2[161];
    assign G[15] = in[160] & in2[160];
    assign P[15] = in[160] ^ in2[160];
    assign G[16] = in[159] & in2[159];
    assign P[16] = in[159] ^ in2[159];
    assign G[17] = in[158] & in2[158];
    assign P[17] = in[158] ^ in2[158];
    assign G[18] = in[157] & in2[157];
    assign P[18] = in[157] ^ in2[157];
    assign G[19] = in[156] & in2[156];
    assign P[19] = in[156] ^ in2[156];
    assign G[20] = in[155] & in2[155];
    assign P[20] = in[155] ^ in2[155];
    assign G[21] = in[154] & in2[154];
    assign P[21] = in[154] ^ in2[154];
    assign G[22] = in[153] & in2[153];
    assign P[22] = in[153] ^ in2[153];
    assign G[23] = in[152] & in2[152];
    assign P[23] = in[152] ^ in2[152];
    assign G[24] = in[151] & in2[151];
    assign P[24] = in[151] ^ in2[151];
    assign G[25] = in[150] & in2[150];
    assign P[25] = in[150] ^ in2[150];
    assign G[26] = in[149] & in2[149];
    assign P[26] = in[149] ^ in2[149];
    assign G[27] = in[148] & in2[148];
    assign P[27] = in[148] ^ in2[148];
    assign G[28] = in[147] & in2[147];
    assign P[28] = in[147] ^ in2[147];
    assign G[29] = in[146] & in2[146];
    assign P[29] = in[146] ^ in2[146];
    assign G[30] = in[145] & in2[145];
    assign P[30] = in[145] ^ in2[145];
    assign G[31] = in[144] & in2[144];
    assign P[31] = in[144] ^ in2[144];
    assign G[32] = in[143] & in2[143];
    assign P[32] = in[143] ^ in2[143];
    assign G[33] = in[142] & in2[142];
    assign P[33] = in[142] ^ in2[142];
    assign G[34] = in[141] & in2[141];
    assign P[34] = in[141] ^ in2[141];
    assign G[35] = in[140] & in2[140];
    assign P[35] = in[140] ^ in2[140];
    assign G[36] = in[139] & in2[139];
    assign P[36] = in[139] ^ in2[139];
    assign G[37] = in[138] & in2[138];
    assign P[37] = in[138] ^ in2[138];
    assign G[38] = in[137] & in2[137];
    assign P[38] = in[137] ^ in2[137];
    assign G[39] = in[136] & in2[136];
    assign P[39] = in[136] ^ in2[136];
    assign G[40] = in[135] & in2[135];
    assign P[40] = in[135] ^ in2[135];
    assign G[41] = in[134] & in2[134];
    assign P[41] = in[134] ^ in2[134];
    assign G[42] = in[133] & in2[133];
    assign P[42] = in[133] ^ in2[133];
    assign G[43] = in[132] & in2[132];
    assign P[43] = in[132] ^ in2[132];
    assign G[44] = in[131] & in2[131];
    assign P[44] = in[131] ^ in2[131];
    assign G[45] = in[130] & in2[130];
    assign P[45] = in[130] ^ in2[130];
    assign G[46] = in[129] & in2[129];
    assign P[46] = in[129] ^ in2[129];
    assign G[47] = in[128] & in2[128];
    assign P[47] = in[128] ^ in2[128];
    assign G[48] = in[127] & in2[127];
    assign P[48] = in[127] ^ in2[127];
    assign G[49] = in[126] & in2[126];
    assign P[49] = in[126] ^ in2[126];
    assign G[50] = in[125] & in2[125];
    assign P[50] = in[125] ^ in2[125];
    assign G[51] = in[124] & in2[124];
    assign P[51] = in[124] ^ in2[124];
    assign G[52] = in[123] & in2[123];
    assign P[52] = in[123] ^ in2[123];
    assign G[53] = in[122] & in2[122];
    assign P[53] = in[122] ^ in2[122];
    assign G[54] = in[121] & in2[121];
    assign P[54] = in[121] ^ in2[121];
    assign G[55] = in[120] & in2[120];
    assign P[55] = in[120] ^ in2[120];
    assign G[56] = in[119] & in2[119];
    assign P[56] = in[119] ^ in2[119];
    assign G[57] = in[118] & in2[118];
    assign P[57] = in[118] ^ in2[118];
    assign G[58] = in[117] & in2[117];
    assign P[58] = in[117] ^ in2[117];
    assign G[59] = in[116] & in2[116];
    assign P[59] = in[116] ^ in2[116];
    assign G[60] = in[115] & in2[115];
    assign P[60] = in[115] ^ in2[115];
    assign G[61] = in[114] & in2[114];
    assign P[61] = in[114] ^ in2[114];
    assign G[62] = in[113] & in2[113];
    assign P[62] = in[113] ^ in2[113];
    assign G[63] = in[112] & in2[112];
    assign P[63] = in[112] ^ in2[112];
    assign G[64] = in[111] & in2[111];
    assign P[64] = in[111] ^ in2[111];
    assign G[65] = in[110] & in2[110];
    assign P[65] = in[110] ^ in2[110];
    assign G[66] = in[109] & in2[109];
    assign P[66] = in[109] ^ in2[109];
    assign G[67] = in[108] & in2[108];
    assign P[67] = in[108] ^ in2[108];
    assign G[68] = in[107] & in2[107];
    assign P[68] = in[107] ^ in2[107];
    assign G[69] = in[106] & in2[106];
    assign P[69] = in[106] ^ in2[106];
    assign G[70] = in[105] & in2[105];
    assign P[70] = in[105] ^ in2[105];
    assign G[71] = in[104] & in2[104];
    assign P[71] = in[104] ^ in2[104];
    assign G[72] = in[103] & in2[103];
    assign P[72] = in[103] ^ in2[103];
    assign G[73] = in[102] & in2[102];
    assign P[73] = in[102] ^ in2[102];
    assign G[74] = in[101] & in2[101];
    assign P[74] = in[101] ^ in2[101];
    assign G[75] = in[100] & in2[100];
    assign P[75] = in[100] ^ in2[100];
    assign G[76] = in[99] & in2[99];
    assign P[76] = in[99] ^ in2[99];
    assign G[77] = in[98] & in2[98];
    assign P[77] = in[98] ^ in2[98];
    assign G[78] = in[97] & in2[97];
    assign P[78] = in[97] ^ in2[97];
    assign G[79] = in[96] & in2[96];
    assign P[79] = in[96] ^ in2[96];
    assign G[80] = in[95] & in2[95];
    assign P[80] = in[95] ^ in2[95];
    assign G[81] = in[94] & in2[94];
    assign P[81] = in[94] ^ in2[94];
    assign G[82] = in[93] & in2[93];
    assign P[82] = in[93] ^ in2[93];
    assign G[83] = in[92] & in2[92];
    assign P[83] = in[92] ^ in2[92];
    assign G[84] = in[91] & in2[91];
    assign P[84] = in[91] ^ in2[91];
    assign G[85] = in[90] & in2[90];
    assign P[85] = in[90] ^ in2[90];
    assign G[86] = in[89] & in2[89];
    assign P[86] = in[89] ^ in2[89];
    assign G[87] = in[88] & in2[88];
    assign P[87] = in[88] ^ in2[88];
    assign G[88] = in[87] & in2[87];
    assign P[88] = in[87] ^ in2[87];
    assign G[89] = in[86] & in2[86];
    assign P[89] = in[86] ^ in2[86];
    assign G[90] = in[85] & in2[85];
    assign P[90] = in[85] ^ in2[85];
    assign G[91] = in[84] & in2[84];
    assign P[91] = in[84] ^ in2[84];
    assign G[92] = in[83] & in2[83];
    assign P[92] = in[83] ^ in2[83];
    assign G[93] = in[82] & in2[82];
    assign P[93] = in[82] ^ in2[82];
    assign G[94] = in[81] & in2[81];
    assign P[94] = in[81] ^ in2[81];
    assign G[95] = in[80] & in2[80];
    assign P[95] = in[80] ^ in2[80];
    assign G[96] = in[79] & in2[79];
    assign P[96] = in[79] ^ in2[79];
    assign G[97] = in[78] & in2[78];
    assign P[97] = in[78] ^ in2[78];
    assign G[98] = in[77] & in2[77];
    assign P[98] = in[77] ^ in2[77];
    assign G[99] = in[76] & in2[76];
    assign P[99] = in[76] ^ in2[76];
    assign G[100] = in[75] & in2[75];
    assign P[100] = in[75] ^ in2[75];
    assign G[101] = in[74] & in2[74];
    assign P[101] = in[74] ^ in2[74];
    assign G[102] = in[73] & in2[73];
    assign P[102] = in[73] ^ in2[73];
    assign G[103] = in[72] & in2[72];
    assign P[103] = in[72] ^ in2[72];
    assign G[104] = in[71] & in2[71];
    assign P[104] = in[71] ^ in2[71];
    assign G[105] = in[70] & in2[70];
    assign P[105] = in[70] ^ in2[70];
    assign G[106] = in[69] & in2[69];
    assign P[106] = in[69] ^ in2[69];
    assign G[107] = in[68] & in2[68];
    assign P[107] = in[68] ^ in2[68];
    assign G[108] = in[67] & in2[67];
    assign P[108] = in[67] ^ in2[67];
    assign G[109] = in[66] & in2[66];
    assign P[109] = in[66] ^ in2[66];
    assign G[110] = in[65] & in2[65];
    assign P[110] = in[65] ^ in2[65];
    assign G[111] = in[64] & in2[64];
    assign P[111] = in[64] ^ in2[64];
    assign G[112] = in[63] & in2[63];
    assign P[112] = in[63] ^ in2[63];
    assign G[113] = in[62] & in2[62];
    assign P[113] = in[62] ^ in2[62];
    assign G[114] = in[61] & in2[61];
    assign P[114] = in[61] ^ in2[61];
    assign G[115] = in[60] & in2[60];
    assign P[115] = in[60] ^ in2[60];
    assign G[116] = in[59] & in2[59];
    assign P[116] = in[59] ^ in2[59];
    assign G[117] = in[58] & in2[58];
    assign P[117] = in[58] ^ in2[58];
    assign G[118] = in[57] & in2[57];
    assign P[118] = in[57] ^ in2[57];
    assign G[119] = in[56] & in2[56];
    assign P[119] = in[56] ^ in2[56];
    assign G[120] = in[55] & in2[55];
    assign P[120] = in[55] ^ in2[55];
    assign G[121] = in[54] & in2[54];
    assign P[121] = in[54] ^ in2[54];
    assign G[122] = in[53] & in2[53];
    assign P[122] = in[53] ^ in2[53];
    assign G[123] = in[52] & in2[52];
    assign P[123] = in[52] ^ in2[52];
    assign G[124] = in[51] & in2[51];
    assign P[124] = in[51] ^ in2[51];
    assign G[125] = in[50] & in2[50];
    assign P[125] = in[50] ^ in2[50];
    assign G[126] = in[49] & in2[49];
    assign P[126] = in[49] ^ in2[49];
    assign G[127] = in[48] & in2[48];
    assign P[127] = in[48] ^ in2[48];
    assign G[128] = in[47] & in2[47];
    assign P[128] = in[47] ^ in2[47];
    assign G[129] = in[46] & in2[46];
    assign P[129] = in[46] ^ in2[46];
    assign G[130] = in[45] & in2[45];
    assign P[130] = in[45] ^ in2[45];
    assign G[131] = in[44] & in2[44];
    assign P[131] = in[44] ^ in2[44];
    assign G[132] = in[43] & in2[43];
    assign P[132] = in[43] ^ in2[43];
    assign G[133] = in[42] & in2[42];
    assign P[133] = in[42] ^ in2[42];
    assign G[134] = in[41] & in2[41];
    assign P[134] = in[41] ^ in2[41];
    assign G[135] = in[40] & in2[40];
    assign P[135] = in[40] ^ in2[40];
    assign G[136] = in[39] & in2[39];
    assign P[136] = in[39] ^ in2[39];
    assign G[137] = in[38] & in2[38];
    assign P[137] = in[38] ^ in2[38];
    assign G[138] = in[37] & in2[37];
    assign P[138] = in[37] ^ in2[37];
    assign G[139] = in[36] & in2[36];
    assign P[139] = in[36] ^ in2[36];
    assign G[140] = in[35] & in2[35];
    assign P[140] = in[35] ^ in2[35];
    assign G[141] = in[34] & in2[34];
    assign P[141] = in[34] ^ in2[34];
    assign G[142] = in[33] & in2[33];
    assign P[142] = in[33] ^ in2[33];
    assign G[143] = in[32] & in2[32];
    assign P[143] = in[32] ^ in2[32];
    assign G[144] = in[31] & in2[31];
    assign P[144] = in[31] ^ in2[31];
    assign G[145] = in[30] & in2[30];
    assign P[145] = in[30] ^ in2[30];
    assign G[146] = in[29] & in2[29];
    assign P[146] = in[29] ^ in2[29];
    assign G[147] = in[28] & in2[28];
    assign P[147] = in[28] ^ in2[28];
    assign G[148] = in[27] & in2[27];
    assign P[148] = in[27] ^ in2[27];
    assign G[149] = in[26] & in2[26];
    assign P[149] = in[26] ^ in2[26];
    assign G[150] = in[25] & in2[25];
    assign P[150] = in[25] ^ in2[25];
    assign G[151] = in[24] & in2[24];
    assign P[151] = in[24] ^ in2[24];
    assign G[152] = in[23] & in2[23];
    assign P[152] = in[23] ^ in2[23];
    assign G[153] = in[22] & in2[22];
    assign P[153] = in[22] ^ in2[22];
    assign G[154] = in[21] & in2[21];
    assign P[154] = in[21] ^ in2[21];
    assign G[155] = in[20] & in2[20];
    assign P[155] = in[20] ^ in2[20];
    assign G[156] = in[19] & in2[19];
    assign P[156] = in[19] ^ in2[19];
    assign G[157] = in[18] & in2[18];
    assign P[157] = in[18] ^ in2[18];
    assign G[158] = in[17] & in2[17];
    assign P[158] = in[17] ^ in2[17];
    assign G[159] = in[16] & in2[16];
    assign P[159] = in[16] ^ in2[16];
    assign G[160] = in[15] & in2[15];
    assign P[160] = in[15] ^ in2[15];
    assign G[161] = in[14] & in2[14];
    assign P[161] = in[14] ^ in2[14];
    assign G[162] = in[13] & in2[13];
    assign P[162] = in[13] ^ in2[13];
    assign G[163] = in[12] & in2[12];
    assign P[163] = in[12] ^ in2[12];
    assign G[164] = in[11] & in2[11];
    assign P[164] = in[11] ^ in2[11];
    assign G[165] = in[10] & in2[10];
    assign P[165] = in[10] ^ in2[10];
    assign G[166] = in[9] & in2[9];
    assign P[166] = in[9] ^ in2[9];
    assign G[167] = in[8] & in2[8];
    assign P[167] = in[8] ^ in2[8];
    assign G[168] = in[7] & in2[7];
    assign P[168] = in[7] ^ in2[7];
    assign G[169] = in[6] & in2[6];
    assign P[169] = in[6] ^ in2[6];
    assign G[170] = in[5] & in2[5];
    assign P[170] = in[5] ^ in2[5];
    assign G[171] = in[4] & in2[4];
    assign P[171] = in[4] ^ in2[4];
    assign G[172] = in[3] & in2[3];
    assign P[172] = in[3] ^ in2[3];
    assign G[173] = in[2] & in2[2];
    assign P[173] = in[2] ^ in2[2];
    assign G[174] = in[1] & in2[1];
    assign P[174] = in[1] ^ in2[1];
    assign G[175] = in[0] & in2[0];
    assign P[175] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign C[175] = G[174] | (P[174] & C[174]);
    assign cout = G[175] | (P[175] & C[175]);
    assign sum = P ^ C;
endmodule

module CLA175(output [174:0] sum, output cout, input [174:0] in1, input [174:0] in2;

    wire[174:0] G;
    wire[174:0] C;
    wire[174:0] P;

    assign G[0] = in[174] & in2[174];
    assign P[0] = in[174] ^ in2[174];
    assign G[1] = in[173] & in2[173];
    assign P[1] = in[173] ^ in2[173];
    assign G[2] = in[172] & in2[172];
    assign P[2] = in[172] ^ in2[172];
    assign G[3] = in[171] & in2[171];
    assign P[3] = in[171] ^ in2[171];
    assign G[4] = in[170] & in2[170];
    assign P[4] = in[170] ^ in2[170];
    assign G[5] = in[169] & in2[169];
    assign P[5] = in[169] ^ in2[169];
    assign G[6] = in[168] & in2[168];
    assign P[6] = in[168] ^ in2[168];
    assign G[7] = in[167] & in2[167];
    assign P[7] = in[167] ^ in2[167];
    assign G[8] = in[166] & in2[166];
    assign P[8] = in[166] ^ in2[166];
    assign G[9] = in[165] & in2[165];
    assign P[9] = in[165] ^ in2[165];
    assign G[10] = in[164] & in2[164];
    assign P[10] = in[164] ^ in2[164];
    assign G[11] = in[163] & in2[163];
    assign P[11] = in[163] ^ in2[163];
    assign G[12] = in[162] & in2[162];
    assign P[12] = in[162] ^ in2[162];
    assign G[13] = in[161] & in2[161];
    assign P[13] = in[161] ^ in2[161];
    assign G[14] = in[160] & in2[160];
    assign P[14] = in[160] ^ in2[160];
    assign G[15] = in[159] & in2[159];
    assign P[15] = in[159] ^ in2[159];
    assign G[16] = in[158] & in2[158];
    assign P[16] = in[158] ^ in2[158];
    assign G[17] = in[157] & in2[157];
    assign P[17] = in[157] ^ in2[157];
    assign G[18] = in[156] & in2[156];
    assign P[18] = in[156] ^ in2[156];
    assign G[19] = in[155] & in2[155];
    assign P[19] = in[155] ^ in2[155];
    assign G[20] = in[154] & in2[154];
    assign P[20] = in[154] ^ in2[154];
    assign G[21] = in[153] & in2[153];
    assign P[21] = in[153] ^ in2[153];
    assign G[22] = in[152] & in2[152];
    assign P[22] = in[152] ^ in2[152];
    assign G[23] = in[151] & in2[151];
    assign P[23] = in[151] ^ in2[151];
    assign G[24] = in[150] & in2[150];
    assign P[24] = in[150] ^ in2[150];
    assign G[25] = in[149] & in2[149];
    assign P[25] = in[149] ^ in2[149];
    assign G[26] = in[148] & in2[148];
    assign P[26] = in[148] ^ in2[148];
    assign G[27] = in[147] & in2[147];
    assign P[27] = in[147] ^ in2[147];
    assign G[28] = in[146] & in2[146];
    assign P[28] = in[146] ^ in2[146];
    assign G[29] = in[145] & in2[145];
    assign P[29] = in[145] ^ in2[145];
    assign G[30] = in[144] & in2[144];
    assign P[30] = in[144] ^ in2[144];
    assign G[31] = in[143] & in2[143];
    assign P[31] = in[143] ^ in2[143];
    assign G[32] = in[142] & in2[142];
    assign P[32] = in[142] ^ in2[142];
    assign G[33] = in[141] & in2[141];
    assign P[33] = in[141] ^ in2[141];
    assign G[34] = in[140] & in2[140];
    assign P[34] = in[140] ^ in2[140];
    assign G[35] = in[139] & in2[139];
    assign P[35] = in[139] ^ in2[139];
    assign G[36] = in[138] & in2[138];
    assign P[36] = in[138] ^ in2[138];
    assign G[37] = in[137] & in2[137];
    assign P[37] = in[137] ^ in2[137];
    assign G[38] = in[136] & in2[136];
    assign P[38] = in[136] ^ in2[136];
    assign G[39] = in[135] & in2[135];
    assign P[39] = in[135] ^ in2[135];
    assign G[40] = in[134] & in2[134];
    assign P[40] = in[134] ^ in2[134];
    assign G[41] = in[133] & in2[133];
    assign P[41] = in[133] ^ in2[133];
    assign G[42] = in[132] & in2[132];
    assign P[42] = in[132] ^ in2[132];
    assign G[43] = in[131] & in2[131];
    assign P[43] = in[131] ^ in2[131];
    assign G[44] = in[130] & in2[130];
    assign P[44] = in[130] ^ in2[130];
    assign G[45] = in[129] & in2[129];
    assign P[45] = in[129] ^ in2[129];
    assign G[46] = in[128] & in2[128];
    assign P[46] = in[128] ^ in2[128];
    assign G[47] = in[127] & in2[127];
    assign P[47] = in[127] ^ in2[127];
    assign G[48] = in[126] & in2[126];
    assign P[48] = in[126] ^ in2[126];
    assign G[49] = in[125] & in2[125];
    assign P[49] = in[125] ^ in2[125];
    assign G[50] = in[124] & in2[124];
    assign P[50] = in[124] ^ in2[124];
    assign G[51] = in[123] & in2[123];
    assign P[51] = in[123] ^ in2[123];
    assign G[52] = in[122] & in2[122];
    assign P[52] = in[122] ^ in2[122];
    assign G[53] = in[121] & in2[121];
    assign P[53] = in[121] ^ in2[121];
    assign G[54] = in[120] & in2[120];
    assign P[54] = in[120] ^ in2[120];
    assign G[55] = in[119] & in2[119];
    assign P[55] = in[119] ^ in2[119];
    assign G[56] = in[118] & in2[118];
    assign P[56] = in[118] ^ in2[118];
    assign G[57] = in[117] & in2[117];
    assign P[57] = in[117] ^ in2[117];
    assign G[58] = in[116] & in2[116];
    assign P[58] = in[116] ^ in2[116];
    assign G[59] = in[115] & in2[115];
    assign P[59] = in[115] ^ in2[115];
    assign G[60] = in[114] & in2[114];
    assign P[60] = in[114] ^ in2[114];
    assign G[61] = in[113] & in2[113];
    assign P[61] = in[113] ^ in2[113];
    assign G[62] = in[112] & in2[112];
    assign P[62] = in[112] ^ in2[112];
    assign G[63] = in[111] & in2[111];
    assign P[63] = in[111] ^ in2[111];
    assign G[64] = in[110] & in2[110];
    assign P[64] = in[110] ^ in2[110];
    assign G[65] = in[109] & in2[109];
    assign P[65] = in[109] ^ in2[109];
    assign G[66] = in[108] & in2[108];
    assign P[66] = in[108] ^ in2[108];
    assign G[67] = in[107] & in2[107];
    assign P[67] = in[107] ^ in2[107];
    assign G[68] = in[106] & in2[106];
    assign P[68] = in[106] ^ in2[106];
    assign G[69] = in[105] & in2[105];
    assign P[69] = in[105] ^ in2[105];
    assign G[70] = in[104] & in2[104];
    assign P[70] = in[104] ^ in2[104];
    assign G[71] = in[103] & in2[103];
    assign P[71] = in[103] ^ in2[103];
    assign G[72] = in[102] & in2[102];
    assign P[72] = in[102] ^ in2[102];
    assign G[73] = in[101] & in2[101];
    assign P[73] = in[101] ^ in2[101];
    assign G[74] = in[100] & in2[100];
    assign P[74] = in[100] ^ in2[100];
    assign G[75] = in[99] & in2[99];
    assign P[75] = in[99] ^ in2[99];
    assign G[76] = in[98] & in2[98];
    assign P[76] = in[98] ^ in2[98];
    assign G[77] = in[97] & in2[97];
    assign P[77] = in[97] ^ in2[97];
    assign G[78] = in[96] & in2[96];
    assign P[78] = in[96] ^ in2[96];
    assign G[79] = in[95] & in2[95];
    assign P[79] = in[95] ^ in2[95];
    assign G[80] = in[94] & in2[94];
    assign P[80] = in[94] ^ in2[94];
    assign G[81] = in[93] & in2[93];
    assign P[81] = in[93] ^ in2[93];
    assign G[82] = in[92] & in2[92];
    assign P[82] = in[92] ^ in2[92];
    assign G[83] = in[91] & in2[91];
    assign P[83] = in[91] ^ in2[91];
    assign G[84] = in[90] & in2[90];
    assign P[84] = in[90] ^ in2[90];
    assign G[85] = in[89] & in2[89];
    assign P[85] = in[89] ^ in2[89];
    assign G[86] = in[88] & in2[88];
    assign P[86] = in[88] ^ in2[88];
    assign G[87] = in[87] & in2[87];
    assign P[87] = in[87] ^ in2[87];
    assign G[88] = in[86] & in2[86];
    assign P[88] = in[86] ^ in2[86];
    assign G[89] = in[85] & in2[85];
    assign P[89] = in[85] ^ in2[85];
    assign G[90] = in[84] & in2[84];
    assign P[90] = in[84] ^ in2[84];
    assign G[91] = in[83] & in2[83];
    assign P[91] = in[83] ^ in2[83];
    assign G[92] = in[82] & in2[82];
    assign P[92] = in[82] ^ in2[82];
    assign G[93] = in[81] & in2[81];
    assign P[93] = in[81] ^ in2[81];
    assign G[94] = in[80] & in2[80];
    assign P[94] = in[80] ^ in2[80];
    assign G[95] = in[79] & in2[79];
    assign P[95] = in[79] ^ in2[79];
    assign G[96] = in[78] & in2[78];
    assign P[96] = in[78] ^ in2[78];
    assign G[97] = in[77] & in2[77];
    assign P[97] = in[77] ^ in2[77];
    assign G[98] = in[76] & in2[76];
    assign P[98] = in[76] ^ in2[76];
    assign G[99] = in[75] & in2[75];
    assign P[99] = in[75] ^ in2[75];
    assign G[100] = in[74] & in2[74];
    assign P[100] = in[74] ^ in2[74];
    assign G[101] = in[73] & in2[73];
    assign P[101] = in[73] ^ in2[73];
    assign G[102] = in[72] & in2[72];
    assign P[102] = in[72] ^ in2[72];
    assign G[103] = in[71] & in2[71];
    assign P[103] = in[71] ^ in2[71];
    assign G[104] = in[70] & in2[70];
    assign P[104] = in[70] ^ in2[70];
    assign G[105] = in[69] & in2[69];
    assign P[105] = in[69] ^ in2[69];
    assign G[106] = in[68] & in2[68];
    assign P[106] = in[68] ^ in2[68];
    assign G[107] = in[67] & in2[67];
    assign P[107] = in[67] ^ in2[67];
    assign G[108] = in[66] & in2[66];
    assign P[108] = in[66] ^ in2[66];
    assign G[109] = in[65] & in2[65];
    assign P[109] = in[65] ^ in2[65];
    assign G[110] = in[64] & in2[64];
    assign P[110] = in[64] ^ in2[64];
    assign G[111] = in[63] & in2[63];
    assign P[111] = in[63] ^ in2[63];
    assign G[112] = in[62] & in2[62];
    assign P[112] = in[62] ^ in2[62];
    assign G[113] = in[61] & in2[61];
    assign P[113] = in[61] ^ in2[61];
    assign G[114] = in[60] & in2[60];
    assign P[114] = in[60] ^ in2[60];
    assign G[115] = in[59] & in2[59];
    assign P[115] = in[59] ^ in2[59];
    assign G[116] = in[58] & in2[58];
    assign P[116] = in[58] ^ in2[58];
    assign G[117] = in[57] & in2[57];
    assign P[117] = in[57] ^ in2[57];
    assign G[118] = in[56] & in2[56];
    assign P[118] = in[56] ^ in2[56];
    assign G[119] = in[55] & in2[55];
    assign P[119] = in[55] ^ in2[55];
    assign G[120] = in[54] & in2[54];
    assign P[120] = in[54] ^ in2[54];
    assign G[121] = in[53] & in2[53];
    assign P[121] = in[53] ^ in2[53];
    assign G[122] = in[52] & in2[52];
    assign P[122] = in[52] ^ in2[52];
    assign G[123] = in[51] & in2[51];
    assign P[123] = in[51] ^ in2[51];
    assign G[124] = in[50] & in2[50];
    assign P[124] = in[50] ^ in2[50];
    assign G[125] = in[49] & in2[49];
    assign P[125] = in[49] ^ in2[49];
    assign G[126] = in[48] & in2[48];
    assign P[126] = in[48] ^ in2[48];
    assign G[127] = in[47] & in2[47];
    assign P[127] = in[47] ^ in2[47];
    assign G[128] = in[46] & in2[46];
    assign P[128] = in[46] ^ in2[46];
    assign G[129] = in[45] & in2[45];
    assign P[129] = in[45] ^ in2[45];
    assign G[130] = in[44] & in2[44];
    assign P[130] = in[44] ^ in2[44];
    assign G[131] = in[43] & in2[43];
    assign P[131] = in[43] ^ in2[43];
    assign G[132] = in[42] & in2[42];
    assign P[132] = in[42] ^ in2[42];
    assign G[133] = in[41] & in2[41];
    assign P[133] = in[41] ^ in2[41];
    assign G[134] = in[40] & in2[40];
    assign P[134] = in[40] ^ in2[40];
    assign G[135] = in[39] & in2[39];
    assign P[135] = in[39] ^ in2[39];
    assign G[136] = in[38] & in2[38];
    assign P[136] = in[38] ^ in2[38];
    assign G[137] = in[37] & in2[37];
    assign P[137] = in[37] ^ in2[37];
    assign G[138] = in[36] & in2[36];
    assign P[138] = in[36] ^ in2[36];
    assign G[139] = in[35] & in2[35];
    assign P[139] = in[35] ^ in2[35];
    assign G[140] = in[34] & in2[34];
    assign P[140] = in[34] ^ in2[34];
    assign G[141] = in[33] & in2[33];
    assign P[141] = in[33] ^ in2[33];
    assign G[142] = in[32] & in2[32];
    assign P[142] = in[32] ^ in2[32];
    assign G[143] = in[31] & in2[31];
    assign P[143] = in[31] ^ in2[31];
    assign G[144] = in[30] & in2[30];
    assign P[144] = in[30] ^ in2[30];
    assign G[145] = in[29] & in2[29];
    assign P[145] = in[29] ^ in2[29];
    assign G[146] = in[28] & in2[28];
    assign P[146] = in[28] ^ in2[28];
    assign G[147] = in[27] & in2[27];
    assign P[147] = in[27] ^ in2[27];
    assign G[148] = in[26] & in2[26];
    assign P[148] = in[26] ^ in2[26];
    assign G[149] = in[25] & in2[25];
    assign P[149] = in[25] ^ in2[25];
    assign G[150] = in[24] & in2[24];
    assign P[150] = in[24] ^ in2[24];
    assign G[151] = in[23] & in2[23];
    assign P[151] = in[23] ^ in2[23];
    assign G[152] = in[22] & in2[22];
    assign P[152] = in[22] ^ in2[22];
    assign G[153] = in[21] & in2[21];
    assign P[153] = in[21] ^ in2[21];
    assign G[154] = in[20] & in2[20];
    assign P[154] = in[20] ^ in2[20];
    assign G[155] = in[19] & in2[19];
    assign P[155] = in[19] ^ in2[19];
    assign G[156] = in[18] & in2[18];
    assign P[156] = in[18] ^ in2[18];
    assign G[157] = in[17] & in2[17];
    assign P[157] = in[17] ^ in2[17];
    assign G[158] = in[16] & in2[16];
    assign P[158] = in[16] ^ in2[16];
    assign G[159] = in[15] & in2[15];
    assign P[159] = in[15] ^ in2[15];
    assign G[160] = in[14] & in2[14];
    assign P[160] = in[14] ^ in2[14];
    assign G[161] = in[13] & in2[13];
    assign P[161] = in[13] ^ in2[13];
    assign G[162] = in[12] & in2[12];
    assign P[162] = in[12] ^ in2[12];
    assign G[163] = in[11] & in2[11];
    assign P[163] = in[11] ^ in2[11];
    assign G[164] = in[10] & in2[10];
    assign P[164] = in[10] ^ in2[10];
    assign G[165] = in[9] & in2[9];
    assign P[165] = in[9] ^ in2[9];
    assign G[166] = in[8] & in2[8];
    assign P[166] = in[8] ^ in2[8];
    assign G[167] = in[7] & in2[7];
    assign P[167] = in[7] ^ in2[7];
    assign G[168] = in[6] & in2[6];
    assign P[168] = in[6] ^ in2[6];
    assign G[169] = in[5] & in2[5];
    assign P[169] = in[5] ^ in2[5];
    assign G[170] = in[4] & in2[4];
    assign P[170] = in[4] ^ in2[4];
    assign G[171] = in[3] & in2[3];
    assign P[171] = in[3] ^ in2[3];
    assign G[172] = in[2] & in2[2];
    assign P[172] = in[2] ^ in2[2];
    assign G[173] = in[1] & in2[1];
    assign P[173] = in[1] ^ in2[1];
    assign G[174] = in[0] & in2[0];
    assign P[174] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign C[174] = G[173] | (P[173] & C[173]);
    assign cout = G[174] | (P[174] & C[174]);
    assign sum = P ^ C;
endmodule

module CLA174(output [173:0] sum, output cout, input [173:0] in1, input [173:0] in2;

    wire[173:0] G;
    wire[173:0] C;
    wire[173:0] P;

    assign G[0] = in[173] & in2[173];
    assign P[0] = in[173] ^ in2[173];
    assign G[1] = in[172] & in2[172];
    assign P[1] = in[172] ^ in2[172];
    assign G[2] = in[171] & in2[171];
    assign P[2] = in[171] ^ in2[171];
    assign G[3] = in[170] & in2[170];
    assign P[3] = in[170] ^ in2[170];
    assign G[4] = in[169] & in2[169];
    assign P[4] = in[169] ^ in2[169];
    assign G[5] = in[168] & in2[168];
    assign P[5] = in[168] ^ in2[168];
    assign G[6] = in[167] & in2[167];
    assign P[6] = in[167] ^ in2[167];
    assign G[7] = in[166] & in2[166];
    assign P[7] = in[166] ^ in2[166];
    assign G[8] = in[165] & in2[165];
    assign P[8] = in[165] ^ in2[165];
    assign G[9] = in[164] & in2[164];
    assign P[9] = in[164] ^ in2[164];
    assign G[10] = in[163] & in2[163];
    assign P[10] = in[163] ^ in2[163];
    assign G[11] = in[162] & in2[162];
    assign P[11] = in[162] ^ in2[162];
    assign G[12] = in[161] & in2[161];
    assign P[12] = in[161] ^ in2[161];
    assign G[13] = in[160] & in2[160];
    assign P[13] = in[160] ^ in2[160];
    assign G[14] = in[159] & in2[159];
    assign P[14] = in[159] ^ in2[159];
    assign G[15] = in[158] & in2[158];
    assign P[15] = in[158] ^ in2[158];
    assign G[16] = in[157] & in2[157];
    assign P[16] = in[157] ^ in2[157];
    assign G[17] = in[156] & in2[156];
    assign P[17] = in[156] ^ in2[156];
    assign G[18] = in[155] & in2[155];
    assign P[18] = in[155] ^ in2[155];
    assign G[19] = in[154] & in2[154];
    assign P[19] = in[154] ^ in2[154];
    assign G[20] = in[153] & in2[153];
    assign P[20] = in[153] ^ in2[153];
    assign G[21] = in[152] & in2[152];
    assign P[21] = in[152] ^ in2[152];
    assign G[22] = in[151] & in2[151];
    assign P[22] = in[151] ^ in2[151];
    assign G[23] = in[150] & in2[150];
    assign P[23] = in[150] ^ in2[150];
    assign G[24] = in[149] & in2[149];
    assign P[24] = in[149] ^ in2[149];
    assign G[25] = in[148] & in2[148];
    assign P[25] = in[148] ^ in2[148];
    assign G[26] = in[147] & in2[147];
    assign P[26] = in[147] ^ in2[147];
    assign G[27] = in[146] & in2[146];
    assign P[27] = in[146] ^ in2[146];
    assign G[28] = in[145] & in2[145];
    assign P[28] = in[145] ^ in2[145];
    assign G[29] = in[144] & in2[144];
    assign P[29] = in[144] ^ in2[144];
    assign G[30] = in[143] & in2[143];
    assign P[30] = in[143] ^ in2[143];
    assign G[31] = in[142] & in2[142];
    assign P[31] = in[142] ^ in2[142];
    assign G[32] = in[141] & in2[141];
    assign P[32] = in[141] ^ in2[141];
    assign G[33] = in[140] & in2[140];
    assign P[33] = in[140] ^ in2[140];
    assign G[34] = in[139] & in2[139];
    assign P[34] = in[139] ^ in2[139];
    assign G[35] = in[138] & in2[138];
    assign P[35] = in[138] ^ in2[138];
    assign G[36] = in[137] & in2[137];
    assign P[36] = in[137] ^ in2[137];
    assign G[37] = in[136] & in2[136];
    assign P[37] = in[136] ^ in2[136];
    assign G[38] = in[135] & in2[135];
    assign P[38] = in[135] ^ in2[135];
    assign G[39] = in[134] & in2[134];
    assign P[39] = in[134] ^ in2[134];
    assign G[40] = in[133] & in2[133];
    assign P[40] = in[133] ^ in2[133];
    assign G[41] = in[132] & in2[132];
    assign P[41] = in[132] ^ in2[132];
    assign G[42] = in[131] & in2[131];
    assign P[42] = in[131] ^ in2[131];
    assign G[43] = in[130] & in2[130];
    assign P[43] = in[130] ^ in2[130];
    assign G[44] = in[129] & in2[129];
    assign P[44] = in[129] ^ in2[129];
    assign G[45] = in[128] & in2[128];
    assign P[45] = in[128] ^ in2[128];
    assign G[46] = in[127] & in2[127];
    assign P[46] = in[127] ^ in2[127];
    assign G[47] = in[126] & in2[126];
    assign P[47] = in[126] ^ in2[126];
    assign G[48] = in[125] & in2[125];
    assign P[48] = in[125] ^ in2[125];
    assign G[49] = in[124] & in2[124];
    assign P[49] = in[124] ^ in2[124];
    assign G[50] = in[123] & in2[123];
    assign P[50] = in[123] ^ in2[123];
    assign G[51] = in[122] & in2[122];
    assign P[51] = in[122] ^ in2[122];
    assign G[52] = in[121] & in2[121];
    assign P[52] = in[121] ^ in2[121];
    assign G[53] = in[120] & in2[120];
    assign P[53] = in[120] ^ in2[120];
    assign G[54] = in[119] & in2[119];
    assign P[54] = in[119] ^ in2[119];
    assign G[55] = in[118] & in2[118];
    assign P[55] = in[118] ^ in2[118];
    assign G[56] = in[117] & in2[117];
    assign P[56] = in[117] ^ in2[117];
    assign G[57] = in[116] & in2[116];
    assign P[57] = in[116] ^ in2[116];
    assign G[58] = in[115] & in2[115];
    assign P[58] = in[115] ^ in2[115];
    assign G[59] = in[114] & in2[114];
    assign P[59] = in[114] ^ in2[114];
    assign G[60] = in[113] & in2[113];
    assign P[60] = in[113] ^ in2[113];
    assign G[61] = in[112] & in2[112];
    assign P[61] = in[112] ^ in2[112];
    assign G[62] = in[111] & in2[111];
    assign P[62] = in[111] ^ in2[111];
    assign G[63] = in[110] & in2[110];
    assign P[63] = in[110] ^ in2[110];
    assign G[64] = in[109] & in2[109];
    assign P[64] = in[109] ^ in2[109];
    assign G[65] = in[108] & in2[108];
    assign P[65] = in[108] ^ in2[108];
    assign G[66] = in[107] & in2[107];
    assign P[66] = in[107] ^ in2[107];
    assign G[67] = in[106] & in2[106];
    assign P[67] = in[106] ^ in2[106];
    assign G[68] = in[105] & in2[105];
    assign P[68] = in[105] ^ in2[105];
    assign G[69] = in[104] & in2[104];
    assign P[69] = in[104] ^ in2[104];
    assign G[70] = in[103] & in2[103];
    assign P[70] = in[103] ^ in2[103];
    assign G[71] = in[102] & in2[102];
    assign P[71] = in[102] ^ in2[102];
    assign G[72] = in[101] & in2[101];
    assign P[72] = in[101] ^ in2[101];
    assign G[73] = in[100] & in2[100];
    assign P[73] = in[100] ^ in2[100];
    assign G[74] = in[99] & in2[99];
    assign P[74] = in[99] ^ in2[99];
    assign G[75] = in[98] & in2[98];
    assign P[75] = in[98] ^ in2[98];
    assign G[76] = in[97] & in2[97];
    assign P[76] = in[97] ^ in2[97];
    assign G[77] = in[96] & in2[96];
    assign P[77] = in[96] ^ in2[96];
    assign G[78] = in[95] & in2[95];
    assign P[78] = in[95] ^ in2[95];
    assign G[79] = in[94] & in2[94];
    assign P[79] = in[94] ^ in2[94];
    assign G[80] = in[93] & in2[93];
    assign P[80] = in[93] ^ in2[93];
    assign G[81] = in[92] & in2[92];
    assign P[81] = in[92] ^ in2[92];
    assign G[82] = in[91] & in2[91];
    assign P[82] = in[91] ^ in2[91];
    assign G[83] = in[90] & in2[90];
    assign P[83] = in[90] ^ in2[90];
    assign G[84] = in[89] & in2[89];
    assign P[84] = in[89] ^ in2[89];
    assign G[85] = in[88] & in2[88];
    assign P[85] = in[88] ^ in2[88];
    assign G[86] = in[87] & in2[87];
    assign P[86] = in[87] ^ in2[87];
    assign G[87] = in[86] & in2[86];
    assign P[87] = in[86] ^ in2[86];
    assign G[88] = in[85] & in2[85];
    assign P[88] = in[85] ^ in2[85];
    assign G[89] = in[84] & in2[84];
    assign P[89] = in[84] ^ in2[84];
    assign G[90] = in[83] & in2[83];
    assign P[90] = in[83] ^ in2[83];
    assign G[91] = in[82] & in2[82];
    assign P[91] = in[82] ^ in2[82];
    assign G[92] = in[81] & in2[81];
    assign P[92] = in[81] ^ in2[81];
    assign G[93] = in[80] & in2[80];
    assign P[93] = in[80] ^ in2[80];
    assign G[94] = in[79] & in2[79];
    assign P[94] = in[79] ^ in2[79];
    assign G[95] = in[78] & in2[78];
    assign P[95] = in[78] ^ in2[78];
    assign G[96] = in[77] & in2[77];
    assign P[96] = in[77] ^ in2[77];
    assign G[97] = in[76] & in2[76];
    assign P[97] = in[76] ^ in2[76];
    assign G[98] = in[75] & in2[75];
    assign P[98] = in[75] ^ in2[75];
    assign G[99] = in[74] & in2[74];
    assign P[99] = in[74] ^ in2[74];
    assign G[100] = in[73] & in2[73];
    assign P[100] = in[73] ^ in2[73];
    assign G[101] = in[72] & in2[72];
    assign P[101] = in[72] ^ in2[72];
    assign G[102] = in[71] & in2[71];
    assign P[102] = in[71] ^ in2[71];
    assign G[103] = in[70] & in2[70];
    assign P[103] = in[70] ^ in2[70];
    assign G[104] = in[69] & in2[69];
    assign P[104] = in[69] ^ in2[69];
    assign G[105] = in[68] & in2[68];
    assign P[105] = in[68] ^ in2[68];
    assign G[106] = in[67] & in2[67];
    assign P[106] = in[67] ^ in2[67];
    assign G[107] = in[66] & in2[66];
    assign P[107] = in[66] ^ in2[66];
    assign G[108] = in[65] & in2[65];
    assign P[108] = in[65] ^ in2[65];
    assign G[109] = in[64] & in2[64];
    assign P[109] = in[64] ^ in2[64];
    assign G[110] = in[63] & in2[63];
    assign P[110] = in[63] ^ in2[63];
    assign G[111] = in[62] & in2[62];
    assign P[111] = in[62] ^ in2[62];
    assign G[112] = in[61] & in2[61];
    assign P[112] = in[61] ^ in2[61];
    assign G[113] = in[60] & in2[60];
    assign P[113] = in[60] ^ in2[60];
    assign G[114] = in[59] & in2[59];
    assign P[114] = in[59] ^ in2[59];
    assign G[115] = in[58] & in2[58];
    assign P[115] = in[58] ^ in2[58];
    assign G[116] = in[57] & in2[57];
    assign P[116] = in[57] ^ in2[57];
    assign G[117] = in[56] & in2[56];
    assign P[117] = in[56] ^ in2[56];
    assign G[118] = in[55] & in2[55];
    assign P[118] = in[55] ^ in2[55];
    assign G[119] = in[54] & in2[54];
    assign P[119] = in[54] ^ in2[54];
    assign G[120] = in[53] & in2[53];
    assign P[120] = in[53] ^ in2[53];
    assign G[121] = in[52] & in2[52];
    assign P[121] = in[52] ^ in2[52];
    assign G[122] = in[51] & in2[51];
    assign P[122] = in[51] ^ in2[51];
    assign G[123] = in[50] & in2[50];
    assign P[123] = in[50] ^ in2[50];
    assign G[124] = in[49] & in2[49];
    assign P[124] = in[49] ^ in2[49];
    assign G[125] = in[48] & in2[48];
    assign P[125] = in[48] ^ in2[48];
    assign G[126] = in[47] & in2[47];
    assign P[126] = in[47] ^ in2[47];
    assign G[127] = in[46] & in2[46];
    assign P[127] = in[46] ^ in2[46];
    assign G[128] = in[45] & in2[45];
    assign P[128] = in[45] ^ in2[45];
    assign G[129] = in[44] & in2[44];
    assign P[129] = in[44] ^ in2[44];
    assign G[130] = in[43] & in2[43];
    assign P[130] = in[43] ^ in2[43];
    assign G[131] = in[42] & in2[42];
    assign P[131] = in[42] ^ in2[42];
    assign G[132] = in[41] & in2[41];
    assign P[132] = in[41] ^ in2[41];
    assign G[133] = in[40] & in2[40];
    assign P[133] = in[40] ^ in2[40];
    assign G[134] = in[39] & in2[39];
    assign P[134] = in[39] ^ in2[39];
    assign G[135] = in[38] & in2[38];
    assign P[135] = in[38] ^ in2[38];
    assign G[136] = in[37] & in2[37];
    assign P[136] = in[37] ^ in2[37];
    assign G[137] = in[36] & in2[36];
    assign P[137] = in[36] ^ in2[36];
    assign G[138] = in[35] & in2[35];
    assign P[138] = in[35] ^ in2[35];
    assign G[139] = in[34] & in2[34];
    assign P[139] = in[34] ^ in2[34];
    assign G[140] = in[33] & in2[33];
    assign P[140] = in[33] ^ in2[33];
    assign G[141] = in[32] & in2[32];
    assign P[141] = in[32] ^ in2[32];
    assign G[142] = in[31] & in2[31];
    assign P[142] = in[31] ^ in2[31];
    assign G[143] = in[30] & in2[30];
    assign P[143] = in[30] ^ in2[30];
    assign G[144] = in[29] & in2[29];
    assign P[144] = in[29] ^ in2[29];
    assign G[145] = in[28] & in2[28];
    assign P[145] = in[28] ^ in2[28];
    assign G[146] = in[27] & in2[27];
    assign P[146] = in[27] ^ in2[27];
    assign G[147] = in[26] & in2[26];
    assign P[147] = in[26] ^ in2[26];
    assign G[148] = in[25] & in2[25];
    assign P[148] = in[25] ^ in2[25];
    assign G[149] = in[24] & in2[24];
    assign P[149] = in[24] ^ in2[24];
    assign G[150] = in[23] & in2[23];
    assign P[150] = in[23] ^ in2[23];
    assign G[151] = in[22] & in2[22];
    assign P[151] = in[22] ^ in2[22];
    assign G[152] = in[21] & in2[21];
    assign P[152] = in[21] ^ in2[21];
    assign G[153] = in[20] & in2[20];
    assign P[153] = in[20] ^ in2[20];
    assign G[154] = in[19] & in2[19];
    assign P[154] = in[19] ^ in2[19];
    assign G[155] = in[18] & in2[18];
    assign P[155] = in[18] ^ in2[18];
    assign G[156] = in[17] & in2[17];
    assign P[156] = in[17] ^ in2[17];
    assign G[157] = in[16] & in2[16];
    assign P[157] = in[16] ^ in2[16];
    assign G[158] = in[15] & in2[15];
    assign P[158] = in[15] ^ in2[15];
    assign G[159] = in[14] & in2[14];
    assign P[159] = in[14] ^ in2[14];
    assign G[160] = in[13] & in2[13];
    assign P[160] = in[13] ^ in2[13];
    assign G[161] = in[12] & in2[12];
    assign P[161] = in[12] ^ in2[12];
    assign G[162] = in[11] & in2[11];
    assign P[162] = in[11] ^ in2[11];
    assign G[163] = in[10] & in2[10];
    assign P[163] = in[10] ^ in2[10];
    assign G[164] = in[9] & in2[9];
    assign P[164] = in[9] ^ in2[9];
    assign G[165] = in[8] & in2[8];
    assign P[165] = in[8] ^ in2[8];
    assign G[166] = in[7] & in2[7];
    assign P[166] = in[7] ^ in2[7];
    assign G[167] = in[6] & in2[6];
    assign P[167] = in[6] ^ in2[6];
    assign G[168] = in[5] & in2[5];
    assign P[168] = in[5] ^ in2[5];
    assign G[169] = in[4] & in2[4];
    assign P[169] = in[4] ^ in2[4];
    assign G[170] = in[3] & in2[3];
    assign P[170] = in[3] ^ in2[3];
    assign G[171] = in[2] & in2[2];
    assign P[171] = in[2] ^ in2[2];
    assign G[172] = in[1] & in2[1];
    assign P[172] = in[1] ^ in2[1];
    assign G[173] = in[0] & in2[0];
    assign P[173] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign C[173] = G[172] | (P[172] & C[172]);
    assign cout = G[173] | (P[173] & C[173]);
    assign sum = P ^ C;
endmodule

module CLA173(output [172:0] sum, output cout, input [172:0] in1, input [172:0] in2;

    wire[172:0] G;
    wire[172:0] C;
    wire[172:0] P;

    assign G[0] = in[172] & in2[172];
    assign P[0] = in[172] ^ in2[172];
    assign G[1] = in[171] & in2[171];
    assign P[1] = in[171] ^ in2[171];
    assign G[2] = in[170] & in2[170];
    assign P[2] = in[170] ^ in2[170];
    assign G[3] = in[169] & in2[169];
    assign P[3] = in[169] ^ in2[169];
    assign G[4] = in[168] & in2[168];
    assign P[4] = in[168] ^ in2[168];
    assign G[5] = in[167] & in2[167];
    assign P[5] = in[167] ^ in2[167];
    assign G[6] = in[166] & in2[166];
    assign P[6] = in[166] ^ in2[166];
    assign G[7] = in[165] & in2[165];
    assign P[7] = in[165] ^ in2[165];
    assign G[8] = in[164] & in2[164];
    assign P[8] = in[164] ^ in2[164];
    assign G[9] = in[163] & in2[163];
    assign P[9] = in[163] ^ in2[163];
    assign G[10] = in[162] & in2[162];
    assign P[10] = in[162] ^ in2[162];
    assign G[11] = in[161] & in2[161];
    assign P[11] = in[161] ^ in2[161];
    assign G[12] = in[160] & in2[160];
    assign P[12] = in[160] ^ in2[160];
    assign G[13] = in[159] & in2[159];
    assign P[13] = in[159] ^ in2[159];
    assign G[14] = in[158] & in2[158];
    assign P[14] = in[158] ^ in2[158];
    assign G[15] = in[157] & in2[157];
    assign P[15] = in[157] ^ in2[157];
    assign G[16] = in[156] & in2[156];
    assign P[16] = in[156] ^ in2[156];
    assign G[17] = in[155] & in2[155];
    assign P[17] = in[155] ^ in2[155];
    assign G[18] = in[154] & in2[154];
    assign P[18] = in[154] ^ in2[154];
    assign G[19] = in[153] & in2[153];
    assign P[19] = in[153] ^ in2[153];
    assign G[20] = in[152] & in2[152];
    assign P[20] = in[152] ^ in2[152];
    assign G[21] = in[151] & in2[151];
    assign P[21] = in[151] ^ in2[151];
    assign G[22] = in[150] & in2[150];
    assign P[22] = in[150] ^ in2[150];
    assign G[23] = in[149] & in2[149];
    assign P[23] = in[149] ^ in2[149];
    assign G[24] = in[148] & in2[148];
    assign P[24] = in[148] ^ in2[148];
    assign G[25] = in[147] & in2[147];
    assign P[25] = in[147] ^ in2[147];
    assign G[26] = in[146] & in2[146];
    assign P[26] = in[146] ^ in2[146];
    assign G[27] = in[145] & in2[145];
    assign P[27] = in[145] ^ in2[145];
    assign G[28] = in[144] & in2[144];
    assign P[28] = in[144] ^ in2[144];
    assign G[29] = in[143] & in2[143];
    assign P[29] = in[143] ^ in2[143];
    assign G[30] = in[142] & in2[142];
    assign P[30] = in[142] ^ in2[142];
    assign G[31] = in[141] & in2[141];
    assign P[31] = in[141] ^ in2[141];
    assign G[32] = in[140] & in2[140];
    assign P[32] = in[140] ^ in2[140];
    assign G[33] = in[139] & in2[139];
    assign P[33] = in[139] ^ in2[139];
    assign G[34] = in[138] & in2[138];
    assign P[34] = in[138] ^ in2[138];
    assign G[35] = in[137] & in2[137];
    assign P[35] = in[137] ^ in2[137];
    assign G[36] = in[136] & in2[136];
    assign P[36] = in[136] ^ in2[136];
    assign G[37] = in[135] & in2[135];
    assign P[37] = in[135] ^ in2[135];
    assign G[38] = in[134] & in2[134];
    assign P[38] = in[134] ^ in2[134];
    assign G[39] = in[133] & in2[133];
    assign P[39] = in[133] ^ in2[133];
    assign G[40] = in[132] & in2[132];
    assign P[40] = in[132] ^ in2[132];
    assign G[41] = in[131] & in2[131];
    assign P[41] = in[131] ^ in2[131];
    assign G[42] = in[130] & in2[130];
    assign P[42] = in[130] ^ in2[130];
    assign G[43] = in[129] & in2[129];
    assign P[43] = in[129] ^ in2[129];
    assign G[44] = in[128] & in2[128];
    assign P[44] = in[128] ^ in2[128];
    assign G[45] = in[127] & in2[127];
    assign P[45] = in[127] ^ in2[127];
    assign G[46] = in[126] & in2[126];
    assign P[46] = in[126] ^ in2[126];
    assign G[47] = in[125] & in2[125];
    assign P[47] = in[125] ^ in2[125];
    assign G[48] = in[124] & in2[124];
    assign P[48] = in[124] ^ in2[124];
    assign G[49] = in[123] & in2[123];
    assign P[49] = in[123] ^ in2[123];
    assign G[50] = in[122] & in2[122];
    assign P[50] = in[122] ^ in2[122];
    assign G[51] = in[121] & in2[121];
    assign P[51] = in[121] ^ in2[121];
    assign G[52] = in[120] & in2[120];
    assign P[52] = in[120] ^ in2[120];
    assign G[53] = in[119] & in2[119];
    assign P[53] = in[119] ^ in2[119];
    assign G[54] = in[118] & in2[118];
    assign P[54] = in[118] ^ in2[118];
    assign G[55] = in[117] & in2[117];
    assign P[55] = in[117] ^ in2[117];
    assign G[56] = in[116] & in2[116];
    assign P[56] = in[116] ^ in2[116];
    assign G[57] = in[115] & in2[115];
    assign P[57] = in[115] ^ in2[115];
    assign G[58] = in[114] & in2[114];
    assign P[58] = in[114] ^ in2[114];
    assign G[59] = in[113] & in2[113];
    assign P[59] = in[113] ^ in2[113];
    assign G[60] = in[112] & in2[112];
    assign P[60] = in[112] ^ in2[112];
    assign G[61] = in[111] & in2[111];
    assign P[61] = in[111] ^ in2[111];
    assign G[62] = in[110] & in2[110];
    assign P[62] = in[110] ^ in2[110];
    assign G[63] = in[109] & in2[109];
    assign P[63] = in[109] ^ in2[109];
    assign G[64] = in[108] & in2[108];
    assign P[64] = in[108] ^ in2[108];
    assign G[65] = in[107] & in2[107];
    assign P[65] = in[107] ^ in2[107];
    assign G[66] = in[106] & in2[106];
    assign P[66] = in[106] ^ in2[106];
    assign G[67] = in[105] & in2[105];
    assign P[67] = in[105] ^ in2[105];
    assign G[68] = in[104] & in2[104];
    assign P[68] = in[104] ^ in2[104];
    assign G[69] = in[103] & in2[103];
    assign P[69] = in[103] ^ in2[103];
    assign G[70] = in[102] & in2[102];
    assign P[70] = in[102] ^ in2[102];
    assign G[71] = in[101] & in2[101];
    assign P[71] = in[101] ^ in2[101];
    assign G[72] = in[100] & in2[100];
    assign P[72] = in[100] ^ in2[100];
    assign G[73] = in[99] & in2[99];
    assign P[73] = in[99] ^ in2[99];
    assign G[74] = in[98] & in2[98];
    assign P[74] = in[98] ^ in2[98];
    assign G[75] = in[97] & in2[97];
    assign P[75] = in[97] ^ in2[97];
    assign G[76] = in[96] & in2[96];
    assign P[76] = in[96] ^ in2[96];
    assign G[77] = in[95] & in2[95];
    assign P[77] = in[95] ^ in2[95];
    assign G[78] = in[94] & in2[94];
    assign P[78] = in[94] ^ in2[94];
    assign G[79] = in[93] & in2[93];
    assign P[79] = in[93] ^ in2[93];
    assign G[80] = in[92] & in2[92];
    assign P[80] = in[92] ^ in2[92];
    assign G[81] = in[91] & in2[91];
    assign P[81] = in[91] ^ in2[91];
    assign G[82] = in[90] & in2[90];
    assign P[82] = in[90] ^ in2[90];
    assign G[83] = in[89] & in2[89];
    assign P[83] = in[89] ^ in2[89];
    assign G[84] = in[88] & in2[88];
    assign P[84] = in[88] ^ in2[88];
    assign G[85] = in[87] & in2[87];
    assign P[85] = in[87] ^ in2[87];
    assign G[86] = in[86] & in2[86];
    assign P[86] = in[86] ^ in2[86];
    assign G[87] = in[85] & in2[85];
    assign P[87] = in[85] ^ in2[85];
    assign G[88] = in[84] & in2[84];
    assign P[88] = in[84] ^ in2[84];
    assign G[89] = in[83] & in2[83];
    assign P[89] = in[83] ^ in2[83];
    assign G[90] = in[82] & in2[82];
    assign P[90] = in[82] ^ in2[82];
    assign G[91] = in[81] & in2[81];
    assign P[91] = in[81] ^ in2[81];
    assign G[92] = in[80] & in2[80];
    assign P[92] = in[80] ^ in2[80];
    assign G[93] = in[79] & in2[79];
    assign P[93] = in[79] ^ in2[79];
    assign G[94] = in[78] & in2[78];
    assign P[94] = in[78] ^ in2[78];
    assign G[95] = in[77] & in2[77];
    assign P[95] = in[77] ^ in2[77];
    assign G[96] = in[76] & in2[76];
    assign P[96] = in[76] ^ in2[76];
    assign G[97] = in[75] & in2[75];
    assign P[97] = in[75] ^ in2[75];
    assign G[98] = in[74] & in2[74];
    assign P[98] = in[74] ^ in2[74];
    assign G[99] = in[73] & in2[73];
    assign P[99] = in[73] ^ in2[73];
    assign G[100] = in[72] & in2[72];
    assign P[100] = in[72] ^ in2[72];
    assign G[101] = in[71] & in2[71];
    assign P[101] = in[71] ^ in2[71];
    assign G[102] = in[70] & in2[70];
    assign P[102] = in[70] ^ in2[70];
    assign G[103] = in[69] & in2[69];
    assign P[103] = in[69] ^ in2[69];
    assign G[104] = in[68] & in2[68];
    assign P[104] = in[68] ^ in2[68];
    assign G[105] = in[67] & in2[67];
    assign P[105] = in[67] ^ in2[67];
    assign G[106] = in[66] & in2[66];
    assign P[106] = in[66] ^ in2[66];
    assign G[107] = in[65] & in2[65];
    assign P[107] = in[65] ^ in2[65];
    assign G[108] = in[64] & in2[64];
    assign P[108] = in[64] ^ in2[64];
    assign G[109] = in[63] & in2[63];
    assign P[109] = in[63] ^ in2[63];
    assign G[110] = in[62] & in2[62];
    assign P[110] = in[62] ^ in2[62];
    assign G[111] = in[61] & in2[61];
    assign P[111] = in[61] ^ in2[61];
    assign G[112] = in[60] & in2[60];
    assign P[112] = in[60] ^ in2[60];
    assign G[113] = in[59] & in2[59];
    assign P[113] = in[59] ^ in2[59];
    assign G[114] = in[58] & in2[58];
    assign P[114] = in[58] ^ in2[58];
    assign G[115] = in[57] & in2[57];
    assign P[115] = in[57] ^ in2[57];
    assign G[116] = in[56] & in2[56];
    assign P[116] = in[56] ^ in2[56];
    assign G[117] = in[55] & in2[55];
    assign P[117] = in[55] ^ in2[55];
    assign G[118] = in[54] & in2[54];
    assign P[118] = in[54] ^ in2[54];
    assign G[119] = in[53] & in2[53];
    assign P[119] = in[53] ^ in2[53];
    assign G[120] = in[52] & in2[52];
    assign P[120] = in[52] ^ in2[52];
    assign G[121] = in[51] & in2[51];
    assign P[121] = in[51] ^ in2[51];
    assign G[122] = in[50] & in2[50];
    assign P[122] = in[50] ^ in2[50];
    assign G[123] = in[49] & in2[49];
    assign P[123] = in[49] ^ in2[49];
    assign G[124] = in[48] & in2[48];
    assign P[124] = in[48] ^ in2[48];
    assign G[125] = in[47] & in2[47];
    assign P[125] = in[47] ^ in2[47];
    assign G[126] = in[46] & in2[46];
    assign P[126] = in[46] ^ in2[46];
    assign G[127] = in[45] & in2[45];
    assign P[127] = in[45] ^ in2[45];
    assign G[128] = in[44] & in2[44];
    assign P[128] = in[44] ^ in2[44];
    assign G[129] = in[43] & in2[43];
    assign P[129] = in[43] ^ in2[43];
    assign G[130] = in[42] & in2[42];
    assign P[130] = in[42] ^ in2[42];
    assign G[131] = in[41] & in2[41];
    assign P[131] = in[41] ^ in2[41];
    assign G[132] = in[40] & in2[40];
    assign P[132] = in[40] ^ in2[40];
    assign G[133] = in[39] & in2[39];
    assign P[133] = in[39] ^ in2[39];
    assign G[134] = in[38] & in2[38];
    assign P[134] = in[38] ^ in2[38];
    assign G[135] = in[37] & in2[37];
    assign P[135] = in[37] ^ in2[37];
    assign G[136] = in[36] & in2[36];
    assign P[136] = in[36] ^ in2[36];
    assign G[137] = in[35] & in2[35];
    assign P[137] = in[35] ^ in2[35];
    assign G[138] = in[34] & in2[34];
    assign P[138] = in[34] ^ in2[34];
    assign G[139] = in[33] & in2[33];
    assign P[139] = in[33] ^ in2[33];
    assign G[140] = in[32] & in2[32];
    assign P[140] = in[32] ^ in2[32];
    assign G[141] = in[31] & in2[31];
    assign P[141] = in[31] ^ in2[31];
    assign G[142] = in[30] & in2[30];
    assign P[142] = in[30] ^ in2[30];
    assign G[143] = in[29] & in2[29];
    assign P[143] = in[29] ^ in2[29];
    assign G[144] = in[28] & in2[28];
    assign P[144] = in[28] ^ in2[28];
    assign G[145] = in[27] & in2[27];
    assign P[145] = in[27] ^ in2[27];
    assign G[146] = in[26] & in2[26];
    assign P[146] = in[26] ^ in2[26];
    assign G[147] = in[25] & in2[25];
    assign P[147] = in[25] ^ in2[25];
    assign G[148] = in[24] & in2[24];
    assign P[148] = in[24] ^ in2[24];
    assign G[149] = in[23] & in2[23];
    assign P[149] = in[23] ^ in2[23];
    assign G[150] = in[22] & in2[22];
    assign P[150] = in[22] ^ in2[22];
    assign G[151] = in[21] & in2[21];
    assign P[151] = in[21] ^ in2[21];
    assign G[152] = in[20] & in2[20];
    assign P[152] = in[20] ^ in2[20];
    assign G[153] = in[19] & in2[19];
    assign P[153] = in[19] ^ in2[19];
    assign G[154] = in[18] & in2[18];
    assign P[154] = in[18] ^ in2[18];
    assign G[155] = in[17] & in2[17];
    assign P[155] = in[17] ^ in2[17];
    assign G[156] = in[16] & in2[16];
    assign P[156] = in[16] ^ in2[16];
    assign G[157] = in[15] & in2[15];
    assign P[157] = in[15] ^ in2[15];
    assign G[158] = in[14] & in2[14];
    assign P[158] = in[14] ^ in2[14];
    assign G[159] = in[13] & in2[13];
    assign P[159] = in[13] ^ in2[13];
    assign G[160] = in[12] & in2[12];
    assign P[160] = in[12] ^ in2[12];
    assign G[161] = in[11] & in2[11];
    assign P[161] = in[11] ^ in2[11];
    assign G[162] = in[10] & in2[10];
    assign P[162] = in[10] ^ in2[10];
    assign G[163] = in[9] & in2[9];
    assign P[163] = in[9] ^ in2[9];
    assign G[164] = in[8] & in2[8];
    assign P[164] = in[8] ^ in2[8];
    assign G[165] = in[7] & in2[7];
    assign P[165] = in[7] ^ in2[7];
    assign G[166] = in[6] & in2[6];
    assign P[166] = in[6] ^ in2[6];
    assign G[167] = in[5] & in2[5];
    assign P[167] = in[5] ^ in2[5];
    assign G[168] = in[4] & in2[4];
    assign P[168] = in[4] ^ in2[4];
    assign G[169] = in[3] & in2[3];
    assign P[169] = in[3] ^ in2[3];
    assign G[170] = in[2] & in2[2];
    assign P[170] = in[2] ^ in2[2];
    assign G[171] = in[1] & in2[1];
    assign P[171] = in[1] ^ in2[1];
    assign G[172] = in[0] & in2[0];
    assign P[172] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign C[172] = G[171] | (P[171] & C[171]);
    assign cout = G[172] | (P[172] & C[172]);
    assign sum = P ^ C;
endmodule

module CLA172(output [171:0] sum, output cout, input [171:0] in1, input [171:0] in2;

    wire[171:0] G;
    wire[171:0] C;
    wire[171:0] P;

    assign G[0] = in[171] & in2[171];
    assign P[0] = in[171] ^ in2[171];
    assign G[1] = in[170] & in2[170];
    assign P[1] = in[170] ^ in2[170];
    assign G[2] = in[169] & in2[169];
    assign P[2] = in[169] ^ in2[169];
    assign G[3] = in[168] & in2[168];
    assign P[3] = in[168] ^ in2[168];
    assign G[4] = in[167] & in2[167];
    assign P[4] = in[167] ^ in2[167];
    assign G[5] = in[166] & in2[166];
    assign P[5] = in[166] ^ in2[166];
    assign G[6] = in[165] & in2[165];
    assign P[6] = in[165] ^ in2[165];
    assign G[7] = in[164] & in2[164];
    assign P[7] = in[164] ^ in2[164];
    assign G[8] = in[163] & in2[163];
    assign P[8] = in[163] ^ in2[163];
    assign G[9] = in[162] & in2[162];
    assign P[9] = in[162] ^ in2[162];
    assign G[10] = in[161] & in2[161];
    assign P[10] = in[161] ^ in2[161];
    assign G[11] = in[160] & in2[160];
    assign P[11] = in[160] ^ in2[160];
    assign G[12] = in[159] & in2[159];
    assign P[12] = in[159] ^ in2[159];
    assign G[13] = in[158] & in2[158];
    assign P[13] = in[158] ^ in2[158];
    assign G[14] = in[157] & in2[157];
    assign P[14] = in[157] ^ in2[157];
    assign G[15] = in[156] & in2[156];
    assign P[15] = in[156] ^ in2[156];
    assign G[16] = in[155] & in2[155];
    assign P[16] = in[155] ^ in2[155];
    assign G[17] = in[154] & in2[154];
    assign P[17] = in[154] ^ in2[154];
    assign G[18] = in[153] & in2[153];
    assign P[18] = in[153] ^ in2[153];
    assign G[19] = in[152] & in2[152];
    assign P[19] = in[152] ^ in2[152];
    assign G[20] = in[151] & in2[151];
    assign P[20] = in[151] ^ in2[151];
    assign G[21] = in[150] & in2[150];
    assign P[21] = in[150] ^ in2[150];
    assign G[22] = in[149] & in2[149];
    assign P[22] = in[149] ^ in2[149];
    assign G[23] = in[148] & in2[148];
    assign P[23] = in[148] ^ in2[148];
    assign G[24] = in[147] & in2[147];
    assign P[24] = in[147] ^ in2[147];
    assign G[25] = in[146] & in2[146];
    assign P[25] = in[146] ^ in2[146];
    assign G[26] = in[145] & in2[145];
    assign P[26] = in[145] ^ in2[145];
    assign G[27] = in[144] & in2[144];
    assign P[27] = in[144] ^ in2[144];
    assign G[28] = in[143] & in2[143];
    assign P[28] = in[143] ^ in2[143];
    assign G[29] = in[142] & in2[142];
    assign P[29] = in[142] ^ in2[142];
    assign G[30] = in[141] & in2[141];
    assign P[30] = in[141] ^ in2[141];
    assign G[31] = in[140] & in2[140];
    assign P[31] = in[140] ^ in2[140];
    assign G[32] = in[139] & in2[139];
    assign P[32] = in[139] ^ in2[139];
    assign G[33] = in[138] & in2[138];
    assign P[33] = in[138] ^ in2[138];
    assign G[34] = in[137] & in2[137];
    assign P[34] = in[137] ^ in2[137];
    assign G[35] = in[136] & in2[136];
    assign P[35] = in[136] ^ in2[136];
    assign G[36] = in[135] & in2[135];
    assign P[36] = in[135] ^ in2[135];
    assign G[37] = in[134] & in2[134];
    assign P[37] = in[134] ^ in2[134];
    assign G[38] = in[133] & in2[133];
    assign P[38] = in[133] ^ in2[133];
    assign G[39] = in[132] & in2[132];
    assign P[39] = in[132] ^ in2[132];
    assign G[40] = in[131] & in2[131];
    assign P[40] = in[131] ^ in2[131];
    assign G[41] = in[130] & in2[130];
    assign P[41] = in[130] ^ in2[130];
    assign G[42] = in[129] & in2[129];
    assign P[42] = in[129] ^ in2[129];
    assign G[43] = in[128] & in2[128];
    assign P[43] = in[128] ^ in2[128];
    assign G[44] = in[127] & in2[127];
    assign P[44] = in[127] ^ in2[127];
    assign G[45] = in[126] & in2[126];
    assign P[45] = in[126] ^ in2[126];
    assign G[46] = in[125] & in2[125];
    assign P[46] = in[125] ^ in2[125];
    assign G[47] = in[124] & in2[124];
    assign P[47] = in[124] ^ in2[124];
    assign G[48] = in[123] & in2[123];
    assign P[48] = in[123] ^ in2[123];
    assign G[49] = in[122] & in2[122];
    assign P[49] = in[122] ^ in2[122];
    assign G[50] = in[121] & in2[121];
    assign P[50] = in[121] ^ in2[121];
    assign G[51] = in[120] & in2[120];
    assign P[51] = in[120] ^ in2[120];
    assign G[52] = in[119] & in2[119];
    assign P[52] = in[119] ^ in2[119];
    assign G[53] = in[118] & in2[118];
    assign P[53] = in[118] ^ in2[118];
    assign G[54] = in[117] & in2[117];
    assign P[54] = in[117] ^ in2[117];
    assign G[55] = in[116] & in2[116];
    assign P[55] = in[116] ^ in2[116];
    assign G[56] = in[115] & in2[115];
    assign P[56] = in[115] ^ in2[115];
    assign G[57] = in[114] & in2[114];
    assign P[57] = in[114] ^ in2[114];
    assign G[58] = in[113] & in2[113];
    assign P[58] = in[113] ^ in2[113];
    assign G[59] = in[112] & in2[112];
    assign P[59] = in[112] ^ in2[112];
    assign G[60] = in[111] & in2[111];
    assign P[60] = in[111] ^ in2[111];
    assign G[61] = in[110] & in2[110];
    assign P[61] = in[110] ^ in2[110];
    assign G[62] = in[109] & in2[109];
    assign P[62] = in[109] ^ in2[109];
    assign G[63] = in[108] & in2[108];
    assign P[63] = in[108] ^ in2[108];
    assign G[64] = in[107] & in2[107];
    assign P[64] = in[107] ^ in2[107];
    assign G[65] = in[106] & in2[106];
    assign P[65] = in[106] ^ in2[106];
    assign G[66] = in[105] & in2[105];
    assign P[66] = in[105] ^ in2[105];
    assign G[67] = in[104] & in2[104];
    assign P[67] = in[104] ^ in2[104];
    assign G[68] = in[103] & in2[103];
    assign P[68] = in[103] ^ in2[103];
    assign G[69] = in[102] & in2[102];
    assign P[69] = in[102] ^ in2[102];
    assign G[70] = in[101] & in2[101];
    assign P[70] = in[101] ^ in2[101];
    assign G[71] = in[100] & in2[100];
    assign P[71] = in[100] ^ in2[100];
    assign G[72] = in[99] & in2[99];
    assign P[72] = in[99] ^ in2[99];
    assign G[73] = in[98] & in2[98];
    assign P[73] = in[98] ^ in2[98];
    assign G[74] = in[97] & in2[97];
    assign P[74] = in[97] ^ in2[97];
    assign G[75] = in[96] & in2[96];
    assign P[75] = in[96] ^ in2[96];
    assign G[76] = in[95] & in2[95];
    assign P[76] = in[95] ^ in2[95];
    assign G[77] = in[94] & in2[94];
    assign P[77] = in[94] ^ in2[94];
    assign G[78] = in[93] & in2[93];
    assign P[78] = in[93] ^ in2[93];
    assign G[79] = in[92] & in2[92];
    assign P[79] = in[92] ^ in2[92];
    assign G[80] = in[91] & in2[91];
    assign P[80] = in[91] ^ in2[91];
    assign G[81] = in[90] & in2[90];
    assign P[81] = in[90] ^ in2[90];
    assign G[82] = in[89] & in2[89];
    assign P[82] = in[89] ^ in2[89];
    assign G[83] = in[88] & in2[88];
    assign P[83] = in[88] ^ in2[88];
    assign G[84] = in[87] & in2[87];
    assign P[84] = in[87] ^ in2[87];
    assign G[85] = in[86] & in2[86];
    assign P[85] = in[86] ^ in2[86];
    assign G[86] = in[85] & in2[85];
    assign P[86] = in[85] ^ in2[85];
    assign G[87] = in[84] & in2[84];
    assign P[87] = in[84] ^ in2[84];
    assign G[88] = in[83] & in2[83];
    assign P[88] = in[83] ^ in2[83];
    assign G[89] = in[82] & in2[82];
    assign P[89] = in[82] ^ in2[82];
    assign G[90] = in[81] & in2[81];
    assign P[90] = in[81] ^ in2[81];
    assign G[91] = in[80] & in2[80];
    assign P[91] = in[80] ^ in2[80];
    assign G[92] = in[79] & in2[79];
    assign P[92] = in[79] ^ in2[79];
    assign G[93] = in[78] & in2[78];
    assign P[93] = in[78] ^ in2[78];
    assign G[94] = in[77] & in2[77];
    assign P[94] = in[77] ^ in2[77];
    assign G[95] = in[76] & in2[76];
    assign P[95] = in[76] ^ in2[76];
    assign G[96] = in[75] & in2[75];
    assign P[96] = in[75] ^ in2[75];
    assign G[97] = in[74] & in2[74];
    assign P[97] = in[74] ^ in2[74];
    assign G[98] = in[73] & in2[73];
    assign P[98] = in[73] ^ in2[73];
    assign G[99] = in[72] & in2[72];
    assign P[99] = in[72] ^ in2[72];
    assign G[100] = in[71] & in2[71];
    assign P[100] = in[71] ^ in2[71];
    assign G[101] = in[70] & in2[70];
    assign P[101] = in[70] ^ in2[70];
    assign G[102] = in[69] & in2[69];
    assign P[102] = in[69] ^ in2[69];
    assign G[103] = in[68] & in2[68];
    assign P[103] = in[68] ^ in2[68];
    assign G[104] = in[67] & in2[67];
    assign P[104] = in[67] ^ in2[67];
    assign G[105] = in[66] & in2[66];
    assign P[105] = in[66] ^ in2[66];
    assign G[106] = in[65] & in2[65];
    assign P[106] = in[65] ^ in2[65];
    assign G[107] = in[64] & in2[64];
    assign P[107] = in[64] ^ in2[64];
    assign G[108] = in[63] & in2[63];
    assign P[108] = in[63] ^ in2[63];
    assign G[109] = in[62] & in2[62];
    assign P[109] = in[62] ^ in2[62];
    assign G[110] = in[61] & in2[61];
    assign P[110] = in[61] ^ in2[61];
    assign G[111] = in[60] & in2[60];
    assign P[111] = in[60] ^ in2[60];
    assign G[112] = in[59] & in2[59];
    assign P[112] = in[59] ^ in2[59];
    assign G[113] = in[58] & in2[58];
    assign P[113] = in[58] ^ in2[58];
    assign G[114] = in[57] & in2[57];
    assign P[114] = in[57] ^ in2[57];
    assign G[115] = in[56] & in2[56];
    assign P[115] = in[56] ^ in2[56];
    assign G[116] = in[55] & in2[55];
    assign P[116] = in[55] ^ in2[55];
    assign G[117] = in[54] & in2[54];
    assign P[117] = in[54] ^ in2[54];
    assign G[118] = in[53] & in2[53];
    assign P[118] = in[53] ^ in2[53];
    assign G[119] = in[52] & in2[52];
    assign P[119] = in[52] ^ in2[52];
    assign G[120] = in[51] & in2[51];
    assign P[120] = in[51] ^ in2[51];
    assign G[121] = in[50] & in2[50];
    assign P[121] = in[50] ^ in2[50];
    assign G[122] = in[49] & in2[49];
    assign P[122] = in[49] ^ in2[49];
    assign G[123] = in[48] & in2[48];
    assign P[123] = in[48] ^ in2[48];
    assign G[124] = in[47] & in2[47];
    assign P[124] = in[47] ^ in2[47];
    assign G[125] = in[46] & in2[46];
    assign P[125] = in[46] ^ in2[46];
    assign G[126] = in[45] & in2[45];
    assign P[126] = in[45] ^ in2[45];
    assign G[127] = in[44] & in2[44];
    assign P[127] = in[44] ^ in2[44];
    assign G[128] = in[43] & in2[43];
    assign P[128] = in[43] ^ in2[43];
    assign G[129] = in[42] & in2[42];
    assign P[129] = in[42] ^ in2[42];
    assign G[130] = in[41] & in2[41];
    assign P[130] = in[41] ^ in2[41];
    assign G[131] = in[40] & in2[40];
    assign P[131] = in[40] ^ in2[40];
    assign G[132] = in[39] & in2[39];
    assign P[132] = in[39] ^ in2[39];
    assign G[133] = in[38] & in2[38];
    assign P[133] = in[38] ^ in2[38];
    assign G[134] = in[37] & in2[37];
    assign P[134] = in[37] ^ in2[37];
    assign G[135] = in[36] & in2[36];
    assign P[135] = in[36] ^ in2[36];
    assign G[136] = in[35] & in2[35];
    assign P[136] = in[35] ^ in2[35];
    assign G[137] = in[34] & in2[34];
    assign P[137] = in[34] ^ in2[34];
    assign G[138] = in[33] & in2[33];
    assign P[138] = in[33] ^ in2[33];
    assign G[139] = in[32] & in2[32];
    assign P[139] = in[32] ^ in2[32];
    assign G[140] = in[31] & in2[31];
    assign P[140] = in[31] ^ in2[31];
    assign G[141] = in[30] & in2[30];
    assign P[141] = in[30] ^ in2[30];
    assign G[142] = in[29] & in2[29];
    assign P[142] = in[29] ^ in2[29];
    assign G[143] = in[28] & in2[28];
    assign P[143] = in[28] ^ in2[28];
    assign G[144] = in[27] & in2[27];
    assign P[144] = in[27] ^ in2[27];
    assign G[145] = in[26] & in2[26];
    assign P[145] = in[26] ^ in2[26];
    assign G[146] = in[25] & in2[25];
    assign P[146] = in[25] ^ in2[25];
    assign G[147] = in[24] & in2[24];
    assign P[147] = in[24] ^ in2[24];
    assign G[148] = in[23] & in2[23];
    assign P[148] = in[23] ^ in2[23];
    assign G[149] = in[22] & in2[22];
    assign P[149] = in[22] ^ in2[22];
    assign G[150] = in[21] & in2[21];
    assign P[150] = in[21] ^ in2[21];
    assign G[151] = in[20] & in2[20];
    assign P[151] = in[20] ^ in2[20];
    assign G[152] = in[19] & in2[19];
    assign P[152] = in[19] ^ in2[19];
    assign G[153] = in[18] & in2[18];
    assign P[153] = in[18] ^ in2[18];
    assign G[154] = in[17] & in2[17];
    assign P[154] = in[17] ^ in2[17];
    assign G[155] = in[16] & in2[16];
    assign P[155] = in[16] ^ in2[16];
    assign G[156] = in[15] & in2[15];
    assign P[156] = in[15] ^ in2[15];
    assign G[157] = in[14] & in2[14];
    assign P[157] = in[14] ^ in2[14];
    assign G[158] = in[13] & in2[13];
    assign P[158] = in[13] ^ in2[13];
    assign G[159] = in[12] & in2[12];
    assign P[159] = in[12] ^ in2[12];
    assign G[160] = in[11] & in2[11];
    assign P[160] = in[11] ^ in2[11];
    assign G[161] = in[10] & in2[10];
    assign P[161] = in[10] ^ in2[10];
    assign G[162] = in[9] & in2[9];
    assign P[162] = in[9] ^ in2[9];
    assign G[163] = in[8] & in2[8];
    assign P[163] = in[8] ^ in2[8];
    assign G[164] = in[7] & in2[7];
    assign P[164] = in[7] ^ in2[7];
    assign G[165] = in[6] & in2[6];
    assign P[165] = in[6] ^ in2[6];
    assign G[166] = in[5] & in2[5];
    assign P[166] = in[5] ^ in2[5];
    assign G[167] = in[4] & in2[4];
    assign P[167] = in[4] ^ in2[4];
    assign G[168] = in[3] & in2[3];
    assign P[168] = in[3] ^ in2[3];
    assign G[169] = in[2] & in2[2];
    assign P[169] = in[2] ^ in2[2];
    assign G[170] = in[1] & in2[1];
    assign P[170] = in[1] ^ in2[1];
    assign G[171] = in[0] & in2[0];
    assign P[171] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign C[171] = G[170] | (P[170] & C[170]);
    assign cout = G[171] | (P[171] & C[171]);
    assign sum = P ^ C;
endmodule

module CLA171(output [170:0] sum, output cout, input [170:0] in1, input [170:0] in2;

    wire[170:0] G;
    wire[170:0] C;
    wire[170:0] P;

    assign G[0] = in[170] & in2[170];
    assign P[0] = in[170] ^ in2[170];
    assign G[1] = in[169] & in2[169];
    assign P[1] = in[169] ^ in2[169];
    assign G[2] = in[168] & in2[168];
    assign P[2] = in[168] ^ in2[168];
    assign G[3] = in[167] & in2[167];
    assign P[3] = in[167] ^ in2[167];
    assign G[4] = in[166] & in2[166];
    assign P[4] = in[166] ^ in2[166];
    assign G[5] = in[165] & in2[165];
    assign P[5] = in[165] ^ in2[165];
    assign G[6] = in[164] & in2[164];
    assign P[6] = in[164] ^ in2[164];
    assign G[7] = in[163] & in2[163];
    assign P[7] = in[163] ^ in2[163];
    assign G[8] = in[162] & in2[162];
    assign P[8] = in[162] ^ in2[162];
    assign G[9] = in[161] & in2[161];
    assign P[9] = in[161] ^ in2[161];
    assign G[10] = in[160] & in2[160];
    assign P[10] = in[160] ^ in2[160];
    assign G[11] = in[159] & in2[159];
    assign P[11] = in[159] ^ in2[159];
    assign G[12] = in[158] & in2[158];
    assign P[12] = in[158] ^ in2[158];
    assign G[13] = in[157] & in2[157];
    assign P[13] = in[157] ^ in2[157];
    assign G[14] = in[156] & in2[156];
    assign P[14] = in[156] ^ in2[156];
    assign G[15] = in[155] & in2[155];
    assign P[15] = in[155] ^ in2[155];
    assign G[16] = in[154] & in2[154];
    assign P[16] = in[154] ^ in2[154];
    assign G[17] = in[153] & in2[153];
    assign P[17] = in[153] ^ in2[153];
    assign G[18] = in[152] & in2[152];
    assign P[18] = in[152] ^ in2[152];
    assign G[19] = in[151] & in2[151];
    assign P[19] = in[151] ^ in2[151];
    assign G[20] = in[150] & in2[150];
    assign P[20] = in[150] ^ in2[150];
    assign G[21] = in[149] & in2[149];
    assign P[21] = in[149] ^ in2[149];
    assign G[22] = in[148] & in2[148];
    assign P[22] = in[148] ^ in2[148];
    assign G[23] = in[147] & in2[147];
    assign P[23] = in[147] ^ in2[147];
    assign G[24] = in[146] & in2[146];
    assign P[24] = in[146] ^ in2[146];
    assign G[25] = in[145] & in2[145];
    assign P[25] = in[145] ^ in2[145];
    assign G[26] = in[144] & in2[144];
    assign P[26] = in[144] ^ in2[144];
    assign G[27] = in[143] & in2[143];
    assign P[27] = in[143] ^ in2[143];
    assign G[28] = in[142] & in2[142];
    assign P[28] = in[142] ^ in2[142];
    assign G[29] = in[141] & in2[141];
    assign P[29] = in[141] ^ in2[141];
    assign G[30] = in[140] & in2[140];
    assign P[30] = in[140] ^ in2[140];
    assign G[31] = in[139] & in2[139];
    assign P[31] = in[139] ^ in2[139];
    assign G[32] = in[138] & in2[138];
    assign P[32] = in[138] ^ in2[138];
    assign G[33] = in[137] & in2[137];
    assign P[33] = in[137] ^ in2[137];
    assign G[34] = in[136] & in2[136];
    assign P[34] = in[136] ^ in2[136];
    assign G[35] = in[135] & in2[135];
    assign P[35] = in[135] ^ in2[135];
    assign G[36] = in[134] & in2[134];
    assign P[36] = in[134] ^ in2[134];
    assign G[37] = in[133] & in2[133];
    assign P[37] = in[133] ^ in2[133];
    assign G[38] = in[132] & in2[132];
    assign P[38] = in[132] ^ in2[132];
    assign G[39] = in[131] & in2[131];
    assign P[39] = in[131] ^ in2[131];
    assign G[40] = in[130] & in2[130];
    assign P[40] = in[130] ^ in2[130];
    assign G[41] = in[129] & in2[129];
    assign P[41] = in[129] ^ in2[129];
    assign G[42] = in[128] & in2[128];
    assign P[42] = in[128] ^ in2[128];
    assign G[43] = in[127] & in2[127];
    assign P[43] = in[127] ^ in2[127];
    assign G[44] = in[126] & in2[126];
    assign P[44] = in[126] ^ in2[126];
    assign G[45] = in[125] & in2[125];
    assign P[45] = in[125] ^ in2[125];
    assign G[46] = in[124] & in2[124];
    assign P[46] = in[124] ^ in2[124];
    assign G[47] = in[123] & in2[123];
    assign P[47] = in[123] ^ in2[123];
    assign G[48] = in[122] & in2[122];
    assign P[48] = in[122] ^ in2[122];
    assign G[49] = in[121] & in2[121];
    assign P[49] = in[121] ^ in2[121];
    assign G[50] = in[120] & in2[120];
    assign P[50] = in[120] ^ in2[120];
    assign G[51] = in[119] & in2[119];
    assign P[51] = in[119] ^ in2[119];
    assign G[52] = in[118] & in2[118];
    assign P[52] = in[118] ^ in2[118];
    assign G[53] = in[117] & in2[117];
    assign P[53] = in[117] ^ in2[117];
    assign G[54] = in[116] & in2[116];
    assign P[54] = in[116] ^ in2[116];
    assign G[55] = in[115] & in2[115];
    assign P[55] = in[115] ^ in2[115];
    assign G[56] = in[114] & in2[114];
    assign P[56] = in[114] ^ in2[114];
    assign G[57] = in[113] & in2[113];
    assign P[57] = in[113] ^ in2[113];
    assign G[58] = in[112] & in2[112];
    assign P[58] = in[112] ^ in2[112];
    assign G[59] = in[111] & in2[111];
    assign P[59] = in[111] ^ in2[111];
    assign G[60] = in[110] & in2[110];
    assign P[60] = in[110] ^ in2[110];
    assign G[61] = in[109] & in2[109];
    assign P[61] = in[109] ^ in2[109];
    assign G[62] = in[108] & in2[108];
    assign P[62] = in[108] ^ in2[108];
    assign G[63] = in[107] & in2[107];
    assign P[63] = in[107] ^ in2[107];
    assign G[64] = in[106] & in2[106];
    assign P[64] = in[106] ^ in2[106];
    assign G[65] = in[105] & in2[105];
    assign P[65] = in[105] ^ in2[105];
    assign G[66] = in[104] & in2[104];
    assign P[66] = in[104] ^ in2[104];
    assign G[67] = in[103] & in2[103];
    assign P[67] = in[103] ^ in2[103];
    assign G[68] = in[102] & in2[102];
    assign P[68] = in[102] ^ in2[102];
    assign G[69] = in[101] & in2[101];
    assign P[69] = in[101] ^ in2[101];
    assign G[70] = in[100] & in2[100];
    assign P[70] = in[100] ^ in2[100];
    assign G[71] = in[99] & in2[99];
    assign P[71] = in[99] ^ in2[99];
    assign G[72] = in[98] & in2[98];
    assign P[72] = in[98] ^ in2[98];
    assign G[73] = in[97] & in2[97];
    assign P[73] = in[97] ^ in2[97];
    assign G[74] = in[96] & in2[96];
    assign P[74] = in[96] ^ in2[96];
    assign G[75] = in[95] & in2[95];
    assign P[75] = in[95] ^ in2[95];
    assign G[76] = in[94] & in2[94];
    assign P[76] = in[94] ^ in2[94];
    assign G[77] = in[93] & in2[93];
    assign P[77] = in[93] ^ in2[93];
    assign G[78] = in[92] & in2[92];
    assign P[78] = in[92] ^ in2[92];
    assign G[79] = in[91] & in2[91];
    assign P[79] = in[91] ^ in2[91];
    assign G[80] = in[90] & in2[90];
    assign P[80] = in[90] ^ in2[90];
    assign G[81] = in[89] & in2[89];
    assign P[81] = in[89] ^ in2[89];
    assign G[82] = in[88] & in2[88];
    assign P[82] = in[88] ^ in2[88];
    assign G[83] = in[87] & in2[87];
    assign P[83] = in[87] ^ in2[87];
    assign G[84] = in[86] & in2[86];
    assign P[84] = in[86] ^ in2[86];
    assign G[85] = in[85] & in2[85];
    assign P[85] = in[85] ^ in2[85];
    assign G[86] = in[84] & in2[84];
    assign P[86] = in[84] ^ in2[84];
    assign G[87] = in[83] & in2[83];
    assign P[87] = in[83] ^ in2[83];
    assign G[88] = in[82] & in2[82];
    assign P[88] = in[82] ^ in2[82];
    assign G[89] = in[81] & in2[81];
    assign P[89] = in[81] ^ in2[81];
    assign G[90] = in[80] & in2[80];
    assign P[90] = in[80] ^ in2[80];
    assign G[91] = in[79] & in2[79];
    assign P[91] = in[79] ^ in2[79];
    assign G[92] = in[78] & in2[78];
    assign P[92] = in[78] ^ in2[78];
    assign G[93] = in[77] & in2[77];
    assign P[93] = in[77] ^ in2[77];
    assign G[94] = in[76] & in2[76];
    assign P[94] = in[76] ^ in2[76];
    assign G[95] = in[75] & in2[75];
    assign P[95] = in[75] ^ in2[75];
    assign G[96] = in[74] & in2[74];
    assign P[96] = in[74] ^ in2[74];
    assign G[97] = in[73] & in2[73];
    assign P[97] = in[73] ^ in2[73];
    assign G[98] = in[72] & in2[72];
    assign P[98] = in[72] ^ in2[72];
    assign G[99] = in[71] & in2[71];
    assign P[99] = in[71] ^ in2[71];
    assign G[100] = in[70] & in2[70];
    assign P[100] = in[70] ^ in2[70];
    assign G[101] = in[69] & in2[69];
    assign P[101] = in[69] ^ in2[69];
    assign G[102] = in[68] & in2[68];
    assign P[102] = in[68] ^ in2[68];
    assign G[103] = in[67] & in2[67];
    assign P[103] = in[67] ^ in2[67];
    assign G[104] = in[66] & in2[66];
    assign P[104] = in[66] ^ in2[66];
    assign G[105] = in[65] & in2[65];
    assign P[105] = in[65] ^ in2[65];
    assign G[106] = in[64] & in2[64];
    assign P[106] = in[64] ^ in2[64];
    assign G[107] = in[63] & in2[63];
    assign P[107] = in[63] ^ in2[63];
    assign G[108] = in[62] & in2[62];
    assign P[108] = in[62] ^ in2[62];
    assign G[109] = in[61] & in2[61];
    assign P[109] = in[61] ^ in2[61];
    assign G[110] = in[60] & in2[60];
    assign P[110] = in[60] ^ in2[60];
    assign G[111] = in[59] & in2[59];
    assign P[111] = in[59] ^ in2[59];
    assign G[112] = in[58] & in2[58];
    assign P[112] = in[58] ^ in2[58];
    assign G[113] = in[57] & in2[57];
    assign P[113] = in[57] ^ in2[57];
    assign G[114] = in[56] & in2[56];
    assign P[114] = in[56] ^ in2[56];
    assign G[115] = in[55] & in2[55];
    assign P[115] = in[55] ^ in2[55];
    assign G[116] = in[54] & in2[54];
    assign P[116] = in[54] ^ in2[54];
    assign G[117] = in[53] & in2[53];
    assign P[117] = in[53] ^ in2[53];
    assign G[118] = in[52] & in2[52];
    assign P[118] = in[52] ^ in2[52];
    assign G[119] = in[51] & in2[51];
    assign P[119] = in[51] ^ in2[51];
    assign G[120] = in[50] & in2[50];
    assign P[120] = in[50] ^ in2[50];
    assign G[121] = in[49] & in2[49];
    assign P[121] = in[49] ^ in2[49];
    assign G[122] = in[48] & in2[48];
    assign P[122] = in[48] ^ in2[48];
    assign G[123] = in[47] & in2[47];
    assign P[123] = in[47] ^ in2[47];
    assign G[124] = in[46] & in2[46];
    assign P[124] = in[46] ^ in2[46];
    assign G[125] = in[45] & in2[45];
    assign P[125] = in[45] ^ in2[45];
    assign G[126] = in[44] & in2[44];
    assign P[126] = in[44] ^ in2[44];
    assign G[127] = in[43] & in2[43];
    assign P[127] = in[43] ^ in2[43];
    assign G[128] = in[42] & in2[42];
    assign P[128] = in[42] ^ in2[42];
    assign G[129] = in[41] & in2[41];
    assign P[129] = in[41] ^ in2[41];
    assign G[130] = in[40] & in2[40];
    assign P[130] = in[40] ^ in2[40];
    assign G[131] = in[39] & in2[39];
    assign P[131] = in[39] ^ in2[39];
    assign G[132] = in[38] & in2[38];
    assign P[132] = in[38] ^ in2[38];
    assign G[133] = in[37] & in2[37];
    assign P[133] = in[37] ^ in2[37];
    assign G[134] = in[36] & in2[36];
    assign P[134] = in[36] ^ in2[36];
    assign G[135] = in[35] & in2[35];
    assign P[135] = in[35] ^ in2[35];
    assign G[136] = in[34] & in2[34];
    assign P[136] = in[34] ^ in2[34];
    assign G[137] = in[33] & in2[33];
    assign P[137] = in[33] ^ in2[33];
    assign G[138] = in[32] & in2[32];
    assign P[138] = in[32] ^ in2[32];
    assign G[139] = in[31] & in2[31];
    assign P[139] = in[31] ^ in2[31];
    assign G[140] = in[30] & in2[30];
    assign P[140] = in[30] ^ in2[30];
    assign G[141] = in[29] & in2[29];
    assign P[141] = in[29] ^ in2[29];
    assign G[142] = in[28] & in2[28];
    assign P[142] = in[28] ^ in2[28];
    assign G[143] = in[27] & in2[27];
    assign P[143] = in[27] ^ in2[27];
    assign G[144] = in[26] & in2[26];
    assign P[144] = in[26] ^ in2[26];
    assign G[145] = in[25] & in2[25];
    assign P[145] = in[25] ^ in2[25];
    assign G[146] = in[24] & in2[24];
    assign P[146] = in[24] ^ in2[24];
    assign G[147] = in[23] & in2[23];
    assign P[147] = in[23] ^ in2[23];
    assign G[148] = in[22] & in2[22];
    assign P[148] = in[22] ^ in2[22];
    assign G[149] = in[21] & in2[21];
    assign P[149] = in[21] ^ in2[21];
    assign G[150] = in[20] & in2[20];
    assign P[150] = in[20] ^ in2[20];
    assign G[151] = in[19] & in2[19];
    assign P[151] = in[19] ^ in2[19];
    assign G[152] = in[18] & in2[18];
    assign P[152] = in[18] ^ in2[18];
    assign G[153] = in[17] & in2[17];
    assign P[153] = in[17] ^ in2[17];
    assign G[154] = in[16] & in2[16];
    assign P[154] = in[16] ^ in2[16];
    assign G[155] = in[15] & in2[15];
    assign P[155] = in[15] ^ in2[15];
    assign G[156] = in[14] & in2[14];
    assign P[156] = in[14] ^ in2[14];
    assign G[157] = in[13] & in2[13];
    assign P[157] = in[13] ^ in2[13];
    assign G[158] = in[12] & in2[12];
    assign P[158] = in[12] ^ in2[12];
    assign G[159] = in[11] & in2[11];
    assign P[159] = in[11] ^ in2[11];
    assign G[160] = in[10] & in2[10];
    assign P[160] = in[10] ^ in2[10];
    assign G[161] = in[9] & in2[9];
    assign P[161] = in[9] ^ in2[9];
    assign G[162] = in[8] & in2[8];
    assign P[162] = in[8] ^ in2[8];
    assign G[163] = in[7] & in2[7];
    assign P[163] = in[7] ^ in2[7];
    assign G[164] = in[6] & in2[6];
    assign P[164] = in[6] ^ in2[6];
    assign G[165] = in[5] & in2[5];
    assign P[165] = in[5] ^ in2[5];
    assign G[166] = in[4] & in2[4];
    assign P[166] = in[4] ^ in2[4];
    assign G[167] = in[3] & in2[3];
    assign P[167] = in[3] ^ in2[3];
    assign G[168] = in[2] & in2[2];
    assign P[168] = in[2] ^ in2[2];
    assign G[169] = in[1] & in2[1];
    assign P[169] = in[1] ^ in2[1];
    assign G[170] = in[0] & in2[0];
    assign P[170] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign C[170] = G[169] | (P[169] & C[169]);
    assign cout = G[170] | (P[170] & C[170]);
    assign sum = P ^ C;
endmodule

module CLA170(output [169:0] sum, output cout, input [169:0] in1, input [169:0] in2;

    wire[169:0] G;
    wire[169:0] C;
    wire[169:0] P;

    assign G[0] = in[169] & in2[169];
    assign P[0] = in[169] ^ in2[169];
    assign G[1] = in[168] & in2[168];
    assign P[1] = in[168] ^ in2[168];
    assign G[2] = in[167] & in2[167];
    assign P[2] = in[167] ^ in2[167];
    assign G[3] = in[166] & in2[166];
    assign P[3] = in[166] ^ in2[166];
    assign G[4] = in[165] & in2[165];
    assign P[4] = in[165] ^ in2[165];
    assign G[5] = in[164] & in2[164];
    assign P[5] = in[164] ^ in2[164];
    assign G[6] = in[163] & in2[163];
    assign P[6] = in[163] ^ in2[163];
    assign G[7] = in[162] & in2[162];
    assign P[7] = in[162] ^ in2[162];
    assign G[8] = in[161] & in2[161];
    assign P[8] = in[161] ^ in2[161];
    assign G[9] = in[160] & in2[160];
    assign P[9] = in[160] ^ in2[160];
    assign G[10] = in[159] & in2[159];
    assign P[10] = in[159] ^ in2[159];
    assign G[11] = in[158] & in2[158];
    assign P[11] = in[158] ^ in2[158];
    assign G[12] = in[157] & in2[157];
    assign P[12] = in[157] ^ in2[157];
    assign G[13] = in[156] & in2[156];
    assign P[13] = in[156] ^ in2[156];
    assign G[14] = in[155] & in2[155];
    assign P[14] = in[155] ^ in2[155];
    assign G[15] = in[154] & in2[154];
    assign P[15] = in[154] ^ in2[154];
    assign G[16] = in[153] & in2[153];
    assign P[16] = in[153] ^ in2[153];
    assign G[17] = in[152] & in2[152];
    assign P[17] = in[152] ^ in2[152];
    assign G[18] = in[151] & in2[151];
    assign P[18] = in[151] ^ in2[151];
    assign G[19] = in[150] & in2[150];
    assign P[19] = in[150] ^ in2[150];
    assign G[20] = in[149] & in2[149];
    assign P[20] = in[149] ^ in2[149];
    assign G[21] = in[148] & in2[148];
    assign P[21] = in[148] ^ in2[148];
    assign G[22] = in[147] & in2[147];
    assign P[22] = in[147] ^ in2[147];
    assign G[23] = in[146] & in2[146];
    assign P[23] = in[146] ^ in2[146];
    assign G[24] = in[145] & in2[145];
    assign P[24] = in[145] ^ in2[145];
    assign G[25] = in[144] & in2[144];
    assign P[25] = in[144] ^ in2[144];
    assign G[26] = in[143] & in2[143];
    assign P[26] = in[143] ^ in2[143];
    assign G[27] = in[142] & in2[142];
    assign P[27] = in[142] ^ in2[142];
    assign G[28] = in[141] & in2[141];
    assign P[28] = in[141] ^ in2[141];
    assign G[29] = in[140] & in2[140];
    assign P[29] = in[140] ^ in2[140];
    assign G[30] = in[139] & in2[139];
    assign P[30] = in[139] ^ in2[139];
    assign G[31] = in[138] & in2[138];
    assign P[31] = in[138] ^ in2[138];
    assign G[32] = in[137] & in2[137];
    assign P[32] = in[137] ^ in2[137];
    assign G[33] = in[136] & in2[136];
    assign P[33] = in[136] ^ in2[136];
    assign G[34] = in[135] & in2[135];
    assign P[34] = in[135] ^ in2[135];
    assign G[35] = in[134] & in2[134];
    assign P[35] = in[134] ^ in2[134];
    assign G[36] = in[133] & in2[133];
    assign P[36] = in[133] ^ in2[133];
    assign G[37] = in[132] & in2[132];
    assign P[37] = in[132] ^ in2[132];
    assign G[38] = in[131] & in2[131];
    assign P[38] = in[131] ^ in2[131];
    assign G[39] = in[130] & in2[130];
    assign P[39] = in[130] ^ in2[130];
    assign G[40] = in[129] & in2[129];
    assign P[40] = in[129] ^ in2[129];
    assign G[41] = in[128] & in2[128];
    assign P[41] = in[128] ^ in2[128];
    assign G[42] = in[127] & in2[127];
    assign P[42] = in[127] ^ in2[127];
    assign G[43] = in[126] & in2[126];
    assign P[43] = in[126] ^ in2[126];
    assign G[44] = in[125] & in2[125];
    assign P[44] = in[125] ^ in2[125];
    assign G[45] = in[124] & in2[124];
    assign P[45] = in[124] ^ in2[124];
    assign G[46] = in[123] & in2[123];
    assign P[46] = in[123] ^ in2[123];
    assign G[47] = in[122] & in2[122];
    assign P[47] = in[122] ^ in2[122];
    assign G[48] = in[121] & in2[121];
    assign P[48] = in[121] ^ in2[121];
    assign G[49] = in[120] & in2[120];
    assign P[49] = in[120] ^ in2[120];
    assign G[50] = in[119] & in2[119];
    assign P[50] = in[119] ^ in2[119];
    assign G[51] = in[118] & in2[118];
    assign P[51] = in[118] ^ in2[118];
    assign G[52] = in[117] & in2[117];
    assign P[52] = in[117] ^ in2[117];
    assign G[53] = in[116] & in2[116];
    assign P[53] = in[116] ^ in2[116];
    assign G[54] = in[115] & in2[115];
    assign P[54] = in[115] ^ in2[115];
    assign G[55] = in[114] & in2[114];
    assign P[55] = in[114] ^ in2[114];
    assign G[56] = in[113] & in2[113];
    assign P[56] = in[113] ^ in2[113];
    assign G[57] = in[112] & in2[112];
    assign P[57] = in[112] ^ in2[112];
    assign G[58] = in[111] & in2[111];
    assign P[58] = in[111] ^ in2[111];
    assign G[59] = in[110] & in2[110];
    assign P[59] = in[110] ^ in2[110];
    assign G[60] = in[109] & in2[109];
    assign P[60] = in[109] ^ in2[109];
    assign G[61] = in[108] & in2[108];
    assign P[61] = in[108] ^ in2[108];
    assign G[62] = in[107] & in2[107];
    assign P[62] = in[107] ^ in2[107];
    assign G[63] = in[106] & in2[106];
    assign P[63] = in[106] ^ in2[106];
    assign G[64] = in[105] & in2[105];
    assign P[64] = in[105] ^ in2[105];
    assign G[65] = in[104] & in2[104];
    assign P[65] = in[104] ^ in2[104];
    assign G[66] = in[103] & in2[103];
    assign P[66] = in[103] ^ in2[103];
    assign G[67] = in[102] & in2[102];
    assign P[67] = in[102] ^ in2[102];
    assign G[68] = in[101] & in2[101];
    assign P[68] = in[101] ^ in2[101];
    assign G[69] = in[100] & in2[100];
    assign P[69] = in[100] ^ in2[100];
    assign G[70] = in[99] & in2[99];
    assign P[70] = in[99] ^ in2[99];
    assign G[71] = in[98] & in2[98];
    assign P[71] = in[98] ^ in2[98];
    assign G[72] = in[97] & in2[97];
    assign P[72] = in[97] ^ in2[97];
    assign G[73] = in[96] & in2[96];
    assign P[73] = in[96] ^ in2[96];
    assign G[74] = in[95] & in2[95];
    assign P[74] = in[95] ^ in2[95];
    assign G[75] = in[94] & in2[94];
    assign P[75] = in[94] ^ in2[94];
    assign G[76] = in[93] & in2[93];
    assign P[76] = in[93] ^ in2[93];
    assign G[77] = in[92] & in2[92];
    assign P[77] = in[92] ^ in2[92];
    assign G[78] = in[91] & in2[91];
    assign P[78] = in[91] ^ in2[91];
    assign G[79] = in[90] & in2[90];
    assign P[79] = in[90] ^ in2[90];
    assign G[80] = in[89] & in2[89];
    assign P[80] = in[89] ^ in2[89];
    assign G[81] = in[88] & in2[88];
    assign P[81] = in[88] ^ in2[88];
    assign G[82] = in[87] & in2[87];
    assign P[82] = in[87] ^ in2[87];
    assign G[83] = in[86] & in2[86];
    assign P[83] = in[86] ^ in2[86];
    assign G[84] = in[85] & in2[85];
    assign P[84] = in[85] ^ in2[85];
    assign G[85] = in[84] & in2[84];
    assign P[85] = in[84] ^ in2[84];
    assign G[86] = in[83] & in2[83];
    assign P[86] = in[83] ^ in2[83];
    assign G[87] = in[82] & in2[82];
    assign P[87] = in[82] ^ in2[82];
    assign G[88] = in[81] & in2[81];
    assign P[88] = in[81] ^ in2[81];
    assign G[89] = in[80] & in2[80];
    assign P[89] = in[80] ^ in2[80];
    assign G[90] = in[79] & in2[79];
    assign P[90] = in[79] ^ in2[79];
    assign G[91] = in[78] & in2[78];
    assign P[91] = in[78] ^ in2[78];
    assign G[92] = in[77] & in2[77];
    assign P[92] = in[77] ^ in2[77];
    assign G[93] = in[76] & in2[76];
    assign P[93] = in[76] ^ in2[76];
    assign G[94] = in[75] & in2[75];
    assign P[94] = in[75] ^ in2[75];
    assign G[95] = in[74] & in2[74];
    assign P[95] = in[74] ^ in2[74];
    assign G[96] = in[73] & in2[73];
    assign P[96] = in[73] ^ in2[73];
    assign G[97] = in[72] & in2[72];
    assign P[97] = in[72] ^ in2[72];
    assign G[98] = in[71] & in2[71];
    assign P[98] = in[71] ^ in2[71];
    assign G[99] = in[70] & in2[70];
    assign P[99] = in[70] ^ in2[70];
    assign G[100] = in[69] & in2[69];
    assign P[100] = in[69] ^ in2[69];
    assign G[101] = in[68] & in2[68];
    assign P[101] = in[68] ^ in2[68];
    assign G[102] = in[67] & in2[67];
    assign P[102] = in[67] ^ in2[67];
    assign G[103] = in[66] & in2[66];
    assign P[103] = in[66] ^ in2[66];
    assign G[104] = in[65] & in2[65];
    assign P[104] = in[65] ^ in2[65];
    assign G[105] = in[64] & in2[64];
    assign P[105] = in[64] ^ in2[64];
    assign G[106] = in[63] & in2[63];
    assign P[106] = in[63] ^ in2[63];
    assign G[107] = in[62] & in2[62];
    assign P[107] = in[62] ^ in2[62];
    assign G[108] = in[61] & in2[61];
    assign P[108] = in[61] ^ in2[61];
    assign G[109] = in[60] & in2[60];
    assign P[109] = in[60] ^ in2[60];
    assign G[110] = in[59] & in2[59];
    assign P[110] = in[59] ^ in2[59];
    assign G[111] = in[58] & in2[58];
    assign P[111] = in[58] ^ in2[58];
    assign G[112] = in[57] & in2[57];
    assign P[112] = in[57] ^ in2[57];
    assign G[113] = in[56] & in2[56];
    assign P[113] = in[56] ^ in2[56];
    assign G[114] = in[55] & in2[55];
    assign P[114] = in[55] ^ in2[55];
    assign G[115] = in[54] & in2[54];
    assign P[115] = in[54] ^ in2[54];
    assign G[116] = in[53] & in2[53];
    assign P[116] = in[53] ^ in2[53];
    assign G[117] = in[52] & in2[52];
    assign P[117] = in[52] ^ in2[52];
    assign G[118] = in[51] & in2[51];
    assign P[118] = in[51] ^ in2[51];
    assign G[119] = in[50] & in2[50];
    assign P[119] = in[50] ^ in2[50];
    assign G[120] = in[49] & in2[49];
    assign P[120] = in[49] ^ in2[49];
    assign G[121] = in[48] & in2[48];
    assign P[121] = in[48] ^ in2[48];
    assign G[122] = in[47] & in2[47];
    assign P[122] = in[47] ^ in2[47];
    assign G[123] = in[46] & in2[46];
    assign P[123] = in[46] ^ in2[46];
    assign G[124] = in[45] & in2[45];
    assign P[124] = in[45] ^ in2[45];
    assign G[125] = in[44] & in2[44];
    assign P[125] = in[44] ^ in2[44];
    assign G[126] = in[43] & in2[43];
    assign P[126] = in[43] ^ in2[43];
    assign G[127] = in[42] & in2[42];
    assign P[127] = in[42] ^ in2[42];
    assign G[128] = in[41] & in2[41];
    assign P[128] = in[41] ^ in2[41];
    assign G[129] = in[40] & in2[40];
    assign P[129] = in[40] ^ in2[40];
    assign G[130] = in[39] & in2[39];
    assign P[130] = in[39] ^ in2[39];
    assign G[131] = in[38] & in2[38];
    assign P[131] = in[38] ^ in2[38];
    assign G[132] = in[37] & in2[37];
    assign P[132] = in[37] ^ in2[37];
    assign G[133] = in[36] & in2[36];
    assign P[133] = in[36] ^ in2[36];
    assign G[134] = in[35] & in2[35];
    assign P[134] = in[35] ^ in2[35];
    assign G[135] = in[34] & in2[34];
    assign P[135] = in[34] ^ in2[34];
    assign G[136] = in[33] & in2[33];
    assign P[136] = in[33] ^ in2[33];
    assign G[137] = in[32] & in2[32];
    assign P[137] = in[32] ^ in2[32];
    assign G[138] = in[31] & in2[31];
    assign P[138] = in[31] ^ in2[31];
    assign G[139] = in[30] & in2[30];
    assign P[139] = in[30] ^ in2[30];
    assign G[140] = in[29] & in2[29];
    assign P[140] = in[29] ^ in2[29];
    assign G[141] = in[28] & in2[28];
    assign P[141] = in[28] ^ in2[28];
    assign G[142] = in[27] & in2[27];
    assign P[142] = in[27] ^ in2[27];
    assign G[143] = in[26] & in2[26];
    assign P[143] = in[26] ^ in2[26];
    assign G[144] = in[25] & in2[25];
    assign P[144] = in[25] ^ in2[25];
    assign G[145] = in[24] & in2[24];
    assign P[145] = in[24] ^ in2[24];
    assign G[146] = in[23] & in2[23];
    assign P[146] = in[23] ^ in2[23];
    assign G[147] = in[22] & in2[22];
    assign P[147] = in[22] ^ in2[22];
    assign G[148] = in[21] & in2[21];
    assign P[148] = in[21] ^ in2[21];
    assign G[149] = in[20] & in2[20];
    assign P[149] = in[20] ^ in2[20];
    assign G[150] = in[19] & in2[19];
    assign P[150] = in[19] ^ in2[19];
    assign G[151] = in[18] & in2[18];
    assign P[151] = in[18] ^ in2[18];
    assign G[152] = in[17] & in2[17];
    assign P[152] = in[17] ^ in2[17];
    assign G[153] = in[16] & in2[16];
    assign P[153] = in[16] ^ in2[16];
    assign G[154] = in[15] & in2[15];
    assign P[154] = in[15] ^ in2[15];
    assign G[155] = in[14] & in2[14];
    assign P[155] = in[14] ^ in2[14];
    assign G[156] = in[13] & in2[13];
    assign P[156] = in[13] ^ in2[13];
    assign G[157] = in[12] & in2[12];
    assign P[157] = in[12] ^ in2[12];
    assign G[158] = in[11] & in2[11];
    assign P[158] = in[11] ^ in2[11];
    assign G[159] = in[10] & in2[10];
    assign P[159] = in[10] ^ in2[10];
    assign G[160] = in[9] & in2[9];
    assign P[160] = in[9] ^ in2[9];
    assign G[161] = in[8] & in2[8];
    assign P[161] = in[8] ^ in2[8];
    assign G[162] = in[7] & in2[7];
    assign P[162] = in[7] ^ in2[7];
    assign G[163] = in[6] & in2[6];
    assign P[163] = in[6] ^ in2[6];
    assign G[164] = in[5] & in2[5];
    assign P[164] = in[5] ^ in2[5];
    assign G[165] = in[4] & in2[4];
    assign P[165] = in[4] ^ in2[4];
    assign G[166] = in[3] & in2[3];
    assign P[166] = in[3] ^ in2[3];
    assign G[167] = in[2] & in2[2];
    assign P[167] = in[2] ^ in2[2];
    assign G[168] = in[1] & in2[1];
    assign P[168] = in[1] ^ in2[1];
    assign G[169] = in[0] & in2[0];
    assign P[169] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign C[169] = G[168] | (P[168] & C[168]);
    assign cout = G[169] | (P[169] & C[169]);
    assign sum = P ^ C;
endmodule

module CLA169(output [168:0] sum, output cout, input [168:0] in1, input [168:0] in2;

    wire[168:0] G;
    wire[168:0] C;
    wire[168:0] P;

    assign G[0] = in[168] & in2[168];
    assign P[0] = in[168] ^ in2[168];
    assign G[1] = in[167] & in2[167];
    assign P[1] = in[167] ^ in2[167];
    assign G[2] = in[166] & in2[166];
    assign P[2] = in[166] ^ in2[166];
    assign G[3] = in[165] & in2[165];
    assign P[3] = in[165] ^ in2[165];
    assign G[4] = in[164] & in2[164];
    assign P[4] = in[164] ^ in2[164];
    assign G[5] = in[163] & in2[163];
    assign P[5] = in[163] ^ in2[163];
    assign G[6] = in[162] & in2[162];
    assign P[6] = in[162] ^ in2[162];
    assign G[7] = in[161] & in2[161];
    assign P[7] = in[161] ^ in2[161];
    assign G[8] = in[160] & in2[160];
    assign P[8] = in[160] ^ in2[160];
    assign G[9] = in[159] & in2[159];
    assign P[9] = in[159] ^ in2[159];
    assign G[10] = in[158] & in2[158];
    assign P[10] = in[158] ^ in2[158];
    assign G[11] = in[157] & in2[157];
    assign P[11] = in[157] ^ in2[157];
    assign G[12] = in[156] & in2[156];
    assign P[12] = in[156] ^ in2[156];
    assign G[13] = in[155] & in2[155];
    assign P[13] = in[155] ^ in2[155];
    assign G[14] = in[154] & in2[154];
    assign P[14] = in[154] ^ in2[154];
    assign G[15] = in[153] & in2[153];
    assign P[15] = in[153] ^ in2[153];
    assign G[16] = in[152] & in2[152];
    assign P[16] = in[152] ^ in2[152];
    assign G[17] = in[151] & in2[151];
    assign P[17] = in[151] ^ in2[151];
    assign G[18] = in[150] & in2[150];
    assign P[18] = in[150] ^ in2[150];
    assign G[19] = in[149] & in2[149];
    assign P[19] = in[149] ^ in2[149];
    assign G[20] = in[148] & in2[148];
    assign P[20] = in[148] ^ in2[148];
    assign G[21] = in[147] & in2[147];
    assign P[21] = in[147] ^ in2[147];
    assign G[22] = in[146] & in2[146];
    assign P[22] = in[146] ^ in2[146];
    assign G[23] = in[145] & in2[145];
    assign P[23] = in[145] ^ in2[145];
    assign G[24] = in[144] & in2[144];
    assign P[24] = in[144] ^ in2[144];
    assign G[25] = in[143] & in2[143];
    assign P[25] = in[143] ^ in2[143];
    assign G[26] = in[142] & in2[142];
    assign P[26] = in[142] ^ in2[142];
    assign G[27] = in[141] & in2[141];
    assign P[27] = in[141] ^ in2[141];
    assign G[28] = in[140] & in2[140];
    assign P[28] = in[140] ^ in2[140];
    assign G[29] = in[139] & in2[139];
    assign P[29] = in[139] ^ in2[139];
    assign G[30] = in[138] & in2[138];
    assign P[30] = in[138] ^ in2[138];
    assign G[31] = in[137] & in2[137];
    assign P[31] = in[137] ^ in2[137];
    assign G[32] = in[136] & in2[136];
    assign P[32] = in[136] ^ in2[136];
    assign G[33] = in[135] & in2[135];
    assign P[33] = in[135] ^ in2[135];
    assign G[34] = in[134] & in2[134];
    assign P[34] = in[134] ^ in2[134];
    assign G[35] = in[133] & in2[133];
    assign P[35] = in[133] ^ in2[133];
    assign G[36] = in[132] & in2[132];
    assign P[36] = in[132] ^ in2[132];
    assign G[37] = in[131] & in2[131];
    assign P[37] = in[131] ^ in2[131];
    assign G[38] = in[130] & in2[130];
    assign P[38] = in[130] ^ in2[130];
    assign G[39] = in[129] & in2[129];
    assign P[39] = in[129] ^ in2[129];
    assign G[40] = in[128] & in2[128];
    assign P[40] = in[128] ^ in2[128];
    assign G[41] = in[127] & in2[127];
    assign P[41] = in[127] ^ in2[127];
    assign G[42] = in[126] & in2[126];
    assign P[42] = in[126] ^ in2[126];
    assign G[43] = in[125] & in2[125];
    assign P[43] = in[125] ^ in2[125];
    assign G[44] = in[124] & in2[124];
    assign P[44] = in[124] ^ in2[124];
    assign G[45] = in[123] & in2[123];
    assign P[45] = in[123] ^ in2[123];
    assign G[46] = in[122] & in2[122];
    assign P[46] = in[122] ^ in2[122];
    assign G[47] = in[121] & in2[121];
    assign P[47] = in[121] ^ in2[121];
    assign G[48] = in[120] & in2[120];
    assign P[48] = in[120] ^ in2[120];
    assign G[49] = in[119] & in2[119];
    assign P[49] = in[119] ^ in2[119];
    assign G[50] = in[118] & in2[118];
    assign P[50] = in[118] ^ in2[118];
    assign G[51] = in[117] & in2[117];
    assign P[51] = in[117] ^ in2[117];
    assign G[52] = in[116] & in2[116];
    assign P[52] = in[116] ^ in2[116];
    assign G[53] = in[115] & in2[115];
    assign P[53] = in[115] ^ in2[115];
    assign G[54] = in[114] & in2[114];
    assign P[54] = in[114] ^ in2[114];
    assign G[55] = in[113] & in2[113];
    assign P[55] = in[113] ^ in2[113];
    assign G[56] = in[112] & in2[112];
    assign P[56] = in[112] ^ in2[112];
    assign G[57] = in[111] & in2[111];
    assign P[57] = in[111] ^ in2[111];
    assign G[58] = in[110] & in2[110];
    assign P[58] = in[110] ^ in2[110];
    assign G[59] = in[109] & in2[109];
    assign P[59] = in[109] ^ in2[109];
    assign G[60] = in[108] & in2[108];
    assign P[60] = in[108] ^ in2[108];
    assign G[61] = in[107] & in2[107];
    assign P[61] = in[107] ^ in2[107];
    assign G[62] = in[106] & in2[106];
    assign P[62] = in[106] ^ in2[106];
    assign G[63] = in[105] & in2[105];
    assign P[63] = in[105] ^ in2[105];
    assign G[64] = in[104] & in2[104];
    assign P[64] = in[104] ^ in2[104];
    assign G[65] = in[103] & in2[103];
    assign P[65] = in[103] ^ in2[103];
    assign G[66] = in[102] & in2[102];
    assign P[66] = in[102] ^ in2[102];
    assign G[67] = in[101] & in2[101];
    assign P[67] = in[101] ^ in2[101];
    assign G[68] = in[100] & in2[100];
    assign P[68] = in[100] ^ in2[100];
    assign G[69] = in[99] & in2[99];
    assign P[69] = in[99] ^ in2[99];
    assign G[70] = in[98] & in2[98];
    assign P[70] = in[98] ^ in2[98];
    assign G[71] = in[97] & in2[97];
    assign P[71] = in[97] ^ in2[97];
    assign G[72] = in[96] & in2[96];
    assign P[72] = in[96] ^ in2[96];
    assign G[73] = in[95] & in2[95];
    assign P[73] = in[95] ^ in2[95];
    assign G[74] = in[94] & in2[94];
    assign P[74] = in[94] ^ in2[94];
    assign G[75] = in[93] & in2[93];
    assign P[75] = in[93] ^ in2[93];
    assign G[76] = in[92] & in2[92];
    assign P[76] = in[92] ^ in2[92];
    assign G[77] = in[91] & in2[91];
    assign P[77] = in[91] ^ in2[91];
    assign G[78] = in[90] & in2[90];
    assign P[78] = in[90] ^ in2[90];
    assign G[79] = in[89] & in2[89];
    assign P[79] = in[89] ^ in2[89];
    assign G[80] = in[88] & in2[88];
    assign P[80] = in[88] ^ in2[88];
    assign G[81] = in[87] & in2[87];
    assign P[81] = in[87] ^ in2[87];
    assign G[82] = in[86] & in2[86];
    assign P[82] = in[86] ^ in2[86];
    assign G[83] = in[85] & in2[85];
    assign P[83] = in[85] ^ in2[85];
    assign G[84] = in[84] & in2[84];
    assign P[84] = in[84] ^ in2[84];
    assign G[85] = in[83] & in2[83];
    assign P[85] = in[83] ^ in2[83];
    assign G[86] = in[82] & in2[82];
    assign P[86] = in[82] ^ in2[82];
    assign G[87] = in[81] & in2[81];
    assign P[87] = in[81] ^ in2[81];
    assign G[88] = in[80] & in2[80];
    assign P[88] = in[80] ^ in2[80];
    assign G[89] = in[79] & in2[79];
    assign P[89] = in[79] ^ in2[79];
    assign G[90] = in[78] & in2[78];
    assign P[90] = in[78] ^ in2[78];
    assign G[91] = in[77] & in2[77];
    assign P[91] = in[77] ^ in2[77];
    assign G[92] = in[76] & in2[76];
    assign P[92] = in[76] ^ in2[76];
    assign G[93] = in[75] & in2[75];
    assign P[93] = in[75] ^ in2[75];
    assign G[94] = in[74] & in2[74];
    assign P[94] = in[74] ^ in2[74];
    assign G[95] = in[73] & in2[73];
    assign P[95] = in[73] ^ in2[73];
    assign G[96] = in[72] & in2[72];
    assign P[96] = in[72] ^ in2[72];
    assign G[97] = in[71] & in2[71];
    assign P[97] = in[71] ^ in2[71];
    assign G[98] = in[70] & in2[70];
    assign P[98] = in[70] ^ in2[70];
    assign G[99] = in[69] & in2[69];
    assign P[99] = in[69] ^ in2[69];
    assign G[100] = in[68] & in2[68];
    assign P[100] = in[68] ^ in2[68];
    assign G[101] = in[67] & in2[67];
    assign P[101] = in[67] ^ in2[67];
    assign G[102] = in[66] & in2[66];
    assign P[102] = in[66] ^ in2[66];
    assign G[103] = in[65] & in2[65];
    assign P[103] = in[65] ^ in2[65];
    assign G[104] = in[64] & in2[64];
    assign P[104] = in[64] ^ in2[64];
    assign G[105] = in[63] & in2[63];
    assign P[105] = in[63] ^ in2[63];
    assign G[106] = in[62] & in2[62];
    assign P[106] = in[62] ^ in2[62];
    assign G[107] = in[61] & in2[61];
    assign P[107] = in[61] ^ in2[61];
    assign G[108] = in[60] & in2[60];
    assign P[108] = in[60] ^ in2[60];
    assign G[109] = in[59] & in2[59];
    assign P[109] = in[59] ^ in2[59];
    assign G[110] = in[58] & in2[58];
    assign P[110] = in[58] ^ in2[58];
    assign G[111] = in[57] & in2[57];
    assign P[111] = in[57] ^ in2[57];
    assign G[112] = in[56] & in2[56];
    assign P[112] = in[56] ^ in2[56];
    assign G[113] = in[55] & in2[55];
    assign P[113] = in[55] ^ in2[55];
    assign G[114] = in[54] & in2[54];
    assign P[114] = in[54] ^ in2[54];
    assign G[115] = in[53] & in2[53];
    assign P[115] = in[53] ^ in2[53];
    assign G[116] = in[52] & in2[52];
    assign P[116] = in[52] ^ in2[52];
    assign G[117] = in[51] & in2[51];
    assign P[117] = in[51] ^ in2[51];
    assign G[118] = in[50] & in2[50];
    assign P[118] = in[50] ^ in2[50];
    assign G[119] = in[49] & in2[49];
    assign P[119] = in[49] ^ in2[49];
    assign G[120] = in[48] & in2[48];
    assign P[120] = in[48] ^ in2[48];
    assign G[121] = in[47] & in2[47];
    assign P[121] = in[47] ^ in2[47];
    assign G[122] = in[46] & in2[46];
    assign P[122] = in[46] ^ in2[46];
    assign G[123] = in[45] & in2[45];
    assign P[123] = in[45] ^ in2[45];
    assign G[124] = in[44] & in2[44];
    assign P[124] = in[44] ^ in2[44];
    assign G[125] = in[43] & in2[43];
    assign P[125] = in[43] ^ in2[43];
    assign G[126] = in[42] & in2[42];
    assign P[126] = in[42] ^ in2[42];
    assign G[127] = in[41] & in2[41];
    assign P[127] = in[41] ^ in2[41];
    assign G[128] = in[40] & in2[40];
    assign P[128] = in[40] ^ in2[40];
    assign G[129] = in[39] & in2[39];
    assign P[129] = in[39] ^ in2[39];
    assign G[130] = in[38] & in2[38];
    assign P[130] = in[38] ^ in2[38];
    assign G[131] = in[37] & in2[37];
    assign P[131] = in[37] ^ in2[37];
    assign G[132] = in[36] & in2[36];
    assign P[132] = in[36] ^ in2[36];
    assign G[133] = in[35] & in2[35];
    assign P[133] = in[35] ^ in2[35];
    assign G[134] = in[34] & in2[34];
    assign P[134] = in[34] ^ in2[34];
    assign G[135] = in[33] & in2[33];
    assign P[135] = in[33] ^ in2[33];
    assign G[136] = in[32] & in2[32];
    assign P[136] = in[32] ^ in2[32];
    assign G[137] = in[31] & in2[31];
    assign P[137] = in[31] ^ in2[31];
    assign G[138] = in[30] & in2[30];
    assign P[138] = in[30] ^ in2[30];
    assign G[139] = in[29] & in2[29];
    assign P[139] = in[29] ^ in2[29];
    assign G[140] = in[28] & in2[28];
    assign P[140] = in[28] ^ in2[28];
    assign G[141] = in[27] & in2[27];
    assign P[141] = in[27] ^ in2[27];
    assign G[142] = in[26] & in2[26];
    assign P[142] = in[26] ^ in2[26];
    assign G[143] = in[25] & in2[25];
    assign P[143] = in[25] ^ in2[25];
    assign G[144] = in[24] & in2[24];
    assign P[144] = in[24] ^ in2[24];
    assign G[145] = in[23] & in2[23];
    assign P[145] = in[23] ^ in2[23];
    assign G[146] = in[22] & in2[22];
    assign P[146] = in[22] ^ in2[22];
    assign G[147] = in[21] & in2[21];
    assign P[147] = in[21] ^ in2[21];
    assign G[148] = in[20] & in2[20];
    assign P[148] = in[20] ^ in2[20];
    assign G[149] = in[19] & in2[19];
    assign P[149] = in[19] ^ in2[19];
    assign G[150] = in[18] & in2[18];
    assign P[150] = in[18] ^ in2[18];
    assign G[151] = in[17] & in2[17];
    assign P[151] = in[17] ^ in2[17];
    assign G[152] = in[16] & in2[16];
    assign P[152] = in[16] ^ in2[16];
    assign G[153] = in[15] & in2[15];
    assign P[153] = in[15] ^ in2[15];
    assign G[154] = in[14] & in2[14];
    assign P[154] = in[14] ^ in2[14];
    assign G[155] = in[13] & in2[13];
    assign P[155] = in[13] ^ in2[13];
    assign G[156] = in[12] & in2[12];
    assign P[156] = in[12] ^ in2[12];
    assign G[157] = in[11] & in2[11];
    assign P[157] = in[11] ^ in2[11];
    assign G[158] = in[10] & in2[10];
    assign P[158] = in[10] ^ in2[10];
    assign G[159] = in[9] & in2[9];
    assign P[159] = in[9] ^ in2[9];
    assign G[160] = in[8] & in2[8];
    assign P[160] = in[8] ^ in2[8];
    assign G[161] = in[7] & in2[7];
    assign P[161] = in[7] ^ in2[7];
    assign G[162] = in[6] & in2[6];
    assign P[162] = in[6] ^ in2[6];
    assign G[163] = in[5] & in2[5];
    assign P[163] = in[5] ^ in2[5];
    assign G[164] = in[4] & in2[4];
    assign P[164] = in[4] ^ in2[4];
    assign G[165] = in[3] & in2[3];
    assign P[165] = in[3] ^ in2[3];
    assign G[166] = in[2] & in2[2];
    assign P[166] = in[2] ^ in2[2];
    assign G[167] = in[1] & in2[1];
    assign P[167] = in[1] ^ in2[1];
    assign G[168] = in[0] & in2[0];
    assign P[168] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign C[168] = G[167] | (P[167] & C[167]);
    assign cout = G[168] | (P[168] & C[168]);
    assign sum = P ^ C;
endmodule

module CLA168(output [167:0] sum, output cout, input [167:0] in1, input [167:0] in2;

    wire[167:0] G;
    wire[167:0] C;
    wire[167:0] P;

    assign G[0] = in[167] & in2[167];
    assign P[0] = in[167] ^ in2[167];
    assign G[1] = in[166] & in2[166];
    assign P[1] = in[166] ^ in2[166];
    assign G[2] = in[165] & in2[165];
    assign P[2] = in[165] ^ in2[165];
    assign G[3] = in[164] & in2[164];
    assign P[3] = in[164] ^ in2[164];
    assign G[4] = in[163] & in2[163];
    assign P[4] = in[163] ^ in2[163];
    assign G[5] = in[162] & in2[162];
    assign P[5] = in[162] ^ in2[162];
    assign G[6] = in[161] & in2[161];
    assign P[6] = in[161] ^ in2[161];
    assign G[7] = in[160] & in2[160];
    assign P[7] = in[160] ^ in2[160];
    assign G[8] = in[159] & in2[159];
    assign P[8] = in[159] ^ in2[159];
    assign G[9] = in[158] & in2[158];
    assign P[9] = in[158] ^ in2[158];
    assign G[10] = in[157] & in2[157];
    assign P[10] = in[157] ^ in2[157];
    assign G[11] = in[156] & in2[156];
    assign P[11] = in[156] ^ in2[156];
    assign G[12] = in[155] & in2[155];
    assign P[12] = in[155] ^ in2[155];
    assign G[13] = in[154] & in2[154];
    assign P[13] = in[154] ^ in2[154];
    assign G[14] = in[153] & in2[153];
    assign P[14] = in[153] ^ in2[153];
    assign G[15] = in[152] & in2[152];
    assign P[15] = in[152] ^ in2[152];
    assign G[16] = in[151] & in2[151];
    assign P[16] = in[151] ^ in2[151];
    assign G[17] = in[150] & in2[150];
    assign P[17] = in[150] ^ in2[150];
    assign G[18] = in[149] & in2[149];
    assign P[18] = in[149] ^ in2[149];
    assign G[19] = in[148] & in2[148];
    assign P[19] = in[148] ^ in2[148];
    assign G[20] = in[147] & in2[147];
    assign P[20] = in[147] ^ in2[147];
    assign G[21] = in[146] & in2[146];
    assign P[21] = in[146] ^ in2[146];
    assign G[22] = in[145] & in2[145];
    assign P[22] = in[145] ^ in2[145];
    assign G[23] = in[144] & in2[144];
    assign P[23] = in[144] ^ in2[144];
    assign G[24] = in[143] & in2[143];
    assign P[24] = in[143] ^ in2[143];
    assign G[25] = in[142] & in2[142];
    assign P[25] = in[142] ^ in2[142];
    assign G[26] = in[141] & in2[141];
    assign P[26] = in[141] ^ in2[141];
    assign G[27] = in[140] & in2[140];
    assign P[27] = in[140] ^ in2[140];
    assign G[28] = in[139] & in2[139];
    assign P[28] = in[139] ^ in2[139];
    assign G[29] = in[138] & in2[138];
    assign P[29] = in[138] ^ in2[138];
    assign G[30] = in[137] & in2[137];
    assign P[30] = in[137] ^ in2[137];
    assign G[31] = in[136] & in2[136];
    assign P[31] = in[136] ^ in2[136];
    assign G[32] = in[135] & in2[135];
    assign P[32] = in[135] ^ in2[135];
    assign G[33] = in[134] & in2[134];
    assign P[33] = in[134] ^ in2[134];
    assign G[34] = in[133] & in2[133];
    assign P[34] = in[133] ^ in2[133];
    assign G[35] = in[132] & in2[132];
    assign P[35] = in[132] ^ in2[132];
    assign G[36] = in[131] & in2[131];
    assign P[36] = in[131] ^ in2[131];
    assign G[37] = in[130] & in2[130];
    assign P[37] = in[130] ^ in2[130];
    assign G[38] = in[129] & in2[129];
    assign P[38] = in[129] ^ in2[129];
    assign G[39] = in[128] & in2[128];
    assign P[39] = in[128] ^ in2[128];
    assign G[40] = in[127] & in2[127];
    assign P[40] = in[127] ^ in2[127];
    assign G[41] = in[126] & in2[126];
    assign P[41] = in[126] ^ in2[126];
    assign G[42] = in[125] & in2[125];
    assign P[42] = in[125] ^ in2[125];
    assign G[43] = in[124] & in2[124];
    assign P[43] = in[124] ^ in2[124];
    assign G[44] = in[123] & in2[123];
    assign P[44] = in[123] ^ in2[123];
    assign G[45] = in[122] & in2[122];
    assign P[45] = in[122] ^ in2[122];
    assign G[46] = in[121] & in2[121];
    assign P[46] = in[121] ^ in2[121];
    assign G[47] = in[120] & in2[120];
    assign P[47] = in[120] ^ in2[120];
    assign G[48] = in[119] & in2[119];
    assign P[48] = in[119] ^ in2[119];
    assign G[49] = in[118] & in2[118];
    assign P[49] = in[118] ^ in2[118];
    assign G[50] = in[117] & in2[117];
    assign P[50] = in[117] ^ in2[117];
    assign G[51] = in[116] & in2[116];
    assign P[51] = in[116] ^ in2[116];
    assign G[52] = in[115] & in2[115];
    assign P[52] = in[115] ^ in2[115];
    assign G[53] = in[114] & in2[114];
    assign P[53] = in[114] ^ in2[114];
    assign G[54] = in[113] & in2[113];
    assign P[54] = in[113] ^ in2[113];
    assign G[55] = in[112] & in2[112];
    assign P[55] = in[112] ^ in2[112];
    assign G[56] = in[111] & in2[111];
    assign P[56] = in[111] ^ in2[111];
    assign G[57] = in[110] & in2[110];
    assign P[57] = in[110] ^ in2[110];
    assign G[58] = in[109] & in2[109];
    assign P[58] = in[109] ^ in2[109];
    assign G[59] = in[108] & in2[108];
    assign P[59] = in[108] ^ in2[108];
    assign G[60] = in[107] & in2[107];
    assign P[60] = in[107] ^ in2[107];
    assign G[61] = in[106] & in2[106];
    assign P[61] = in[106] ^ in2[106];
    assign G[62] = in[105] & in2[105];
    assign P[62] = in[105] ^ in2[105];
    assign G[63] = in[104] & in2[104];
    assign P[63] = in[104] ^ in2[104];
    assign G[64] = in[103] & in2[103];
    assign P[64] = in[103] ^ in2[103];
    assign G[65] = in[102] & in2[102];
    assign P[65] = in[102] ^ in2[102];
    assign G[66] = in[101] & in2[101];
    assign P[66] = in[101] ^ in2[101];
    assign G[67] = in[100] & in2[100];
    assign P[67] = in[100] ^ in2[100];
    assign G[68] = in[99] & in2[99];
    assign P[68] = in[99] ^ in2[99];
    assign G[69] = in[98] & in2[98];
    assign P[69] = in[98] ^ in2[98];
    assign G[70] = in[97] & in2[97];
    assign P[70] = in[97] ^ in2[97];
    assign G[71] = in[96] & in2[96];
    assign P[71] = in[96] ^ in2[96];
    assign G[72] = in[95] & in2[95];
    assign P[72] = in[95] ^ in2[95];
    assign G[73] = in[94] & in2[94];
    assign P[73] = in[94] ^ in2[94];
    assign G[74] = in[93] & in2[93];
    assign P[74] = in[93] ^ in2[93];
    assign G[75] = in[92] & in2[92];
    assign P[75] = in[92] ^ in2[92];
    assign G[76] = in[91] & in2[91];
    assign P[76] = in[91] ^ in2[91];
    assign G[77] = in[90] & in2[90];
    assign P[77] = in[90] ^ in2[90];
    assign G[78] = in[89] & in2[89];
    assign P[78] = in[89] ^ in2[89];
    assign G[79] = in[88] & in2[88];
    assign P[79] = in[88] ^ in2[88];
    assign G[80] = in[87] & in2[87];
    assign P[80] = in[87] ^ in2[87];
    assign G[81] = in[86] & in2[86];
    assign P[81] = in[86] ^ in2[86];
    assign G[82] = in[85] & in2[85];
    assign P[82] = in[85] ^ in2[85];
    assign G[83] = in[84] & in2[84];
    assign P[83] = in[84] ^ in2[84];
    assign G[84] = in[83] & in2[83];
    assign P[84] = in[83] ^ in2[83];
    assign G[85] = in[82] & in2[82];
    assign P[85] = in[82] ^ in2[82];
    assign G[86] = in[81] & in2[81];
    assign P[86] = in[81] ^ in2[81];
    assign G[87] = in[80] & in2[80];
    assign P[87] = in[80] ^ in2[80];
    assign G[88] = in[79] & in2[79];
    assign P[88] = in[79] ^ in2[79];
    assign G[89] = in[78] & in2[78];
    assign P[89] = in[78] ^ in2[78];
    assign G[90] = in[77] & in2[77];
    assign P[90] = in[77] ^ in2[77];
    assign G[91] = in[76] & in2[76];
    assign P[91] = in[76] ^ in2[76];
    assign G[92] = in[75] & in2[75];
    assign P[92] = in[75] ^ in2[75];
    assign G[93] = in[74] & in2[74];
    assign P[93] = in[74] ^ in2[74];
    assign G[94] = in[73] & in2[73];
    assign P[94] = in[73] ^ in2[73];
    assign G[95] = in[72] & in2[72];
    assign P[95] = in[72] ^ in2[72];
    assign G[96] = in[71] & in2[71];
    assign P[96] = in[71] ^ in2[71];
    assign G[97] = in[70] & in2[70];
    assign P[97] = in[70] ^ in2[70];
    assign G[98] = in[69] & in2[69];
    assign P[98] = in[69] ^ in2[69];
    assign G[99] = in[68] & in2[68];
    assign P[99] = in[68] ^ in2[68];
    assign G[100] = in[67] & in2[67];
    assign P[100] = in[67] ^ in2[67];
    assign G[101] = in[66] & in2[66];
    assign P[101] = in[66] ^ in2[66];
    assign G[102] = in[65] & in2[65];
    assign P[102] = in[65] ^ in2[65];
    assign G[103] = in[64] & in2[64];
    assign P[103] = in[64] ^ in2[64];
    assign G[104] = in[63] & in2[63];
    assign P[104] = in[63] ^ in2[63];
    assign G[105] = in[62] & in2[62];
    assign P[105] = in[62] ^ in2[62];
    assign G[106] = in[61] & in2[61];
    assign P[106] = in[61] ^ in2[61];
    assign G[107] = in[60] & in2[60];
    assign P[107] = in[60] ^ in2[60];
    assign G[108] = in[59] & in2[59];
    assign P[108] = in[59] ^ in2[59];
    assign G[109] = in[58] & in2[58];
    assign P[109] = in[58] ^ in2[58];
    assign G[110] = in[57] & in2[57];
    assign P[110] = in[57] ^ in2[57];
    assign G[111] = in[56] & in2[56];
    assign P[111] = in[56] ^ in2[56];
    assign G[112] = in[55] & in2[55];
    assign P[112] = in[55] ^ in2[55];
    assign G[113] = in[54] & in2[54];
    assign P[113] = in[54] ^ in2[54];
    assign G[114] = in[53] & in2[53];
    assign P[114] = in[53] ^ in2[53];
    assign G[115] = in[52] & in2[52];
    assign P[115] = in[52] ^ in2[52];
    assign G[116] = in[51] & in2[51];
    assign P[116] = in[51] ^ in2[51];
    assign G[117] = in[50] & in2[50];
    assign P[117] = in[50] ^ in2[50];
    assign G[118] = in[49] & in2[49];
    assign P[118] = in[49] ^ in2[49];
    assign G[119] = in[48] & in2[48];
    assign P[119] = in[48] ^ in2[48];
    assign G[120] = in[47] & in2[47];
    assign P[120] = in[47] ^ in2[47];
    assign G[121] = in[46] & in2[46];
    assign P[121] = in[46] ^ in2[46];
    assign G[122] = in[45] & in2[45];
    assign P[122] = in[45] ^ in2[45];
    assign G[123] = in[44] & in2[44];
    assign P[123] = in[44] ^ in2[44];
    assign G[124] = in[43] & in2[43];
    assign P[124] = in[43] ^ in2[43];
    assign G[125] = in[42] & in2[42];
    assign P[125] = in[42] ^ in2[42];
    assign G[126] = in[41] & in2[41];
    assign P[126] = in[41] ^ in2[41];
    assign G[127] = in[40] & in2[40];
    assign P[127] = in[40] ^ in2[40];
    assign G[128] = in[39] & in2[39];
    assign P[128] = in[39] ^ in2[39];
    assign G[129] = in[38] & in2[38];
    assign P[129] = in[38] ^ in2[38];
    assign G[130] = in[37] & in2[37];
    assign P[130] = in[37] ^ in2[37];
    assign G[131] = in[36] & in2[36];
    assign P[131] = in[36] ^ in2[36];
    assign G[132] = in[35] & in2[35];
    assign P[132] = in[35] ^ in2[35];
    assign G[133] = in[34] & in2[34];
    assign P[133] = in[34] ^ in2[34];
    assign G[134] = in[33] & in2[33];
    assign P[134] = in[33] ^ in2[33];
    assign G[135] = in[32] & in2[32];
    assign P[135] = in[32] ^ in2[32];
    assign G[136] = in[31] & in2[31];
    assign P[136] = in[31] ^ in2[31];
    assign G[137] = in[30] & in2[30];
    assign P[137] = in[30] ^ in2[30];
    assign G[138] = in[29] & in2[29];
    assign P[138] = in[29] ^ in2[29];
    assign G[139] = in[28] & in2[28];
    assign P[139] = in[28] ^ in2[28];
    assign G[140] = in[27] & in2[27];
    assign P[140] = in[27] ^ in2[27];
    assign G[141] = in[26] & in2[26];
    assign P[141] = in[26] ^ in2[26];
    assign G[142] = in[25] & in2[25];
    assign P[142] = in[25] ^ in2[25];
    assign G[143] = in[24] & in2[24];
    assign P[143] = in[24] ^ in2[24];
    assign G[144] = in[23] & in2[23];
    assign P[144] = in[23] ^ in2[23];
    assign G[145] = in[22] & in2[22];
    assign P[145] = in[22] ^ in2[22];
    assign G[146] = in[21] & in2[21];
    assign P[146] = in[21] ^ in2[21];
    assign G[147] = in[20] & in2[20];
    assign P[147] = in[20] ^ in2[20];
    assign G[148] = in[19] & in2[19];
    assign P[148] = in[19] ^ in2[19];
    assign G[149] = in[18] & in2[18];
    assign P[149] = in[18] ^ in2[18];
    assign G[150] = in[17] & in2[17];
    assign P[150] = in[17] ^ in2[17];
    assign G[151] = in[16] & in2[16];
    assign P[151] = in[16] ^ in2[16];
    assign G[152] = in[15] & in2[15];
    assign P[152] = in[15] ^ in2[15];
    assign G[153] = in[14] & in2[14];
    assign P[153] = in[14] ^ in2[14];
    assign G[154] = in[13] & in2[13];
    assign P[154] = in[13] ^ in2[13];
    assign G[155] = in[12] & in2[12];
    assign P[155] = in[12] ^ in2[12];
    assign G[156] = in[11] & in2[11];
    assign P[156] = in[11] ^ in2[11];
    assign G[157] = in[10] & in2[10];
    assign P[157] = in[10] ^ in2[10];
    assign G[158] = in[9] & in2[9];
    assign P[158] = in[9] ^ in2[9];
    assign G[159] = in[8] & in2[8];
    assign P[159] = in[8] ^ in2[8];
    assign G[160] = in[7] & in2[7];
    assign P[160] = in[7] ^ in2[7];
    assign G[161] = in[6] & in2[6];
    assign P[161] = in[6] ^ in2[6];
    assign G[162] = in[5] & in2[5];
    assign P[162] = in[5] ^ in2[5];
    assign G[163] = in[4] & in2[4];
    assign P[163] = in[4] ^ in2[4];
    assign G[164] = in[3] & in2[3];
    assign P[164] = in[3] ^ in2[3];
    assign G[165] = in[2] & in2[2];
    assign P[165] = in[2] ^ in2[2];
    assign G[166] = in[1] & in2[1];
    assign P[166] = in[1] ^ in2[1];
    assign G[167] = in[0] & in2[0];
    assign P[167] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign C[167] = G[166] | (P[166] & C[166]);
    assign cout = G[167] | (P[167] & C[167]);
    assign sum = P ^ C;
endmodule

module CLA167(output [166:0] sum, output cout, input [166:0] in1, input [166:0] in2;

    wire[166:0] G;
    wire[166:0] C;
    wire[166:0] P;

    assign G[0] = in[166] & in2[166];
    assign P[0] = in[166] ^ in2[166];
    assign G[1] = in[165] & in2[165];
    assign P[1] = in[165] ^ in2[165];
    assign G[2] = in[164] & in2[164];
    assign P[2] = in[164] ^ in2[164];
    assign G[3] = in[163] & in2[163];
    assign P[3] = in[163] ^ in2[163];
    assign G[4] = in[162] & in2[162];
    assign P[4] = in[162] ^ in2[162];
    assign G[5] = in[161] & in2[161];
    assign P[5] = in[161] ^ in2[161];
    assign G[6] = in[160] & in2[160];
    assign P[6] = in[160] ^ in2[160];
    assign G[7] = in[159] & in2[159];
    assign P[7] = in[159] ^ in2[159];
    assign G[8] = in[158] & in2[158];
    assign P[8] = in[158] ^ in2[158];
    assign G[9] = in[157] & in2[157];
    assign P[9] = in[157] ^ in2[157];
    assign G[10] = in[156] & in2[156];
    assign P[10] = in[156] ^ in2[156];
    assign G[11] = in[155] & in2[155];
    assign P[11] = in[155] ^ in2[155];
    assign G[12] = in[154] & in2[154];
    assign P[12] = in[154] ^ in2[154];
    assign G[13] = in[153] & in2[153];
    assign P[13] = in[153] ^ in2[153];
    assign G[14] = in[152] & in2[152];
    assign P[14] = in[152] ^ in2[152];
    assign G[15] = in[151] & in2[151];
    assign P[15] = in[151] ^ in2[151];
    assign G[16] = in[150] & in2[150];
    assign P[16] = in[150] ^ in2[150];
    assign G[17] = in[149] & in2[149];
    assign P[17] = in[149] ^ in2[149];
    assign G[18] = in[148] & in2[148];
    assign P[18] = in[148] ^ in2[148];
    assign G[19] = in[147] & in2[147];
    assign P[19] = in[147] ^ in2[147];
    assign G[20] = in[146] & in2[146];
    assign P[20] = in[146] ^ in2[146];
    assign G[21] = in[145] & in2[145];
    assign P[21] = in[145] ^ in2[145];
    assign G[22] = in[144] & in2[144];
    assign P[22] = in[144] ^ in2[144];
    assign G[23] = in[143] & in2[143];
    assign P[23] = in[143] ^ in2[143];
    assign G[24] = in[142] & in2[142];
    assign P[24] = in[142] ^ in2[142];
    assign G[25] = in[141] & in2[141];
    assign P[25] = in[141] ^ in2[141];
    assign G[26] = in[140] & in2[140];
    assign P[26] = in[140] ^ in2[140];
    assign G[27] = in[139] & in2[139];
    assign P[27] = in[139] ^ in2[139];
    assign G[28] = in[138] & in2[138];
    assign P[28] = in[138] ^ in2[138];
    assign G[29] = in[137] & in2[137];
    assign P[29] = in[137] ^ in2[137];
    assign G[30] = in[136] & in2[136];
    assign P[30] = in[136] ^ in2[136];
    assign G[31] = in[135] & in2[135];
    assign P[31] = in[135] ^ in2[135];
    assign G[32] = in[134] & in2[134];
    assign P[32] = in[134] ^ in2[134];
    assign G[33] = in[133] & in2[133];
    assign P[33] = in[133] ^ in2[133];
    assign G[34] = in[132] & in2[132];
    assign P[34] = in[132] ^ in2[132];
    assign G[35] = in[131] & in2[131];
    assign P[35] = in[131] ^ in2[131];
    assign G[36] = in[130] & in2[130];
    assign P[36] = in[130] ^ in2[130];
    assign G[37] = in[129] & in2[129];
    assign P[37] = in[129] ^ in2[129];
    assign G[38] = in[128] & in2[128];
    assign P[38] = in[128] ^ in2[128];
    assign G[39] = in[127] & in2[127];
    assign P[39] = in[127] ^ in2[127];
    assign G[40] = in[126] & in2[126];
    assign P[40] = in[126] ^ in2[126];
    assign G[41] = in[125] & in2[125];
    assign P[41] = in[125] ^ in2[125];
    assign G[42] = in[124] & in2[124];
    assign P[42] = in[124] ^ in2[124];
    assign G[43] = in[123] & in2[123];
    assign P[43] = in[123] ^ in2[123];
    assign G[44] = in[122] & in2[122];
    assign P[44] = in[122] ^ in2[122];
    assign G[45] = in[121] & in2[121];
    assign P[45] = in[121] ^ in2[121];
    assign G[46] = in[120] & in2[120];
    assign P[46] = in[120] ^ in2[120];
    assign G[47] = in[119] & in2[119];
    assign P[47] = in[119] ^ in2[119];
    assign G[48] = in[118] & in2[118];
    assign P[48] = in[118] ^ in2[118];
    assign G[49] = in[117] & in2[117];
    assign P[49] = in[117] ^ in2[117];
    assign G[50] = in[116] & in2[116];
    assign P[50] = in[116] ^ in2[116];
    assign G[51] = in[115] & in2[115];
    assign P[51] = in[115] ^ in2[115];
    assign G[52] = in[114] & in2[114];
    assign P[52] = in[114] ^ in2[114];
    assign G[53] = in[113] & in2[113];
    assign P[53] = in[113] ^ in2[113];
    assign G[54] = in[112] & in2[112];
    assign P[54] = in[112] ^ in2[112];
    assign G[55] = in[111] & in2[111];
    assign P[55] = in[111] ^ in2[111];
    assign G[56] = in[110] & in2[110];
    assign P[56] = in[110] ^ in2[110];
    assign G[57] = in[109] & in2[109];
    assign P[57] = in[109] ^ in2[109];
    assign G[58] = in[108] & in2[108];
    assign P[58] = in[108] ^ in2[108];
    assign G[59] = in[107] & in2[107];
    assign P[59] = in[107] ^ in2[107];
    assign G[60] = in[106] & in2[106];
    assign P[60] = in[106] ^ in2[106];
    assign G[61] = in[105] & in2[105];
    assign P[61] = in[105] ^ in2[105];
    assign G[62] = in[104] & in2[104];
    assign P[62] = in[104] ^ in2[104];
    assign G[63] = in[103] & in2[103];
    assign P[63] = in[103] ^ in2[103];
    assign G[64] = in[102] & in2[102];
    assign P[64] = in[102] ^ in2[102];
    assign G[65] = in[101] & in2[101];
    assign P[65] = in[101] ^ in2[101];
    assign G[66] = in[100] & in2[100];
    assign P[66] = in[100] ^ in2[100];
    assign G[67] = in[99] & in2[99];
    assign P[67] = in[99] ^ in2[99];
    assign G[68] = in[98] & in2[98];
    assign P[68] = in[98] ^ in2[98];
    assign G[69] = in[97] & in2[97];
    assign P[69] = in[97] ^ in2[97];
    assign G[70] = in[96] & in2[96];
    assign P[70] = in[96] ^ in2[96];
    assign G[71] = in[95] & in2[95];
    assign P[71] = in[95] ^ in2[95];
    assign G[72] = in[94] & in2[94];
    assign P[72] = in[94] ^ in2[94];
    assign G[73] = in[93] & in2[93];
    assign P[73] = in[93] ^ in2[93];
    assign G[74] = in[92] & in2[92];
    assign P[74] = in[92] ^ in2[92];
    assign G[75] = in[91] & in2[91];
    assign P[75] = in[91] ^ in2[91];
    assign G[76] = in[90] & in2[90];
    assign P[76] = in[90] ^ in2[90];
    assign G[77] = in[89] & in2[89];
    assign P[77] = in[89] ^ in2[89];
    assign G[78] = in[88] & in2[88];
    assign P[78] = in[88] ^ in2[88];
    assign G[79] = in[87] & in2[87];
    assign P[79] = in[87] ^ in2[87];
    assign G[80] = in[86] & in2[86];
    assign P[80] = in[86] ^ in2[86];
    assign G[81] = in[85] & in2[85];
    assign P[81] = in[85] ^ in2[85];
    assign G[82] = in[84] & in2[84];
    assign P[82] = in[84] ^ in2[84];
    assign G[83] = in[83] & in2[83];
    assign P[83] = in[83] ^ in2[83];
    assign G[84] = in[82] & in2[82];
    assign P[84] = in[82] ^ in2[82];
    assign G[85] = in[81] & in2[81];
    assign P[85] = in[81] ^ in2[81];
    assign G[86] = in[80] & in2[80];
    assign P[86] = in[80] ^ in2[80];
    assign G[87] = in[79] & in2[79];
    assign P[87] = in[79] ^ in2[79];
    assign G[88] = in[78] & in2[78];
    assign P[88] = in[78] ^ in2[78];
    assign G[89] = in[77] & in2[77];
    assign P[89] = in[77] ^ in2[77];
    assign G[90] = in[76] & in2[76];
    assign P[90] = in[76] ^ in2[76];
    assign G[91] = in[75] & in2[75];
    assign P[91] = in[75] ^ in2[75];
    assign G[92] = in[74] & in2[74];
    assign P[92] = in[74] ^ in2[74];
    assign G[93] = in[73] & in2[73];
    assign P[93] = in[73] ^ in2[73];
    assign G[94] = in[72] & in2[72];
    assign P[94] = in[72] ^ in2[72];
    assign G[95] = in[71] & in2[71];
    assign P[95] = in[71] ^ in2[71];
    assign G[96] = in[70] & in2[70];
    assign P[96] = in[70] ^ in2[70];
    assign G[97] = in[69] & in2[69];
    assign P[97] = in[69] ^ in2[69];
    assign G[98] = in[68] & in2[68];
    assign P[98] = in[68] ^ in2[68];
    assign G[99] = in[67] & in2[67];
    assign P[99] = in[67] ^ in2[67];
    assign G[100] = in[66] & in2[66];
    assign P[100] = in[66] ^ in2[66];
    assign G[101] = in[65] & in2[65];
    assign P[101] = in[65] ^ in2[65];
    assign G[102] = in[64] & in2[64];
    assign P[102] = in[64] ^ in2[64];
    assign G[103] = in[63] & in2[63];
    assign P[103] = in[63] ^ in2[63];
    assign G[104] = in[62] & in2[62];
    assign P[104] = in[62] ^ in2[62];
    assign G[105] = in[61] & in2[61];
    assign P[105] = in[61] ^ in2[61];
    assign G[106] = in[60] & in2[60];
    assign P[106] = in[60] ^ in2[60];
    assign G[107] = in[59] & in2[59];
    assign P[107] = in[59] ^ in2[59];
    assign G[108] = in[58] & in2[58];
    assign P[108] = in[58] ^ in2[58];
    assign G[109] = in[57] & in2[57];
    assign P[109] = in[57] ^ in2[57];
    assign G[110] = in[56] & in2[56];
    assign P[110] = in[56] ^ in2[56];
    assign G[111] = in[55] & in2[55];
    assign P[111] = in[55] ^ in2[55];
    assign G[112] = in[54] & in2[54];
    assign P[112] = in[54] ^ in2[54];
    assign G[113] = in[53] & in2[53];
    assign P[113] = in[53] ^ in2[53];
    assign G[114] = in[52] & in2[52];
    assign P[114] = in[52] ^ in2[52];
    assign G[115] = in[51] & in2[51];
    assign P[115] = in[51] ^ in2[51];
    assign G[116] = in[50] & in2[50];
    assign P[116] = in[50] ^ in2[50];
    assign G[117] = in[49] & in2[49];
    assign P[117] = in[49] ^ in2[49];
    assign G[118] = in[48] & in2[48];
    assign P[118] = in[48] ^ in2[48];
    assign G[119] = in[47] & in2[47];
    assign P[119] = in[47] ^ in2[47];
    assign G[120] = in[46] & in2[46];
    assign P[120] = in[46] ^ in2[46];
    assign G[121] = in[45] & in2[45];
    assign P[121] = in[45] ^ in2[45];
    assign G[122] = in[44] & in2[44];
    assign P[122] = in[44] ^ in2[44];
    assign G[123] = in[43] & in2[43];
    assign P[123] = in[43] ^ in2[43];
    assign G[124] = in[42] & in2[42];
    assign P[124] = in[42] ^ in2[42];
    assign G[125] = in[41] & in2[41];
    assign P[125] = in[41] ^ in2[41];
    assign G[126] = in[40] & in2[40];
    assign P[126] = in[40] ^ in2[40];
    assign G[127] = in[39] & in2[39];
    assign P[127] = in[39] ^ in2[39];
    assign G[128] = in[38] & in2[38];
    assign P[128] = in[38] ^ in2[38];
    assign G[129] = in[37] & in2[37];
    assign P[129] = in[37] ^ in2[37];
    assign G[130] = in[36] & in2[36];
    assign P[130] = in[36] ^ in2[36];
    assign G[131] = in[35] & in2[35];
    assign P[131] = in[35] ^ in2[35];
    assign G[132] = in[34] & in2[34];
    assign P[132] = in[34] ^ in2[34];
    assign G[133] = in[33] & in2[33];
    assign P[133] = in[33] ^ in2[33];
    assign G[134] = in[32] & in2[32];
    assign P[134] = in[32] ^ in2[32];
    assign G[135] = in[31] & in2[31];
    assign P[135] = in[31] ^ in2[31];
    assign G[136] = in[30] & in2[30];
    assign P[136] = in[30] ^ in2[30];
    assign G[137] = in[29] & in2[29];
    assign P[137] = in[29] ^ in2[29];
    assign G[138] = in[28] & in2[28];
    assign P[138] = in[28] ^ in2[28];
    assign G[139] = in[27] & in2[27];
    assign P[139] = in[27] ^ in2[27];
    assign G[140] = in[26] & in2[26];
    assign P[140] = in[26] ^ in2[26];
    assign G[141] = in[25] & in2[25];
    assign P[141] = in[25] ^ in2[25];
    assign G[142] = in[24] & in2[24];
    assign P[142] = in[24] ^ in2[24];
    assign G[143] = in[23] & in2[23];
    assign P[143] = in[23] ^ in2[23];
    assign G[144] = in[22] & in2[22];
    assign P[144] = in[22] ^ in2[22];
    assign G[145] = in[21] & in2[21];
    assign P[145] = in[21] ^ in2[21];
    assign G[146] = in[20] & in2[20];
    assign P[146] = in[20] ^ in2[20];
    assign G[147] = in[19] & in2[19];
    assign P[147] = in[19] ^ in2[19];
    assign G[148] = in[18] & in2[18];
    assign P[148] = in[18] ^ in2[18];
    assign G[149] = in[17] & in2[17];
    assign P[149] = in[17] ^ in2[17];
    assign G[150] = in[16] & in2[16];
    assign P[150] = in[16] ^ in2[16];
    assign G[151] = in[15] & in2[15];
    assign P[151] = in[15] ^ in2[15];
    assign G[152] = in[14] & in2[14];
    assign P[152] = in[14] ^ in2[14];
    assign G[153] = in[13] & in2[13];
    assign P[153] = in[13] ^ in2[13];
    assign G[154] = in[12] & in2[12];
    assign P[154] = in[12] ^ in2[12];
    assign G[155] = in[11] & in2[11];
    assign P[155] = in[11] ^ in2[11];
    assign G[156] = in[10] & in2[10];
    assign P[156] = in[10] ^ in2[10];
    assign G[157] = in[9] & in2[9];
    assign P[157] = in[9] ^ in2[9];
    assign G[158] = in[8] & in2[8];
    assign P[158] = in[8] ^ in2[8];
    assign G[159] = in[7] & in2[7];
    assign P[159] = in[7] ^ in2[7];
    assign G[160] = in[6] & in2[6];
    assign P[160] = in[6] ^ in2[6];
    assign G[161] = in[5] & in2[5];
    assign P[161] = in[5] ^ in2[5];
    assign G[162] = in[4] & in2[4];
    assign P[162] = in[4] ^ in2[4];
    assign G[163] = in[3] & in2[3];
    assign P[163] = in[3] ^ in2[3];
    assign G[164] = in[2] & in2[2];
    assign P[164] = in[2] ^ in2[2];
    assign G[165] = in[1] & in2[1];
    assign P[165] = in[1] ^ in2[1];
    assign G[166] = in[0] & in2[0];
    assign P[166] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign C[166] = G[165] | (P[165] & C[165]);
    assign cout = G[166] | (P[166] & C[166]);
    assign sum = P ^ C;
endmodule

module CLA166(output [165:0] sum, output cout, input [165:0] in1, input [165:0] in2;

    wire[165:0] G;
    wire[165:0] C;
    wire[165:0] P;

    assign G[0] = in[165] & in2[165];
    assign P[0] = in[165] ^ in2[165];
    assign G[1] = in[164] & in2[164];
    assign P[1] = in[164] ^ in2[164];
    assign G[2] = in[163] & in2[163];
    assign P[2] = in[163] ^ in2[163];
    assign G[3] = in[162] & in2[162];
    assign P[3] = in[162] ^ in2[162];
    assign G[4] = in[161] & in2[161];
    assign P[4] = in[161] ^ in2[161];
    assign G[5] = in[160] & in2[160];
    assign P[5] = in[160] ^ in2[160];
    assign G[6] = in[159] & in2[159];
    assign P[6] = in[159] ^ in2[159];
    assign G[7] = in[158] & in2[158];
    assign P[7] = in[158] ^ in2[158];
    assign G[8] = in[157] & in2[157];
    assign P[8] = in[157] ^ in2[157];
    assign G[9] = in[156] & in2[156];
    assign P[9] = in[156] ^ in2[156];
    assign G[10] = in[155] & in2[155];
    assign P[10] = in[155] ^ in2[155];
    assign G[11] = in[154] & in2[154];
    assign P[11] = in[154] ^ in2[154];
    assign G[12] = in[153] & in2[153];
    assign P[12] = in[153] ^ in2[153];
    assign G[13] = in[152] & in2[152];
    assign P[13] = in[152] ^ in2[152];
    assign G[14] = in[151] & in2[151];
    assign P[14] = in[151] ^ in2[151];
    assign G[15] = in[150] & in2[150];
    assign P[15] = in[150] ^ in2[150];
    assign G[16] = in[149] & in2[149];
    assign P[16] = in[149] ^ in2[149];
    assign G[17] = in[148] & in2[148];
    assign P[17] = in[148] ^ in2[148];
    assign G[18] = in[147] & in2[147];
    assign P[18] = in[147] ^ in2[147];
    assign G[19] = in[146] & in2[146];
    assign P[19] = in[146] ^ in2[146];
    assign G[20] = in[145] & in2[145];
    assign P[20] = in[145] ^ in2[145];
    assign G[21] = in[144] & in2[144];
    assign P[21] = in[144] ^ in2[144];
    assign G[22] = in[143] & in2[143];
    assign P[22] = in[143] ^ in2[143];
    assign G[23] = in[142] & in2[142];
    assign P[23] = in[142] ^ in2[142];
    assign G[24] = in[141] & in2[141];
    assign P[24] = in[141] ^ in2[141];
    assign G[25] = in[140] & in2[140];
    assign P[25] = in[140] ^ in2[140];
    assign G[26] = in[139] & in2[139];
    assign P[26] = in[139] ^ in2[139];
    assign G[27] = in[138] & in2[138];
    assign P[27] = in[138] ^ in2[138];
    assign G[28] = in[137] & in2[137];
    assign P[28] = in[137] ^ in2[137];
    assign G[29] = in[136] & in2[136];
    assign P[29] = in[136] ^ in2[136];
    assign G[30] = in[135] & in2[135];
    assign P[30] = in[135] ^ in2[135];
    assign G[31] = in[134] & in2[134];
    assign P[31] = in[134] ^ in2[134];
    assign G[32] = in[133] & in2[133];
    assign P[32] = in[133] ^ in2[133];
    assign G[33] = in[132] & in2[132];
    assign P[33] = in[132] ^ in2[132];
    assign G[34] = in[131] & in2[131];
    assign P[34] = in[131] ^ in2[131];
    assign G[35] = in[130] & in2[130];
    assign P[35] = in[130] ^ in2[130];
    assign G[36] = in[129] & in2[129];
    assign P[36] = in[129] ^ in2[129];
    assign G[37] = in[128] & in2[128];
    assign P[37] = in[128] ^ in2[128];
    assign G[38] = in[127] & in2[127];
    assign P[38] = in[127] ^ in2[127];
    assign G[39] = in[126] & in2[126];
    assign P[39] = in[126] ^ in2[126];
    assign G[40] = in[125] & in2[125];
    assign P[40] = in[125] ^ in2[125];
    assign G[41] = in[124] & in2[124];
    assign P[41] = in[124] ^ in2[124];
    assign G[42] = in[123] & in2[123];
    assign P[42] = in[123] ^ in2[123];
    assign G[43] = in[122] & in2[122];
    assign P[43] = in[122] ^ in2[122];
    assign G[44] = in[121] & in2[121];
    assign P[44] = in[121] ^ in2[121];
    assign G[45] = in[120] & in2[120];
    assign P[45] = in[120] ^ in2[120];
    assign G[46] = in[119] & in2[119];
    assign P[46] = in[119] ^ in2[119];
    assign G[47] = in[118] & in2[118];
    assign P[47] = in[118] ^ in2[118];
    assign G[48] = in[117] & in2[117];
    assign P[48] = in[117] ^ in2[117];
    assign G[49] = in[116] & in2[116];
    assign P[49] = in[116] ^ in2[116];
    assign G[50] = in[115] & in2[115];
    assign P[50] = in[115] ^ in2[115];
    assign G[51] = in[114] & in2[114];
    assign P[51] = in[114] ^ in2[114];
    assign G[52] = in[113] & in2[113];
    assign P[52] = in[113] ^ in2[113];
    assign G[53] = in[112] & in2[112];
    assign P[53] = in[112] ^ in2[112];
    assign G[54] = in[111] & in2[111];
    assign P[54] = in[111] ^ in2[111];
    assign G[55] = in[110] & in2[110];
    assign P[55] = in[110] ^ in2[110];
    assign G[56] = in[109] & in2[109];
    assign P[56] = in[109] ^ in2[109];
    assign G[57] = in[108] & in2[108];
    assign P[57] = in[108] ^ in2[108];
    assign G[58] = in[107] & in2[107];
    assign P[58] = in[107] ^ in2[107];
    assign G[59] = in[106] & in2[106];
    assign P[59] = in[106] ^ in2[106];
    assign G[60] = in[105] & in2[105];
    assign P[60] = in[105] ^ in2[105];
    assign G[61] = in[104] & in2[104];
    assign P[61] = in[104] ^ in2[104];
    assign G[62] = in[103] & in2[103];
    assign P[62] = in[103] ^ in2[103];
    assign G[63] = in[102] & in2[102];
    assign P[63] = in[102] ^ in2[102];
    assign G[64] = in[101] & in2[101];
    assign P[64] = in[101] ^ in2[101];
    assign G[65] = in[100] & in2[100];
    assign P[65] = in[100] ^ in2[100];
    assign G[66] = in[99] & in2[99];
    assign P[66] = in[99] ^ in2[99];
    assign G[67] = in[98] & in2[98];
    assign P[67] = in[98] ^ in2[98];
    assign G[68] = in[97] & in2[97];
    assign P[68] = in[97] ^ in2[97];
    assign G[69] = in[96] & in2[96];
    assign P[69] = in[96] ^ in2[96];
    assign G[70] = in[95] & in2[95];
    assign P[70] = in[95] ^ in2[95];
    assign G[71] = in[94] & in2[94];
    assign P[71] = in[94] ^ in2[94];
    assign G[72] = in[93] & in2[93];
    assign P[72] = in[93] ^ in2[93];
    assign G[73] = in[92] & in2[92];
    assign P[73] = in[92] ^ in2[92];
    assign G[74] = in[91] & in2[91];
    assign P[74] = in[91] ^ in2[91];
    assign G[75] = in[90] & in2[90];
    assign P[75] = in[90] ^ in2[90];
    assign G[76] = in[89] & in2[89];
    assign P[76] = in[89] ^ in2[89];
    assign G[77] = in[88] & in2[88];
    assign P[77] = in[88] ^ in2[88];
    assign G[78] = in[87] & in2[87];
    assign P[78] = in[87] ^ in2[87];
    assign G[79] = in[86] & in2[86];
    assign P[79] = in[86] ^ in2[86];
    assign G[80] = in[85] & in2[85];
    assign P[80] = in[85] ^ in2[85];
    assign G[81] = in[84] & in2[84];
    assign P[81] = in[84] ^ in2[84];
    assign G[82] = in[83] & in2[83];
    assign P[82] = in[83] ^ in2[83];
    assign G[83] = in[82] & in2[82];
    assign P[83] = in[82] ^ in2[82];
    assign G[84] = in[81] & in2[81];
    assign P[84] = in[81] ^ in2[81];
    assign G[85] = in[80] & in2[80];
    assign P[85] = in[80] ^ in2[80];
    assign G[86] = in[79] & in2[79];
    assign P[86] = in[79] ^ in2[79];
    assign G[87] = in[78] & in2[78];
    assign P[87] = in[78] ^ in2[78];
    assign G[88] = in[77] & in2[77];
    assign P[88] = in[77] ^ in2[77];
    assign G[89] = in[76] & in2[76];
    assign P[89] = in[76] ^ in2[76];
    assign G[90] = in[75] & in2[75];
    assign P[90] = in[75] ^ in2[75];
    assign G[91] = in[74] & in2[74];
    assign P[91] = in[74] ^ in2[74];
    assign G[92] = in[73] & in2[73];
    assign P[92] = in[73] ^ in2[73];
    assign G[93] = in[72] & in2[72];
    assign P[93] = in[72] ^ in2[72];
    assign G[94] = in[71] & in2[71];
    assign P[94] = in[71] ^ in2[71];
    assign G[95] = in[70] & in2[70];
    assign P[95] = in[70] ^ in2[70];
    assign G[96] = in[69] & in2[69];
    assign P[96] = in[69] ^ in2[69];
    assign G[97] = in[68] & in2[68];
    assign P[97] = in[68] ^ in2[68];
    assign G[98] = in[67] & in2[67];
    assign P[98] = in[67] ^ in2[67];
    assign G[99] = in[66] & in2[66];
    assign P[99] = in[66] ^ in2[66];
    assign G[100] = in[65] & in2[65];
    assign P[100] = in[65] ^ in2[65];
    assign G[101] = in[64] & in2[64];
    assign P[101] = in[64] ^ in2[64];
    assign G[102] = in[63] & in2[63];
    assign P[102] = in[63] ^ in2[63];
    assign G[103] = in[62] & in2[62];
    assign P[103] = in[62] ^ in2[62];
    assign G[104] = in[61] & in2[61];
    assign P[104] = in[61] ^ in2[61];
    assign G[105] = in[60] & in2[60];
    assign P[105] = in[60] ^ in2[60];
    assign G[106] = in[59] & in2[59];
    assign P[106] = in[59] ^ in2[59];
    assign G[107] = in[58] & in2[58];
    assign P[107] = in[58] ^ in2[58];
    assign G[108] = in[57] & in2[57];
    assign P[108] = in[57] ^ in2[57];
    assign G[109] = in[56] & in2[56];
    assign P[109] = in[56] ^ in2[56];
    assign G[110] = in[55] & in2[55];
    assign P[110] = in[55] ^ in2[55];
    assign G[111] = in[54] & in2[54];
    assign P[111] = in[54] ^ in2[54];
    assign G[112] = in[53] & in2[53];
    assign P[112] = in[53] ^ in2[53];
    assign G[113] = in[52] & in2[52];
    assign P[113] = in[52] ^ in2[52];
    assign G[114] = in[51] & in2[51];
    assign P[114] = in[51] ^ in2[51];
    assign G[115] = in[50] & in2[50];
    assign P[115] = in[50] ^ in2[50];
    assign G[116] = in[49] & in2[49];
    assign P[116] = in[49] ^ in2[49];
    assign G[117] = in[48] & in2[48];
    assign P[117] = in[48] ^ in2[48];
    assign G[118] = in[47] & in2[47];
    assign P[118] = in[47] ^ in2[47];
    assign G[119] = in[46] & in2[46];
    assign P[119] = in[46] ^ in2[46];
    assign G[120] = in[45] & in2[45];
    assign P[120] = in[45] ^ in2[45];
    assign G[121] = in[44] & in2[44];
    assign P[121] = in[44] ^ in2[44];
    assign G[122] = in[43] & in2[43];
    assign P[122] = in[43] ^ in2[43];
    assign G[123] = in[42] & in2[42];
    assign P[123] = in[42] ^ in2[42];
    assign G[124] = in[41] & in2[41];
    assign P[124] = in[41] ^ in2[41];
    assign G[125] = in[40] & in2[40];
    assign P[125] = in[40] ^ in2[40];
    assign G[126] = in[39] & in2[39];
    assign P[126] = in[39] ^ in2[39];
    assign G[127] = in[38] & in2[38];
    assign P[127] = in[38] ^ in2[38];
    assign G[128] = in[37] & in2[37];
    assign P[128] = in[37] ^ in2[37];
    assign G[129] = in[36] & in2[36];
    assign P[129] = in[36] ^ in2[36];
    assign G[130] = in[35] & in2[35];
    assign P[130] = in[35] ^ in2[35];
    assign G[131] = in[34] & in2[34];
    assign P[131] = in[34] ^ in2[34];
    assign G[132] = in[33] & in2[33];
    assign P[132] = in[33] ^ in2[33];
    assign G[133] = in[32] & in2[32];
    assign P[133] = in[32] ^ in2[32];
    assign G[134] = in[31] & in2[31];
    assign P[134] = in[31] ^ in2[31];
    assign G[135] = in[30] & in2[30];
    assign P[135] = in[30] ^ in2[30];
    assign G[136] = in[29] & in2[29];
    assign P[136] = in[29] ^ in2[29];
    assign G[137] = in[28] & in2[28];
    assign P[137] = in[28] ^ in2[28];
    assign G[138] = in[27] & in2[27];
    assign P[138] = in[27] ^ in2[27];
    assign G[139] = in[26] & in2[26];
    assign P[139] = in[26] ^ in2[26];
    assign G[140] = in[25] & in2[25];
    assign P[140] = in[25] ^ in2[25];
    assign G[141] = in[24] & in2[24];
    assign P[141] = in[24] ^ in2[24];
    assign G[142] = in[23] & in2[23];
    assign P[142] = in[23] ^ in2[23];
    assign G[143] = in[22] & in2[22];
    assign P[143] = in[22] ^ in2[22];
    assign G[144] = in[21] & in2[21];
    assign P[144] = in[21] ^ in2[21];
    assign G[145] = in[20] & in2[20];
    assign P[145] = in[20] ^ in2[20];
    assign G[146] = in[19] & in2[19];
    assign P[146] = in[19] ^ in2[19];
    assign G[147] = in[18] & in2[18];
    assign P[147] = in[18] ^ in2[18];
    assign G[148] = in[17] & in2[17];
    assign P[148] = in[17] ^ in2[17];
    assign G[149] = in[16] & in2[16];
    assign P[149] = in[16] ^ in2[16];
    assign G[150] = in[15] & in2[15];
    assign P[150] = in[15] ^ in2[15];
    assign G[151] = in[14] & in2[14];
    assign P[151] = in[14] ^ in2[14];
    assign G[152] = in[13] & in2[13];
    assign P[152] = in[13] ^ in2[13];
    assign G[153] = in[12] & in2[12];
    assign P[153] = in[12] ^ in2[12];
    assign G[154] = in[11] & in2[11];
    assign P[154] = in[11] ^ in2[11];
    assign G[155] = in[10] & in2[10];
    assign P[155] = in[10] ^ in2[10];
    assign G[156] = in[9] & in2[9];
    assign P[156] = in[9] ^ in2[9];
    assign G[157] = in[8] & in2[8];
    assign P[157] = in[8] ^ in2[8];
    assign G[158] = in[7] & in2[7];
    assign P[158] = in[7] ^ in2[7];
    assign G[159] = in[6] & in2[6];
    assign P[159] = in[6] ^ in2[6];
    assign G[160] = in[5] & in2[5];
    assign P[160] = in[5] ^ in2[5];
    assign G[161] = in[4] & in2[4];
    assign P[161] = in[4] ^ in2[4];
    assign G[162] = in[3] & in2[3];
    assign P[162] = in[3] ^ in2[3];
    assign G[163] = in[2] & in2[2];
    assign P[163] = in[2] ^ in2[2];
    assign G[164] = in[1] & in2[1];
    assign P[164] = in[1] ^ in2[1];
    assign G[165] = in[0] & in2[0];
    assign P[165] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign C[165] = G[164] | (P[164] & C[164]);
    assign cout = G[165] | (P[165] & C[165]);
    assign sum = P ^ C;
endmodule

module CLA165(output [164:0] sum, output cout, input [164:0] in1, input [164:0] in2;

    wire[164:0] G;
    wire[164:0] C;
    wire[164:0] P;

    assign G[0] = in[164] & in2[164];
    assign P[0] = in[164] ^ in2[164];
    assign G[1] = in[163] & in2[163];
    assign P[1] = in[163] ^ in2[163];
    assign G[2] = in[162] & in2[162];
    assign P[2] = in[162] ^ in2[162];
    assign G[3] = in[161] & in2[161];
    assign P[3] = in[161] ^ in2[161];
    assign G[4] = in[160] & in2[160];
    assign P[4] = in[160] ^ in2[160];
    assign G[5] = in[159] & in2[159];
    assign P[5] = in[159] ^ in2[159];
    assign G[6] = in[158] & in2[158];
    assign P[6] = in[158] ^ in2[158];
    assign G[7] = in[157] & in2[157];
    assign P[7] = in[157] ^ in2[157];
    assign G[8] = in[156] & in2[156];
    assign P[8] = in[156] ^ in2[156];
    assign G[9] = in[155] & in2[155];
    assign P[9] = in[155] ^ in2[155];
    assign G[10] = in[154] & in2[154];
    assign P[10] = in[154] ^ in2[154];
    assign G[11] = in[153] & in2[153];
    assign P[11] = in[153] ^ in2[153];
    assign G[12] = in[152] & in2[152];
    assign P[12] = in[152] ^ in2[152];
    assign G[13] = in[151] & in2[151];
    assign P[13] = in[151] ^ in2[151];
    assign G[14] = in[150] & in2[150];
    assign P[14] = in[150] ^ in2[150];
    assign G[15] = in[149] & in2[149];
    assign P[15] = in[149] ^ in2[149];
    assign G[16] = in[148] & in2[148];
    assign P[16] = in[148] ^ in2[148];
    assign G[17] = in[147] & in2[147];
    assign P[17] = in[147] ^ in2[147];
    assign G[18] = in[146] & in2[146];
    assign P[18] = in[146] ^ in2[146];
    assign G[19] = in[145] & in2[145];
    assign P[19] = in[145] ^ in2[145];
    assign G[20] = in[144] & in2[144];
    assign P[20] = in[144] ^ in2[144];
    assign G[21] = in[143] & in2[143];
    assign P[21] = in[143] ^ in2[143];
    assign G[22] = in[142] & in2[142];
    assign P[22] = in[142] ^ in2[142];
    assign G[23] = in[141] & in2[141];
    assign P[23] = in[141] ^ in2[141];
    assign G[24] = in[140] & in2[140];
    assign P[24] = in[140] ^ in2[140];
    assign G[25] = in[139] & in2[139];
    assign P[25] = in[139] ^ in2[139];
    assign G[26] = in[138] & in2[138];
    assign P[26] = in[138] ^ in2[138];
    assign G[27] = in[137] & in2[137];
    assign P[27] = in[137] ^ in2[137];
    assign G[28] = in[136] & in2[136];
    assign P[28] = in[136] ^ in2[136];
    assign G[29] = in[135] & in2[135];
    assign P[29] = in[135] ^ in2[135];
    assign G[30] = in[134] & in2[134];
    assign P[30] = in[134] ^ in2[134];
    assign G[31] = in[133] & in2[133];
    assign P[31] = in[133] ^ in2[133];
    assign G[32] = in[132] & in2[132];
    assign P[32] = in[132] ^ in2[132];
    assign G[33] = in[131] & in2[131];
    assign P[33] = in[131] ^ in2[131];
    assign G[34] = in[130] & in2[130];
    assign P[34] = in[130] ^ in2[130];
    assign G[35] = in[129] & in2[129];
    assign P[35] = in[129] ^ in2[129];
    assign G[36] = in[128] & in2[128];
    assign P[36] = in[128] ^ in2[128];
    assign G[37] = in[127] & in2[127];
    assign P[37] = in[127] ^ in2[127];
    assign G[38] = in[126] & in2[126];
    assign P[38] = in[126] ^ in2[126];
    assign G[39] = in[125] & in2[125];
    assign P[39] = in[125] ^ in2[125];
    assign G[40] = in[124] & in2[124];
    assign P[40] = in[124] ^ in2[124];
    assign G[41] = in[123] & in2[123];
    assign P[41] = in[123] ^ in2[123];
    assign G[42] = in[122] & in2[122];
    assign P[42] = in[122] ^ in2[122];
    assign G[43] = in[121] & in2[121];
    assign P[43] = in[121] ^ in2[121];
    assign G[44] = in[120] & in2[120];
    assign P[44] = in[120] ^ in2[120];
    assign G[45] = in[119] & in2[119];
    assign P[45] = in[119] ^ in2[119];
    assign G[46] = in[118] & in2[118];
    assign P[46] = in[118] ^ in2[118];
    assign G[47] = in[117] & in2[117];
    assign P[47] = in[117] ^ in2[117];
    assign G[48] = in[116] & in2[116];
    assign P[48] = in[116] ^ in2[116];
    assign G[49] = in[115] & in2[115];
    assign P[49] = in[115] ^ in2[115];
    assign G[50] = in[114] & in2[114];
    assign P[50] = in[114] ^ in2[114];
    assign G[51] = in[113] & in2[113];
    assign P[51] = in[113] ^ in2[113];
    assign G[52] = in[112] & in2[112];
    assign P[52] = in[112] ^ in2[112];
    assign G[53] = in[111] & in2[111];
    assign P[53] = in[111] ^ in2[111];
    assign G[54] = in[110] & in2[110];
    assign P[54] = in[110] ^ in2[110];
    assign G[55] = in[109] & in2[109];
    assign P[55] = in[109] ^ in2[109];
    assign G[56] = in[108] & in2[108];
    assign P[56] = in[108] ^ in2[108];
    assign G[57] = in[107] & in2[107];
    assign P[57] = in[107] ^ in2[107];
    assign G[58] = in[106] & in2[106];
    assign P[58] = in[106] ^ in2[106];
    assign G[59] = in[105] & in2[105];
    assign P[59] = in[105] ^ in2[105];
    assign G[60] = in[104] & in2[104];
    assign P[60] = in[104] ^ in2[104];
    assign G[61] = in[103] & in2[103];
    assign P[61] = in[103] ^ in2[103];
    assign G[62] = in[102] & in2[102];
    assign P[62] = in[102] ^ in2[102];
    assign G[63] = in[101] & in2[101];
    assign P[63] = in[101] ^ in2[101];
    assign G[64] = in[100] & in2[100];
    assign P[64] = in[100] ^ in2[100];
    assign G[65] = in[99] & in2[99];
    assign P[65] = in[99] ^ in2[99];
    assign G[66] = in[98] & in2[98];
    assign P[66] = in[98] ^ in2[98];
    assign G[67] = in[97] & in2[97];
    assign P[67] = in[97] ^ in2[97];
    assign G[68] = in[96] & in2[96];
    assign P[68] = in[96] ^ in2[96];
    assign G[69] = in[95] & in2[95];
    assign P[69] = in[95] ^ in2[95];
    assign G[70] = in[94] & in2[94];
    assign P[70] = in[94] ^ in2[94];
    assign G[71] = in[93] & in2[93];
    assign P[71] = in[93] ^ in2[93];
    assign G[72] = in[92] & in2[92];
    assign P[72] = in[92] ^ in2[92];
    assign G[73] = in[91] & in2[91];
    assign P[73] = in[91] ^ in2[91];
    assign G[74] = in[90] & in2[90];
    assign P[74] = in[90] ^ in2[90];
    assign G[75] = in[89] & in2[89];
    assign P[75] = in[89] ^ in2[89];
    assign G[76] = in[88] & in2[88];
    assign P[76] = in[88] ^ in2[88];
    assign G[77] = in[87] & in2[87];
    assign P[77] = in[87] ^ in2[87];
    assign G[78] = in[86] & in2[86];
    assign P[78] = in[86] ^ in2[86];
    assign G[79] = in[85] & in2[85];
    assign P[79] = in[85] ^ in2[85];
    assign G[80] = in[84] & in2[84];
    assign P[80] = in[84] ^ in2[84];
    assign G[81] = in[83] & in2[83];
    assign P[81] = in[83] ^ in2[83];
    assign G[82] = in[82] & in2[82];
    assign P[82] = in[82] ^ in2[82];
    assign G[83] = in[81] & in2[81];
    assign P[83] = in[81] ^ in2[81];
    assign G[84] = in[80] & in2[80];
    assign P[84] = in[80] ^ in2[80];
    assign G[85] = in[79] & in2[79];
    assign P[85] = in[79] ^ in2[79];
    assign G[86] = in[78] & in2[78];
    assign P[86] = in[78] ^ in2[78];
    assign G[87] = in[77] & in2[77];
    assign P[87] = in[77] ^ in2[77];
    assign G[88] = in[76] & in2[76];
    assign P[88] = in[76] ^ in2[76];
    assign G[89] = in[75] & in2[75];
    assign P[89] = in[75] ^ in2[75];
    assign G[90] = in[74] & in2[74];
    assign P[90] = in[74] ^ in2[74];
    assign G[91] = in[73] & in2[73];
    assign P[91] = in[73] ^ in2[73];
    assign G[92] = in[72] & in2[72];
    assign P[92] = in[72] ^ in2[72];
    assign G[93] = in[71] & in2[71];
    assign P[93] = in[71] ^ in2[71];
    assign G[94] = in[70] & in2[70];
    assign P[94] = in[70] ^ in2[70];
    assign G[95] = in[69] & in2[69];
    assign P[95] = in[69] ^ in2[69];
    assign G[96] = in[68] & in2[68];
    assign P[96] = in[68] ^ in2[68];
    assign G[97] = in[67] & in2[67];
    assign P[97] = in[67] ^ in2[67];
    assign G[98] = in[66] & in2[66];
    assign P[98] = in[66] ^ in2[66];
    assign G[99] = in[65] & in2[65];
    assign P[99] = in[65] ^ in2[65];
    assign G[100] = in[64] & in2[64];
    assign P[100] = in[64] ^ in2[64];
    assign G[101] = in[63] & in2[63];
    assign P[101] = in[63] ^ in2[63];
    assign G[102] = in[62] & in2[62];
    assign P[102] = in[62] ^ in2[62];
    assign G[103] = in[61] & in2[61];
    assign P[103] = in[61] ^ in2[61];
    assign G[104] = in[60] & in2[60];
    assign P[104] = in[60] ^ in2[60];
    assign G[105] = in[59] & in2[59];
    assign P[105] = in[59] ^ in2[59];
    assign G[106] = in[58] & in2[58];
    assign P[106] = in[58] ^ in2[58];
    assign G[107] = in[57] & in2[57];
    assign P[107] = in[57] ^ in2[57];
    assign G[108] = in[56] & in2[56];
    assign P[108] = in[56] ^ in2[56];
    assign G[109] = in[55] & in2[55];
    assign P[109] = in[55] ^ in2[55];
    assign G[110] = in[54] & in2[54];
    assign P[110] = in[54] ^ in2[54];
    assign G[111] = in[53] & in2[53];
    assign P[111] = in[53] ^ in2[53];
    assign G[112] = in[52] & in2[52];
    assign P[112] = in[52] ^ in2[52];
    assign G[113] = in[51] & in2[51];
    assign P[113] = in[51] ^ in2[51];
    assign G[114] = in[50] & in2[50];
    assign P[114] = in[50] ^ in2[50];
    assign G[115] = in[49] & in2[49];
    assign P[115] = in[49] ^ in2[49];
    assign G[116] = in[48] & in2[48];
    assign P[116] = in[48] ^ in2[48];
    assign G[117] = in[47] & in2[47];
    assign P[117] = in[47] ^ in2[47];
    assign G[118] = in[46] & in2[46];
    assign P[118] = in[46] ^ in2[46];
    assign G[119] = in[45] & in2[45];
    assign P[119] = in[45] ^ in2[45];
    assign G[120] = in[44] & in2[44];
    assign P[120] = in[44] ^ in2[44];
    assign G[121] = in[43] & in2[43];
    assign P[121] = in[43] ^ in2[43];
    assign G[122] = in[42] & in2[42];
    assign P[122] = in[42] ^ in2[42];
    assign G[123] = in[41] & in2[41];
    assign P[123] = in[41] ^ in2[41];
    assign G[124] = in[40] & in2[40];
    assign P[124] = in[40] ^ in2[40];
    assign G[125] = in[39] & in2[39];
    assign P[125] = in[39] ^ in2[39];
    assign G[126] = in[38] & in2[38];
    assign P[126] = in[38] ^ in2[38];
    assign G[127] = in[37] & in2[37];
    assign P[127] = in[37] ^ in2[37];
    assign G[128] = in[36] & in2[36];
    assign P[128] = in[36] ^ in2[36];
    assign G[129] = in[35] & in2[35];
    assign P[129] = in[35] ^ in2[35];
    assign G[130] = in[34] & in2[34];
    assign P[130] = in[34] ^ in2[34];
    assign G[131] = in[33] & in2[33];
    assign P[131] = in[33] ^ in2[33];
    assign G[132] = in[32] & in2[32];
    assign P[132] = in[32] ^ in2[32];
    assign G[133] = in[31] & in2[31];
    assign P[133] = in[31] ^ in2[31];
    assign G[134] = in[30] & in2[30];
    assign P[134] = in[30] ^ in2[30];
    assign G[135] = in[29] & in2[29];
    assign P[135] = in[29] ^ in2[29];
    assign G[136] = in[28] & in2[28];
    assign P[136] = in[28] ^ in2[28];
    assign G[137] = in[27] & in2[27];
    assign P[137] = in[27] ^ in2[27];
    assign G[138] = in[26] & in2[26];
    assign P[138] = in[26] ^ in2[26];
    assign G[139] = in[25] & in2[25];
    assign P[139] = in[25] ^ in2[25];
    assign G[140] = in[24] & in2[24];
    assign P[140] = in[24] ^ in2[24];
    assign G[141] = in[23] & in2[23];
    assign P[141] = in[23] ^ in2[23];
    assign G[142] = in[22] & in2[22];
    assign P[142] = in[22] ^ in2[22];
    assign G[143] = in[21] & in2[21];
    assign P[143] = in[21] ^ in2[21];
    assign G[144] = in[20] & in2[20];
    assign P[144] = in[20] ^ in2[20];
    assign G[145] = in[19] & in2[19];
    assign P[145] = in[19] ^ in2[19];
    assign G[146] = in[18] & in2[18];
    assign P[146] = in[18] ^ in2[18];
    assign G[147] = in[17] & in2[17];
    assign P[147] = in[17] ^ in2[17];
    assign G[148] = in[16] & in2[16];
    assign P[148] = in[16] ^ in2[16];
    assign G[149] = in[15] & in2[15];
    assign P[149] = in[15] ^ in2[15];
    assign G[150] = in[14] & in2[14];
    assign P[150] = in[14] ^ in2[14];
    assign G[151] = in[13] & in2[13];
    assign P[151] = in[13] ^ in2[13];
    assign G[152] = in[12] & in2[12];
    assign P[152] = in[12] ^ in2[12];
    assign G[153] = in[11] & in2[11];
    assign P[153] = in[11] ^ in2[11];
    assign G[154] = in[10] & in2[10];
    assign P[154] = in[10] ^ in2[10];
    assign G[155] = in[9] & in2[9];
    assign P[155] = in[9] ^ in2[9];
    assign G[156] = in[8] & in2[8];
    assign P[156] = in[8] ^ in2[8];
    assign G[157] = in[7] & in2[7];
    assign P[157] = in[7] ^ in2[7];
    assign G[158] = in[6] & in2[6];
    assign P[158] = in[6] ^ in2[6];
    assign G[159] = in[5] & in2[5];
    assign P[159] = in[5] ^ in2[5];
    assign G[160] = in[4] & in2[4];
    assign P[160] = in[4] ^ in2[4];
    assign G[161] = in[3] & in2[3];
    assign P[161] = in[3] ^ in2[3];
    assign G[162] = in[2] & in2[2];
    assign P[162] = in[2] ^ in2[2];
    assign G[163] = in[1] & in2[1];
    assign P[163] = in[1] ^ in2[1];
    assign G[164] = in[0] & in2[0];
    assign P[164] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign C[164] = G[163] | (P[163] & C[163]);
    assign cout = G[164] | (P[164] & C[164]);
    assign sum = P ^ C;
endmodule

module CLA164(output [163:0] sum, output cout, input [163:0] in1, input [163:0] in2;

    wire[163:0] G;
    wire[163:0] C;
    wire[163:0] P;

    assign G[0] = in[163] & in2[163];
    assign P[0] = in[163] ^ in2[163];
    assign G[1] = in[162] & in2[162];
    assign P[1] = in[162] ^ in2[162];
    assign G[2] = in[161] & in2[161];
    assign P[2] = in[161] ^ in2[161];
    assign G[3] = in[160] & in2[160];
    assign P[3] = in[160] ^ in2[160];
    assign G[4] = in[159] & in2[159];
    assign P[4] = in[159] ^ in2[159];
    assign G[5] = in[158] & in2[158];
    assign P[5] = in[158] ^ in2[158];
    assign G[6] = in[157] & in2[157];
    assign P[6] = in[157] ^ in2[157];
    assign G[7] = in[156] & in2[156];
    assign P[7] = in[156] ^ in2[156];
    assign G[8] = in[155] & in2[155];
    assign P[8] = in[155] ^ in2[155];
    assign G[9] = in[154] & in2[154];
    assign P[9] = in[154] ^ in2[154];
    assign G[10] = in[153] & in2[153];
    assign P[10] = in[153] ^ in2[153];
    assign G[11] = in[152] & in2[152];
    assign P[11] = in[152] ^ in2[152];
    assign G[12] = in[151] & in2[151];
    assign P[12] = in[151] ^ in2[151];
    assign G[13] = in[150] & in2[150];
    assign P[13] = in[150] ^ in2[150];
    assign G[14] = in[149] & in2[149];
    assign P[14] = in[149] ^ in2[149];
    assign G[15] = in[148] & in2[148];
    assign P[15] = in[148] ^ in2[148];
    assign G[16] = in[147] & in2[147];
    assign P[16] = in[147] ^ in2[147];
    assign G[17] = in[146] & in2[146];
    assign P[17] = in[146] ^ in2[146];
    assign G[18] = in[145] & in2[145];
    assign P[18] = in[145] ^ in2[145];
    assign G[19] = in[144] & in2[144];
    assign P[19] = in[144] ^ in2[144];
    assign G[20] = in[143] & in2[143];
    assign P[20] = in[143] ^ in2[143];
    assign G[21] = in[142] & in2[142];
    assign P[21] = in[142] ^ in2[142];
    assign G[22] = in[141] & in2[141];
    assign P[22] = in[141] ^ in2[141];
    assign G[23] = in[140] & in2[140];
    assign P[23] = in[140] ^ in2[140];
    assign G[24] = in[139] & in2[139];
    assign P[24] = in[139] ^ in2[139];
    assign G[25] = in[138] & in2[138];
    assign P[25] = in[138] ^ in2[138];
    assign G[26] = in[137] & in2[137];
    assign P[26] = in[137] ^ in2[137];
    assign G[27] = in[136] & in2[136];
    assign P[27] = in[136] ^ in2[136];
    assign G[28] = in[135] & in2[135];
    assign P[28] = in[135] ^ in2[135];
    assign G[29] = in[134] & in2[134];
    assign P[29] = in[134] ^ in2[134];
    assign G[30] = in[133] & in2[133];
    assign P[30] = in[133] ^ in2[133];
    assign G[31] = in[132] & in2[132];
    assign P[31] = in[132] ^ in2[132];
    assign G[32] = in[131] & in2[131];
    assign P[32] = in[131] ^ in2[131];
    assign G[33] = in[130] & in2[130];
    assign P[33] = in[130] ^ in2[130];
    assign G[34] = in[129] & in2[129];
    assign P[34] = in[129] ^ in2[129];
    assign G[35] = in[128] & in2[128];
    assign P[35] = in[128] ^ in2[128];
    assign G[36] = in[127] & in2[127];
    assign P[36] = in[127] ^ in2[127];
    assign G[37] = in[126] & in2[126];
    assign P[37] = in[126] ^ in2[126];
    assign G[38] = in[125] & in2[125];
    assign P[38] = in[125] ^ in2[125];
    assign G[39] = in[124] & in2[124];
    assign P[39] = in[124] ^ in2[124];
    assign G[40] = in[123] & in2[123];
    assign P[40] = in[123] ^ in2[123];
    assign G[41] = in[122] & in2[122];
    assign P[41] = in[122] ^ in2[122];
    assign G[42] = in[121] & in2[121];
    assign P[42] = in[121] ^ in2[121];
    assign G[43] = in[120] & in2[120];
    assign P[43] = in[120] ^ in2[120];
    assign G[44] = in[119] & in2[119];
    assign P[44] = in[119] ^ in2[119];
    assign G[45] = in[118] & in2[118];
    assign P[45] = in[118] ^ in2[118];
    assign G[46] = in[117] & in2[117];
    assign P[46] = in[117] ^ in2[117];
    assign G[47] = in[116] & in2[116];
    assign P[47] = in[116] ^ in2[116];
    assign G[48] = in[115] & in2[115];
    assign P[48] = in[115] ^ in2[115];
    assign G[49] = in[114] & in2[114];
    assign P[49] = in[114] ^ in2[114];
    assign G[50] = in[113] & in2[113];
    assign P[50] = in[113] ^ in2[113];
    assign G[51] = in[112] & in2[112];
    assign P[51] = in[112] ^ in2[112];
    assign G[52] = in[111] & in2[111];
    assign P[52] = in[111] ^ in2[111];
    assign G[53] = in[110] & in2[110];
    assign P[53] = in[110] ^ in2[110];
    assign G[54] = in[109] & in2[109];
    assign P[54] = in[109] ^ in2[109];
    assign G[55] = in[108] & in2[108];
    assign P[55] = in[108] ^ in2[108];
    assign G[56] = in[107] & in2[107];
    assign P[56] = in[107] ^ in2[107];
    assign G[57] = in[106] & in2[106];
    assign P[57] = in[106] ^ in2[106];
    assign G[58] = in[105] & in2[105];
    assign P[58] = in[105] ^ in2[105];
    assign G[59] = in[104] & in2[104];
    assign P[59] = in[104] ^ in2[104];
    assign G[60] = in[103] & in2[103];
    assign P[60] = in[103] ^ in2[103];
    assign G[61] = in[102] & in2[102];
    assign P[61] = in[102] ^ in2[102];
    assign G[62] = in[101] & in2[101];
    assign P[62] = in[101] ^ in2[101];
    assign G[63] = in[100] & in2[100];
    assign P[63] = in[100] ^ in2[100];
    assign G[64] = in[99] & in2[99];
    assign P[64] = in[99] ^ in2[99];
    assign G[65] = in[98] & in2[98];
    assign P[65] = in[98] ^ in2[98];
    assign G[66] = in[97] & in2[97];
    assign P[66] = in[97] ^ in2[97];
    assign G[67] = in[96] & in2[96];
    assign P[67] = in[96] ^ in2[96];
    assign G[68] = in[95] & in2[95];
    assign P[68] = in[95] ^ in2[95];
    assign G[69] = in[94] & in2[94];
    assign P[69] = in[94] ^ in2[94];
    assign G[70] = in[93] & in2[93];
    assign P[70] = in[93] ^ in2[93];
    assign G[71] = in[92] & in2[92];
    assign P[71] = in[92] ^ in2[92];
    assign G[72] = in[91] & in2[91];
    assign P[72] = in[91] ^ in2[91];
    assign G[73] = in[90] & in2[90];
    assign P[73] = in[90] ^ in2[90];
    assign G[74] = in[89] & in2[89];
    assign P[74] = in[89] ^ in2[89];
    assign G[75] = in[88] & in2[88];
    assign P[75] = in[88] ^ in2[88];
    assign G[76] = in[87] & in2[87];
    assign P[76] = in[87] ^ in2[87];
    assign G[77] = in[86] & in2[86];
    assign P[77] = in[86] ^ in2[86];
    assign G[78] = in[85] & in2[85];
    assign P[78] = in[85] ^ in2[85];
    assign G[79] = in[84] & in2[84];
    assign P[79] = in[84] ^ in2[84];
    assign G[80] = in[83] & in2[83];
    assign P[80] = in[83] ^ in2[83];
    assign G[81] = in[82] & in2[82];
    assign P[81] = in[82] ^ in2[82];
    assign G[82] = in[81] & in2[81];
    assign P[82] = in[81] ^ in2[81];
    assign G[83] = in[80] & in2[80];
    assign P[83] = in[80] ^ in2[80];
    assign G[84] = in[79] & in2[79];
    assign P[84] = in[79] ^ in2[79];
    assign G[85] = in[78] & in2[78];
    assign P[85] = in[78] ^ in2[78];
    assign G[86] = in[77] & in2[77];
    assign P[86] = in[77] ^ in2[77];
    assign G[87] = in[76] & in2[76];
    assign P[87] = in[76] ^ in2[76];
    assign G[88] = in[75] & in2[75];
    assign P[88] = in[75] ^ in2[75];
    assign G[89] = in[74] & in2[74];
    assign P[89] = in[74] ^ in2[74];
    assign G[90] = in[73] & in2[73];
    assign P[90] = in[73] ^ in2[73];
    assign G[91] = in[72] & in2[72];
    assign P[91] = in[72] ^ in2[72];
    assign G[92] = in[71] & in2[71];
    assign P[92] = in[71] ^ in2[71];
    assign G[93] = in[70] & in2[70];
    assign P[93] = in[70] ^ in2[70];
    assign G[94] = in[69] & in2[69];
    assign P[94] = in[69] ^ in2[69];
    assign G[95] = in[68] & in2[68];
    assign P[95] = in[68] ^ in2[68];
    assign G[96] = in[67] & in2[67];
    assign P[96] = in[67] ^ in2[67];
    assign G[97] = in[66] & in2[66];
    assign P[97] = in[66] ^ in2[66];
    assign G[98] = in[65] & in2[65];
    assign P[98] = in[65] ^ in2[65];
    assign G[99] = in[64] & in2[64];
    assign P[99] = in[64] ^ in2[64];
    assign G[100] = in[63] & in2[63];
    assign P[100] = in[63] ^ in2[63];
    assign G[101] = in[62] & in2[62];
    assign P[101] = in[62] ^ in2[62];
    assign G[102] = in[61] & in2[61];
    assign P[102] = in[61] ^ in2[61];
    assign G[103] = in[60] & in2[60];
    assign P[103] = in[60] ^ in2[60];
    assign G[104] = in[59] & in2[59];
    assign P[104] = in[59] ^ in2[59];
    assign G[105] = in[58] & in2[58];
    assign P[105] = in[58] ^ in2[58];
    assign G[106] = in[57] & in2[57];
    assign P[106] = in[57] ^ in2[57];
    assign G[107] = in[56] & in2[56];
    assign P[107] = in[56] ^ in2[56];
    assign G[108] = in[55] & in2[55];
    assign P[108] = in[55] ^ in2[55];
    assign G[109] = in[54] & in2[54];
    assign P[109] = in[54] ^ in2[54];
    assign G[110] = in[53] & in2[53];
    assign P[110] = in[53] ^ in2[53];
    assign G[111] = in[52] & in2[52];
    assign P[111] = in[52] ^ in2[52];
    assign G[112] = in[51] & in2[51];
    assign P[112] = in[51] ^ in2[51];
    assign G[113] = in[50] & in2[50];
    assign P[113] = in[50] ^ in2[50];
    assign G[114] = in[49] & in2[49];
    assign P[114] = in[49] ^ in2[49];
    assign G[115] = in[48] & in2[48];
    assign P[115] = in[48] ^ in2[48];
    assign G[116] = in[47] & in2[47];
    assign P[116] = in[47] ^ in2[47];
    assign G[117] = in[46] & in2[46];
    assign P[117] = in[46] ^ in2[46];
    assign G[118] = in[45] & in2[45];
    assign P[118] = in[45] ^ in2[45];
    assign G[119] = in[44] & in2[44];
    assign P[119] = in[44] ^ in2[44];
    assign G[120] = in[43] & in2[43];
    assign P[120] = in[43] ^ in2[43];
    assign G[121] = in[42] & in2[42];
    assign P[121] = in[42] ^ in2[42];
    assign G[122] = in[41] & in2[41];
    assign P[122] = in[41] ^ in2[41];
    assign G[123] = in[40] & in2[40];
    assign P[123] = in[40] ^ in2[40];
    assign G[124] = in[39] & in2[39];
    assign P[124] = in[39] ^ in2[39];
    assign G[125] = in[38] & in2[38];
    assign P[125] = in[38] ^ in2[38];
    assign G[126] = in[37] & in2[37];
    assign P[126] = in[37] ^ in2[37];
    assign G[127] = in[36] & in2[36];
    assign P[127] = in[36] ^ in2[36];
    assign G[128] = in[35] & in2[35];
    assign P[128] = in[35] ^ in2[35];
    assign G[129] = in[34] & in2[34];
    assign P[129] = in[34] ^ in2[34];
    assign G[130] = in[33] & in2[33];
    assign P[130] = in[33] ^ in2[33];
    assign G[131] = in[32] & in2[32];
    assign P[131] = in[32] ^ in2[32];
    assign G[132] = in[31] & in2[31];
    assign P[132] = in[31] ^ in2[31];
    assign G[133] = in[30] & in2[30];
    assign P[133] = in[30] ^ in2[30];
    assign G[134] = in[29] & in2[29];
    assign P[134] = in[29] ^ in2[29];
    assign G[135] = in[28] & in2[28];
    assign P[135] = in[28] ^ in2[28];
    assign G[136] = in[27] & in2[27];
    assign P[136] = in[27] ^ in2[27];
    assign G[137] = in[26] & in2[26];
    assign P[137] = in[26] ^ in2[26];
    assign G[138] = in[25] & in2[25];
    assign P[138] = in[25] ^ in2[25];
    assign G[139] = in[24] & in2[24];
    assign P[139] = in[24] ^ in2[24];
    assign G[140] = in[23] & in2[23];
    assign P[140] = in[23] ^ in2[23];
    assign G[141] = in[22] & in2[22];
    assign P[141] = in[22] ^ in2[22];
    assign G[142] = in[21] & in2[21];
    assign P[142] = in[21] ^ in2[21];
    assign G[143] = in[20] & in2[20];
    assign P[143] = in[20] ^ in2[20];
    assign G[144] = in[19] & in2[19];
    assign P[144] = in[19] ^ in2[19];
    assign G[145] = in[18] & in2[18];
    assign P[145] = in[18] ^ in2[18];
    assign G[146] = in[17] & in2[17];
    assign P[146] = in[17] ^ in2[17];
    assign G[147] = in[16] & in2[16];
    assign P[147] = in[16] ^ in2[16];
    assign G[148] = in[15] & in2[15];
    assign P[148] = in[15] ^ in2[15];
    assign G[149] = in[14] & in2[14];
    assign P[149] = in[14] ^ in2[14];
    assign G[150] = in[13] & in2[13];
    assign P[150] = in[13] ^ in2[13];
    assign G[151] = in[12] & in2[12];
    assign P[151] = in[12] ^ in2[12];
    assign G[152] = in[11] & in2[11];
    assign P[152] = in[11] ^ in2[11];
    assign G[153] = in[10] & in2[10];
    assign P[153] = in[10] ^ in2[10];
    assign G[154] = in[9] & in2[9];
    assign P[154] = in[9] ^ in2[9];
    assign G[155] = in[8] & in2[8];
    assign P[155] = in[8] ^ in2[8];
    assign G[156] = in[7] & in2[7];
    assign P[156] = in[7] ^ in2[7];
    assign G[157] = in[6] & in2[6];
    assign P[157] = in[6] ^ in2[6];
    assign G[158] = in[5] & in2[5];
    assign P[158] = in[5] ^ in2[5];
    assign G[159] = in[4] & in2[4];
    assign P[159] = in[4] ^ in2[4];
    assign G[160] = in[3] & in2[3];
    assign P[160] = in[3] ^ in2[3];
    assign G[161] = in[2] & in2[2];
    assign P[161] = in[2] ^ in2[2];
    assign G[162] = in[1] & in2[1];
    assign P[162] = in[1] ^ in2[1];
    assign G[163] = in[0] & in2[0];
    assign P[163] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign C[163] = G[162] | (P[162] & C[162]);
    assign cout = G[163] | (P[163] & C[163]);
    assign sum = P ^ C;
endmodule

module CLA163(output [162:0] sum, output cout, input [162:0] in1, input [162:0] in2;

    wire[162:0] G;
    wire[162:0] C;
    wire[162:0] P;

    assign G[0] = in[162] & in2[162];
    assign P[0] = in[162] ^ in2[162];
    assign G[1] = in[161] & in2[161];
    assign P[1] = in[161] ^ in2[161];
    assign G[2] = in[160] & in2[160];
    assign P[2] = in[160] ^ in2[160];
    assign G[3] = in[159] & in2[159];
    assign P[3] = in[159] ^ in2[159];
    assign G[4] = in[158] & in2[158];
    assign P[4] = in[158] ^ in2[158];
    assign G[5] = in[157] & in2[157];
    assign P[5] = in[157] ^ in2[157];
    assign G[6] = in[156] & in2[156];
    assign P[6] = in[156] ^ in2[156];
    assign G[7] = in[155] & in2[155];
    assign P[7] = in[155] ^ in2[155];
    assign G[8] = in[154] & in2[154];
    assign P[8] = in[154] ^ in2[154];
    assign G[9] = in[153] & in2[153];
    assign P[9] = in[153] ^ in2[153];
    assign G[10] = in[152] & in2[152];
    assign P[10] = in[152] ^ in2[152];
    assign G[11] = in[151] & in2[151];
    assign P[11] = in[151] ^ in2[151];
    assign G[12] = in[150] & in2[150];
    assign P[12] = in[150] ^ in2[150];
    assign G[13] = in[149] & in2[149];
    assign P[13] = in[149] ^ in2[149];
    assign G[14] = in[148] & in2[148];
    assign P[14] = in[148] ^ in2[148];
    assign G[15] = in[147] & in2[147];
    assign P[15] = in[147] ^ in2[147];
    assign G[16] = in[146] & in2[146];
    assign P[16] = in[146] ^ in2[146];
    assign G[17] = in[145] & in2[145];
    assign P[17] = in[145] ^ in2[145];
    assign G[18] = in[144] & in2[144];
    assign P[18] = in[144] ^ in2[144];
    assign G[19] = in[143] & in2[143];
    assign P[19] = in[143] ^ in2[143];
    assign G[20] = in[142] & in2[142];
    assign P[20] = in[142] ^ in2[142];
    assign G[21] = in[141] & in2[141];
    assign P[21] = in[141] ^ in2[141];
    assign G[22] = in[140] & in2[140];
    assign P[22] = in[140] ^ in2[140];
    assign G[23] = in[139] & in2[139];
    assign P[23] = in[139] ^ in2[139];
    assign G[24] = in[138] & in2[138];
    assign P[24] = in[138] ^ in2[138];
    assign G[25] = in[137] & in2[137];
    assign P[25] = in[137] ^ in2[137];
    assign G[26] = in[136] & in2[136];
    assign P[26] = in[136] ^ in2[136];
    assign G[27] = in[135] & in2[135];
    assign P[27] = in[135] ^ in2[135];
    assign G[28] = in[134] & in2[134];
    assign P[28] = in[134] ^ in2[134];
    assign G[29] = in[133] & in2[133];
    assign P[29] = in[133] ^ in2[133];
    assign G[30] = in[132] & in2[132];
    assign P[30] = in[132] ^ in2[132];
    assign G[31] = in[131] & in2[131];
    assign P[31] = in[131] ^ in2[131];
    assign G[32] = in[130] & in2[130];
    assign P[32] = in[130] ^ in2[130];
    assign G[33] = in[129] & in2[129];
    assign P[33] = in[129] ^ in2[129];
    assign G[34] = in[128] & in2[128];
    assign P[34] = in[128] ^ in2[128];
    assign G[35] = in[127] & in2[127];
    assign P[35] = in[127] ^ in2[127];
    assign G[36] = in[126] & in2[126];
    assign P[36] = in[126] ^ in2[126];
    assign G[37] = in[125] & in2[125];
    assign P[37] = in[125] ^ in2[125];
    assign G[38] = in[124] & in2[124];
    assign P[38] = in[124] ^ in2[124];
    assign G[39] = in[123] & in2[123];
    assign P[39] = in[123] ^ in2[123];
    assign G[40] = in[122] & in2[122];
    assign P[40] = in[122] ^ in2[122];
    assign G[41] = in[121] & in2[121];
    assign P[41] = in[121] ^ in2[121];
    assign G[42] = in[120] & in2[120];
    assign P[42] = in[120] ^ in2[120];
    assign G[43] = in[119] & in2[119];
    assign P[43] = in[119] ^ in2[119];
    assign G[44] = in[118] & in2[118];
    assign P[44] = in[118] ^ in2[118];
    assign G[45] = in[117] & in2[117];
    assign P[45] = in[117] ^ in2[117];
    assign G[46] = in[116] & in2[116];
    assign P[46] = in[116] ^ in2[116];
    assign G[47] = in[115] & in2[115];
    assign P[47] = in[115] ^ in2[115];
    assign G[48] = in[114] & in2[114];
    assign P[48] = in[114] ^ in2[114];
    assign G[49] = in[113] & in2[113];
    assign P[49] = in[113] ^ in2[113];
    assign G[50] = in[112] & in2[112];
    assign P[50] = in[112] ^ in2[112];
    assign G[51] = in[111] & in2[111];
    assign P[51] = in[111] ^ in2[111];
    assign G[52] = in[110] & in2[110];
    assign P[52] = in[110] ^ in2[110];
    assign G[53] = in[109] & in2[109];
    assign P[53] = in[109] ^ in2[109];
    assign G[54] = in[108] & in2[108];
    assign P[54] = in[108] ^ in2[108];
    assign G[55] = in[107] & in2[107];
    assign P[55] = in[107] ^ in2[107];
    assign G[56] = in[106] & in2[106];
    assign P[56] = in[106] ^ in2[106];
    assign G[57] = in[105] & in2[105];
    assign P[57] = in[105] ^ in2[105];
    assign G[58] = in[104] & in2[104];
    assign P[58] = in[104] ^ in2[104];
    assign G[59] = in[103] & in2[103];
    assign P[59] = in[103] ^ in2[103];
    assign G[60] = in[102] & in2[102];
    assign P[60] = in[102] ^ in2[102];
    assign G[61] = in[101] & in2[101];
    assign P[61] = in[101] ^ in2[101];
    assign G[62] = in[100] & in2[100];
    assign P[62] = in[100] ^ in2[100];
    assign G[63] = in[99] & in2[99];
    assign P[63] = in[99] ^ in2[99];
    assign G[64] = in[98] & in2[98];
    assign P[64] = in[98] ^ in2[98];
    assign G[65] = in[97] & in2[97];
    assign P[65] = in[97] ^ in2[97];
    assign G[66] = in[96] & in2[96];
    assign P[66] = in[96] ^ in2[96];
    assign G[67] = in[95] & in2[95];
    assign P[67] = in[95] ^ in2[95];
    assign G[68] = in[94] & in2[94];
    assign P[68] = in[94] ^ in2[94];
    assign G[69] = in[93] & in2[93];
    assign P[69] = in[93] ^ in2[93];
    assign G[70] = in[92] & in2[92];
    assign P[70] = in[92] ^ in2[92];
    assign G[71] = in[91] & in2[91];
    assign P[71] = in[91] ^ in2[91];
    assign G[72] = in[90] & in2[90];
    assign P[72] = in[90] ^ in2[90];
    assign G[73] = in[89] & in2[89];
    assign P[73] = in[89] ^ in2[89];
    assign G[74] = in[88] & in2[88];
    assign P[74] = in[88] ^ in2[88];
    assign G[75] = in[87] & in2[87];
    assign P[75] = in[87] ^ in2[87];
    assign G[76] = in[86] & in2[86];
    assign P[76] = in[86] ^ in2[86];
    assign G[77] = in[85] & in2[85];
    assign P[77] = in[85] ^ in2[85];
    assign G[78] = in[84] & in2[84];
    assign P[78] = in[84] ^ in2[84];
    assign G[79] = in[83] & in2[83];
    assign P[79] = in[83] ^ in2[83];
    assign G[80] = in[82] & in2[82];
    assign P[80] = in[82] ^ in2[82];
    assign G[81] = in[81] & in2[81];
    assign P[81] = in[81] ^ in2[81];
    assign G[82] = in[80] & in2[80];
    assign P[82] = in[80] ^ in2[80];
    assign G[83] = in[79] & in2[79];
    assign P[83] = in[79] ^ in2[79];
    assign G[84] = in[78] & in2[78];
    assign P[84] = in[78] ^ in2[78];
    assign G[85] = in[77] & in2[77];
    assign P[85] = in[77] ^ in2[77];
    assign G[86] = in[76] & in2[76];
    assign P[86] = in[76] ^ in2[76];
    assign G[87] = in[75] & in2[75];
    assign P[87] = in[75] ^ in2[75];
    assign G[88] = in[74] & in2[74];
    assign P[88] = in[74] ^ in2[74];
    assign G[89] = in[73] & in2[73];
    assign P[89] = in[73] ^ in2[73];
    assign G[90] = in[72] & in2[72];
    assign P[90] = in[72] ^ in2[72];
    assign G[91] = in[71] & in2[71];
    assign P[91] = in[71] ^ in2[71];
    assign G[92] = in[70] & in2[70];
    assign P[92] = in[70] ^ in2[70];
    assign G[93] = in[69] & in2[69];
    assign P[93] = in[69] ^ in2[69];
    assign G[94] = in[68] & in2[68];
    assign P[94] = in[68] ^ in2[68];
    assign G[95] = in[67] & in2[67];
    assign P[95] = in[67] ^ in2[67];
    assign G[96] = in[66] & in2[66];
    assign P[96] = in[66] ^ in2[66];
    assign G[97] = in[65] & in2[65];
    assign P[97] = in[65] ^ in2[65];
    assign G[98] = in[64] & in2[64];
    assign P[98] = in[64] ^ in2[64];
    assign G[99] = in[63] & in2[63];
    assign P[99] = in[63] ^ in2[63];
    assign G[100] = in[62] & in2[62];
    assign P[100] = in[62] ^ in2[62];
    assign G[101] = in[61] & in2[61];
    assign P[101] = in[61] ^ in2[61];
    assign G[102] = in[60] & in2[60];
    assign P[102] = in[60] ^ in2[60];
    assign G[103] = in[59] & in2[59];
    assign P[103] = in[59] ^ in2[59];
    assign G[104] = in[58] & in2[58];
    assign P[104] = in[58] ^ in2[58];
    assign G[105] = in[57] & in2[57];
    assign P[105] = in[57] ^ in2[57];
    assign G[106] = in[56] & in2[56];
    assign P[106] = in[56] ^ in2[56];
    assign G[107] = in[55] & in2[55];
    assign P[107] = in[55] ^ in2[55];
    assign G[108] = in[54] & in2[54];
    assign P[108] = in[54] ^ in2[54];
    assign G[109] = in[53] & in2[53];
    assign P[109] = in[53] ^ in2[53];
    assign G[110] = in[52] & in2[52];
    assign P[110] = in[52] ^ in2[52];
    assign G[111] = in[51] & in2[51];
    assign P[111] = in[51] ^ in2[51];
    assign G[112] = in[50] & in2[50];
    assign P[112] = in[50] ^ in2[50];
    assign G[113] = in[49] & in2[49];
    assign P[113] = in[49] ^ in2[49];
    assign G[114] = in[48] & in2[48];
    assign P[114] = in[48] ^ in2[48];
    assign G[115] = in[47] & in2[47];
    assign P[115] = in[47] ^ in2[47];
    assign G[116] = in[46] & in2[46];
    assign P[116] = in[46] ^ in2[46];
    assign G[117] = in[45] & in2[45];
    assign P[117] = in[45] ^ in2[45];
    assign G[118] = in[44] & in2[44];
    assign P[118] = in[44] ^ in2[44];
    assign G[119] = in[43] & in2[43];
    assign P[119] = in[43] ^ in2[43];
    assign G[120] = in[42] & in2[42];
    assign P[120] = in[42] ^ in2[42];
    assign G[121] = in[41] & in2[41];
    assign P[121] = in[41] ^ in2[41];
    assign G[122] = in[40] & in2[40];
    assign P[122] = in[40] ^ in2[40];
    assign G[123] = in[39] & in2[39];
    assign P[123] = in[39] ^ in2[39];
    assign G[124] = in[38] & in2[38];
    assign P[124] = in[38] ^ in2[38];
    assign G[125] = in[37] & in2[37];
    assign P[125] = in[37] ^ in2[37];
    assign G[126] = in[36] & in2[36];
    assign P[126] = in[36] ^ in2[36];
    assign G[127] = in[35] & in2[35];
    assign P[127] = in[35] ^ in2[35];
    assign G[128] = in[34] & in2[34];
    assign P[128] = in[34] ^ in2[34];
    assign G[129] = in[33] & in2[33];
    assign P[129] = in[33] ^ in2[33];
    assign G[130] = in[32] & in2[32];
    assign P[130] = in[32] ^ in2[32];
    assign G[131] = in[31] & in2[31];
    assign P[131] = in[31] ^ in2[31];
    assign G[132] = in[30] & in2[30];
    assign P[132] = in[30] ^ in2[30];
    assign G[133] = in[29] & in2[29];
    assign P[133] = in[29] ^ in2[29];
    assign G[134] = in[28] & in2[28];
    assign P[134] = in[28] ^ in2[28];
    assign G[135] = in[27] & in2[27];
    assign P[135] = in[27] ^ in2[27];
    assign G[136] = in[26] & in2[26];
    assign P[136] = in[26] ^ in2[26];
    assign G[137] = in[25] & in2[25];
    assign P[137] = in[25] ^ in2[25];
    assign G[138] = in[24] & in2[24];
    assign P[138] = in[24] ^ in2[24];
    assign G[139] = in[23] & in2[23];
    assign P[139] = in[23] ^ in2[23];
    assign G[140] = in[22] & in2[22];
    assign P[140] = in[22] ^ in2[22];
    assign G[141] = in[21] & in2[21];
    assign P[141] = in[21] ^ in2[21];
    assign G[142] = in[20] & in2[20];
    assign P[142] = in[20] ^ in2[20];
    assign G[143] = in[19] & in2[19];
    assign P[143] = in[19] ^ in2[19];
    assign G[144] = in[18] & in2[18];
    assign P[144] = in[18] ^ in2[18];
    assign G[145] = in[17] & in2[17];
    assign P[145] = in[17] ^ in2[17];
    assign G[146] = in[16] & in2[16];
    assign P[146] = in[16] ^ in2[16];
    assign G[147] = in[15] & in2[15];
    assign P[147] = in[15] ^ in2[15];
    assign G[148] = in[14] & in2[14];
    assign P[148] = in[14] ^ in2[14];
    assign G[149] = in[13] & in2[13];
    assign P[149] = in[13] ^ in2[13];
    assign G[150] = in[12] & in2[12];
    assign P[150] = in[12] ^ in2[12];
    assign G[151] = in[11] & in2[11];
    assign P[151] = in[11] ^ in2[11];
    assign G[152] = in[10] & in2[10];
    assign P[152] = in[10] ^ in2[10];
    assign G[153] = in[9] & in2[9];
    assign P[153] = in[9] ^ in2[9];
    assign G[154] = in[8] & in2[8];
    assign P[154] = in[8] ^ in2[8];
    assign G[155] = in[7] & in2[7];
    assign P[155] = in[7] ^ in2[7];
    assign G[156] = in[6] & in2[6];
    assign P[156] = in[6] ^ in2[6];
    assign G[157] = in[5] & in2[5];
    assign P[157] = in[5] ^ in2[5];
    assign G[158] = in[4] & in2[4];
    assign P[158] = in[4] ^ in2[4];
    assign G[159] = in[3] & in2[3];
    assign P[159] = in[3] ^ in2[3];
    assign G[160] = in[2] & in2[2];
    assign P[160] = in[2] ^ in2[2];
    assign G[161] = in[1] & in2[1];
    assign P[161] = in[1] ^ in2[1];
    assign G[162] = in[0] & in2[0];
    assign P[162] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign C[162] = G[161] | (P[161] & C[161]);
    assign cout = G[162] | (P[162] & C[162]);
    assign sum = P ^ C;
endmodule

module CLA162(output [161:0] sum, output cout, input [161:0] in1, input [161:0] in2;

    wire[161:0] G;
    wire[161:0] C;
    wire[161:0] P;

    assign G[0] = in[161] & in2[161];
    assign P[0] = in[161] ^ in2[161];
    assign G[1] = in[160] & in2[160];
    assign P[1] = in[160] ^ in2[160];
    assign G[2] = in[159] & in2[159];
    assign P[2] = in[159] ^ in2[159];
    assign G[3] = in[158] & in2[158];
    assign P[3] = in[158] ^ in2[158];
    assign G[4] = in[157] & in2[157];
    assign P[4] = in[157] ^ in2[157];
    assign G[5] = in[156] & in2[156];
    assign P[5] = in[156] ^ in2[156];
    assign G[6] = in[155] & in2[155];
    assign P[6] = in[155] ^ in2[155];
    assign G[7] = in[154] & in2[154];
    assign P[7] = in[154] ^ in2[154];
    assign G[8] = in[153] & in2[153];
    assign P[8] = in[153] ^ in2[153];
    assign G[9] = in[152] & in2[152];
    assign P[9] = in[152] ^ in2[152];
    assign G[10] = in[151] & in2[151];
    assign P[10] = in[151] ^ in2[151];
    assign G[11] = in[150] & in2[150];
    assign P[11] = in[150] ^ in2[150];
    assign G[12] = in[149] & in2[149];
    assign P[12] = in[149] ^ in2[149];
    assign G[13] = in[148] & in2[148];
    assign P[13] = in[148] ^ in2[148];
    assign G[14] = in[147] & in2[147];
    assign P[14] = in[147] ^ in2[147];
    assign G[15] = in[146] & in2[146];
    assign P[15] = in[146] ^ in2[146];
    assign G[16] = in[145] & in2[145];
    assign P[16] = in[145] ^ in2[145];
    assign G[17] = in[144] & in2[144];
    assign P[17] = in[144] ^ in2[144];
    assign G[18] = in[143] & in2[143];
    assign P[18] = in[143] ^ in2[143];
    assign G[19] = in[142] & in2[142];
    assign P[19] = in[142] ^ in2[142];
    assign G[20] = in[141] & in2[141];
    assign P[20] = in[141] ^ in2[141];
    assign G[21] = in[140] & in2[140];
    assign P[21] = in[140] ^ in2[140];
    assign G[22] = in[139] & in2[139];
    assign P[22] = in[139] ^ in2[139];
    assign G[23] = in[138] & in2[138];
    assign P[23] = in[138] ^ in2[138];
    assign G[24] = in[137] & in2[137];
    assign P[24] = in[137] ^ in2[137];
    assign G[25] = in[136] & in2[136];
    assign P[25] = in[136] ^ in2[136];
    assign G[26] = in[135] & in2[135];
    assign P[26] = in[135] ^ in2[135];
    assign G[27] = in[134] & in2[134];
    assign P[27] = in[134] ^ in2[134];
    assign G[28] = in[133] & in2[133];
    assign P[28] = in[133] ^ in2[133];
    assign G[29] = in[132] & in2[132];
    assign P[29] = in[132] ^ in2[132];
    assign G[30] = in[131] & in2[131];
    assign P[30] = in[131] ^ in2[131];
    assign G[31] = in[130] & in2[130];
    assign P[31] = in[130] ^ in2[130];
    assign G[32] = in[129] & in2[129];
    assign P[32] = in[129] ^ in2[129];
    assign G[33] = in[128] & in2[128];
    assign P[33] = in[128] ^ in2[128];
    assign G[34] = in[127] & in2[127];
    assign P[34] = in[127] ^ in2[127];
    assign G[35] = in[126] & in2[126];
    assign P[35] = in[126] ^ in2[126];
    assign G[36] = in[125] & in2[125];
    assign P[36] = in[125] ^ in2[125];
    assign G[37] = in[124] & in2[124];
    assign P[37] = in[124] ^ in2[124];
    assign G[38] = in[123] & in2[123];
    assign P[38] = in[123] ^ in2[123];
    assign G[39] = in[122] & in2[122];
    assign P[39] = in[122] ^ in2[122];
    assign G[40] = in[121] & in2[121];
    assign P[40] = in[121] ^ in2[121];
    assign G[41] = in[120] & in2[120];
    assign P[41] = in[120] ^ in2[120];
    assign G[42] = in[119] & in2[119];
    assign P[42] = in[119] ^ in2[119];
    assign G[43] = in[118] & in2[118];
    assign P[43] = in[118] ^ in2[118];
    assign G[44] = in[117] & in2[117];
    assign P[44] = in[117] ^ in2[117];
    assign G[45] = in[116] & in2[116];
    assign P[45] = in[116] ^ in2[116];
    assign G[46] = in[115] & in2[115];
    assign P[46] = in[115] ^ in2[115];
    assign G[47] = in[114] & in2[114];
    assign P[47] = in[114] ^ in2[114];
    assign G[48] = in[113] & in2[113];
    assign P[48] = in[113] ^ in2[113];
    assign G[49] = in[112] & in2[112];
    assign P[49] = in[112] ^ in2[112];
    assign G[50] = in[111] & in2[111];
    assign P[50] = in[111] ^ in2[111];
    assign G[51] = in[110] & in2[110];
    assign P[51] = in[110] ^ in2[110];
    assign G[52] = in[109] & in2[109];
    assign P[52] = in[109] ^ in2[109];
    assign G[53] = in[108] & in2[108];
    assign P[53] = in[108] ^ in2[108];
    assign G[54] = in[107] & in2[107];
    assign P[54] = in[107] ^ in2[107];
    assign G[55] = in[106] & in2[106];
    assign P[55] = in[106] ^ in2[106];
    assign G[56] = in[105] & in2[105];
    assign P[56] = in[105] ^ in2[105];
    assign G[57] = in[104] & in2[104];
    assign P[57] = in[104] ^ in2[104];
    assign G[58] = in[103] & in2[103];
    assign P[58] = in[103] ^ in2[103];
    assign G[59] = in[102] & in2[102];
    assign P[59] = in[102] ^ in2[102];
    assign G[60] = in[101] & in2[101];
    assign P[60] = in[101] ^ in2[101];
    assign G[61] = in[100] & in2[100];
    assign P[61] = in[100] ^ in2[100];
    assign G[62] = in[99] & in2[99];
    assign P[62] = in[99] ^ in2[99];
    assign G[63] = in[98] & in2[98];
    assign P[63] = in[98] ^ in2[98];
    assign G[64] = in[97] & in2[97];
    assign P[64] = in[97] ^ in2[97];
    assign G[65] = in[96] & in2[96];
    assign P[65] = in[96] ^ in2[96];
    assign G[66] = in[95] & in2[95];
    assign P[66] = in[95] ^ in2[95];
    assign G[67] = in[94] & in2[94];
    assign P[67] = in[94] ^ in2[94];
    assign G[68] = in[93] & in2[93];
    assign P[68] = in[93] ^ in2[93];
    assign G[69] = in[92] & in2[92];
    assign P[69] = in[92] ^ in2[92];
    assign G[70] = in[91] & in2[91];
    assign P[70] = in[91] ^ in2[91];
    assign G[71] = in[90] & in2[90];
    assign P[71] = in[90] ^ in2[90];
    assign G[72] = in[89] & in2[89];
    assign P[72] = in[89] ^ in2[89];
    assign G[73] = in[88] & in2[88];
    assign P[73] = in[88] ^ in2[88];
    assign G[74] = in[87] & in2[87];
    assign P[74] = in[87] ^ in2[87];
    assign G[75] = in[86] & in2[86];
    assign P[75] = in[86] ^ in2[86];
    assign G[76] = in[85] & in2[85];
    assign P[76] = in[85] ^ in2[85];
    assign G[77] = in[84] & in2[84];
    assign P[77] = in[84] ^ in2[84];
    assign G[78] = in[83] & in2[83];
    assign P[78] = in[83] ^ in2[83];
    assign G[79] = in[82] & in2[82];
    assign P[79] = in[82] ^ in2[82];
    assign G[80] = in[81] & in2[81];
    assign P[80] = in[81] ^ in2[81];
    assign G[81] = in[80] & in2[80];
    assign P[81] = in[80] ^ in2[80];
    assign G[82] = in[79] & in2[79];
    assign P[82] = in[79] ^ in2[79];
    assign G[83] = in[78] & in2[78];
    assign P[83] = in[78] ^ in2[78];
    assign G[84] = in[77] & in2[77];
    assign P[84] = in[77] ^ in2[77];
    assign G[85] = in[76] & in2[76];
    assign P[85] = in[76] ^ in2[76];
    assign G[86] = in[75] & in2[75];
    assign P[86] = in[75] ^ in2[75];
    assign G[87] = in[74] & in2[74];
    assign P[87] = in[74] ^ in2[74];
    assign G[88] = in[73] & in2[73];
    assign P[88] = in[73] ^ in2[73];
    assign G[89] = in[72] & in2[72];
    assign P[89] = in[72] ^ in2[72];
    assign G[90] = in[71] & in2[71];
    assign P[90] = in[71] ^ in2[71];
    assign G[91] = in[70] & in2[70];
    assign P[91] = in[70] ^ in2[70];
    assign G[92] = in[69] & in2[69];
    assign P[92] = in[69] ^ in2[69];
    assign G[93] = in[68] & in2[68];
    assign P[93] = in[68] ^ in2[68];
    assign G[94] = in[67] & in2[67];
    assign P[94] = in[67] ^ in2[67];
    assign G[95] = in[66] & in2[66];
    assign P[95] = in[66] ^ in2[66];
    assign G[96] = in[65] & in2[65];
    assign P[96] = in[65] ^ in2[65];
    assign G[97] = in[64] & in2[64];
    assign P[97] = in[64] ^ in2[64];
    assign G[98] = in[63] & in2[63];
    assign P[98] = in[63] ^ in2[63];
    assign G[99] = in[62] & in2[62];
    assign P[99] = in[62] ^ in2[62];
    assign G[100] = in[61] & in2[61];
    assign P[100] = in[61] ^ in2[61];
    assign G[101] = in[60] & in2[60];
    assign P[101] = in[60] ^ in2[60];
    assign G[102] = in[59] & in2[59];
    assign P[102] = in[59] ^ in2[59];
    assign G[103] = in[58] & in2[58];
    assign P[103] = in[58] ^ in2[58];
    assign G[104] = in[57] & in2[57];
    assign P[104] = in[57] ^ in2[57];
    assign G[105] = in[56] & in2[56];
    assign P[105] = in[56] ^ in2[56];
    assign G[106] = in[55] & in2[55];
    assign P[106] = in[55] ^ in2[55];
    assign G[107] = in[54] & in2[54];
    assign P[107] = in[54] ^ in2[54];
    assign G[108] = in[53] & in2[53];
    assign P[108] = in[53] ^ in2[53];
    assign G[109] = in[52] & in2[52];
    assign P[109] = in[52] ^ in2[52];
    assign G[110] = in[51] & in2[51];
    assign P[110] = in[51] ^ in2[51];
    assign G[111] = in[50] & in2[50];
    assign P[111] = in[50] ^ in2[50];
    assign G[112] = in[49] & in2[49];
    assign P[112] = in[49] ^ in2[49];
    assign G[113] = in[48] & in2[48];
    assign P[113] = in[48] ^ in2[48];
    assign G[114] = in[47] & in2[47];
    assign P[114] = in[47] ^ in2[47];
    assign G[115] = in[46] & in2[46];
    assign P[115] = in[46] ^ in2[46];
    assign G[116] = in[45] & in2[45];
    assign P[116] = in[45] ^ in2[45];
    assign G[117] = in[44] & in2[44];
    assign P[117] = in[44] ^ in2[44];
    assign G[118] = in[43] & in2[43];
    assign P[118] = in[43] ^ in2[43];
    assign G[119] = in[42] & in2[42];
    assign P[119] = in[42] ^ in2[42];
    assign G[120] = in[41] & in2[41];
    assign P[120] = in[41] ^ in2[41];
    assign G[121] = in[40] & in2[40];
    assign P[121] = in[40] ^ in2[40];
    assign G[122] = in[39] & in2[39];
    assign P[122] = in[39] ^ in2[39];
    assign G[123] = in[38] & in2[38];
    assign P[123] = in[38] ^ in2[38];
    assign G[124] = in[37] & in2[37];
    assign P[124] = in[37] ^ in2[37];
    assign G[125] = in[36] & in2[36];
    assign P[125] = in[36] ^ in2[36];
    assign G[126] = in[35] & in2[35];
    assign P[126] = in[35] ^ in2[35];
    assign G[127] = in[34] & in2[34];
    assign P[127] = in[34] ^ in2[34];
    assign G[128] = in[33] & in2[33];
    assign P[128] = in[33] ^ in2[33];
    assign G[129] = in[32] & in2[32];
    assign P[129] = in[32] ^ in2[32];
    assign G[130] = in[31] & in2[31];
    assign P[130] = in[31] ^ in2[31];
    assign G[131] = in[30] & in2[30];
    assign P[131] = in[30] ^ in2[30];
    assign G[132] = in[29] & in2[29];
    assign P[132] = in[29] ^ in2[29];
    assign G[133] = in[28] & in2[28];
    assign P[133] = in[28] ^ in2[28];
    assign G[134] = in[27] & in2[27];
    assign P[134] = in[27] ^ in2[27];
    assign G[135] = in[26] & in2[26];
    assign P[135] = in[26] ^ in2[26];
    assign G[136] = in[25] & in2[25];
    assign P[136] = in[25] ^ in2[25];
    assign G[137] = in[24] & in2[24];
    assign P[137] = in[24] ^ in2[24];
    assign G[138] = in[23] & in2[23];
    assign P[138] = in[23] ^ in2[23];
    assign G[139] = in[22] & in2[22];
    assign P[139] = in[22] ^ in2[22];
    assign G[140] = in[21] & in2[21];
    assign P[140] = in[21] ^ in2[21];
    assign G[141] = in[20] & in2[20];
    assign P[141] = in[20] ^ in2[20];
    assign G[142] = in[19] & in2[19];
    assign P[142] = in[19] ^ in2[19];
    assign G[143] = in[18] & in2[18];
    assign P[143] = in[18] ^ in2[18];
    assign G[144] = in[17] & in2[17];
    assign P[144] = in[17] ^ in2[17];
    assign G[145] = in[16] & in2[16];
    assign P[145] = in[16] ^ in2[16];
    assign G[146] = in[15] & in2[15];
    assign P[146] = in[15] ^ in2[15];
    assign G[147] = in[14] & in2[14];
    assign P[147] = in[14] ^ in2[14];
    assign G[148] = in[13] & in2[13];
    assign P[148] = in[13] ^ in2[13];
    assign G[149] = in[12] & in2[12];
    assign P[149] = in[12] ^ in2[12];
    assign G[150] = in[11] & in2[11];
    assign P[150] = in[11] ^ in2[11];
    assign G[151] = in[10] & in2[10];
    assign P[151] = in[10] ^ in2[10];
    assign G[152] = in[9] & in2[9];
    assign P[152] = in[9] ^ in2[9];
    assign G[153] = in[8] & in2[8];
    assign P[153] = in[8] ^ in2[8];
    assign G[154] = in[7] & in2[7];
    assign P[154] = in[7] ^ in2[7];
    assign G[155] = in[6] & in2[6];
    assign P[155] = in[6] ^ in2[6];
    assign G[156] = in[5] & in2[5];
    assign P[156] = in[5] ^ in2[5];
    assign G[157] = in[4] & in2[4];
    assign P[157] = in[4] ^ in2[4];
    assign G[158] = in[3] & in2[3];
    assign P[158] = in[3] ^ in2[3];
    assign G[159] = in[2] & in2[2];
    assign P[159] = in[2] ^ in2[2];
    assign G[160] = in[1] & in2[1];
    assign P[160] = in[1] ^ in2[1];
    assign G[161] = in[0] & in2[0];
    assign P[161] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign C[161] = G[160] | (P[160] & C[160]);
    assign cout = G[161] | (P[161] & C[161]);
    assign sum = P ^ C;
endmodule

module CLA161(output [160:0] sum, output cout, input [160:0] in1, input [160:0] in2;

    wire[160:0] G;
    wire[160:0] C;
    wire[160:0] P;

    assign G[0] = in[160] & in2[160];
    assign P[0] = in[160] ^ in2[160];
    assign G[1] = in[159] & in2[159];
    assign P[1] = in[159] ^ in2[159];
    assign G[2] = in[158] & in2[158];
    assign P[2] = in[158] ^ in2[158];
    assign G[3] = in[157] & in2[157];
    assign P[3] = in[157] ^ in2[157];
    assign G[4] = in[156] & in2[156];
    assign P[4] = in[156] ^ in2[156];
    assign G[5] = in[155] & in2[155];
    assign P[5] = in[155] ^ in2[155];
    assign G[6] = in[154] & in2[154];
    assign P[6] = in[154] ^ in2[154];
    assign G[7] = in[153] & in2[153];
    assign P[7] = in[153] ^ in2[153];
    assign G[8] = in[152] & in2[152];
    assign P[8] = in[152] ^ in2[152];
    assign G[9] = in[151] & in2[151];
    assign P[9] = in[151] ^ in2[151];
    assign G[10] = in[150] & in2[150];
    assign P[10] = in[150] ^ in2[150];
    assign G[11] = in[149] & in2[149];
    assign P[11] = in[149] ^ in2[149];
    assign G[12] = in[148] & in2[148];
    assign P[12] = in[148] ^ in2[148];
    assign G[13] = in[147] & in2[147];
    assign P[13] = in[147] ^ in2[147];
    assign G[14] = in[146] & in2[146];
    assign P[14] = in[146] ^ in2[146];
    assign G[15] = in[145] & in2[145];
    assign P[15] = in[145] ^ in2[145];
    assign G[16] = in[144] & in2[144];
    assign P[16] = in[144] ^ in2[144];
    assign G[17] = in[143] & in2[143];
    assign P[17] = in[143] ^ in2[143];
    assign G[18] = in[142] & in2[142];
    assign P[18] = in[142] ^ in2[142];
    assign G[19] = in[141] & in2[141];
    assign P[19] = in[141] ^ in2[141];
    assign G[20] = in[140] & in2[140];
    assign P[20] = in[140] ^ in2[140];
    assign G[21] = in[139] & in2[139];
    assign P[21] = in[139] ^ in2[139];
    assign G[22] = in[138] & in2[138];
    assign P[22] = in[138] ^ in2[138];
    assign G[23] = in[137] & in2[137];
    assign P[23] = in[137] ^ in2[137];
    assign G[24] = in[136] & in2[136];
    assign P[24] = in[136] ^ in2[136];
    assign G[25] = in[135] & in2[135];
    assign P[25] = in[135] ^ in2[135];
    assign G[26] = in[134] & in2[134];
    assign P[26] = in[134] ^ in2[134];
    assign G[27] = in[133] & in2[133];
    assign P[27] = in[133] ^ in2[133];
    assign G[28] = in[132] & in2[132];
    assign P[28] = in[132] ^ in2[132];
    assign G[29] = in[131] & in2[131];
    assign P[29] = in[131] ^ in2[131];
    assign G[30] = in[130] & in2[130];
    assign P[30] = in[130] ^ in2[130];
    assign G[31] = in[129] & in2[129];
    assign P[31] = in[129] ^ in2[129];
    assign G[32] = in[128] & in2[128];
    assign P[32] = in[128] ^ in2[128];
    assign G[33] = in[127] & in2[127];
    assign P[33] = in[127] ^ in2[127];
    assign G[34] = in[126] & in2[126];
    assign P[34] = in[126] ^ in2[126];
    assign G[35] = in[125] & in2[125];
    assign P[35] = in[125] ^ in2[125];
    assign G[36] = in[124] & in2[124];
    assign P[36] = in[124] ^ in2[124];
    assign G[37] = in[123] & in2[123];
    assign P[37] = in[123] ^ in2[123];
    assign G[38] = in[122] & in2[122];
    assign P[38] = in[122] ^ in2[122];
    assign G[39] = in[121] & in2[121];
    assign P[39] = in[121] ^ in2[121];
    assign G[40] = in[120] & in2[120];
    assign P[40] = in[120] ^ in2[120];
    assign G[41] = in[119] & in2[119];
    assign P[41] = in[119] ^ in2[119];
    assign G[42] = in[118] & in2[118];
    assign P[42] = in[118] ^ in2[118];
    assign G[43] = in[117] & in2[117];
    assign P[43] = in[117] ^ in2[117];
    assign G[44] = in[116] & in2[116];
    assign P[44] = in[116] ^ in2[116];
    assign G[45] = in[115] & in2[115];
    assign P[45] = in[115] ^ in2[115];
    assign G[46] = in[114] & in2[114];
    assign P[46] = in[114] ^ in2[114];
    assign G[47] = in[113] & in2[113];
    assign P[47] = in[113] ^ in2[113];
    assign G[48] = in[112] & in2[112];
    assign P[48] = in[112] ^ in2[112];
    assign G[49] = in[111] & in2[111];
    assign P[49] = in[111] ^ in2[111];
    assign G[50] = in[110] & in2[110];
    assign P[50] = in[110] ^ in2[110];
    assign G[51] = in[109] & in2[109];
    assign P[51] = in[109] ^ in2[109];
    assign G[52] = in[108] & in2[108];
    assign P[52] = in[108] ^ in2[108];
    assign G[53] = in[107] & in2[107];
    assign P[53] = in[107] ^ in2[107];
    assign G[54] = in[106] & in2[106];
    assign P[54] = in[106] ^ in2[106];
    assign G[55] = in[105] & in2[105];
    assign P[55] = in[105] ^ in2[105];
    assign G[56] = in[104] & in2[104];
    assign P[56] = in[104] ^ in2[104];
    assign G[57] = in[103] & in2[103];
    assign P[57] = in[103] ^ in2[103];
    assign G[58] = in[102] & in2[102];
    assign P[58] = in[102] ^ in2[102];
    assign G[59] = in[101] & in2[101];
    assign P[59] = in[101] ^ in2[101];
    assign G[60] = in[100] & in2[100];
    assign P[60] = in[100] ^ in2[100];
    assign G[61] = in[99] & in2[99];
    assign P[61] = in[99] ^ in2[99];
    assign G[62] = in[98] & in2[98];
    assign P[62] = in[98] ^ in2[98];
    assign G[63] = in[97] & in2[97];
    assign P[63] = in[97] ^ in2[97];
    assign G[64] = in[96] & in2[96];
    assign P[64] = in[96] ^ in2[96];
    assign G[65] = in[95] & in2[95];
    assign P[65] = in[95] ^ in2[95];
    assign G[66] = in[94] & in2[94];
    assign P[66] = in[94] ^ in2[94];
    assign G[67] = in[93] & in2[93];
    assign P[67] = in[93] ^ in2[93];
    assign G[68] = in[92] & in2[92];
    assign P[68] = in[92] ^ in2[92];
    assign G[69] = in[91] & in2[91];
    assign P[69] = in[91] ^ in2[91];
    assign G[70] = in[90] & in2[90];
    assign P[70] = in[90] ^ in2[90];
    assign G[71] = in[89] & in2[89];
    assign P[71] = in[89] ^ in2[89];
    assign G[72] = in[88] & in2[88];
    assign P[72] = in[88] ^ in2[88];
    assign G[73] = in[87] & in2[87];
    assign P[73] = in[87] ^ in2[87];
    assign G[74] = in[86] & in2[86];
    assign P[74] = in[86] ^ in2[86];
    assign G[75] = in[85] & in2[85];
    assign P[75] = in[85] ^ in2[85];
    assign G[76] = in[84] & in2[84];
    assign P[76] = in[84] ^ in2[84];
    assign G[77] = in[83] & in2[83];
    assign P[77] = in[83] ^ in2[83];
    assign G[78] = in[82] & in2[82];
    assign P[78] = in[82] ^ in2[82];
    assign G[79] = in[81] & in2[81];
    assign P[79] = in[81] ^ in2[81];
    assign G[80] = in[80] & in2[80];
    assign P[80] = in[80] ^ in2[80];
    assign G[81] = in[79] & in2[79];
    assign P[81] = in[79] ^ in2[79];
    assign G[82] = in[78] & in2[78];
    assign P[82] = in[78] ^ in2[78];
    assign G[83] = in[77] & in2[77];
    assign P[83] = in[77] ^ in2[77];
    assign G[84] = in[76] & in2[76];
    assign P[84] = in[76] ^ in2[76];
    assign G[85] = in[75] & in2[75];
    assign P[85] = in[75] ^ in2[75];
    assign G[86] = in[74] & in2[74];
    assign P[86] = in[74] ^ in2[74];
    assign G[87] = in[73] & in2[73];
    assign P[87] = in[73] ^ in2[73];
    assign G[88] = in[72] & in2[72];
    assign P[88] = in[72] ^ in2[72];
    assign G[89] = in[71] & in2[71];
    assign P[89] = in[71] ^ in2[71];
    assign G[90] = in[70] & in2[70];
    assign P[90] = in[70] ^ in2[70];
    assign G[91] = in[69] & in2[69];
    assign P[91] = in[69] ^ in2[69];
    assign G[92] = in[68] & in2[68];
    assign P[92] = in[68] ^ in2[68];
    assign G[93] = in[67] & in2[67];
    assign P[93] = in[67] ^ in2[67];
    assign G[94] = in[66] & in2[66];
    assign P[94] = in[66] ^ in2[66];
    assign G[95] = in[65] & in2[65];
    assign P[95] = in[65] ^ in2[65];
    assign G[96] = in[64] & in2[64];
    assign P[96] = in[64] ^ in2[64];
    assign G[97] = in[63] & in2[63];
    assign P[97] = in[63] ^ in2[63];
    assign G[98] = in[62] & in2[62];
    assign P[98] = in[62] ^ in2[62];
    assign G[99] = in[61] & in2[61];
    assign P[99] = in[61] ^ in2[61];
    assign G[100] = in[60] & in2[60];
    assign P[100] = in[60] ^ in2[60];
    assign G[101] = in[59] & in2[59];
    assign P[101] = in[59] ^ in2[59];
    assign G[102] = in[58] & in2[58];
    assign P[102] = in[58] ^ in2[58];
    assign G[103] = in[57] & in2[57];
    assign P[103] = in[57] ^ in2[57];
    assign G[104] = in[56] & in2[56];
    assign P[104] = in[56] ^ in2[56];
    assign G[105] = in[55] & in2[55];
    assign P[105] = in[55] ^ in2[55];
    assign G[106] = in[54] & in2[54];
    assign P[106] = in[54] ^ in2[54];
    assign G[107] = in[53] & in2[53];
    assign P[107] = in[53] ^ in2[53];
    assign G[108] = in[52] & in2[52];
    assign P[108] = in[52] ^ in2[52];
    assign G[109] = in[51] & in2[51];
    assign P[109] = in[51] ^ in2[51];
    assign G[110] = in[50] & in2[50];
    assign P[110] = in[50] ^ in2[50];
    assign G[111] = in[49] & in2[49];
    assign P[111] = in[49] ^ in2[49];
    assign G[112] = in[48] & in2[48];
    assign P[112] = in[48] ^ in2[48];
    assign G[113] = in[47] & in2[47];
    assign P[113] = in[47] ^ in2[47];
    assign G[114] = in[46] & in2[46];
    assign P[114] = in[46] ^ in2[46];
    assign G[115] = in[45] & in2[45];
    assign P[115] = in[45] ^ in2[45];
    assign G[116] = in[44] & in2[44];
    assign P[116] = in[44] ^ in2[44];
    assign G[117] = in[43] & in2[43];
    assign P[117] = in[43] ^ in2[43];
    assign G[118] = in[42] & in2[42];
    assign P[118] = in[42] ^ in2[42];
    assign G[119] = in[41] & in2[41];
    assign P[119] = in[41] ^ in2[41];
    assign G[120] = in[40] & in2[40];
    assign P[120] = in[40] ^ in2[40];
    assign G[121] = in[39] & in2[39];
    assign P[121] = in[39] ^ in2[39];
    assign G[122] = in[38] & in2[38];
    assign P[122] = in[38] ^ in2[38];
    assign G[123] = in[37] & in2[37];
    assign P[123] = in[37] ^ in2[37];
    assign G[124] = in[36] & in2[36];
    assign P[124] = in[36] ^ in2[36];
    assign G[125] = in[35] & in2[35];
    assign P[125] = in[35] ^ in2[35];
    assign G[126] = in[34] & in2[34];
    assign P[126] = in[34] ^ in2[34];
    assign G[127] = in[33] & in2[33];
    assign P[127] = in[33] ^ in2[33];
    assign G[128] = in[32] & in2[32];
    assign P[128] = in[32] ^ in2[32];
    assign G[129] = in[31] & in2[31];
    assign P[129] = in[31] ^ in2[31];
    assign G[130] = in[30] & in2[30];
    assign P[130] = in[30] ^ in2[30];
    assign G[131] = in[29] & in2[29];
    assign P[131] = in[29] ^ in2[29];
    assign G[132] = in[28] & in2[28];
    assign P[132] = in[28] ^ in2[28];
    assign G[133] = in[27] & in2[27];
    assign P[133] = in[27] ^ in2[27];
    assign G[134] = in[26] & in2[26];
    assign P[134] = in[26] ^ in2[26];
    assign G[135] = in[25] & in2[25];
    assign P[135] = in[25] ^ in2[25];
    assign G[136] = in[24] & in2[24];
    assign P[136] = in[24] ^ in2[24];
    assign G[137] = in[23] & in2[23];
    assign P[137] = in[23] ^ in2[23];
    assign G[138] = in[22] & in2[22];
    assign P[138] = in[22] ^ in2[22];
    assign G[139] = in[21] & in2[21];
    assign P[139] = in[21] ^ in2[21];
    assign G[140] = in[20] & in2[20];
    assign P[140] = in[20] ^ in2[20];
    assign G[141] = in[19] & in2[19];
    assign P[141] = in[19] ^ in2[19];
    assign G[142] = in[18] & in2[18];
    assign P[142] = in[18] ^ in2[18];
    assign G[143] = in[17] & in2[17];
    assign P[143] = in[17] ^ in2[17];
    assign G[144] = in[16] & in2[16];
    assign P[144] = in[16] ^ in2[16];
    assign G[145] = in[15] & in2[15];
    assign P[145] = in[15] ^ in2[15];
    assign G[146] = in[14] & in2[14];
    assign P[146] = in[14] ^ in2[14];
    assign G[147] = in[13] & in2[13];
    assign P[147] = in[13] ^ in2[13];
    assign G[148] = in[12] & in2[12];
    assign P[148] = in[12] ^ in2[12];
    assign G[149] = in[11] & in2[11];
    assign P[149] = in[11] ^ in2[11];
    assign G[150] = in[10] & in2[10];
    assign P[150] = in[10] ^ in2[10];
    assign G[151] = in[9] & in2[9];
    assign P[151] = in[9] ^ in2[9];
    assign G[152] = in[8] & in2[8];
    assign P[152] = in[8] ^ in2[8];
    assign G[153] = in[7] & in2[7];
    assign P[153] = in[7] ^ in2[7];
    assign G[154] = in[6] & in2[6];
    assign P[154] = in[6] ^ in2[6];
    assign G[155] = in[5] & in2[5];
    assign P[155] = in[5] ^ in2[5];
    assign G[156] = in[4] & in2[4];
    assign P[156] = in[4] ^ in2[4];
    assign G[157] = in[3] & in2[3];
    assign P[157] = in[3] ^ in2[3];
    assign G[158] = in[2] & in2[2];
    assign P[158] = in[2] ^ in2[2];
    assign G[159] = in[1] & in2[1];
    assign P[159] = in[1] ^ in2[1];
    assign G[160] = in[0] & in2[0];
    assign P[160] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign C[160] = G[159] | (P[159] & C[159]);
    assign cout = G[160] | (P[160] & C[160]);
    assign sum = P ^ C;
endmodule

module CLA160(output [159:0] sum, output cout, input [159:0] in1, input [159:0] in2;

    wire[159:0] G;
    wire[159:0] C;
    wire[159:0] P;

    assign G[0] = in[159] & in2[159];
    assign P[0] = in[159] ^ in2[159];
    assign G[1] = in[158] & in2[158];
    assign P[1] = in[158] ^ in2[158];
    assign G[2] = in[157] & in2[157];
    assign P[2] = in[157] ^ in2[157];
    assign G[3] = in[156] & in2[156];
    assign P[3] = in[156] ^ in2[156];
    assign G[4] = in[155] & in2[155];
    assign P[4] = in[155] ^ in2[155];
    assign G[5] = in[154] & in2[154];
    assign P[5] = in[154] ^ in2[154];
    assign G[6] = in[153] & in2[153];
    assign P[6] = in[153] ^ in2[153];
    assign G[7] = in[152] & in2[152];
    assign P[7] = in[152] ^ in2[152];
    assign G[8] = in[151] & in2[151];
    assign P[8] = in[151] ^ in2[151];
    assign G[9] = in[150] & in2[150];
    assign P[9] = in[150] ^ in2[150];
    assign G[10] = in[149] & in2[149];
    assign P[10] = in[149] ^ in2[149];
    assign G[11] = in[148] & in2[148];
    assign P[11] = in[148] ^ in2[148];
    assign G[12] = in[147] & in2[147];
    assign P[12] = in[147] ^ in2[147];
    assign G[13] = in[146] & in2[146];
    assign P[13] = in[146] ^ in2[146];
    assign G[14] = in[145] & in2[145];
    assign P[14] = in[145] ^ in2[145];
    assign G[15] = in[144] & in2[144];
    assign P[15] = in[144] ^ in2[144];
    assign G[16] = in[143] & in2[143];
    assign P[16] = in[143] ^ in2[143];
    assign G[17] = in[142] & in2[142];
    assign P[17] = in[142] ^ in2[142];
    assign G[18] = in[141] & in2[141];
    assign P[18] = in[141] ^ in2[141];
    assign G[19] = in[140] & in2[140];
    assign P[19] = in[140] ^ in2[140];
    assign G[20] = in[139] & in2[139];
    assign P[20] = in[139] ^ in2[139];
    assign G[21] = in[138] & in2[138];
    assign P[21] = in[138] ^ in2[138];
    assign G[22] = in[137] & in2[137];
    assign P[22] = in[137] ^ in2[137];
    assign G[23] = in[136] & in2[136];
    assign P[23] = in[136] ^ in2[136];
    assign G[24] = in[135] & in2[135];
    assign P[24] = in[135] ^ in2[135];
    assign G[25] = in[134] & in2[134];
    assign P[25] = in[134] ^ in2[134];
    assign G[26] = in[133] & in2[133];
    assign P[26] = in[133] ^ in2[133];
    assign G[27] = in[132] & in2[132];
    assign P[27] = in[132] ^ in2[132];
    assign G[28] = in[131] & in2[131];
    assign P[28] = in[131] ^ in2[131];
    assign G[29] = in[130] & in2[130];
    assign P[29] = in[130] ^ in2[130];
    assign G[30] = in[129] & in2[129];
    assign P[30] = in[129] ^ in2[129];
    assign G[31] = in[128] & in2[128];
    assign P[31] = in[128] ^ in2[128];
    assign G[32] = in[127] & in2[127];
    assign P[32] = in[127] ^ in2[127];
    assign G[33] = in[126] & in2[126];
    assign P[33] = in[126] ^ in2[126];
    assign G[34] = in[125] & in2[125];
    assign P[34] = in[125] ^ in2[125];
    assign G[35] = in[124] & in2[124];
    assign P[35] = in[124] ^ in2[124];
    assign G[36] = in[123] & in2[123];
    assign P[36] = in[123] ^ in2[123];
    assign G[37] = in[122] & in2[122];
    assign P[37] = in[122] ^ in2[122];
    assign G[38] = in[121] & in2[121];
    assign P[38] = in[121] ^ in2[121];
    assign G[39] = in[120] & in2[120];
    assign P[39] = in[120] ^ in2[120];
    assign G[40] = in[119] & in2[119];
    assign P[40] = in[119] ^ in2[119];
    assign G[41] = in[118] & in2[118];
    assign P[41] = in[118] ^ in2[118];
    assign G[42] = in[117] & in2[117];
    assign P[42] = in[117] ^ in2[117];
    assign G[43] = in[116] & in2[116];
    assign P[43] = in[116] ^ in2[116];
    assign G[44] = in[115] & in2[115];
    assign P[44] = in[115] ^ in2[115];
    assign G[45] = in[114] & in2[114];
    assign P[45] = in[114] ^ in2[114];
    assign G[46] = in[113] & in2[113];
    assign P[46] = in[113] ^ in2[113];
    assign G[47] = in[112] & in2[112];
    assign P[47] = in[112] ^ in2[112];
    assign G[48] = in[111] & in2[111];
    assign P[48] = in[111] ^ in2[111];
    assign G[49] = in[110] & in2[110];
    assign P[49] = in[110] ^ in2[110];
    assign G[50] = in[109] & in2[109];
    assign P[50] = in[109] ^ in2[109];
    assign G[51] = in[108] & in2[108];
    assign P[51] = in[108] ^ in2[108];
    assign G[52] = in[107] & in2[107];
    assign P[52] = in[107] ^ in2[107];
    assign G[53] = in[106] & in2[106];
    assign P[53] = in[106] ^ in2[106];
    assign G[54] = in[105] & in2[105];
    assign P[54] = in[105] ^ in2[105];
    assign G[55] = in[104] & in2[104];
    assign P[55] = in[104] ^ in2[104];
    assign G[56] = in[103] & in2[103];
    assign P[56] = in[103] ^ in2[103];
    assign G[57] = in[102] & in2[102];
    assign P[57] = in[102] ^ in2[102];
    assign G[58] = in[101] & in2[101];
    assign P[58] = in[101] ^ in2[101];
    assign G[59] = in[100] & in2[100];
    assign P[59] = in[100] ^ in2[100];
    assign G[60] = in[99] & in2[99];
    assign P[60] = in[99] ^ in2[99];
    assign G[61] = in[98] & in2[98];
    assign P[61] = in[98] ^ in2[98];
    assign G[62] = in[97] & in2[97];
    assign P[62] = in[97] ^ in2[97];
    assign G[63] = in[96] & in2[96];
    assign P[63] = in[96] ^ in2[96];
    assign G[64] = in[95] & in2[95];
    assign P[64] = in[95] ^ in2[95];
    assign G[65] = in[94] & in2[94];
    assign P[65] = in[94] ^ in2[94];
    assign G[66] = in[93] & in2[93];
    assign P[66] = in[93] ^ in2[93];
    assign G[67] = in[92] & in2[92];
    assign P[67] = in[92] ^ in2[92];
    assign G[68] = in[91] & in2[91];
    assign P[68] = in[91] ^ in2[91];
    assign G[69] = in[90] & in2[90];
    assign P[69] = in[90] ^ in2[90];
    assign G[70] = in[89] & in2[89];
    assign P[70] = in[89] ^ in2[89];
    assign G[71] = in[88] & in2[88];
    assign P[71] = in[88] ^ in2[88];
    assign G[72] = in[87] & in2[87];
    assign P[72] = in[87] ^ in2[87];
    assign G[73] = in[86] & in2[86];
    assign P[73] = in[86] ^ in2[86];
    assign G[74] = in[85] & in2[85];
    assign P[74] = in[85] ^ in2[85];
    assign G[75] = in[84] & in2[84];
    assign P[75] = in[84] ^ in2[84];
    assign G[76] = in[83] & in2[83];
    assign P[76] = in[83] ^ in2[83];
    assign G[77] = in[82] & in2[82];
    assign P[77] = in[82] ^ in2[82];
    assign G[78] = in[81] & in2[81];
    assign P[78] = in[81] ^ in2[81];
    assign G[79] = in[80] & in2[80];
    assign P[79] = in[80] ^ in2[80];
    assign G[80] = in[79] & in2[79];
    assign P[80] = in[79] ^ in2[79];
    assign G[81] = in[78] & in2[78];
    assign P[81] = in[78] ^ in2[78];
    assign G[82] = in[77] & in2[77];
    assign P[82] = in[77] ^ in2[77];
    assign G[83] = in[76] & in2[76];
    assign P[83] = in[76] ^ in2[76];
    assign G[84] = in[75] & in2[75];
    assign P[84] = in[75] ^ in2[75];
    assign G[85] = in[74] & in2[74];
    assign P[85] = in[74] ^ in2[74];
    assign G[86] = in[73] & in2[73];
    assign P[86] = in[73] ^ in2[73];
    assign G[87] = in[72] & in2[72];
    assign P[87] = in[72] ^ in2[72];
    assign G[88] = in[71] & in2[71];
    assign P[88] = in[71] ^ in2[71];
    assign G[89] = in[70] & in2[70];
    assign P[89] = in[70] ^ in2[70];
    assign G[90] = in[69] & in2[69];
    assign P[90] = in[69] ^ in2[69];
    assign G[91] = in[68] & in2[68];
    assign P[91] = in[68] ^ in2[68];
    assign G[92] = in[67] & in2[67];
    assign P[92] = in[67] ^ in2[67];
    assign G[93] = in[66] & in2[66];
    assign P[93] = in[66] ^ in2[66];
    assign G[94] = in[65] & in2[65];
    assign P[94] = in[65] ^ in2[65];
    assign G[95] = in[64] & in2[64];
    assign P[95] = in[64] ^ in2[64];
    assign G[96] = in[63] & in2[63];
    assign P[96] = in[63] ^ in2[63];
    assign G[97] = in[62] & in2[62];
    assign P[97] = in[62] ^ in2[62];
    assign G[98] = in[61] & in2[61];
    assign P[98] = in[61] ^ in2[61];
    assign G[99] = in[60] & in2[60];
    assign P[99] = in[60] ^ in2[60];
    assign G[100] = in[59] & in2[59];
    assign P[100] = in[59] ^ in2[59];
    assign G[101] = in[58] & in2[58];
    assign P[101] = in[58] ^ in2[58];
    assign G[102] = in[57] & in2[57];
    assign P[102] = in[57] ^ in2[57];
    assign G[103] = in[56] & in2[56];
    assign P[103] = in[56] ^ in2[56];
    assign G[104] = in[55] & in2[55];
    assign P[104] = in[55] ^ in2[55];
    assign G[105] = in[54] & in2[54];
    assign P[105] = in[54] ^ in2[54];
    assign G[106] = in[53] & in2[53];
    assign P[106] = in[53] ^ in2[53];
    assign G[107] = in[52] & in2[52];
    assign P[107] = in[52] ^ in2[52];
    assign G[108] = in[51] & in2[51];
    assign P[108] = in[51] ^ in2[51];
    assign G[109] = in[50] & in2[50];
    assign P[109] = in[50] ^ in2[50];
    assign G[110] = in[49] & in2[49];
    assign P[110] = in[49] ^ in2[49];
    assign G[111] = in[48] & in2[48];
    assign P[111] = in[48] ^ in2[48];
    assign G[112] = in[47] & in2[47];
    assign P[112] = in[47] ^ in2[47];
    assign G[113] = in[46] & in2[46];
    assign P[113] = in[46] ^ in2[46];
    assign G[114] = in[45] & in2[45];
    assign P[114] = in[45] ^ in2[45];
    assign G[115] = in[44] & in2[44];
    assign P[115] = in[44] ^ in2[44];
    assign G[116] = in[43] & in2[43];
    assign P[116] = in[43] ^ in2[43];
    assign G[117] = in[42] & in2[42];
    assign P[117] = in[42] ^ in2[42];
    assign G[118] = in[41] & in2[41];
    assign P[118] = in[41] ^ in2[41];
    assign G[119] = in[40] & in2[40];
    assign P[119] = in[40] ^ in2[40];
    assign G[120] = in[39] & in2[39];
    assign P[120] = in[39] ^ in2[39];
    assign G[121] = in[38] & in2[38];
    assign P[121] = in[38] ^ in2[38];
    assign G[122] = in[37] & in2[37];
    assign P[122] = in[37] ^ in2[37];
    assign G[123] = in[36] & in2[36];
    assign P[123] = in[36] ^ in2[36];
    assign G[124] = in[35] & in2[35];
    assign P[124] = in[35] ^ in2[35];
    assign G[125] = in[34] & in2[34];
    assign P[125] = in[34] ^ in2[34];
    assign G[126] = in[33] & in2[33];
    assign P[126] = in[33] ^ in2[33];
    assign G[127] = in[32] & in2[32];
    assign P[127] = in[32] ^ in2[32];
    assign G[128] = in[31] & in2[31];
    assign P[128] = in[31] ^ in2[31];
    assign G[129] = in[30] & in2[30];
    assign P[129] = in[30] ^ in2[30];
    assign G[130] = in[29] & in2[29];
    assign P[130] = in[29] ^ in2[29];
    assign G[131] = in[28] & in2[28];
    assign P[131] = in[28] ^ in2[28];
    assign G[132] = in[27] & in2[27];
    assign P[132] = in[27] ^ in2[27];
    assign G[133] = in[26] & in2[26];
    assign P[133] = in[26] ^ in2[26];
    assign G[134] = in[25] & in2[25];
    assign P[134] = in[25] ^ in2[25];
    assign G[135] = in[24] & in2[24];
    assign P[135] = in[24] ^ in2[24];
    assign G[136] = in[23] & in2[23];
    assign P[136] = in[23] ^ in2[23];
    assign G[137] = in[22] & in2[22];
    assign P[137] = in[22] ^ in2[22];
    assign G[138] = in[21] & in2[21];
    assign P[138] = in[21] ^ in2[21];
    assign G[139] = in[20] & in2[20];
    assign P[139] = in[20] ^ in2[20];
    assign G[140] = in[19] & in2[19];
    assign P[140] = in[19] ^ in2[19];
    assign G[141] = in[18] & in2[18];
    assign P[141] = in[18] ^ in2[18];
    assign G[142] = in[17] & in2[17];
    assign P[142] = in[17] ^ in2[17];
    assign G[143] = in[16] & in2[16];
    assign P[143] = in[16] ^ in2[16];
    assign G[144] = in[15] & in2[15];
    assign P[144] = in[15] ^ in2[15];
    assign G[145] = in[14] & in2[14];
    assign P[145] = in[14] ^ in2[14];
    assign G[146] = in[13] & in2[13];
    assign P[146] = in[13] ^ in2[13];
    assign G[147] = in[12] & in2[12];
    assign P[147] = in[12] ^ in2[12];
    assign G[148] = in[11] & in2[11];
    assign P[148] = in[11] ^ in2[11];
    assign G[149] = in[10] & in2[10];
    assign P[149] = in[10] ^ in2[10];
    assign G[150] = in[9] & in2[9];
    assign P[150] = in[9] ^ in2[9];
    assign G[151] = in[8] & in2[8];
    assign P[151] = in[8] ^ in2[8];
    assign G[152] = in[7] & in2[7];
    assign P[152] = in[7] ^ in2[7];
    assign G[153] = in[6] & in2[6];
    assign P[153] = in[6] ^ in2[6];
    assign G[154] = in[5] & in2[5];
    assign P[154] = in[5] ^ in2[5];
    assign G[155] = in[4] & in2[4];
    assign P[155] = in[4] ^ in2[4];
    assign G[156] = in[3] & in2[3];
    assign P[156] = in[3] ^ in2[3];
    assign G[157] = in[2] & in2[2];
    assign P[157] = in[2] ^ in2[2];
    assign G[158] = in[1] & in2[1];
    assign P[158] = in[1] ^ in2[1];
    assign G[159] = in[0] & in2[0];
    assign P[159] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign C[159] = G[158] | (P[158] & C[158]);
    assign cout = G[159] | (P[159] & C[159]);
    assign sum = P ^ C;
endmodule

module CLA159(output [158:0] sum, output cout, input [158:0] in1, input [158:0] in2;

    wire[158:0] G;
    wire[158:0] C;
    wire[158:0] P;

    assign G[0] = in[158] & in2[158];
    assign P[0] = in[158] ^ in2[158];
    assign G[1] = in[157] & in2[157];
    assign P[1] = in[157] ^ in2[157];
    assign G[2] = in[156] & in2[156];
    assign P[2] = in[156] ^ in2[156];
    assign G[3] = in[155] & in2[155];
    assign P[3] = in[155] ^ in2[155];
    assign G[4] = in[154] & in2[154];
    assign P[4] = in[154] ^ in2[154];
    assign G[5] = in[153] & in2[153];
    assign P[5] = in[153] ^ in2[153];
    assign G[6] = in[152] & in2[152];
    assign P[6] = in[152] ^ in2[152];
    assign G[7] = in[151] & in2[151];
    assign P[7] = in[151] ^ in2[151];
    assign G[8] = in[150] & in2[150];
    assign P[8] = in[150] ^ in2[150];
    assign G[9] = in[149] & in2[149];
    assign P[9] = in[149] ^ in2[149];
    assign G[10] = in[148] & in2[148];
    assign P[10] = in[148] ^ in2[148];
    assign G[11] = in[147] & in2[147];
    assign P[11] = in[147] ^ in2[147];
    assign G[12] = in[146] & in2[146];
    assign P[12] = in[146] ^ in2[146];
    assign G[13] = in[145] & in2[145];
    assign P[13] = in[145] ^ in2[145];
    assign G[14] = in[144] & in2[144];
    assign P[14] = in[144] ^ in2[144];
    assign G[15] = in[143] & in2[143];
    assign P[15] = in[143] ^ in2[143];
    assign G[16] = in[142] & in2[142];
    assign P[16] = in[142] ^ in2[142];
    assign G[17] = in[141] & in2[141];
    assign P[17] = in[141] ^ in2[141];
    assign G[18] = in[140] & in2[140];
    assign P[18] = in[140] ^ in2[140];
    assign G[19] = in[139] & in2[139];
    assign P[19] = in[139] ^ in2[139];
    assign G[20] = in[138] & in2[138];
    assign P[20] = in[138] ^ in2[138];
    assign G[21] = in[137] & in2[137];
    assign P[21] = in[137] ^ in2[137];
    assign G[22] = in[136] & in2[136];
    assign P[22] = in[136] ^ in2[136];
    assign G[23] = in[135] & in2[135];
    assign P[23] = in[135] ^ in2[135];
    assign G[24] = in[134] & in2[134];
    assign P[24] = in[134] ^ in2[134];
    assign G[25] = in[133] & in2[133];
    assign P[25] = in[133] ^ in2[133];
    assign G[26] = in[132] & in2[132];
    assign P[26] = in[132] ^ in2[132];
    assign G[27] = in[131] & in2[131];
    assign P[27] = in[131] ^ in2[131];
    assign G[28] = in[130] & in2[130];
    assign P[28] = in[130] ^ in2[130];
    assign G[29] = in[129] & in2[129];
    assign P[29] = in[129] ^ in2[129];
    assign G[30] = in[128] & in2[128];
    assign P[30] = in[128] ^ in2[128];
    assign G[31] = in[127] & in2[127];
    assign P[31] = in[127] ^ in2[127];
    assign G[32] = in[126] & in2[126];
    assign P[32] = in[126] ^ in2[126];
    assign G[33] = in[125] & in2[125];
    assign P[33] = in[125] ^ in2[125];
    assign G[34] = in[124] & in2[124];
    assign P[34] = in[124] ^ in2[124];
    assign G[35] = in[123] & in2[123];
    assign P[35] = in[123] ^ in2[123];
    assign G[36] = in[122] & in2[122];
    assign P[36] = in[122] ^ in2[122];
    assign G[37] = in[121] & in2[121];
    assign P[37] = in[121] ^ in2[121];
    assign G[38] = in[120] & in2[120];
    assign P[38] = in[120] ^ in2[120];
    assign G[39] = in[119] & in2[119];
    assign P[39] = in[119] ^ in2[119];
    assign G[40] = in[118] & in2[118];
    assign P[40] = in[118] ^ in2[118];
    assign G[41] = in[117] & in2[117];
    assign P[41] = in[117] ^ in2[117];
    assign G[42] = in[116] & in2[116];
    assign P[42] = in[116] ^ in2[116];
    assign G[43] = in[115] & in2[115];
    assign P[43] = in[115] ^ in2[115];
    assign G[44] = in[114] & in2[114];
    assign P[44] = in[114] ^ in2[114];
    assign G[45] = in[113] & in2[113];
    assign P[45] = in[113] ^ in2[113];
    assign G[46] = in[112] & in2[112];
    assign P[46] = in[112] ^ in2[112];
    assign G[47] = in[111] & in2[111];
    assign P[47] = in[111] ^ in2[111];
    assign G[48] = in[110] & in2[110];
    assign P[48] = in[110] ^ in2[110];
    assign G[49] = in[109] & in2[109];
    assign P[49] = in[109] ^ in2[109];
    assign G[50] = in[108] & in2[108];
    assign P[50] = in[108] ^ in2[108];
    assign G[51] = in[107] & in2[107];
    assign P[51] = in[107] ^ in2[107];
    assign G[52] = in[106] & in2[106];
    assign P[52] = in[106] ^ in2[106];
    assign G[53] = in[105] & in2[105];
    assign P[53] = in[105] ^ in2[105];
    assign G[54] = in[104] & in2[104];
    assign P[54] = in[104] ^ in2[104];
    assign G[55] = in[103] & in2[103];
    assign P[55] = in[103] ^ in2[103];
    assign G[56] = in[102] & in2[102];
    assign P[56] = in[102] ^ in2[102];
    assign G[57] = in[101] & in2[101];
    assign P[57] = in[101] ^ in2[101];
    assign G[58] = in[100] & in2[100];
    assign P[58] = in[100] ^ in2[100];
    assign G[59] = in[99] & in2[99];
    assign P[59] = in[99] ^ in2[99];
    assign G[60] = in[98] & in2[98];
    assign P[60] = in[98] ^ in2[98];
    assign G[61] = in[97] & in2[97];
    assign P[61] = in[97] ^ in2[97];
    assign G[62] = in[96] & in2[96];
    assign P[62] = in[96] ^ in2[96];
    assign G[63] = in[95] & in2[95];
    assign P[63] = in[95] ^ in2[95];
    assign G[64] = in[94] & in2[94];
    assign P[64] = in[94] ^ in2[94];
    assign G[65] = in[93] & in2[93];
    assign P[65] = in[93] ^ in2[93];
    assign G[66] = in[92] & in2[92];
    assign P[66] = in[92] ^ in2[92];
    assign G[67] = in[91] & in2[91];
    assign P[67] = in[91] ^ in2[91];
    assign G[68] = in[90] & in2[90];
    assign P[68] = in[90] ^ in2[90];
    assign G[69] = in[89] & in2[89];
    assign P[69] = in[89] ^ in2[89];
    assign G[70] = in[88] & in2[88];
    assign P[70] = in[88] ^ in2[88];
    assign G[71] = in[87] & in2[87];
    assign P[71] = in[87] ^ in2[87];
    assign G[72] = in[86] & in2[86];
    assign P[72] = in[86] ^ in2[86];
    assign G[73] = in[85] & in2[85];
    assign P[73] = in[85] ^ in2[85];
    assign G[74] = in[84] & in2[84];
    assign P[74] = in[84] ^ in2[84];
    assign G[75] = in[83] & in2[83];
    assign P[75] = in[83] ^ in2[83];
    assign G[76] = in[82] & in2[82];
    assign P[76] = in[82] ^ in2[82];
    assign G[77] = in[81] & in2[81];
    assign P[77] = in[81] ^ in2[81];
    assign G[78] = in[80] & in2[80];
    assign P[78] = in[80] ^ in2[80];
    assign G[79] = in[79] & in2[79];
    assign P[79] = in[79] ^ in2[79];
    assign G[80] = in[78] & in2[78];
    assign P[80] = in[78] ^ in2[78];
    assign G[81] = in[77] & in2[77];
    assign P[81] = in[77] ^ in2[77];
    assign G[82] = in[76] & in2[76];
    assign P[82] = in[76] ^ in2[76];
    assign G[83] = in[75] & in2[75];
    assign P[83] = in[75] ^ in2[75];
    assign G[84] = in[74] & in2[74];
    assign P[84] = in[74] ^ in2[74];
    assign G[85] = in[73] & in2[73];
    assign P[85] = in[73] ^ in2[73];
    assign G[86] = in[72] & in2[72];
    assign P[86] = in[72] ^ in2[72];
    assign G[87] = in[71] & in2[71];
    assign P[87] = in[71] ^ in2[71];
    assign G[88] = in[70] & in2[70];
    assign P[88] = in[70] ^ in2[70];
    assign G[89] = in[69] & in2[69];
    assign P[89] = in[69] ^ in2[69];
    assign G[90] = in[68] & in2[68];
    assign P[90] = in[68] ^ in2[68];
    assign G[91] = in[67] & in2[67];
    assign P[91] = in[67] ^ in2[67];
    assign G[92] = in[66] & in2[66];
    assign P[92] = in[66] ^ in2[66];
    assign G[93] = in[65] & in2[65];
    assign P[93] = in[65] ^ in2[65];
    assign G[94] = in[64] & in2[64];
    assign P[94] = in[64] ^ in2[64];
    assign G[95] = in[63] & in2[63];
    assign P[95] = in[63] ^ in2[63];
    assign G[96] = in[62] & in2[62];
    assign P[96] = in[62] ^ in2[62];
    assign G[97] = in[61] & in2[61];
    assign P[97] = in[61] ^ in2[61];
    assign G[98] = in[60] & in2[60];
    assign P[98] = in[60] ^ in2[60];
    assign G[99] = in[59] & in2[59];
    assign P[99] = in[59] ^ in2[59];
    assign G[100] = in[58] & in2[58];
    assign P[100] = in[58] ^ in2[58];
    assign G[101] = in[57] & in2[57];
    assign P[101] = in[57] ^ in2[57];
    assign G[102] = in[56] & in2[56];
    assign P[102] = in[56] ^ in2[56];
    assign G[103] = in[55] & in2[55];
    assign P[103] = in[55] ^ in2[55];
    assign G[104] = in[54] & in2[54];
    assign P[104] = in[54] ^ in2[54];
    assign G[105] = in[53] & in2[53];
    assign P[105] = in[53] ^ in2[53];
    assign G[106] = in[52] & in2[52];
    assign P[106] = in[52] ^ in2[52];
    assign G[107] = in[51] & in2[51];
    assign P[107] = in[51] ^ in2[51];
    assign G[108] = in[50] & in2[50];
    assign P[108] = in[50] ^ in2[50];
    assign G[109] = in[49] & in2[49];
    assign P[109] = in[49] ^ in2[49];
    assign G[110] = in[48] & in2[48];
    assign P[110] = in[48] ^ in2[48];
    assign G[111] = in[47] & in2[47];
    assign P[111] = in[47] ^ in2[47];
    assign G[112] = in[46] & in2[46];
    assign P[112] = in[46] ^ in2[46];
    assign G[113] = in[45] & in2[45];
    assign P[113] = in[45] ^ in2[45];
    assign G[114] = in[44] & in2[44];
    assign P[114] = in[44] ^ in2[44];
    assign G[115] = in[43] & in2[43];
    assign P[115] = in[43] ^ in2[43];
    assign G[116] = in[42] & in2[42];
    assign P[116] = in[42] ^ in2[42];
    assign G[117] = in[41] & in2[41];
    assign P[117] = in[41] ^ in2[41];
    assign G[118] = in[40] & in2[40];
    assign P[118] = in[40] ^ in2[40];
    assign G[119] = in[39] & in2[39];
    assign P[119] = in[39] ^ in2[39];
    assign G[120] = in[38] & in2[38];
    assign P[120] = in[38] ^ in2[38];
    assign G[121] = in[37] & in2[37];
    assign P[121] = in[37] ^ in2[37];
    assign G[122] = in[36] & in2[36];
    assign P[122] = in[36] ^ in2[36];
    assign G[123] = in[35] & in2[35];
    assign P[123] = in[35] ^ in2[35];
    assign G[124] = in[34] & in2[34];
    assign P[124] = in[34] ^ in2[34];
    assign G[125] = in[33] & in2[33];
    assign P[125] = in[33] ^ in2[33];
    assign G[126] = in[32] & in2[32];
    assign P[126] = in[32] ^ in2[32];
    assign G[127] = in[31] & in2[31];
    assign P[127] = in[31] ^ in2[31];
    assign G[128] = in[30] & in2[30];
    assign P[128] = in[30] ^ in2[30];
    assign G[129] = in[29] & in2[29];
    assign P[129] = in[29] ^ in2[29];
    assign G[130] = in[28] & in2[28];
    assign P[130] = in[28] ^ in2[28];
    assign G[131] = in[27] & in2[27];
    assign P[131] = in[27] ^ in2[27];
    assign G[132] = in[26] & in2[26];
    assign P[132] = in[26] ^ in2[26];
    assign G[133] = in[25] & in2[25];
    assign P[133] = in[25] ^ in2[25];
    assign G[134] = in[24] & in2[24];
    assign P[134] = in[24] ^ in2[24];
    assign G[135] = in[23] & in2[23];
    assign P[135] = in[23] ^ in2[23];
    assign G[136] = in[22] & in2[22];
    assign P[136] = in[22] ^ in2[22];
    assign G[137] = in[21] & in2[21];
    assign P[137] = in[21] ^ in2[21];
    assign G[138] = in[20] & in2[20];
    assign P[138] = in[20] ^ in2[20];
    assign G[139] = in[19] & in2[19];
    assign P[139] = in[19] ^ in2[19];
    assign G[140] = in[18] & in2[18];
    assign P[140] = in[18] ^ in2[18];
    assign G[141] = in[17] & in2[17];
    assign P[141] = in[17] ^ in2[17];
    assign G[142] = in[16] & in2[16];
    assign P[142] = in[16] ^ in2[16];
    assign G[143] = in[15] & in2[15];
    assign P[143] = in[15] ^ in2[15];
    assign G[144] = in[14] & in2[14];
    assign P[144] = in[14] ^ in2[14];
    assign G[145] = in[13] & in2[13];
    assign P[145] = in[13] ^ in2[13];
    assign G[146] = in[12] & in2[12];
    assign P[146] = in[12] ^ in2[12];
    assign G[147] = in[11] & in2[11];
    assign P[147] = in[11] ^ in2[11];
    assign G[148] = in[10] & in2[10];
    assign P[148] = in[10] ^ in2[10];
    assign G[149] = in[9] & in2[9];
    assign P[149] = in[9] ^ in2[9];
    assign G[150] = in[8] & in2[8];
    assign P[150] = in[8] ^ in2[8];
    assign G[151] = in[7] & in2[7];
    assign P[151] = in[7] ^ in2[7];
    assign G[152] = in[6] & in2[6];
    assign P[152] = in[6] ^ in2[6];
    assign G[153] = in[5] & in2[5];
    assign P[153] = in[5] ^ in2[5];
    assign G[154] = in[4] & in2[4];
    assign P[154] = in[4] ^ in2[4];
    assign G[155] = in[3] & in2[3];
    assign P[155] = in[3] ^ in2[3];
    assign G[156] = in[2] & in2[2];
    assign P[156] = in[2] ^ in2[2];
    assign G[157] = in[1] & in2[1];
    assign P[157] = in[1] ^ in2[1];
    assign G[158] = in[0] & in2[0];
    assign P[158] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign C[158] = G[157] | (P[157] & C[157]);
    assign cout = G[158] | (P[158] & C[158]);
    assign sum = P ^ C;
endmodule

module CLA158(output [157:0] sum, output cout, input [157:0] in1, input [157:0] in2;

    wire[157:0] G;
    wire[157:0] C;
    wire[157:0] P;

    assign G[0] = in[157] & in2[157];
    assign P[0] = in[157] ^ in2[157];
    assign G[1] = in[156] & in2[156];
    assign P[1] = in[156] ^ in2[156];
    assign G[2] = in[155] & in2[155];
    assign P[2] = in[155] ^ in2[155];
    assign G[3] = in[154] & in2[154];
    assign P[3] = in[154] ^ in2[154];
    assign G[4] = in[153] & in2[153];
    assign P[4] = in[153] ^ in2[153];
    assign G[5] = in[152] & in2[152];
    assign P[5] = in[152] ^ in2[152];
    assign G[6] = in[151] & in2[151];
    assign P[6] = in[151] ^ in2[151];
    assign G[7] = in[150] & in2[150];
    assign P[7] = in[150] ^ in2[150];
    assign G[8] = in[149] & in2[149];
    assign P[8] = in[149] ^ in2[149];
    assign G[9] = in[148] & in2[148];
    assign P[9] = in[148] ^ in2[148];
    assign G[10] = in[147] & in2[147];
    assign P[10] = in[147] ^ in2[147];
    assign G[11] = in[146] & in2[146];
    assign P[11] = in[146] ^ in2[146];
    assign G[12] = in[145] & in2[145];
    assign P[12] = in[145] ^ in2[145];
    assign G[13] = in[144] & in2[144];
    assign P[13] = in[144] ^ in2[144];
    assign G[14] = in[143] & in2[143];
    assign P[14] = in[143] ^ in2[143];
    assign G[15] = in[142] & in2[142];
    assign P[15] = in[142] ^ in2[142];
    assign G[16] = in[141] & in2[141];
    assign P[16] = in[141] ^ in2[141];
    assign G[17] = in[140] & in2[140];
    assign P[17] = in[140] ^ in2[140];
    assign G[18] = in[139] & in2[139];
    assign P[18] = in[139] ^ in2[139];
    assign G[19] = in[138] & in2[138];
    assign P[19] = in[138] ^ in2[138];
    assign G[20] = in[137] & in2[137];
    assign P[20] = in[137] ^ in2[137];
    assign G[21] = in[136] & in2[136];
    assign P[21] = in[136] ^ in2[136];
    assign G[22] = in[135] & in2[135];
    assign P[22] = in[135] ^ in2[135];
    assign G[23] = in[134] & in2[134];
    assign P[23] = in[134] ^ in2[134];
    assign G[24] = in[133] & in2[133];
    assign P[24] = in[133] ^ in2[133];
    assign G[25] = in[132] & in2[132];
    assign P[25] = in[132] ^ in2[132];
    assign G[26] = in[131] & in2[131];
    assign P[26] = in[131] ^ in2[131];
    assign G[27] = in[130] & in2[130];
    assign P[27] = in[130] ^ in2[130];
    assign G[28] = in[129] & in2[129];
    assign P[28] = in[129] ^ in2[129];
    assign G[29] = in[128] & in2[128];
    assign P[29] = in[128] ^ in2[128];
    assign G[30] = in[127] & in2[127];
    assign P[30] = in[127] ^ in2[127];
    assign G[31] = in[126] & in2[126];
    assign P[31] = in[126] ^ in2[126];
    assign G[32] = in[125] & in2[125];
    assign P[32] = in[125] ^ in2[125];
    assign G[33] = in[124] & in2[124];
    assign P[33] = in[124] ^ in2[124];
    assign G[34] = in[123] & in2[123];
    assign P[34] = in[123] ^ in2[123];
    assign G[35] = in[122] & in2[122];
    assign P[35] = in[122] ^ in2[122];
    assign G[36] = in[121] & in2[121];
    assign P[36] = in[121] ^ in2[121];
    assign G[37] = in[120] & in2[120];
    assign P[37] = in[120] ^ in2[120];
    assign G[38] = in[119] & in2[119];
    assign P[38] = in[119] ^ in2[119];
    assign G[39] = in[118] & in2[118];
    assign P[39] = in[118] ^ in2[118];
    assign G[40] = in[117] & in2[117];
    assign P[40] = in[117] ^ in2[117];
    assign G[41] = in[116] & in2[116];
    assign P[41] = in[116] ^ in2[116];
    assign G[42] = in[115] & in2[115];
    assign P[42] = in[115] ^ in2[115];
    assign G[43] = in[114] & in2[114];
    assign P[43] = in[114] ^ in2[114];
    assign G[44] = in[113] & in2[113];
    assign P[44] = in[113] ^ in2[113];
    assign G[45] = in[112] & in2[112];
    assign P[45] = in[112] ^ in2[112];
    assign G[46] = in[111] & in2[111];
    assign P[46] = in[111] ^ in2[111];
    assign G[47] = in[110] & in2[110];
    assign P[47] = in[110] ^ in2[110];
    assign G[48] = in[109] & in2[109];
    assign P[48] = in[109] ^ in2[109];
    assign G[49] = in[108] & in2[108];
    assign P[49] = in[108] ^ in2[108];
    assign G[50] = in[107] & in2[107];
    assign P[50] = in[107] ^ in2[107];
    assign G[51] = in[106] & in2[106];
    assign P[51] = in[106] ^ in2[106];
    assign G[52] = in[105] & in2[105];
    assign P[52] = in[105] ^ in2[105];
    assign G[53] = in[104] & in2[104];
    assign P[53] = in[104] ^ in2[104];
    assign G[54] = in[103] & in2[103];
    assign P[54] = in[103] ^ in2[103];
    assign G[55] = in[102] & in2[102];
    assign P[55] = in[102] ^ in2[102];
    assign G[56] = in[101] & in2[101];
    assign P[56] = in[101] ^ in2[101];
    assign G[57] = in[100] & in2[100];
    assign P[57] = in[100] ^ in2[100];
    assign G[58] = in[99] & in2[99];
    assign P[58] = in[99] ^ in2[99];
    assign G[59] = in[98] & in2[98];
    assign P[59] = in[98] ^ in2[98];
    assign G[60] = in[97] & in2[97];
    assign P[60] = in[97] ^ in2[97];
    assign G[61] = in[96] & in2[96];
    assign P[61] = in[96] ^ in2[96];
    assign G[62] = in[95] & in2[95];
    assign P[62] = in[95] ^ in2[95];
    assign G[63] = in[94] & in2[94];
    assign P[63] = in[94] ^ in2[94];
    assign G[64] = in[93] & in2[93];
    assign P[64] = in[93] ^ in2[93];
    assign G[65] = in[92] & in2[92];
    assign P[65] = in[92] ^ in2[92];
    assign G[66] = in[91] & in2[91];
    assign P[66] = in[91] ^ in2[91];
    assign G[67] = in[90] & in2[90];
    assign P[67] = in[90] ^ in2[90];
    assign G[68] = in[89] & in2[89];
    assign P[68] = in[89] ^ in2[89];
    assign G[69] = in[88] & in2[88];
    assign P[69] = in[88] ^ in2[88];
    assign G[70] = in[87] & in2[87];
    assign P[70] = in[87] ^ in2[87];
    assign G[71] = in[86] & in2[86];
    assign P[71] = in[86] ^ in2[86];
    assign G[72] = in[85] & in2[85];
    assign P[72] = in[85] ^ in2[85];
    assign G[73] = in[84] & in2[84];
    assign P[73] = in[84] ^ in2[84];
    assign G[74] = in[83] & in2[83];
    assign P[74] = in[83] ^ in2[83];
    assign G[75] = in[82] & in2[82];
    assign P[75] = in[82] ^ in2[82];
    assign G[76] = in[81] & in2[81];
    assign P[76] = in[81] ^ in2[81];
    assign G[77] = in[80] & in2[80];
    assign P[77] = in[80] ^ in2[80];
    assign G[78] = in[79] & in2[79];
    assign P[78] = in[79] ^ in2[79];
    assign G[79] = in[78] & in2[78];
    assign P[79] = in[78] ^ in2[78];
    assign G[80] = in[77] & in2[77];
    assign P[80] = in[77] ^ in2[77];
    assign G[81] = in[76] & in2[76];
    assign P[81] = in[76] ^ in2[76];
    assign G[82] = in[75] & in2[75];
    assign P[82] = in[75] ^ in2[75];
    assign G[83] = in[74] & in2[74];
    assign P[83] = in[74] ^ in2[74];
    assign G[84] = in[73] & in2[73];
    assign P[84] = in[73] ^ in2[73];
    assign G[85] = in[72] & in2[72];
    assign P[85] = in[72] ^ in2[72];
    assign G[86] = in[71] & in2[71];
    assign P[86] = in[71] ^ in2[71];
    assign G[87] = in[70] & in2[70];
    assign P[87] = in[70] ^ in2[70];
    assign G[88] = in[69] & in2[69];
    assign P[88] = in[69] ^ in2[69];
    assign G[89] = in[68] & in2[68];
    assign P[89] = in[68] ^ in2[68];
    assign G[90] = in[67] & in2[67];
    assign P[90] = in[67] ^ in2[67];
    assign G[91] = in[66] & in2[66];
    assign P[91] = in[66] ^ in2[66];
    assign G[92] = in[65] & in2[65];
    assign P[92] = in[65] ^ in2[65];
    assign G[93] = in[64] & in2[64];
    assign P[93] = in[64] ^ in2[64];
    assign G[94] = in[63] & in2[63];
    assign P[94] = in[63] ^ in2[63];
    assign G[95] = in[62] & in2[62];
    assign P[95] = in[62] ^ in2[62];
    assign G[96] = in[61] & in2[61];
    assign P[96] = in[61] ^ in2[61];
    assign G[97] = in[60] & in2[60];
    assign P[97] = in[60] ^ in2[60];
    assign G[98] = in[59] & in2[59];
    assign P[98] = in[59] ^ in2[59];
    assign G[99] = in[58] & in2[58];
    assign P[99] = in[58] ^ in2[58];
    assign G[100] = in[57] & in2[57];
    assign P[100] = in[57] ^ in2[57];
    assign G[101] = in[56] & in2[56];
    assign P[101] = in[56] ^ in2[56];
    assign G[102] = in[55] & in2[55];
    assign P[102] = in[55] ^ in2[55];
    assign G[103] = in[54] & in2[54];
    assign P[103] = in[54] ^ in2[54];
    assign G[104] = in[53] & in2[53];
    assign P[104] = in[53] ^ in2[53];
    assign G[105] = in[52] & in2[52];
    assign P[105] = in[52] ^ in2[52];
    assign G[106] = in[51] & in2[51];
    assign P[106] = in[51] ^ in2[51];
    assign G[107] = in[50] & in2[50];
    assign P[107] = in[50] ^ in2[50];
    assign G[108] = in[49] & in2[49];
    assign P[108] = in[49] ^ in2[49];
    assign G[109] = in[48] & in2[48];
    assign P[109] = in[48] ^ in2[48];
    assign G[110] = in[47] & in2[47];
    assign P[110] = in[47] ^ in2[47];
    assign G[111] = in[46] & in2[46];
    assign P[111] = in[46] ^ in2[46];
    assign G[112] = in[45] & in2[45];
    assign P[112] = in[45] ^ in2[45];
    assign G[113] = in[44] & in2[44];
    assign P[113] = in[44] ^ in2[44];
    assign G[114] = in[43] & in2[43];
    assign P[114] = in[43] ^ in2[43];
    assign G[115] = in[42] & in2[42];
    assign P[115] = in[42] ^ in2[42];
    assign G[116] = in[41] & in2[41];
    assign P[116] = in[41] ^ in2[41];
    assign G[117] = in[40] & in2[40];
    assign P[117] = in[40] ^ in2[40];
    assign G[118] = in[39] & in2[39];
    assign P[118] = in[39] ^ in2[39];
    assign G[119] = in[38] & in2[38];
    assign P[119] = in[38] ^ in2[38];
    assign G[120] = in[37] & in2[37];
    assign P[120] = in[37] ^ in2[37];
    assign G[121] = in[36] & in2[36];
    assign P[121] = in[36] ^ in2[36];
    assign G[122] = in[35] & in2[35];
    assign P[122] = in[35] ^ in2[35];
    assign G[123] = in[34] & in2[34];
    assign P[123] = in[34] ^ in2[34];
    assign G[124] = in[33] & in2[33];
    assign P[124] = in[33] ^ in2[33];
    assign G[125] = in[32] & in2[32];
    assign P[125] = in[32] ^ in2[32];
    assign G[126] = in[31] & in2[31];
    assign P[126] = in[31] ^ in2[31];
    assign G[127] = in[30] & in2[30];
    assign P[127] = in[30] ^ in2[30];
    assign G[128] = in[29] & in2[29];
    assign P[128] = in[29] ^ in2[29];
    assign G[129] = in[28] & in2[28];
    assign P[129] = in[28] ^ in2[28];
    assign G[130] = in[27] & in2[27];
    assign P[130] = in[27] ^ in2[27];
    assign G[131] = in[26] & in2[26];
    assign P[131] = in[26] ^ in2[26];
    assign G[132] = in[25] & in2[25];
    assign P[132] = in[25] ^ in2[25];
    assign G[133] = in[24] & in2[24];
    assign P[133] = in[24] ^ in2[24];
    assign G[134] = in[23] & in2[23];
    assign P[134] = in[23] ^ in2[23];
    assign G[135] = in[22] & in2[22];
    assign P[135] = in[22] ^ in2[22];
    assign G[136] = in[21] & in2[21];
    assign P[136] = in[21] ^ in2[21];
    assign G[137] = in[20] & in2[20];
    assign P[137] = in[20] ^ in2[20];
    assign G[138] = in[19] & in2[19];
    assign P[138] = in[19] ^ in2[19];
    assign G[139] = in[18] & in2[18];
    assign P[139] = in[18] ^ in2[18];
    assign G[140] = in[17] & in2[17];
    assign P[140] = in[17] ^ in2[17];
    assign G[141] = in[16] & in2[16];
    assign P[141] = in[16] ^ in2[16];
    assign G[142] = in[15] & in2[15];
    assign P[142] = in[15] ^ in2[15];
    assign G[143] = in[14] & in2[14];
    assign P[143] = in[14] ^ in2[14];
    assign G[144] = in[13] & in2[13];
    assign P[144] = in[13] ^ in2[13];
    assign G[145] = in[12] & in2[12];
    assign P[145] = in[12] ^ in2[12];
    assign G[146] = in[11] & in2[11];
    assign P[146] = in[11] ^ in2[11];
    assign G[147] = in[10] & in2[10];
    assign P[147] = in[10] ^ in2[10];
    assign G[148] = in[9] & in2[9];
    assign P[148] = in[9] ^ in2[9];
    assign G[149] = in[8] & in2[8];
    assign P[149] = in[8] ^ in2[8];
    assign G[150] = in[7] & in2[7];
    assign P[150] = in[7] ^ in2[7];
    assign G[151] = in[6] & in2[6];
    assign P[151] = in[6] ^ in2[6];
    assign G[152] = in[5] & in2[5];
    assign P[152] = in[5] ^ in2[5];
    assign G[153] = in[4] & in2[4];
    assign P[153] = in[4] ^ in2[4];
    assign G[154] = in[3] & in2[3];
    assign P[154] = in[3] ^ in2[3];
    assign G[155] = in[2] & in2[2];
    assign P[155] = in[2] ^ in2[2];
    assign G[156] = in[1] & in2[1];
    assign P[156] = in[1] ^ in2[1];
    assign G[157] = in[0] & in2[0];
    assign P[157] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign C[157] = G[156] | (P[156] & C[156]);
    assign cout = G[157] | (P[157] & C[157]);
    assign sum = P ^ C;
endmodule

module CLA157(output [156:0] sum, output cout, input [156:0] in1, input [156:0] in2;

    wire[156:0] G;
    wire[156:0] C;
    wire[156:0] P;

    assign G[0] = in[156] & in2[156];
    assign P[0] = in[156] ^ in2[156];
    assign G[1] = in[155] & in2[155];
    assign P[1] = in[155] ^ in2[155];
    assign G[2] = in[154] & in2[154];
    assign P[2] = in[154] ^ in2[154];
    assign G[3] = in[153] & in2[153];
    assign P[3] = in[153] ^ in2[153];
    assign G[4] = in[152] & in2[152];
    assign P[4] = in[152] ^ in2[152];
    assign G[5] = in[151] & in2[151];
    assign P[5] = in[151] ^ in2[151];
    assign G[6] = in[150] & in2[150];
    assign P[6] = in[150] ^ in2[150];
    assign G[7] = in[149] & in2[149];
    assign P[7] = in[149] ^ in2[149];
    assign G[8] = in[148] & in2[148];
    assign P[8] = in[148] ^ in2[148];
    assign G[9] = in[147] & in2[147];
    assign P[9] = in[147] ^ in2[147];
    assign G[10] = in[146] & in2[146];
    assign P[10] = in[146] ^ in2[146];
    assign G[11] = in[145] & in2[145];
    assign P[11] = in[145] ^ in2[145];
    assign G[12] = in[144] & in2[144];
    assign P[12] = in[144] ^ in2[144];
    assign G[13] = in[143] & in2[143];
    assign P[13] = in[143] ^ in2[143];
    assign G[14] = in[142] & in2[142];
    assign P[14] = in[142] ^ in2[142];
    assign G[15] = in[141] & in2[141];
    assign P[15] = in[141] ^ in2[141];
    assign G[16] = in[140] & in2[140];
    assign P[16] = in[140] ^ in2[140];
    assign G[17] = in[139] & in2[139];
    assign P[17] = in[139] ^ in2[139];
    assign G[18] = in[138] & in2[138];
    assign P[18] = in[138] ^ in2[138];
    assign G[19] = in[137] & in2[137];
    assign P[19] = in[137] ^ in2[137];
    assign G[20] = in[136] & in2[136];
    assign P[20] = in[136] ^ in2[136];
    assign G[21] = in[135] & in2[135];
    assign P[21] = in[135] ^ in2[135];
    assign G[22] = in[134] & in2[134];
    assign P[22] = in[134] ^ in2[134];
    assign G[23] = in[133] & in2[133];
    assign P[23] = in[133] ^ in2[133];
    assign G[24] = in[132] & in2[132];
    assign P[24] = in[132] ^ in2[132];
    assign G[25] = in[131] & in2[131];
    assign P[25] = in[131] ^ in2[131];
    assign G[26] = in[130] & in2[130];
    assign P[26] = in[130] ^ in2[130];
    assign G[27] = in[129] & in2[129];
    assign P[27] = in[129] ^ in2[129];
    assign G[28] = in[128] & in2[128];
    assign P[28] = in[128] ^ in2[128];
    assign G[29] = in[127] & in2[127];
    assign P[29] = in[127] ^ in2[127];
    assign G[30] = in[126] & in2[126];
    assign P[30] = in[126] ^ in2[126];
    assign G[31] = in[125] & in2[125];
    assign P[31] = in[125] ^ in2[125];
    assign G[32] = in[124] & in2[124];
    assign P[32] = in[124] ^ in2[124];
    assign G[33] = in[123] & in2[123];
    assign P[33] = in[123] ^ in2[123];
    assign G[34] = in[122] & in2[122];
    assign P[34] = in[122] ^ in2[122];
    assign G[35] = in[121] & in2[121];
    assign P[35] = in[121] ^ in2[121];
    assign G[36] = in[120] & in2[120];
    assign P[36] = in[120] ^ in2[120];
    assign G[37] = in[119] & in2[119];
    assign P[37] = in[119] ^ in2[119];
    assign G[38] = in[118] & in2[118];
    assign P[38] = in[118] ^ in2[118];
    assign G[39] = in[117] & in2[117];
    assign P[39] = in[117] ^ in2[117];
    assign G[40] = in[116] & in2[116];
    assign P[40] = in[116] ^ in2[116];
    assign G[41] = in[115] & in2[115];
    assign P[41] = in[115] ^ in2[115];
    assign G[42] = in[114] & in2[114];
    assign P[42] = in[114] ^ in2[114];
    assign G[43] = in[113] & in2[113];
    assign P[43] = in[113] ^ in2[113];
    assign G[44] = in[112] & in2[112];
    assign P[44] = in[112] ^ in2[112];
    assign G[45] = in[111] & in2[111];
    assign P[45] = in[111] ^ in2[111];
    assign G[46] = in[110] & in2[110];
    assign P[46] = in[110] ^ in2[110];
    assign G[47] = in[109] & in2[109];
    assign P[47] = in[109] ^ in2[109];
    assign G[48] = in[108] & in2[108];
    assign P[48] = in[108] ^ in2[108];
    assign G[49] = in[107] & in2[107];
    assign P[49] = in[107] ^ in2[107];
    assign G[50] = in[106] & in2[106];
    assign P[50] = in[106] ^ in2[106];
    assign G[51] = in[105] & in2[105];
    assign P[51] = in[105] ^ in2[105];
    assign G[52] = in[104] & in2[104];
    assign P[52] = in[104] ^ in2[104];
    assign G[53] = in[103] & in2[103];
    assign P[53] = in[103] ^ in2[103];
    assign G[54] = in[102] & in2[102];
    assign P[54] = in[102] ^ in2[102];
    assign G[55] = in[101] & in2[101];
    assign P[55] = in[101] ^ in2[101];
    assign G[56] = in[100] & in2[100];
    assign P[56] = in[100] ^ in2[100];
    assign G[57] = in[99] & in2[99];
    assign P[57] = in[99] ^ in2[99];
    assign G[58] = in[98] & in2[98];
    assign P[58] = in[98] ^ in2[98];
    assign G[59] = in[97] & in2[97];
    assign P[59] = in[97] ^ in2[97];
    assign G[60] = in[96] & in2[96];
    assign P[60] = in[96] ^ in2[96];
    assign G[61] = in[95] & in2[95];
    assign P[61] = in[95] ^ in2[95];
    assign G[62] = in[94] & in2[94];
    assign P[62] = in[94] ^ in2[94];
    assign G[63] = in[93] & in2[93];
    assign P[63] = in[93] ^ in2[93];
    assign G[64] = in[92] & in2[92];
    assign P[64] = in[92] ^ in2[92];
    assign G[65] = in[91] & in2[91];
    assign P[65] = in[91] ^ in2[91];
    assign G[66] = in[90] & in2[90];
    assign P[66] = in[90] ^ in2[90];
    assign G[67] = in[89] & in2[89];
    assign P[67] = in[89] ^ in2[89];
    assign G[68] = in[88] & in2[88];
    assign P[68] = in[88] ^ in2[88];
    assign G[69] = in[87] & in2[87];
    assign P[69] = in[87] ^ in2[87];
    assign G[70] = in[86] & in2[86];
    assign P[70] = in[86] ^ in2[86];
    assign G[71] = in[85] & in2[85];
    assign P[71] = in[85] ^ in2[85];
    assign G[72] = in[84] & in2[84];
    assign P[72] = in[84] ^ in2[84];
    assign G[73] = in[83] & in2[83];
    assign P[73] = in[83] ^ in2[83];
    assign G[74] = in[82] & in2[82];
    assign P[74] = in[82] ^ in2[82];
    assign G[75] = in[81] & in2[81];
    assign P[75] = in[81] ^ in2[81];
    assign G[76] = in[80] & in2[80];
    assign P[76] = in[80] ^ in2[80];
    assign G[77] = in[79] & in2[79];
    assign P[77] = in[79] ^ in2[79];
    assign G[78] = in[78] & in2[78];
    assign P[78] = in[78] ^ in2[78];
    assign G[79] = in[77] & in2[77];
    assign P[79] = in[77] ^ in2[77];
    assign G[80] = in[76] & in2[76];
    assign P[80] = in[76] ^ in2[76];
    assign G[81] = in[75] & in2[75];
    assign P[81] = in[75] ^ in2[75];
    assign G[82] = in[74] & in2[74];
    assign P[82] = in[74] ^ in2[74];
    assign G[83] = in[73] & in2[73];
    assign P[83] = in[73] ^ in2[73];
    assign G[84] = in[72] & in2[72];
    assign P[84] = in[72] ^ in2[72];
    assign G[85] = in[71] & in2[71];
    assign P[85] = in[71] ^ in2[71];
    assign G[86] = in[70] & in2[70];
    assign P[86] = in[70] ^ in2[70];
    assign G[87] = in[69] & in2[69];
    assign P[87] = in[69] ^ in2[69];
    assign G[88] = in[68] & in2[68];
    assign P[88] = in[68] ^ in2[68];
    assign G[89] = in[67] & in2[67];
    assign P[89] = in[67] ^ in2[67];
    assign G[90] = in[66] & in2[66];
    assign P[90] = in[66] ^ in2[66];
    assign G[91] = in[65] & in2[65];
    assign P[91] = in[65] ^ in2[65];
    assign G[92] = in[64] & in2[64];
    assign P[92] = in[64] ^ in2[64];
    assign G[93] = in[63] & in2[63];
    assign P[93] = in[63] ^ in2[63];
    assign G[94] = in[62] & in2[62];
    assign P[94] = in[62] ^ in2[62];
    assign G[95] = in[61] & in2[61];
    assign P[95] = in[61] ^ in2[61];
    assign G[96] = in[60] & in2[60];
    assign P[96] = in[60] ^ in2[60];
    assign G[97] = in[59] & in2[59];
    assign P[97] = in[59] ^ in2[59];
    assign G[98] = in[58] & in2[58];
    assign P[98] = in[58] ^ in2[58];
    assign G[99] = in[57] & in2[57];
    assign P[99] = in[57] ^ in2[57];
    assign G[100] = in[56] & in2[56];
    assign P[100] = in[56] ^ in2[56];
    assign G[101] = in[55] & in2[55];
    assign P[101] = in[55] ^ in2[55];
    assign G[102] = in[54] & in2[54];
    assign P[102] = in[54] ^ in2[54];
    assign G[103] = in[53] & in2[53];
    assign P[103] = in[53] ^ in2[53];
    assign G[104] = in[52] & in2[52];
    assign P[104] = in[52] ^ in2[52];
    assign G[105] = in[51] & in2[51];
    assign P[105] = in[51] ^ in2[51];
    assign G[106] = in[50] & in2[50];
    assign P[106] = in[50] ^ in2[50];
    assign G[107] = in[49] & in2[49];
    assign P[107] = in[49] ^ in2[49];
    assign G[108] = in[48] & in2[48];
    assign P[108] = in[48] ^ in2[48];
    assign G[109] = in[47] & in2[47];
    assign P[109] = in[47] ^ in2[47];
    assign G[110] = in[46] & in2[46];
    assign P[110] = in[46] ^ in2[46];
    assign G[111] = in[45] & in2[45];
    assign P[111] = in[45] ^ in2[45];
    assign G[112] = in[44] & in2[44];
    assign P[112] = in[44] ^ in2[44];
    assign G[113] = in[43] & in2[43];
    assign P[113] = in[43] ^ in2[43];
    assign G[114] = in[42] & in2[42];
    assign P[114] = in[42] ^ in2[42];
    assign G[115] = in[41] & in2[41];
    assign P[115] = in[41] ^ in2[41];
    assign G[116] = in[40] & in2[40];
    assign P[116] = in[40] ^ in2[40];
    assign G[117] = in[39] & in2[39];
    assign P[117] = in[39] ^ in2[39];
    assign G[118] = in[38] & in2[38];
    assign P[118] = in[38] ^ in2[38];
    assign G[119] = in[37] & in2[37];
    assign P[119] = in[37] ^ in2[37];
    assign G[120] = in[36] & in2[36];
    assign P[120] = in[36] ^ in2[36];
    assign G[121] = in[35] & in2[35];
    assign P[121] = in[35] ^ in2[35];
    assign G[122] = in[34] & in2[34];
    assign P[122] = in[34] ^ in2[34];
    assign G[123] = in[33] & in2[33];
    assign P[123] = in[33] ^ in2[33];
    assign G[124] = in[32] & in2[32];
    assign P[124] = in[32] ^ in2[32];
    assign G[125] = in[31] & in2[31];
    assign P[125] = in[31] ^ in2[31];
    assign G[126] = in[30] & in2[30];
    assign P[126] = in[30] ^ in2[30];
    assign G[127] = in[29] & in2[29];
    assign P[127] = in[29] ^ in2[29];
    assign G[128] = in[28] & in2[28];
    assign P[128] = in[28] ^ in2[28];
    assign G[129] = in[27] & in2[27];
    assign P[129] = in[27] ^ in2[27];
    assign G[130] = in[26] & in2[26];
    assign P[130] = in[26] ^ in2[26];
    assign G[131] = in[25] & in2[25];
    assign P[131] = in[25] ^ in2[25];
    assign G[132] = in[24] & in2[24];
    assign P[132] = in[24] ^ in2[24];
    assign G[133] = in[23] & in2[23];
    assign P[133] = in[23] ^ in2[23];
    assign G[134] = in[22] & in2[22];
    assign P[134] = in[22] ^ in2[22];
    assign G[135] = in[21] & in2[21];
    assign P[135] = in[21] ^ in2[21];
    assign G[136] = in[20] & in2[20];
    assign P[136] = in[20] ^ in2[20];
    assign G[137] = in[19] & in2[19];
    assign P[137] = in[19] ^ in2[19];
    assign G[138] = in[18] & in2[18];
    assign P[138] = in[18] ^ in2[18];
    assign G[139] = in[17] & in2[17];
    assign P[139] = in[17] ^ in2[17];
    assign G[140] = in[16] & in2[16];
    assign P[140] = in[16] ^ in2[16];
    assign G[141] = in[15] & in2[15];
    assign P[141] = in[15] ^ in2[15];
    assign G[142] = in[14] & in2[14];
    assign P[142] = in[14] ^ in2[14];
    assign G[143] = in[13] & in2[13];
    assign P[143] = in[13] ^ in2[13];
    assign G[144] = in[12] & in2[12];
    assign P[144] = in[12] ^ in2[12];
    assign G[145] = in[11] & in2[11];
    assign P[145] = in[11] ^ in2[11];
    assign G[146] = in[10] & in2[10];
    assign P[146] = in[10] ^ in2[10];
    assign G[147] = in[9] & in2[9];
    assign P[147] = in[9] ^ in2[9];
    assign G[148] = in[8] & in2[8];
    assign P[148] = in[8] ^ in2[8];
    assign G[149] = in[7] & in2[7];
    assign P[149] = in[7] ^ in2[7];
    assign G[150] = in[6] & in2[6];
    assign P[150] = in[6] ^ in2[6];
    assign G[151] = in[5] & in2[5];
    assign P[151] = in[5] ^ in2[5];
    assign G[152] = in[4] & in2[4];
    assign P[152] = in[4] ^ in2[4];
    assign G[153] = in[3] & in2[3];
    assign P[153] = in[3] ^ in2[3];
    assign G[154] = in[2] & in2[2];
    assign P[154] = in[2] ^ in2[2];
    assign G[155] = in[1] & in2[1];
    assign P[155] = in[1] ^ in2[1];
    assign G[156] = in[0] & in2[0];
    assign P[156] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign C[156] = G[155] | (P[155] & C[155]);
    assign cout = G[156] | (P[156] & C[156]);
    assign sum = P ^ C;
endmodule

module CLA156(output [155:0] sum, output cout, input [155:0] in1, input [155:0] in2;

    wire[155:0] G;
    wire[155:0] C;
    wire[155:0] P;

    assign G[0] = in[155] & in2[155];
    assign P[0] = in[155] ^ in2[155];
    assign G[1] = in[154] & in2[154];
    assign P[1] = in[154] ^ in2[154];
    assign G[2] = in[153] & in2[153];
    assign P[2] = in[153] ^ in2[153];
    assign G[3] = in[152] & in2[152];
    assign P[3] = in[152] ^ in2[152];
    assign G[4] = in[151] & in2[151];
    assign P[4] = in[151] ^ in2[151];
    assign G[5] = in[150] & in2[150];
    assign P[5] = in[150] ^ in2[150];
    assign G[6] = in[149] & in2[149];
    assign P[6] = in[149] ^ in2[149];
    assign G[7] = in[148] & in2[148];
    assign P[7] = in[148] ^ in2[148];
    assign G[8] = in[147] & in2[147];
    assign P[8] = in[147] ^ in2[147];
    assign G[9] = in[146] & in2[146];
    assign P[9] = in[146] ^ in2[146];
    assign G[10] = in[145] & in2[145];
    assign P[10] = in[145] ^ in2[145];
    assign G[11] = in[144] & in2[144];
    assign P[11] = in[144] ^ in2[144];
    assign G[12] = in[143] & in2[143];
    assign P[12] = in[143] ^ in2[143];
    assign G[13] = in[142] & in2[142];
    assign P[13] = in[142] ^ in2[142];
    assign G[14] = in[141] & in2[141];
    assign P[14] = in[141] ^ in2[141];
    assign G[15] = in[140] & in2[140];
    assign P[15] = in[140] ^ in2[140];
    assign G[16] = in[139] & in2[139];
    assign P[16] = in[139] ^ in2[139];
    assign G[17] = in[138] & in2[138];
    assign P[17] = in[138] ^ in2[138];
    assign G[18] = in[137] & in2[137];
    assign P[18] = in[137] ^ in2[137];
    assign G[19] = in[136] & in2[136];
    assign P[19] = in[136] ^ in2[136];
    assign G[20] = in[135] & in2[135];
    assign P[20] = in[135] ^ in2[135];
    assign G[21] = in[134] & in2[134];
    assign P[21] = in[134] ^ in2[134];
    assign G[22] = in[133] & in2[133];
    assign P[22] = in[133] ^ in2[133];
    assign G[23] = in[132] & in2[132];
    assign P[23] = in[132] ^ in2[132];
    assign G[24] = in[131] & in2[131];
    assign P[24] = in[131] ^ in2[131];
    assign G[25] = in[130] & in2[130];
    assign P[25] = in[130] ^ in2[130];
    assign G[26] = in[129] & in2[129];
    assign P[26] = in[129] ^ in2[129];
    assign G[27] = in[128] & in2[128];
    assign P[27] = in[128] ^ in2[128];
    assign G[28] = in[127] & in2[127];
    assign P[28] = in[127] ^ in2[127];
    assign G[29] = in[126] & in2[126];
    assign P[29] = in[126] ^ in2[126];
    assign G[30] = in[125] & in2[125];
    assign P[30] = in[125] ^ in2[125];
    assign G[31] = in[124] & in2[124];
    assign P[31] = in[124] ^ in2[124];
    assign G[32] = in[123] & in2[123];
    assign P[32] = in[123] ^ in2[123];
    assign G[33] = in[122] & in2[122];
    assign P[33] = in[122] ^ in2[122];
    assign G[34] = in[121] & in2[121];
    assign P[34] = in[121] ^ in2[121];
    assign G[35] = in[120] & in2[120];
    assign P[35] = in[120] ^ in2[120];
    assign G[36] = in[119] & in2[119];
    assign P[36] = in[119] ^ in2[119];
    assign G[37] = in[118] & in2[118];
    assign P[37] = in[118] ^ in2[118];
    assign G[38] = in[117] & in2[117];
    assign P[38] = in[117] ^ in2[117];
    assign G[39] = in[116] & in2[116];
    assign P[39] = in[116] ^ in2[116];
    assign G[40] = in[115] & in2[115];
    assign P[40] = in[115] ^ in2[115];
    assign G[41] = in[114] & in2[114];
    assign P[41] = in[114] ^ in2[114];
    assign G[42] = in[113] & in2[113];
    assign P[42] = in[113] ^ in2[113];
    assign G[43] = in[112] & in2[112];
    assign P[43] = in[112] ^ in2[112];
    assign G[44] = in[111] & in2[111];
    assign P[44] = in[111] ^ in2[111];
    assign G[45] = in[110] & in2[110];
    assign P[45] = in[110] ^ in2[110];
    assign G[46] = in[109] & in2[109];
    assign P[46] = in[109] ^ in2[109];
    assign G[47] = in[108] & in2[108];
    assign P[47] = in[108] ^ in2[108];
    assign G[48] = in[107] & in2[107];
    assign P[48] = in[107] ^ in2[107];
    assign G[49] = in[106] & in2[106];
    assign P[49] = in[106] ^ in2[106];
    assign G[50] = in[105] & in2[105];
    assign P[50] = in[105] ^ in2[105];
    assign G[51] = in[104] & in2[104];
    assign P[51] = in[104] ^ in2[104];
    assign G[52] = in[103] & in2[103];
    assign P[52] = in[103] ^ in2[103];
    assign G[53] = in[102] & in2[102];
    assign P[53] = in[102] ^ in2[102];
    assign G[54] = in[101] & in2[101];
    assign P[54] = in[101] ^ in2[101];
    assign G[55] = in[100] & in2[100];
    assign P[55] = in[100] ^ in2[100];
    assign G[56] = in[99] & in2[99];
    assign P[56] = in[99] ^ in2[99];
    assign G[57] = in[98] & in2[98];
    assign P[57] = in[98] ^ in2[98];
    assign G[58] = in[97] & in2[97];
    assign P[58] = in[97] ^ in2[97];
    assign G[59] = in[96] & in2[96];
    assign P[59] = in[96] ^ in2[96];
    assign G[60] = in[95] & in2[95];
    assign P[60] = in[95] ^ in2[95];
    assign G[61] = in[94] & in2[94];
    assign P[61] = in[94] ^ in2[94];
    assign G[62] = in[93] & in2[93];
    assign P[62] = in[93] ^ in2[93];
    assign G[63] = in[92] & in2[92];
    assign P[63] = in[92] ^ in2[92];
    assign G[64] = in[91] & in2[91];
    assign P[64] = in[91] ^ in2[91];
    assign G[65] = in[90] & in2[90];
    assign P[65] = in[90] ^ in2[90];
    assign G[66] = in[89] & in2[89];
    assign P[66] = in[89] ^ in2[89];
    assign G[67] = in[88] & in2[88];
    assign P[67] = in[88] ^ in2[88];
    assign G[68] = in[87] & in2[87];
    assign P[68] = in[87] ^ in2[87];
    assign G[69] = in[86] & in2[86];
    assign P[69] = in[86] ^ in2[86];
    assign G[70] = in[85] & in2[85];
    assign P[70] = in[85] ^ in2[85];
    assign G[71] = in[84] & in2[84];
    assign P[71] = in[84] ^ in2[84];
    assign G[72] = in[83] & in2[83];
    assign P[72] = in[83] ^ in2[83];
    assign G[73] = in[82] & in2[82];
    assign P[73] = in[82] ^ in2[82];
    assign G[74] = in[81] & in2[81];
    assign P[74] = in[81] ^ in2[81];
    assign G[75] = in[80] & in2[80];
    assign P[75] = in[80] ^ in2[80];
    assign G[76] = in[79] & in2[79];
    assign P[76] = in[79] ^ in2[79];
    assign G[77] = in[78] & in2[78];
    assign P[77] = in[78] ^ in2[78];
    assign G[78] = in[77] & in2[77];
    assign P[78] = in[77] ^ in2[77];
    assign G[79] = in[76] & in2[76];
    assign P[79] = in[76] ^ in2[76];
    assign G[80] = in[75] & in2[75];
    assign P[80] = in[75] ^ in2[75];
    assign G[81] = in[74] & in2[74];
    assign P[81] = in[74] ^ in2[74];
    assign G[82] = in[73] & in2[73];
    assign P[82] = in[73] ^ in2[73];
    assign G[83] = in[72] & in2[72];
    assign P[83] = in[72] ^ in2[72];
    assign G[84] = in[71] & in2[71];
    assign P[84] = in[71] ^ in2[71];
    assign G[85] = in[70] & in2[70];
    assign P[85] = in[70] ^ in2[70];
    assign G[86] = in[69] & in2[69];
    assign P[86] = in[69] ^ in2[69];
    assign G[87] = in[68] & in2[68];
    assign P[87] = in[68] ^ in2[68];
    assign G[88] = in[67] & in2[67];
    assign P[88] = in[67] ^ in2[67];
    assign G[89] = in[66] & in2[66];
    assign P[89] = in[66] ^ in2[66];
    assign G[90] = in[65] & in2[65];
    assign P[90] = in[65] ^ in2[65];
    assign G[91] = in[64] & in2[64];
    assign P[91] = in[64] ^ in2[64];
    assign G[92] = in[63] & in2[63];
    assign P[92] = in[63] ^ in2[63];
    assign G[93] = in[62] & in2[62];
    assign P[93] = in[62] ^ in2[62];
    assign G[94] = in[61] & in2[61];
    assign P[94] = in[61] ^ in2[61];
    assign G[95] = in[60] & in2[60];
    assign P[95] = in[60] ^ in2[60];
    assign G[96] = in[59] & in2[59];
    assign P[96] = in[59] ^ in2[59];
    assign G[97] = in[58] & in2[58];
    assign P[97] = in[58] ^ in2[58];
    assign G[98] = in[57] & in2[57];
    assign P[98] = in[57] ^ in2[57];
    assign G[99] = in[56] & in2[56];
    assign P[99] = in[56] ^ in2[56];
    assign G[100] = in[55] & in2[55];
    assign P[100] = in[55] ^ in2[55];
    assign G[101] = in[54] & in2[54];
    assign P[101] = in[54] ^ in2[54];
    assign G[102] = in[53] & in2[53];
    assign P[102] = in[53] ^ in2[53];
    assign G[103] = in[52] & in2[52];
    assign P[103] = in[52] ^ in2[52];
    assign G[104] = in[51] & in2[51];
    assign P[104] = in[51] ^ in2[51];
    assign G[105] = in[50] & in2[50];
    assign P[105] = in[50] ^ in2[50];
    assign G[106] = in[49] & in2[49];
    assign P[106] = in[49] ^ in2[49];
    assign G[107] = in[48] & in2[48];
    assign P[107] = in[48] ^ in2[48];
    assign G[108] = in[47] & in2[47];
    assign P[108] = in[47] ^ in2[47];
    assign G[109] = in[46] & in2[46];
    assign P[109] = in[46] ^ in2[46];
    assign G[110] = in[45] & in2[45];
    assign P[110] = in[45] ^ in2[45];
    assign G[111] = in[44] & in2[44];
    assign P[111] = in[44] ^ in2[44];
    assign G[112] = in[43] & in2[43];
    assign P[112] = in[43] ^ in2[43];
    assign G[113] = in[42] & in2[42];
    assign P[113] = in[42] ^ in2[42];
    assign G[114] = in[41] & in2[41];
    assign P[114] = in[41] ^ in2[41];
    assign G[115] = in[40] & in2[40];
    assign P[115] = in[40] ^ in2[40];
    assign G[116] = in[39] & in2[39];
    assign P[116] = in[39] ^ in2[39];
    assign G[117] = in[38] & in2[38];
    assign P[117] = in[38] ^ in2[38];
    assign G[118] = in[37] & in2[37];
    assign P[118] = in[37] ^ in2[37];
    assign G[119] = in[36] & in2[36];
    assign P[119] = in[36] ^ in2[36];
    assign G[120] = in[35] & in2[35];
    assign P[120] = in[35] ^ in2[35];
    assign G[121] = in[34] & in2[34];
    assign P[121] = in[34] ^ in2[34];
    assign G[122] = in[33] & in2[33];
    assign P[122] = in[33] ^ in2[33];
    assign G[123] = in[32] & in2[32];
    assign P[123] = in[32] ^ in2[32];
    assign G[124] = in[31] & in2[31];
    assign P[124] = in[31] ^ in2[31];
    assign G[125] = in[30] & in2[30];
    assign P[125] = in[30] ^ in2[30];
    assign G[126] = in[29] & in2[29];
    assign P[126] = in[29] ^ in2[29];
    assign G[127] = in[28] & in2[28];
    assign P[127] = in[28] ^ in2[28];
    assign G[128] = in[27] & in2[27];
    assign P[128] = in[27] ^ in2[27];
    assign G[129] = in[26] & in2[26];
    assign P[129] = in[26] ^ in2[26];
    assign G[130] = in[25] & in2[25];
    assign P[130] = in[25] ^ in2[25];
    assign G[131] = in[24] & in2[24];
    assign P[131] = in[24] ^ in2[24];
    assign G[132] = in[23] & in2[23];
    assign P[132] = in[23] ^ in2[23];
    assign G[133] = in[22] & in2[22];
    assign P[133] = in[22] ^ in2[22];
    assign G[134] = in[21] & in2[21];
    assign P[134] = in[21] ^ in2[21];
    assign G[135] = in[20] & in2[20];
    assign P[135] = in[20] ^ in2[20];
    assign G[136] = in[19] & in2[19];
    assign P[136] = in[19] ^ in2[19];
    assign G[137] = in[18] & in2[18];
    assign P[137] = in[18] ^ in2[18];
    assign G[138] = in[17] & in2[17];
    assign P[138] = in[17] ^ in2[17];
    assign G[139] = in[16] & in2[16];
    assign P[139] = in[16] ^ in2[16];
    assign G[140] = in[15] & in2[15];
    assign P[140] = in[15] ^ in2[15];
    assign G[141] = in[14] & in2[14];
    assign P[141] = in[14] ^ in2[14];
    assign G[142] = in[13] & in2[13];
    assign P[142] = in[13] ^ in2[13];
    assign G[143] = in[12] & in2[12];
    assign P[143] = in[12] ^ in2[12];
    assign G[144] = in[11] & in2[11];
    assign P[144] = in[11] ^ in2[11];
    assign G[145] = in[10] & in2[10];
    assign P[145] = in[10] ^ in2[10];
    assign G[146] = in[9] & in2[9];
    assign P[146] = in[9] ^ in2[9];
    assign G[147] = in[8] & in2[8];
    assign P[147] = in[8] ^ in2[8];
    assign G[148] = in[7] & in2[7];
    assign P[148] = in[7] ^ in2[7];
    assign G[149] = in[6] & in2[6];
    assign P[149] = in[6] ^ in2[6];
    assign G[150] = in[5] & in2[5];
    assign P[150] = in[5] ^ in2[5];
    assign G[151] = in[4] & in2[4];
    assign P[151] = in[4] ^ in2[4];
    assign G[152] = in[3] & in2[3];
    assign P[152] = in[3] ^ in2[3];
    assign G[153] = in[2] & in2[2];
    assign P[153] = in[2] ^ in2[2];
    assign G[154] = in[1] & in2[1];
    assign P[154] = in[1] ^ in2[1];
    assign G[155] = in[0] & in2[0];
    assign P[155] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign C[155] = G[154] | (P[154] & C[154]);
    assign cout = G[155] | (P[155] & C[155]);
    assign sum = P ^ C;
endmodule

module CLA155(output [154:0] sum, output cout, input [154:0] in1, input [154:0] in2;

    wire[154:0] G;
    wire[154:0] C;
    wire[154:0] P;

    assign G[0] = in[154] & in2[154];
    assign P[0] = in[154] ^ in2[154];
    assign G[1] = in[153] & in2[153];
    assign P[1] = in[153] ^ in2[153];
    assign G[2] = in[152] & in2[152];
    assign P[2] = in[152] ^ in2[152];
    assign G[3] = in[151] & in2[151];
    assign P[3] = in[151] ^ in2[151];
    assign G[4] = in[150] & in2[150];
    assign P[4] = in[150] ^ in2[150];
    assign G[5] = in[149] & in2[149];
    assign P[5] = in[149] ^ in2[149];
    assign G[6] = in[148] & in2[148];
    assign P[6] = in[148] ^ in2[148];
    assign G[7] = in[147] & in2[147];
    assign P[7] = in[147] ^ in2[147];
    assign G[8] = in[146] & in2[146];
    assign P[8] = in[146] ^ in2[146];
    assign G[9] = in[145] & in2[145];
    assign P[9] = in[145] ^ in2[145];
    assign G[10] = in[144] & in2[144];
    assign P[10] = in[144] ^ in2[144];
    assign G[11] = in[143] & in2[143];
    assign P[11] = in[143] ^ in2[143];
    assign G[12] = in[142] & in2[142];
    assign P[12] = in[142] ^ in2[142];
    assign G[13] = in[141] & in2[141];
    assign P[13] = in[141] ^ in2[141];
    assign G[14] = in[140] & in2[140];
    assign P[14] = in[140] ^ in2[140];
    assign G[15] = in[139] & in2[139];
    assign P[15] = in[139] ^ in2[139];
    assign G[16] = in[138] & in2[138];
    assign P[16] = in[138] ^ in2[138];
    assign G[17] = in[137] & in2[137];
    assign P[17] = in[137] ^ in2[137];
    assign G[18] = in[136] & in2[136];
    assign P[18] = in[136] ^ in2[136];
    assign G[19] = in[135] & in2[135];
    assign P[19] = in[135] ^ in2[135];
    assign G[20] = in[134] & in2[134];
    assign P[20] = in[134] ^ in2[134];
    assign G[21] = in[133] & in2[133];
    assign P[21] = in[133] ^ in2[133];
    assign G[22] = in[132] & in2[132];
    assign P[22] = in[132] ^ in2[132];
    assign G[23] = in[131] & in2[131];
    assign P[23] = in[131] ^ in2[131];
    assign G[24] = in[130] & in2[130];
    assign P[24] = in[130] ^ in2[130];
    assign G[25] = in[129] & in2[129];
    assign P[25] = in[129] ^ in2[129];
    assign G[26] = in[128] & in2[128];
    assign P[26] = in[128] ^ in2[128];
    assign G[27] = in[127] & in2[127];
    assign P[27] = in[127] ^ in2[127];
    assign G[28] = in[126] & in2[126];
    assign P[28] = in[126] ^ in2[126];
    assign G[29] = in[125] & in2[125];
    assign P[29] = in[125] ^ in2[125];
    assign G[30] = in[124] & in2[124];
    assign P[30] = in[124] ^ in2[124];
    assign G[31] = in[123] & in2[123];
    assign P[31] = in[123] ^ in2[123];
    assign G[32] = in[122] & in2[122];
    assign P[32] = in[122] ^ in2[122];
    assign G[33] = in[121] & in2[121];
    assign P[33] = in[121] ^ in2[121];
    assign G[34] = in[120] & in2[120];
    assign P[34] = in[120] ^ in2[120];
    assign G[35] = in[119] & in2[119];
    assign P[35] = in[119] ^ in2[119];
    assign G[36] = in[118] & in2[118];
    assign P[36] = in[118] ^ in2[118];
    assign G[37] = in[117] & in2[117];
    assign P[37] = in[117] ^ in2[117];
    assign G[38] = in[116] & in2[116];
    assign P[38] = in[116] ^ in2[116];
    assign G[39] = in[115] & in2[115];
    assign P[39] = in[115] ^ in2[115];
    assign G[40] = in[114] & in2[114];
    assign P[40] = in[114] ^ in2[114];
    assign G[41] = in[113] & in2[113];
    assign P[41] = in[113] ^ in2[113];
    assign G[42] = in[112] & in2[112];
    assign P[42] = in[112] ^ in2[112];
    assign G[43] = in[111] & in2[111];
    assign P[43] = in[111] ^ in2[111];
    assign G[44] = in[110] & in2[110];
    assign P[44] = in[110] ^ in2[110];
    assign G[45] = in[109] & in2[109];
    assign P[45] = in[109] ^ in2[109];
    assign G[46] = in[108] & in2[108];
    assign P[46] = in[108] ^ in2[108];
    assign G[47] = in[107] & in2[107];
    assign P[47] = in[107] ^ in2[107];
    assign G[48] = in[106] & in2[106];
    assign P[48] = in[106] ^ in2[106];
    assign G[49] = in[105] & in2[105];
    assign P[49] = in[105] ^ in2[105];
    assign G[50] = in[104] & in2[104];
    assign P[50] = in[104] ^ in2[104];
    assign G[51] = in[103] & in2[103];
    assign P[51] = in[103] ^ in2[103];
    assign G[52] = in[102] & in2[102];
    assign P[52] = in[102] ^ in2[102];
    assign G[53] = in[101] & in2[101];
    assign P[53] = in[101] ^ in2[101];
    assign G[54] = in[100] & in2[100];
    assign P[54] = in[100] ^ in2[100];
    assign G[55] = in[99] & in2[99];
    assign P[55] = in[99] ^ in2[99];
    assign G[56] = in[98] & in2[98];
    assign P[56] = in[98] ^ in2[98];
    assign G[57] = in[97] & in2[97];
    assign P[57] = in[97] ^ in2[97];
    assign G[58] = in[96] & in2[96];
    assign P[58] = in[96] ^ in2[96];
    assign G[59] = in[95] & in2[95];
    assign P[59] = in[95] ^ in2[95];
    assign G[60] = in[94] & in2[94];
    assign P[60] = in[94] ^ in2[94];
    assign G[61] = in[93] & in2[93];
    assign P[61] = in[93] ^ in2[93];
    assign G[62] = in[92] & in2[92];
    assign P[62] = in[92] ^ in2[92];
    assign G[63] = in[91] & in2[91];
    assign P[63] = in[91] ^ in2[91];
    assign G[64] = in[90] & in2[90];
    assign P[64] = in[90] ^ in2[90];
    assign G[65] = in[89] & in2[89];
    assign P[65] = in[89] ^ in2[89];
    assign G[66] = in[88] & in2[88];
    assign P[66] = in[88] ^ in2[88];
    assign G[67] = in[87] & in2[87];
    assign P[67] = in[87] ^ in2[87];
    assign G[68] = in[86] & in2[86];
    assign P[68] = in[86] ^ in2[86];
    assign G[69] = in[85] & in2[85];
    assign P[69] = in[85] ^ in2[85];
    assign G[70] = in[84] & in2[84];
    assign P[70] = in[84] ^ in2[84];
    assign G[71] = in[83] & in2[83];
    assign P[71] = in[83] ^ in2[83];
    assign G[72] = in[82] & in2[82];
    assign P[72] = in[82] ^ in2[82];
    assign G[73] = in[81] & in2[81];
    assign P[73] = in[81] ^ in2[81];
    assign G[74] = in[80] & in2[80];
    assign P[74] = in[80] ^ in2[80];
    assign G[75] = in[79] & in2[79];
    assign P[75] = in[79] ^ in2[79];
    assign G[76] = in[78] & in2[78];
    assign P[76] = in[78] ^ in2[78];
    assign G[77] = in[77] & in2[77];
    assign P[77] = in[77] ^ in2[77];
    assign G[78] = in[76] & in2[76];
    assign P[78] = in[76] ^ in2[76];
    assign G[79] = in[75] & in2[75];
    assign P[79] = in[75] ^ in2[75];
    assign G[80] = in[74] & in2[74];
    assign P[80] = in[74] ^ in2[74];
    assign G[81] = in[73] & in2[73];
    assign P[81] = in[73] ^ in2[73];
    assign G[82] = in[72] & in2[72];
    assign P[82] = in[72] ^ in2[72];
    assign G[83] = in[71] & in2[71];
    assign P[83] = in[71] ^ in2[71];
    assign G[84] = in[70] & in2[70];
    assign P[84] = in[70] ^ in2[70];
    assign G[85] = in[69] & in2[69];
    assign P[85] = in[69] ^ in2[69];
    assign G[86] = in[68] & in2[68];
    assign P[86] = in[68] ^ in2[68];
    assign G[87] = in[67] & in2[67];
    assign P[87] = in[67] ^ in2[67];
    assign G[88] = in[66] & in2[66];
    assign P[88] = in[66] ^ in2[66];
    assign G[89] = in[65] & in2[65];
    assign P[89] = in[65] ^ in2[65];
    assign G[90] = in[64] & in2[64];
    assign P[90] = in[64] ^ in2[64];
    assign G[91] = in[63] & in2[63];
    assign P[91] = in[63] ^ in2[63];
    assign G[92] = in[62] & in2[62];
    assign P[92] = in[62] ^ in2[62];
    assign G[93] = in[61] & in2[61];
    assign P[93] = in[61] ^ in2[61];
    assign G[94] = in[60] & in2[60];
    assign P[94] = in[60] ^ in2[60];
    assign G[95] = in[59] & in2[59];
    assign P[95] = in[59] ^ in2[59];
    assign G[96] = in[58] & in2[58];
    assign P[96] = in[58] ^ in2[58];
    assign G[97] = in[57] & in2[57];
    assign P[97] = in[57] ^ in2[57];
    assign G[98] = in[56] & in2[56];
    assign P[98] = in[56] ^ in2[56];
    assign G[99] = in[55] & in2[55];
    assign P[99] = in[55] ^ in2[55];
    assign G[100] = in[54] & in2[54];
    assign P[100] = in[54] ^ in2[54];
    assign G[101] = in[53] & in2[53];
    assign P[101] = in[53] ^ in2[53];
    assign G[102] = in[52] & in2[52];
    assign P[102] = in[52] ^ in2[52];
    assign G[103] = in[51] & in2[51];
    assign P[103] = in[51] ^ in2[51];
    assign G[104] = in[50] & in2[50];
    assign P[104] = in[50] ^ in2[50];
    assign G[105] = in[49] & in2[49];
    assign P[105] = in[49] ^ in2[49];
    assign G[106] = in[48] & in2[48];
    assign P[106] = in[48] ^ in2[48];
    assign G[107] = in[47] & in2[47];
    assign P[107] = in[47] ^ in2[47];
    assign G[108] = in[46] & in2[46];
    assign P[108] = in[46] ^ in2[46];
    assign G[109] = in[45] & in2[45];
    assign P[109] = in[45] ^ in2[45];
    assign G[110] = in[44] & in2[44];
    assign P[110] = in[44] ^ in2[44];
    assign G[111] = in[43] & in2[43];
    assign P[111] = in[43] ^ in2[43];
    assign G[112] = in[42] & in2[42];
    assign P[112] = in[42] ^ in2[42];
    assign G[113] = in[41] & in2[41];
    assign P[113] = in[41] ^ in2[41];
    assign G[114] = in[40] & in2[40];
    assign P[114] = in[40] ^ in2[40];
    assign G[115] = in[39] & in2[39];
    assign P[115] = in[39] ^ in2[39];
    assign G[116] = in[38] & in2[38];
    assign P[116] = in[38] ^ in2[38];
    assign G[117] = in[37] & in2[37];
    assign P[117] = in[37] ^ in2[37];
    assign G[118] = in[36] & in2[36];
    assign P[118] = in[36] ^ in2[36];
    assign G[119] = in[35] & in2[35];
    assign P[119] = in[35] ^ in2[35];
    assign G[120] = in[34] & in2[34];
    assign P[120] = in[34] ^ in2[34];
    assign G[121] = in[33] & in2[33];
    assign P[121] = in[33] ^ in2[33];
    assign G[122] = in[32] & in2[32];
    assign P[122] = in[32] ^ in2[32];
    assign G[123] = in[31] & in2[31];
    assign P[123] = in[31] ^ in2[31];
    assign G[124] = in[30] & in2[30];
    assign P[124] = in[30] ^ in2[30];
    assign G[125] = in[29] & in2[29];
    assign P[125] = in[29] ^ in2[29];
    assign G[126] = in[28] & in2[28];
    assign P[126] = in[28] ^ in2[28];
    assign G[127] = in[27] & in2[27];
    assign P[127] = in[27] ^ in2[27];
    assign G[128] = in[26] & in2[26];
    assign P[128] = in[26] ^ in2[26];
    assign G[129] = in[25] & in2[25];
    assign P[129] = in[25] ^ in2[25];
    assign G[130] = in[24] & in2[24];
    assign P[130] = in[24] ^ in2[24];
    assign G[131] = in[23] & in2[23];
    assign P[131] = in[23] ^ in2[23];
    assign G[132] = in[22] & in2[22];
    assign P[132] = in[22] ^ in2[22];
    assign G[133] = in[21] & in2[21];
    assign P[133] = in[21] ^ in2[21];
    assign G[134] = in[20] & in2[20];
    assign P[134] = in[20] ^ in2[20];
    assign G[135] = in[19] & in2[19];
    assign P[135] = in[19] ^ in2[19];
    assign G[136] = in[18] & in2[18];
    assign P[136] = in[18] ^ in2[18];
    assign G[137] = in[17] & in2[17];
    assign P[137] = in[17] ^ in2[17];
    assign G[138] = in[16] & in2[16];
    assign P[138] = in[16] ^ in2[16];
    assign G[139] = in[15] & in2[15];
    assign P[139] = in[15] ^ in2[15];
    assign G[140] = in[14] & in2[14];
    assign P[140] = in[14] ^ in2[14];
    assign G[141] = in[13] & in2[13];
    assign P[141] = in[13] ^ in2[13];
    assign G[142] = in[12] & in2[12];
    assign P[142] = in[12] ^ in2[12];
    assign G[143] = in[11] & in2[11];
    assign P[143] = in[11] ^ in2[11];
    assign G[144] = in[10] & in2[10];
    assign P[144] = in[10] ^ in2[10];
    assign G[145] = in[9] & in2[9];
    assign P[145] = in[9] ^ in2[9];
    assign G[146] = in[8] & in2[8];
    assign P[146] = in[8] ^ in2[8];
    assign G[147] = in[7] & in2[7];
    assign P[147] = in[7] ^ in2[7];
    assign G[148] = in[6] & in2[6];
    assign P[148] = in[6] ^ in2[6];
    assign G[149] = in[5] & in2[5];
    assign P[149] = in[5] ^ in2[5];
    assign G[150] = in[4] & in2[4];
    assign P[150] = in[4] ^ in2[4];
    assign G[151] = in[3] & in2[3];
    assign P[151] = in[3] ^ in2[3];
    assign G[152] = in[2] & in2[2];
    assign P[152] = in[2] ^ in2[2];
    assign G[153] = in[1] & in2[1];
    assign P[153] = in[1] ^ in2[1];
    assign G[154] = in[0] & in2[0];
    assign P[154] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign C[154] = G[153] | (P[153] & C[153]);
    assign cout = G[154] | (P[154] & C[154]);
    assign sum = P ^ C;
endmodule

module CLA154(output [153:0] sum, output cout, input [153:0] in1, input [153:0] in2;

    wire[153:0] G;
    wire[153:0] C;
    wire[153:0] P;

    assign G[0] = in[153] & in2[153];
    assign P[0] = in[153] ^ in2[153];
    assign G[1] = in[152] & in2[152];
    assign P[1] = in[152] ^ in2[152];
    assign G[2] = in[151] & in2[151];
    assign P[2] = in[151] ^ in2[151];
    assign G[3] = in[150] & in2[150];
    assign P[3] = in[150] ^ in2[150];
    assign G[4] = in[149] & in2[149];
    assign P[4] = in[149] ^ in2[149];
    assign G[5] = in[148] & in2[148];
    assign P[5] = in[148] ^ in2[148];
    assign G[6] = in[147] & in2[147];
    assign P[6] = in[147] ^ in2[147];
    assign G[7] = in[146] & in2[146];
    assign P[7] = in[146] ^ in2[146];
    assign G[8] = in[145] & in2[145];
    assign P[8] = in[145] ^ in2[145];
    assign G[9] = in[144] & in2[144];
    assign P[9] = in[144] ^ in2[144];
    assign G[10] = in[143] & in2[143];
    assign P[10] = in[143] ^ in2[143];
    assign G[11] = in[142] & in2[142];
    assign P[11] = in[142] ^ in2[142];
    assign G[12] = in[141] & in2[141];
    assign P[12] = in[141] ^ in2[141];
    assign G[13] = in[140] & in2[140];
    assign P[13] = in[140] ^ in2[140];
    assign G[14] = in[139] & in2[139];
    assign P[14] = in[139] ^ in2[139];
    assign G[15] = in[138] & in2[138];
    assign P[15] = in[138] ^ in2[138];
    assign G[16] = in[137] & in2[137];
    assign P[16] = in[137] ^ in2[137];
    assign G[17] = in[136] & in2[136];
    assign P[17] = in[136] ^ in2[136];
    assign G[18] = in[135] & in2[135];
    assign P[18] = in[135] ^ in2[135];
    assign G[19] = in[134] & in2[134];
    assign P[19] = in[134] ^ in2[134];
    assign G[20] = in[133] & in2[133];
    assign P[20] = in[133] ^ in2[133];
    assign G[21] = in[132] & in2[132];
    assign P[21] = in[132] ^ in2[132];
    assign G[22] = in[131] & in2[131];
    assign P[22] = in[131] ^ in2[131];
    assign G[23] = in[130] & in2[130];
    assign P[23] = in[130] ^ in2[130];
    assign G[24] = in[129] & in2[129];
    assign P[24] = in[129] ^ in2[129];
    assign G[25] = in[128] & in2[128];
    assign P[25] = in[128] ^ in2[128];
    assign G[26] = in[127] & in2[127];
    assign P[26] = in[127] ^ in2[127];
    assign G[27] = in[126] & in2[126];
    assign P[27] = in[126] ^ in2[126];
    assign G[28] = in[125] & in2[125];
    assign P[28] = in[125] ^ in2[125];
    assign G[29] = in[124] & in2[124];
    assign P[29] = in[124] ^ in2[124];
    assign G[30] = in[123] & in2[123];
    assign P[30] = in[123] ^ in2[123];
    assign G[31] = in[122] & in2[122];
    assign P[31] = in[122] ^ in2[122];
    assign G[32] = in[121] & in2[121];
    assign P[32] = in[121] ^ in2[121];
    assign G[33] = in[120] & in2[120];
    assign P[33] = in[120] ^ in2[120];
    assign G[34] = in[119] & in2[119];
    assign P[34] = in[119] ^ in2[119];
    assign G[35] = in[118] & in2[118];
    assign P[35] = in[118] ^ in2[118];
    assign G[36] = in[117] & in2[117];
    assign P[36] = in[117] ^ in2[117];
    assign G[37] = in[116] & in2[116];
    assign P[37] = in[116] ^ in2[116];
    assign G[38] = in[115] & in2[115];
    assign P[38] = in[115] ^ in2[115];
    assign G[39] = in[114] & in2[114];
    assign P[39] = in[114] ^ in2[114];
    assign G[40] = in[113] & in2[113];
    assign P[40] = in[113] ^ in2[113];
    assign G[41] = in[112] & in2[112];
    assign P[41] = in[112] ^ in2[112];
    assign G[42] = in[111] & in2[111];
    assign P[42] = in[111] ^ in2[111];
    assign G[43] = in[110] & in2[110];
    assign P[43] = in[110] ^ in2[110];
    assign G[44] = in[109] & in2[109];
    assign P[44] = in[109] ^ in2[109];
    assign G[45] = in[108] & in2[108];
    assign P[45] = in[108] ^ in2[108];
    assign G[46] = in[107] & in2[107];
    assign P[46] = in[107] ^ in2[107];
    assign G[47] = in[106] & in2[106];
    assign P[47] = in[106] ^ in2[106];
    assign G[48] = in[105] & in2[105];
    assign P[48] = in[105] ^ in2[105];
    assign G[49] = in[104] & in2[104];
    assign P[49] = in[104] ^ in2[104];
    assign G[50] = in[103] & in2[103];
    assign P[50] = in[103] ^ in2[103];
    assign G[51] = in[102] & in2[102];
    assign P[51] = in[102] ^ in2[102];
    assign G[52] = in[101] & in2[101];
    assign P[52] = in[101] ^ in2[101];
    assign G[53] = in[100] & in2[100];
    assign P[53] = in[100] ^ in2[100];
    assign G[54] = in[99] & in2[99];
    assign P[54] = in[99] ^ in2[99];
    assign G[55] = in[98] & in2[98];
    assign P[55] = in[98] ^ in2[98];
    assign G[56] = in[97] & in2[97];
    assign P[56] = in[97] ^ in2[97];
    assign G[57] = in[96] & in2[96];
    assign P[57] = in[96] ^ in2[96];
    assign G[58] = in[95] & in2[95];
    assign P[58] = in[95] ^ in2[95];
    assign G[59] = in[94] & in2[94];
    assign P[59] = in[94] ^ in2[94];
    assign G[60] = in[93] & in2[93];
    assign P[60] = in[93] ^ in2[93];
    assign G[61] = in[92] & in2[92];
    assign P[61] = in[92] ^ in2[92];
    assign G[62] = in[91] & in2[91];
    assign P[62] = in[91] ^ in2[91];
    assign G[63] = in[90] & in2[90];
    assign P[63] = in[90] ^ in2[90];
    assign G[64] = in[89] & in2[89];
    assign P[64] = in[89] ^ in2[89];
    assign G[65] = in[88] & in2[88];
    assign P[65] = in[88] ^ in2[88];
    assign G[66] = in[87] & in2[87];
    assign P[66] = in[87] ^ in2[87];
    assign G[67] = in[86] & in2[86];
    assign P[67] = in[86] ^ in2[86];
    assign G[68] = in[85] & in2[85];
    assign P[68] = in[85] ^ in2[85];
    assign G[69] = in[84] & in2[84];
    assign P[69] = in[84] ^ in2[84];
    assign G[70] = in[83] & in2[83];
    assign P[70] = in[83] ^ in2[83];
    assign G[71] = in[82] & in2[82];
    assign P[71] = in[82] ^ in2[82];
    assign G[72] = in[81] & in2[81];
    assign P[72] = in[81] ^ in2[81];
    assign G[73] = in[80] & in2[80];
    assign P[73] = in[80] ^ in2[80];
    assign G[74] = in[79] & in2[79];
    assign P[74] = in[79] ^ in2[79];
    assign G[75] = in[78] & in2[78];
    assign P[75] = in[78] ^ in2[78];
    assign G[76] = in[77] & in2[77];
    assign P[76] = in[77] ^ in2[77];
    assign G[77] = in[76] & in2[76];
    assign P[77] = in[76] ^ in2[76];
    assign G[78] = in[75] & in2[75];
    assign P[78] = in[75] ^ in2[75];
    assign G[79] = in[74] & in2[74];
    assign P[79] = in[74] ^ in2[74];
    assign G[80] = in[73] & in2[73];
    assign P[80] = in[73] ^ in2[73];
    assign G[81] = in[72] & in2[72];
    assign P[81] = in[72] ^ in2[72];
    assign G[82] = in[71] & in2[71];
    assign P[82] = in[71] ^ in2[71];
    assign G[83] = in[70] & in2[70];
    assign P[83] = in[70] ^ in2[70];
    assign G[84] = in[69] & in2[69];
    assign P[84] = in[69] ^ in2[69];
    assign G[85] = in[68] & in2[68];
    assign P[85] = in[68] ^ in2[68];
    assign G[86] = in[67] & in2[67];
    assign P[86] = in[67] ^ in2[67];
    assign G[87] = in[66] & in2[66];
    assign P[87] = in[66] ^ in2[66];
    assign G[88] = in[65] & in2[65];
    assign P[88] = in[65] ^ in2[65];
    assign G[89] = in[64] & in2[64];
    assign P[89] = in[64] ^ in2[64];
    assign G[90] = in[63] & in2[63];
    assign P[90] = in[63] ^ in2[63];
    assign G[91] = in[62] & in2[62];
    assign P[91] = in[62] ^ in2[62];
    assign G[92] = in[61] & in2[61];
    assign P[92] = in[61] ^ in2[61];
    assign G[93] = in[60] & in2[60];
    assign P[93] = in[60] ^ in2[60];
    assign G[94] = in[59] & in2[59];
    assign P[94] = in[59] ^ in2[59];
    assign G[95] = in[58] & in2[58];
    assign P[95] = in[58] ^ in2[58];
    assign G[96] = in[57] & in2[57];
    assign P[96] = in[57] ^ in2[57];
    assign G[97] = in[56] & in2[56];
    assign P[97] = in[56] ^ in2[56];
    assign G[98] = in[55] & in2[55];
    assign P[98] = in[55] ^ in2[55];
    assign G[99] = in[54] & in2[54];
    assign P[99] = in[54] ^ in2[54];
    assign G[100] = in[53] & in2[53];
    assign P[100] = in[53] ^ in2[53];
    assign G[101] = in[52] & in2[52];
    assign P[101] = in[52] ^ in2[52];
    assign G[102] = in[51] & in2[51];
    assign P[102] = in[51] ^ in2[51];
    assign G[103] = in[50] & in2[50];
    assign P[103] = in[50] ^ in2[50];
    assign G[104] = in[49] & in2[49];
    assign P[104] = in[49] ^ in2[49];
    assign G[105] = in[48] & in2[48];
    assign P[105] = in[48] ^ in2[48];
    assign G[106] = in[47] & in2[47];
    assign P[106] = in[47] ^ in2[47];
    assign G[107] = in[46] & in2[46];
    assign P[107] = in[46] ^ in2[46];
    assign G[108] = in[45] & in2[45];
    assign P[108] = in[45] ^ in2[45];
    assign G[109] = in[44] & in2[44];
    assign P[109] = in[44] ^ in2[44];
    assign G[110] = in[43] & in2[43];
    assign P[110] = in[43] ^ in2[43];
    assign G[111] = in[42] & in2[42];
    assign P[111] = in[42] ^ in2[42];
    assign G[112] = in[41] & in2[41];
    assign P[112] = in[41] ^ in2[41];
    assign G[113] = in[40] & in2[40];
    assign P[113] = in[40] ^ in2[40];
    assign G[114] = in[39] & in2[39];
    assign P[114] = in[39] ^ in2[39];
    assign G[115] = in[38] & in2[38];
    assign P[115] = in[38] ^ in2[38];
    assign G[116] = in[37] & in2[37];
    assign P[116] = in[37] ^ in2[37];
    assign G[117] = in[36] & in2[36];
    assign P[117] = in[36] ^ in2[36];
    assign G[118] = in[35] & in2[35];
    assign P[118] = in[35] ^ in2[35];
    assign G[119] = in[34] & in2[34];
    assign P[119] = in[34] ^ in2[34];
    assign G[120] = in[33] & in2[33];
    assign P[120] = in[33] ^ in2[33];
    assign G[121] = in[32] & in2[32];
    assign P[121] = in[32] ^ in2[32];
    assign G[122] = in[31] & in2[31];
    assign P[122] = in[31] ^ in2[31];
    assign G[123] = in[30] & in2[30];
    assign P[123] = in[30] ^ in2[30];
    assign G[124] = in[29] & in2[29];
    assign P[124] = in[29] ^ in2[29];
    assign G[125] = in[28] & in2[28];
    assign P[125] = in[28] ^ in2[28];
    assign G[126] = in[27] & in2[27];
    assign P[126] = in[27] ^ in2[27];
    assign G[127] = in[26] & in2[26];
    assign P[127] = in[26] ^ in2[26];
    assign G[128] = in[25] & in2[25];
    assign P[128] = in[25] ^ in2[25];
    assign G[129] = in[24] & in2[24];
    assign P[129] = in[24] ^ in2[24];
    assign G[130] = in[23] & in2[23];
    assign P[130] = in[23] ^ in2[23];
    assign G[131] = in[22] & in2[22];
    assign P[131] = in[22] ^ in2[22];
    assign G[132] = in[21] & in2[21];
    assign P[132] = in[21] ^ in2[21];
    assign G[133] = in[20] & in2[20];
    assign P[133] = in[20] ^ in2[20];
    assign G[134] = in[19] & in2[19];
    assign P[134] = in[19] ^ in2[19];
    assign G[135] = in[18] & in2[18];
    assign P[135] = in[18] ^ in2[18];
    assign G[136] = in[17] & in2[17];
    assign P[136] = in[17] ^ in2[17];
    assign G[137] = in[16] & in2[16];
    assign P[137] = in[16] ^ in2[16];
    assign G[138] = in[15] & in2[15];
    assign P[138] = in[15] ^ in2[15];
    assign G[139] = in[14] & in2[14];
    assign P[139] = in[14] ^ in2[14];
    assign G[140] = in[13] & in2[13];
    assign P[140] = in[13] ^ in2[13];
    assign G[141] = in[12] & in2[12];
    assign P[141] = in[12] ^ in2[12];
    assign G[142] = in[11] & in2[11];
    assign P[142] = in[11] ^ in2[11];
    assign G[143] = in[10] & in2[10];
    assign P[143] = in[10] ^ in2[10];
    assign G[144] = in[9] & in2[9];
    assign P[144] = in[9] ^ in2[9];
    assign G[145] = in[8] & in2[8];
    assign P[145] = in[8] ^ in2[8];
    assign G[146] = in[7] & in2[7];
    assign P[146] = in[7] ^ in2[7];
    assign G[147] = in[6] & in2[6];
    assign P[147] = in[6] ^ in2[6];
    assign G[148] = in[5] & in2[5];
    assign P[148] = in[5] ^ in2[5];
    assign G[149] = in[4] & in2[4];
    assign P[149] = in[4] ^ in2[4];
    assign G[150] = in[3] & in2[3];
    assign P[150] = in[3] ^ in2[3];
    assign G[151] = in[2] & in2[2];
    assign P[151] = in[2] ^ in2[2];
    assign G[152] = in[1] & in2[1];
    assign P[152] = in[1] ^ in2[1];
    assign G[153] = in[0] & in2[0];
    assign P[153] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign C[153] = G[152] | (P[152] & C[152]);
    assign cout = G[153] | (P[153] & C[153]);
    assign sum = P ^ C;
endmodule

module CLA153(output [152:0] sum, output cout, input [152:0] in1, input [152:0] in2;

    wire[152:0] G;
    wire[152:0] C;
    wire[152:0] P;

    assign G[0] = in[152] & in2[152];
    assign P[0] = in[152] ^ in2[152];
    assign G[1] = in[151] & in2[151];
    assign P[1] = in[151] ^ in2[151];
    assign G[2] = in[150] & in2[150];
    assign P[2] = in[150] ^ in2[150];
    assign G[3] = in[149] & in2[149];
    assign P[3] = in[149] ^ in2[149];
    assign G[4] = in[148] & in2[148];
    assign P[4] = in[148] ^ in2[148];
    assign G[5] = in[147] & in2[147];
    assign P[5] = in[147] ^ in2[147];
    assign G[6] = in[146] & in2[146];
    assign P[6] = in[146] ^ in2[146];
    assign G[7] = in[145] & in2[145];
    assign P[7] = in[145] ^ in2[145];
    assign G[8] = in[144] & in2[144];
    assign P[8] = in[144] ^ in2[144];
    assign G[9] = in[143] & in2[143];
    assign P[9] = in[143] ^ in2[143];
    assign G[10] = in[142] & in2[142];
    assign P[10] = in[142] ^ in2[142];
    assign G[11] = in[141] & in2[141];
    assign P[11] = in[141] ^ in2[141];
    assign G[12] = in[140] & in2[140];
    assign P[12] = in[140] ^ in2[140];
    assign G[13] = in[139] & in2[139];
    assign P[13] = in[139] ^ in2[139];
    assign G[14] = in[138] & in2[138];
    assign P[14] = in[138] ^ in2[138];
    assign G[15] = in[137] & in2[137];
    assign P[15] = in[137] ^ in2[137];
    assign G[16] = in[136] & in2[136];
    assign P[16] = in[136] ^ in2[136];
    assign G[17] = in[135] & in2[135];
    assign P[17] = in[135] ^ in2[135];
    assign G[18] = in[134] & in2[134];
    assign P[18] = in[134] ^ in2[134];
    assign G[19] = in[133] & in2[133];
    assign P[19] = in[133] ^ in2[133];
    assign G[20] = in[132] & in2[132];
    assign P[20] = in[132] ^ in2[132];
    assign G[21] = in[131] & in2[131];
    assign P[21] = in[131] ^ in2[131];
    assign G[22] = in[130] & in2[130];
    assign P[22] = in[130] ^ in2[130];
    assign G[23] = in[129] & in2[129];
    assign P[23] = in[129] ^ in2[129];
    assign G[24] = in[128] & in2[128];
    assign P[24] = in[128] ^ in2[128];
    assign G[25] = in[127] & in2[127];
    assign P[25] = in[127] ^ in2[127];
    assign G[26] = in[126] & in2[126];
    assign P[26] = in[126] ^ in2[126];
    assign G[27] = in[125] & in2[125];
    assign P[27] = in[125] ^ in2[125];
    assign G[28] = in[124] & in2[124];
    assign P[28] = in[124] ^ in2[124];
    assign G[29] = in[123] & in2[123];
    assign P[29] = in[123] ^ in2[123];
    assign G[30] = in[122] & in2[122];
    assign P[30] = in[122] ^ in2[122];
    assign G[31] = in[121] & in2[121];
    assign P[31] = in[121] ^ in2[121];
    assign G[32] = in[120] & in2[120];
    assign P[32] = in[120] ^ in2[120];
    assign G[33] = in[119] & in2[119];
    assign P[33] = in[119] ^ in2[119];
    assign G[34] = in[118] & in2[118];
    assign P[34] = in[118] ^ in2[118];
    assign G[35] = in[117] & in2[117];
    assign P[35] = in[117] ^ in2[117];
    assign G[36] = in[116] & in2[116];
    assign P[36] = in[116] ^ in2[116];
    assign G[37] = in[115] & in2[115];
    assign P[37] = in[115] ^ in2[115];
    assign G[38] = in[114] & in2[114];
    assign P[38] = in[114] ^ in2[114];
    assign G[39] = in[113] & in2[113];
    assign P[39] = in[113] ^ in2[113];
    assign G[40] = in[112] & in2[112];
    assign P[40] = in[112] ^ in2[112];
    assign G[41] = in[111] & in2[111];
    assign P[41] = in[111] ^ in2[111];
    assign G[42] = in[110] & in2[110];
    assign P[42] = in[110] ^ in2[110];
    assign G[43] = in[109] & in2[109];
    assign P[43] = in[109] ^ in2[109];
    assign G[44] = in[108] & in2[108];
    assign P[44] = in[108] ^ in2[108];
    assign G[45] = in[107] & in2[107];
    assign P[45] = in[107] ^ in2[107];
    assign G[46] = in[106] & in2[106];
    assign P[46] = in[106] ^ in2[106];
    assign G[47] = in[105] & in2[105];
    assign P[47] = in[105] ^ in2[105];
    assign G[48] = in[104] & in2[104];
    assign P[48] = in[104] ^ in2[104];
    assign G[49] = in[103] & in2[103];
    assign P[49] = in[103] ^ in2[103];
    assign G[50] = in[102] & in2[102];
    assign P[50] = in[102] ^ in2[102];
    assign G[51] = in[101] & in2[101];
    assign P[51] = in[101] ^ in2[101];
    assign G[52] = in[100] & in2[100];
    assign P[52] = in[100] ^ in2[100];
    assign G[53] = in[99] & in2[99];
    assign P[53] = in[99] ^ in2[99];
    assign G[54] = in[98] & in2[98];
    assign P[54] = in[98] ^ in2[98];
    assign G[55] = in[97] & in2[97];
    assign P[55] = in[97] ^ in2[97];
    assign G[56] = in[96] & in2[96];
    assign P[56] = in[96] ^ in2[96];
    assign G[57] = in[95] & in2[95];
    assign P[57] = in[95] ^ in2[95];
    assign G[58] = in[94] & in2[94];
    assign P[58] = in[94] ^ in2[94];
    assign G[59] = in[93] & in2[93];
    assign P[59] = in[93] ^ in2[93];
    assign G[60] = in[92] & in2[92];
    assign P[60] = in[92] ^ in2[92];
    assign G[61] = in[91] & in2[91];
    assign P[61] = in[91] ^ in2[91];
    assign G[62] = in[90] & in2[90];
    assign P[62] = in[90] ^ in2[90];
    assign G[63] = in[89] & in2[89];
    assign P[63] = in[89] ^ in2[89];
    assign G[64] = in[88] & in2[88];
    assign P[64] = in[88] ^ in2[88];
    assign G[65] = in[87] & in2[87];
    assign P[65] = in[87] ^ in2[87];
    assign G[66] = in[86] & in2[86];
    assign P[66] = in[86] ^ in2[86];
    assign G[67] = in[85] & in2[85];
    assign P[67] = in[85] ^ in2[85];
    assign G[68] = in[84] & in2[84];
    assign P[68] = in[84] ^ in2[84];
    assign G[69] = in[83] & in2[83];
    assign P[69] = in[83] ^ in2[83];
    assign G[70] = in[82] & in2[82];
    assign P[70] = in[82] ^ in2[82];
    assign G[71] = in[81] & in2[81];
    assign P[71] = in[81] ^ in2[81];
    assign G[72] = in[80] & in2[80];
    assign P[72] = in[80] ^ in2[80];
    assign G[73] = in[79] & in2[79];
    assign P[73] = in[79] ^ in2[79];
    assign G[74] = in[78] & in2[78];
    assign P[74] = in[78] ^ in2[78];
    assign G[75] = in[77] & in2[77];
    assign P[75] = in[77] ^ in2[77];
    assign G[76] = in[76] & in2[76];
    assign P[76] = in[76] ^ in2[76];
    assign G[77] = in[75] & in2[75];
    assign P[77] = in[75] ^ in2[75];
    assign G[78] = in[74] & in2[74];
    assign P[78] = in[74] ^ in2[74];
    assign G[79] = in[73] & in2[73];
    assign P[79] = in[73] ^ in2[73];
    assign G[80] = in[72] & in2[72];
    assign P[80] = in[72] ^ in2[72];
    assign G[81] = in[71] & in2[71];
    assign P[81] = in[71] ^ in2[71];
    assign G[82] = in[70] & in2[70];
    assign P[82] = in[70] ^ in2[70];
    assign G[83] = in[69] & in2[69];
    assign P[83] = in[69] ^ in2[69];
    assign G[84] = in[68] & in2[68];
    assign P[84] = in[68] ^ in2[68];
    assign G[85] = in[67] & in2[67];
    assign P[85] = in[67] ^ in2[67];
    assign G[86] = in[66] & in2[66];
    assign P[86] = in[66] ^ in2[66];
    assign G[87] = in[65] & in2[65];
    assign P[87] = in[65] ^ in2[65];
    assign G[88] = in[64] & in2[64];
    assign P[88] = in[64] ^ in2[64];
    assign G[89] = in[63] & in2[63];
    assign P[89] = in[63] ^ in2[63];
    assign G[90] = in[62] & in2[62];
    assign P[90] = in[62] ^ in2[62];
    assign G[91] = in[61] & in2[61];
    assign P[91] = in[61] ^ in2[61];
    assign G[92] = in[60] & in2[60];
    assign P[92] = in[60] ^ in2[60];
    assign G[93] = in[59] & in2[59];
    assign P[93] = in[59] ^ in2[59];
    assign G[94] = in[58] & in2[58];
    assign P[94] = in[58] ^ in2[58];
    assign G[95] = in[57] & in2[57];
    assign P[95] = in[57] ^ in2[57];
    assign G[96] = in[56] & in2[56];
    assign P[96] = in[56] ^ in2[56];
    assign G[97] = in[55] & in2[55];
    assign P[97] = in[55] ^ in2[55];
    assign G[98] = in[54] & in2[54];
    assign P[98] = in[54] ^ in2[54];
    assign G[99] = in[53] & in2[53];
    assign P[99] = in[53] ^ in2[53];
    assign G[100] = in[52] & in2[52];
    assign P[100] = in[52] ^ in2[52];
    assign G[101] = in[51] & in2[51];
    assign P[101] = in[51] ^ in2[51];
    assign G[102] = in[50] & in2[50];
    assign P[102] = in[50] ^ in2[50];
    assign G[103] = in[49] & in2[49];
    assign P[103] = in[49] ^ in2[49];
    assign G[104] = in[48] & in2[48];
    assign P[104] = in[48] ^ in2[48];
    assign G[105] = in[47] & in2[47];
    assign P[105] = in[47] ^ in2[47];
    assign G[106] = in[46] & in2[46];
    assign P[106] = in[46] ^ in2[46];
    assign G[107] = in[45] & in2[45];
    assign P[107] = in[45] ^ in2[45];
    assign G[108] = in[44] & in2[44];
    assign P[108] = in[44] ^ in2[44];
    assign G[109] = in[43] & in2[43];
    assign P[109] = in[43] ^ in2[43];
    assign G[110] = in[42] & in2[42];
    assign P[110] = in[42] ^ in2[42];
    assign G[111] = in[41] & in2[41];
    assign P[111] = in[41] ^ in2[41];
    assign G[112] = in[40] & in2[40];
    assign P[112] = in[40] ^ in2[40];
    assign G[113] = in[39] & in2[39];
    assign P[113] = in[39] ^ in2[39];
    assign G[114] = in[38] & in2[38];
    assign P[114] = in[38] ^ in2[38];
    assign G[115] = in[37] & in2[37];
    assign P[115] = in[37] ^ in2[37];
    assign G[116] = in[36] & in2[36];
    assign P[116] = in[36] ^ in2[36];
    assign G[117] = in[35] & in2[35];
    assign P[117] = in[35] ^ in2[35];
    assign G[118] = in[34] & in2[34];
    assign P[118] = in[34] ^ in2[34];
    assign G[119] = in[33] & in2[33];
    assign P[119] = in[33] ^ in2[33];
    assign G[120] = in[32] & in2[32];
    assign P[120] = in[32] ^ in2[32];
    assign G[121] = in[31] & in2[31];
    assign P[121] = in[31] ^ in2[31];
    assign G[122] = in[30] & in2[30];
    assign P[122] = in[30] ^ in2[30];
    assign G[123] = in[29] & in2[29];
    assign P[123] = in[29] ^ in2[29];
    assign G[124] = in[28] & in2[28];
    assign P[124] = in[28] ^ in2[28];
    assign G[125] = in[27] & in2[27];
    assign P[125] = in[27] ^ in2[27];
    assign G[126] = in[26] & in2[26];
    assign P[126] = in[26] ^ in2[26];
    assign G[127] = in[25] & in2[25];
    assign P[127] = in[25] ^ in2[25];
    assign G[128] = in[24] & in2[24];
    assign P[128] = in[24] ^ in2[24];
    assign G[129] = in[23] & in2[23];
    assign P[129] = in[23] ^ in2[23];
    assign G[130] = in[22] & in2[22];
    assign P[130] = in[22] ^ in2[22];
    assign G[131] = in[21] & in2[21];
    assign P[131] = in[21] ^ in2[21];
    assign G[132] = in[20] & in2[20];
    assign P[132] = in[20] ^ in2[20];
    assign G[133] = in[19] & in2[19];
    assign P[133] = in[19] ^ in2[19];
    assign G[134] = in[18] & in2[18];
    assign P[134] = in[18] ^ in2[18];
    assign G[135] = in[17] & in2[17];
    assign P[135] = in[17] ^ in2[17];
    assign G[136] = in[16] & in2[16];
    assign P[136] = in[16] ^ in2[16];
    assign G[137] = in[15] & in2[15];
    assign P[137] = in[15] ^ in2[15];
    assign G[138] = in[14] & in2[14];
    assign P[138] = in[14] ^ in2[14];
    assign G[139] = in[13] & in2[13];
    assign P[139] = in[13] ^ in2[13];
    assign G[140] = in[12] & in2[12];
    assign P[140] = in[12] ^ in2[12];
    assign G[141] = in[11] & in2[11];
    assign P[141] = in[11] ^ in2[11];
    assign G[142] = in[10] & in2[10];
    assign P[142] = in[10] ^ in2[10];
    assign G[143] = in[9] & in2[9];
    assign P[143] = in[9] ^ in2[9];
    assign G[144] = in[8] & in2[8];
    assign P[144] = in[8] ^ in2[8];
    assign G[145] = in[7] & in2[7];
    assign P[145] = in[7] ^ in2[7];
    assign G[146] = in[6] & in2[6];
    assign P[146] = in[6] ^ in2[6];
    assign G[147] = in[5] & in2[5];
    assign P[147] = in[5] ^ in2[5];
    assign G[148] = in[4] & in2[4];
    assign P[148] = in[4] ^ in2[4];
    assign G[149] = in[3] & in2[3];
    assign P[149] = in[3] ^ in2[3];
    assign G[150] = in[2] & in2[2];
    assign P[150] = in[2] ^ in2[2];
    assign G[151] = in[1] & in2[1];
    assign P[151] = in[1] ^ in2[1];
    assign G[152] = in[0] & in2[0];
    assign P[152] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign C[152] = G[151] | (P[151] & C[151]);
    assign cout = G[152] | (P[152] & C[152]);
    assign sum = P ^ C;
endmodule

module CLA152(output [151:0] sum, output cout, input [151:0] in1, input [151:0] in2;

    wire[151:0] G;
    wire[151:0] C;
    wire[151:0] P;

    assign G[0] = in[151] & in2[151];
    assign P[0] = in[151] ^ in2[151];
    assign G[1] = in[150] & in2[150];
    assign P[1] = in[150] ^ in2[150];
    assign G[2] = in[149] & in2[149];
    assign P[2] = in[149] ^ in2[149];
    assign G[3] = in[148] & in2[148];
    assign P[3] = in[148] ^ in2[148];
    assign G[4] = in[147] & in2[147];
    assign P[4] = in[147] ^ in2[147];
    assign G[5] = in[146] & in2[146];
    assign P[5] = in[146] ^ in2[146];
    assign G[6] = in[145] & in2[145];
    assign P[6] = in[145] ^ in2[145];
    assign G[7] = in[144] & in2[144];
    assign P[7] = in[144] ^ in2[144];
    assign G[8] = in[143] & in2[143];
    assign P[8] = in[143] ^ in2[143];
    assign G[9] = in[142] & in2[142];
    assign P[9] = in[142] ^ in2[142];
    assign G[10] = in[141] & in2[141];
    assign P[10] = in[141] ^ in2[141];
    assign G[11] = in[140] & in2[140];
    assign P[11] = in[140] ^ in2[140];
    assign G[12] = in[139] & in2[139];
    assign P[12] = in[139] ^ in2[139];
    assign G[13] = in[138] & in2[138];
    assign P[13] = in[138] ^ in2[138];
    assign G[14] = in[137] & in2[137];
    assign P[14] = in[137] ^ in2[137];
    assign G[15] = in[136] & in2[136];
    assign P[15] = in[136] ^ in2[136];
    assign G[16] = in[135] & in2[135];
    assign P[16] = in[135] ^ in2[135];
    assign G[17] = in[134] & in2[134];
    assign P[17] = in[134] ^ in2[134];
    assign G[18] = in[133] & in2[133];
    assign P[18] = in[133] ^ in2[133];
    assign G[19] = in[132] & in2[132];
    assign P[19] = in[132] ^ in2[132];
    assign G[20] = in[131] & in2[131];
    assign P[20] = in[131] ^ in2[131];
    assign G[21] = in[130] & in2[130];
    assign P[21] = in[130] ^ in2[130];
    assign G[22] = in[129] & in2[129];
    assign P[22] = in[129] ^ in2[129];
    assign G[23] = in[128] & in2[128];
    assign P[23] = in[128] ^ in2[128];
    assign G[24] = in[127] & in2[127];
    assign P[24] = in[127] ^ in2[127];
    assign G[25] = in[126] & in2[126];
    assign P[25] = in[126] ^ in2[126];
    assign G[26] = in[125] & in2[125];
    assign P[26] = in[125] ^ in2[125];
    assign G[27] = in[124] & in2[124];
    assign P[27] = in[124] ^ in2[124];
    assign G[28] = in[123] & in2[123];
    assign P[28] = in[123] ^ in2[123];
    assign G[29] = in[122] & in2[122];
    assign P[29] = in[122] ^ in2[122];
    assign G[30] = in[121] & in2[121];
    assign P[30] = in[121] ^ in2[121];
    assign G[31] = in[120] & in2[120];
    assign P[31] = in[120] ^ in2[120];
    assign G[32] = in[119] & in2[119];
    assign P[32] = in[119] ^ in2[119];
    assign G[33] = in[118] & in2[118];
    assign P[33] = in[118] ^ in2[118];
    assign G[34] = in[117] & in2[117];
    assign P[34] = in[117] ^ in2[117];
    assign G[35] = in[116] & in2[116];
    assign P[35] = in[116] ^ in2[116];
    assign G[36] = in[115] & in2[115];
    assign P[36] = in[115] ^ in2[115];
    assign G[37] = in[114] & in2[114];
    assign P[37] = in[114] ^ in2[114];
    assign G[38] = in[113] & in2[113];
    assign P[38] = in[113] ^ in2[113];
    assign G[39] = in[112] & in2[112];
    assign P[39] = in[112] ^ in2[112];
    assign G[40] = in[111] & in2[111];
    assign P[40] = in[111] ^ in2[111];
    assign G[41] = in[110] & in2[110];
    assign P[41] = in[110] ^ in2[110];
    assign G[42] = in[109] & in2[109];
    assign P[42] = in[109] ^ in2[109];
    assign G[43] = in[108] & in2[108];
    assign P[43] = in[108] ^ in2[108];
    assign G[44] = in[107] & in2[107];
    assign P[44] = in[107] ^ in2[107];
    assign G[45] = in[106] & in2[106];
    assign P[45] = in[106] ^ in2[106];
    assign G[46] = in[105] & in2[105];
    assign P[46] = in[105] ^ in2[105];
    assign G[47] = in[104] & in2[104];
    assign P[47] = in[104] ^ in2[104];
    assign G[48] = in[103] & in2[103];
    assign P[48] = in[103] ^ in2[103];
    assign G[49] = in[102] & in2[102];
    assign P[49] = in[102] ^ in2[102];
    assign G[50] = in[101] & in2[101];
    assign P[50] = in[101] ^ in2[101];
    assign G[51] = in[100] & in2[100];
    assign P[51] = in[100] ^ in2[100];
    assign G[52] = in[99] & in2[99];
    assign P[52] = in[99] ^ in2[99];
    assign G[53] = in[98] & in2[98];
    assign P[53] = in[98] ^ in2[98];
    assign G[54] = in[97] & in2[97];
    assign P[54] = in[97] ^ in2[97];
    assign G[55] = in[96] & in2[96];
    assign P[55] = in[96] ^ in2[96];
    assign G[56] = in[95] & in2[95];
    assign P[56] = in[95] ^ in2[95];
    assign G[57] = in[94] & in2[94];
    assign P[57] = in[94] ^ in2[94];
    assign G[58] = in[93] & in2[93];
    assign P[58] = in[93] ^ in2[93];
    assign G[59] = in[92] & in2[92];
    assign P[59] = in[92] ^ in2[92];
    assign G[60] = in[91] & in2[91];
    assign P[60] = in[91] ^ in2[91];
    assign G[61] = in[90] & in2[90];
    assign P[61] = in[90] ^ in2[90];
    assign G[62] = in[89] & in2[89];
    assign P[62] = in[89] ^ in2[89];
    assign G[63] = in[88] & in2[88];
    assign P[63] = in[88] ^ in2[88];
    assign G[64] = in[87] & in2[87];
    assign P[64] = in[87] ^ in2[87];
    assign G[65] = in[86] & in2[86];
    assign P[65] = in[86] ^ in2[86];
    assign G[66] = in[85] & in2[85];
    assign P[66] = in[85] ^ in2[85];
    assign G[67] = in[84] & in2[84];
    assign P[67] = in[84] ^ in2[84];
    assign G[68] = in[83] & in2[83];
    assign P[68] = in[83] ^ in2[83];
    assign G[69] = in[82] & in2[82];
    assign P[69] = in[82] ^ in2[82];
    assign G[70] = in[81] & in2[81];
    assign P[70] = in[81] ^ in2[81];
    assign G[71] = in[80] & in2[80];
    assign P[71] = in[80] ^ in2[80];
    assign G[72] = in[79] & in2[79];
    assign P[72] = in[79] ^ in2[79];
    assign G[73] = in[78] & in2[78];
    assign P[73] = in[78] ^ in2[78];
    assign G[74] = in[77] & in2[77];
    assign P[74] = in[77] ^ in2[77];
    assign G[75] = in[76] & in2[76];
    assign P[75] = in[76] ^ in2[76];
    assign G[76] = in[75] & in2[75];
    assign P[76] = in[75] ^ in2[75];
    assign G[77] = in[74] & in2[74];
    assign P[77] = in[74] ^ in2[74];
    assign G[78] = in[73] & in2[73];
    assign P[78] = in[73] ^ in2[73];
    assign G[79] = in[72] & in2[72];
    assign P[79] = in[72] ^ in2[72];
    assign G[80] = in[71] & in2[71];
    assign P[80] = in[71] ^ in2[71];
    assign G[81] = in[70] & in2[70];
    assign P[81] = in[70] ^ in2[70];
    assign G[82] = in[69] & in2[69];
    assign P[82] = in[69] ^ in2[69];
    assign G[83] = in[68] & in2[68];
    assign P[83] = in[68] ^ in2[68];
    assign G[84] = in[67] & in2[67];
    assign P[84] = in[67] ^ in2[67];
    assign G[85] = in[66] & in2[66];
    assign P[85] = in[66] ^ in2[66];
    assign G[86] = in[65] & in2[65];
    assign P[86] = in[65] ^ in2[65];
    assign G[87] = in[64] & in2[64];
    assign P[87] = in[64] ^ in2[64];
    assign G[88] = in[63] & in2[63];
    assign P[88] = in[63] ^ in2[63];
    assign G[89] = in[62] & in2[62];
    assign P[89] = in[62] ^ in2[62];
    assign G[90] = in[61] & in2[61];
    assign P[90] = in[61] ^ in2[61];
    assign G[91] = in[60] & in2[60];
    assign P[91] = in[60] ^ in2[60];
    assign G[92] = in[59] & in2[59];
    assign P[92] = in[59] ^ in2[59];
    assign G[93] = in[58] & in2[58];
    assign P[93] = in[58] ^ in2[58];
    assign G[94] = in[57] & in2[57];
    assign P[94] = in[57] ^ in2[57];
    assign G[95] = in[56] & in2[56];
    assign P[95] = in[56] ^ in2[56];
    assign G[96] = in[55] & in2[55];
    assign P[96] = in[55] ^ in2[55];
    assign G[97] = in[54] & in2[54];
    assign P[97] = in[54] ^ in2[54];
    assign G[98] = in[53] & in2[53];
    assign P[98] = in[53] ^ in2[53];
    assign G[99] = in[52] & in2[52];
    assign P[99] = in[52] ^ in2[52];
    assign G[100] = in[51] & in2[51];
    assign P[100] = in[51] ^ in2[51];
    assign G[101] = in[50] & in2[50];
    assign P[101] = in[50] ^ in2[50];
    assign G[102] = in[49] & in2[49];
    assign P[102] = in[49] ^ in2[49];
    assign G[103] = in[48] & in2[48];
    assign P[103] = in[48] ^ in2[48];
    assign G[104] = in[47] & in2[47];
    assign P[104] = in[47] ^ in2[47];
    assign G[105] = in[46] & in2[46];
    assign P[105] = in[46] ^ in2[46];
    assign G[106] = in[45] & in2[45];
    assign P[106] = in[45] ^ in2[45];
    assign G[107] = in[44] & in2[44];
    assign P[107] = in[44] ^ in2[44];
    assign G[108] = in[43] & in2[43];
    assign P[108] = in[43] ^ in2[43];
    assign G[109] = in[42] & in2[42];
    assign P[109] = in[42] ^ in2[42];
    assign G[110] = in[41] & in2[41];
    assign P[110] = in[41] ^ in2[41];
    assign G[111] = in[40] & in2[40];
    assign P[111] = in[40] ^ in2[40];
    assign G[112] = in[39] & in2[39];
    assign P[112] = in[39] ^ in2[39];
    assign G[113] = in[38] & in2[38];
    assign P[113] = in[38] ^ in2[38];
    assign G[114] = in[37] & in2[37];
    assign P[114] = in[37] ^ in2[37];
    assign G[115] = in[36] & in2[36];
    assign P[115] = in[36] ^ in2[36];
    assign G[116] = in[35] & in2[35];
    assign P[116] = in[35] ^ in2[35];
    assign G[117] = in[34] & in2[34];
    assign P[117] = in[34] ^ in2[34];
    assign G[118] = in[33] & in2[33];
    assign P[118] = in[33] ^ in2[33];
    assign G[119] = in[32] & in2[32];
    assign P[119] = in[32] ^ in2[32];
    assign G[120] = in[31] & in2[31];
    assign P[120] = in[31] ^ in2[31];
    assign G[121] = in[30] & in2[30];
    assign P[121] = in[30] ^ in2[30];
    assign G[122] = in[29] & in2[29];
    assign P[122] = in[29] ^ in2[29];
    assign G[123] = in[28] & in2[28];
    assign P[123] = in[28] ^ in2[28];
    assign G[124] = in[27] & in2[27];
    assign P[124] = in[27] ^ in2[27];
    assign G[125] = in[26] & in2[26];
    assign P[125] = in[26] ^ in2[26];
    assign G[126] = in[25] & in2[25];
    assign P[126] = in[25] ^ in2[25];
    assign G[127] = in[24] & in2[24];
    assign P[127] = in[24] ^ in2[24];
    assign G[128] = in[23] & in2[23];
    assign P[128] = in[23] ^ in2[23];
    assign G[129] = in[22] & in2[22];
    assign P[129] = in[22] ^ in2[22];
    assign G[130] = in[21] & in2[21];
    assign P[130] = in[21] ^ in2[21];
    assign G[131] = in[20] & in2[20];
    assign P[131] = in[20] ^ in2[20];
    assign G[132] = in[19] & in2[19];
    assign P[132] = in[19] ^ in2[19];
    assign G[133] = in[18] & in2[18];
    assign P[133] = in[18] ^ in2[18];
    assign G[134] = in[17] & in2[17];
    assign P[134] = in[17] ^ in2[17];
    assign G[135] = in[16] & in2[16];
    assign P[135] = in[16] ^ in2[16];
    assign G[136] = in[15] & in2[15];
    assign P[136] = in[15] ^ in2[15];
    assign G[137] = in[14] & in2[14];
    assign P[137] = in[14] ^ in2[14];
    assign G[138] = in[13] & in2[13];
    assign P[138] = in[13] ^ in2[13];
    assign G[139] = in[12] & in2[12];
    assign P[139] = in[12] ^ in2[12];
    assign G[140] = in[11] & in2[11];
    assign P[140] = in[11] ^ in2[11];
    assign G[141] = in[10] & in2[10];
    assign P[141] = in[10] ^ in2[10];
    assign G[142] = in[9] & in2[9];
    assign P[142] = in[9] ^ in2[9];
    assign G[143] = in[8] & in2[8];
    assign P[143] = in[8] ^ in2[8];
    assign G[144] = in[7] & in2[7];
    assign P[144] = in[7] ^ in2[7];
    assign G[145] = in[6] & in2[6];
    assign P[145] = in[6] ^ in2[6];
    assign G[146] = in[5] & in2[5];
    assign P[146] = in[5] ^ in2[5];
    assign G[147] = in[4] & in2[4];
    assign P[147] = in[4] ^ in2[4];
    assign G[148] = in[3] & in2[3];
    assign P[148] = in[3] ^ in2[3];
    assign G[149] = in[2] & in2[2];
    assign P[149] = in[2] ^ in2[2];
    assign G[150] = in[1] & in2[1];
    assign P[150] = in[1] ^ in2[1];
    assign G[151] = in[0] & in2[0];
    assign P[151] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign C[151] = G[150] | (P[150] & C[150]);
    assign cout = G[151] | (P[151] & C[151]);
    assign sum = P ^ C;
endmodule

module CLA151(output [150:0] sum, output cout, input [150:0] in1, input [150:0] in2;

    wire[150:0] G;
    wire[150:0] C;
    wire[150:0] P;

    assign G[0] = in[150] & in2[150];
    assign P[0] = in[150] ^ in2[150];
    assign G[1] = in[149] & in2[149];
    assign P[1] = in[149] ^ in2[149];
    assign G[2] = in[148] & in2[148];
    assign P[2] = in[148] ^ in2[148];
    assign G[3] = in[147] & in2[147];
    assign P[3] = in[147] ^ in2[147];
    assign G[4] = in[146] & in2[146];
    assign P[4] = in[146] ^ in2[146];
    assign G[5] = in[145] & in2[145];
    assign P[5] = in[145] ^ in2[145];
    assign G[6] = in[144] & in2[144];
    assign P[6] = in[144] ^ in2[144];
    assign G[7] = in[143] & in2[143];
    assign P[7] = in[143] ^ in2[143];
    assign G[8] = in[142] & in2[142];
    assign P[8] = in[142] ^ in2[142];
    assign G[9] = in[141] & in2[141];
    assign P[9] = in[141] ^ in2[141];
    assign G[10] = in[140] & in2[140];
    assign P[10] = in[140] ^ in2[140];
    assign G[11] = in[139] & in2[139];
    assign P[11] = in[139] ^ in2[139];
    assign G[12] = in[138] & in2[138];
    assign P[12] = in[138] ^ in2[138];
    assign G[13] = in[137] & in2[137];
    assign P[13] = in[137] ^ in2[137];
    assign G[14] = in[136] & in2[136];
    assign P[14] = in[136] ^ in2[136];
    assign G[15] = in[135] & in2[135];
    assign P[15] = in[135] ^ in2[135];
    assign G[16] = in[134] & in2[134];
    assign P[16] = in[134] ^ in2[134];
    assign G[17] = in[133] & in2[133];
    assign P[17] = in[133] ^ in2[133];
    assign G[18] = in[132] & in2[132];
    assign P[18] = in[132] ^ in2[132];
    assign G[19] = in[131] & in2[131];
    assign P[19] = in[131] ^ in2[131];
    assign G[20] = in[130] & in2[130];
    assign P[20] = in[130] ^ in2[130];
    assign G[21] = in[129] & in2[129];
    assign P[21] = in[129] ^ in2[129];
    assign G[22] = in[128] & in2[128];
    assign P[22] = in[128] ^ in2[128];
    assign G[23] = in[127] & in2[127];
    assign P[23] = in[127] ^ in2[127];
    assign G[24] = in[126] & in2[126];
    assign P[24] = in[126] ^ in2[126];
    assign G[25] = in[125] & in2[125];
    assign P[25] = in[125] ^ in2[125];
    assign G[26] = in[124] & in2[124];
    assign P[26] = in[124] ^ in2[124];
    assign G[27] = in[123] & in2[123];
    assign P[27] = in[123] ^ in2[123];
    assign G[28] = in[122] & in2[122];
    assign P[28] = in[122] ^ in2[122];
    assign G[29] = in[121] & in2[121];
    assign P[29] = in[121] ^ in2[121];
    assign G[30] = in[120] & in2[120];
    assign P[30] = in[120] ^ in2[120];
    assign G[31] = in[119] & in2[119];
    assign P[31] = in[119] ^ in2[119];
    assign G[32] = in[118] & in2[118];
    assign P[32] = in[118] ^ in2[118];
    assign G[33] = in[117] & in2[117];
    assign P[33] = in[117] ^ in2[117];
    assign G[34] = in[116] & in2[116];
    assign P[34] = in[116] ^ in2[116];
    assign G[35] = in[115] & in2[115];
    assign P[35] = in[115] ^ in2[115];
    assign G[36] = in[114] & in2[114];
    assign P[36] = in[114] ^ in2[114];
    assign G[37] = in[113] & in2[113];
    assign P[37] = in[113] ^ in2[113];
    assign G[38] = in[112] & in2[112];
    assign P[38] = in[112] ^ in2[112];
    assign G[39] = in[111] & in2[111];
    assign P[39] = in[111] ^ in2[111];
    assign G[40] = in[110] & in2[110];
    assign P[40] = in[110] ^ in2[110];
    assign G[41] = in[109] & in2[109];
    assign P[41] = in[109] ^ in2[109];
    assign G[42] = in[108] & in2[108];
    assign P[42] = in[108] ^ in2[108];
    assign G[43] = in[107] & in2[107];
    assign P[43] = in[107] ^ in2[107];
    assign G[44] = in[106] & in2[106];
    assign P[44] = in[106] ^ in2[106];
    assign G[45] = in[105] & in2[105];
    assign P[45] = in[105] ^ in2[105];
    assign G[46] = in[104] & in2[104];
    assign P[46] = in[104] ^ in2[104];
    assign G[47] = in[103] & in2[103];
    assign P[47] = in[103] ^ in2[103];
    assign G[48] = in[102] & in2[102];
    assign P[48] = in[102] ^ in2[102];
    assign G[49] = in[101] & in2[101];
    assign P[49] = in[101] ^ in2[101];
    assign G[50] = in[100] & in2[100];
    assign P[50] = in[100] ^ in2[100];
    assign G[51] = in[99] & in2[99];
    assign P[51] = in[99] ^ in2[99];
    assign G[52] = in[98] & in2[98];
    assign P[52] = in[98] ^ in2[98];
    assign G[53] = in[97] & in2[97];
    assign P[53] = in[97] ^ in2[97];
    assign G[54] = in[96] & in2[96];
    assign P[54] = in[96] ^ in2[96];
    assign G[55] = in[95] & in2[95];
    assign P[55] = in[95] ^ in2[95];
    assign G[56] = in[94] & in2[94];
    assign P[56] = in[94] ^ in2[94];
    assign G[57] = in[93] & in2[93];
    assign P[57] = in[93] ^ in2[93];
    assign G[58] = in[92] & in2[92];
    assign P[58] = in[92] ^ in2[92];
    assign G[59] = in[91] & in2[91];
    assign P[59] = in[91] ^ in2[91];
    assign G[60] = in[90] & in2[90];
    assign P[60] = in[90] ^ in2[90];
    assign G[61] = in[89] & in2[89];
    assign P[61] = in[89] ^ in2[89];
    assign G[62] = in[88] & in2[88];
    assign P[62] = in[88] ^ in2[88];
    assign G[63] = in[87] & in2[87];
    assign P[63] = in[87] ^ in2[87];
    assign G[64] = in[86] & in2[86];
    assign P[64] = in[86] ^ in2[86];
    assign G[65] = in[85] & in2[85];
    assign P[65] = in[85] ^ in2[85];
    assign G[66] = in[84] & in2[84];
    assign P[66] = in[84] ^ in2[84];
    assign G[67] = in[83] & in2[83];
    assign P[67] = in[83] ^ in2[83];
    assign G[68] = in[82] & in2[82];
    assign P[68] = in[82] ^ in2[82];
    assign G[69] = in[81] & in2[81];
    assign P[69] = in[81] ^ in2[81];
    assign G[70] = in[80] & in2[80];
    assign P[70] = in[80] ^ in2[80];
    assign G[71] = in[79] & in2[79];
    assign P[71] = in[79] ^ in2[79];
    assign G[72] = in[78] & in2[78];
    assign P[72] = in[78] ^ in2[78];
    assign G[73] = in[77] & in2[77];
    assign P[73] = in[77] ^ in2[77];
    assign G[74] = in[76] & in2[76];
    assign P[74] = in[76] ^ in2[76];
    assign G[75] = in[75] & in2[75];
    assign P[75] = in[75] ^ in2[75];
    assign G[76] = in[74] & in2[74];
    assign P[76] = in[74] ^ in2[74];
    assign G[77] = in[73] & in2[73];
    assign P[77] = in[73] ^ in2[73];
    assign G[78] = in[72] & in2[72];
    assign P[78] = in[72] ^ in2[72];
    assign G[79] = in[71] & in2[71];
    assign P[79] = in[71] ^ in2[71];
    assign G[80] = in[70] & in2[70];
    assign P[80] = in[70] ^ in2[70];
    assign G[81] = in[69] & in2[69];
    assign P[81] = in[69] ^ in2[69];
    assign G[82] = in[68] & in2[68];
    assign P[82] = in[68] ^ in2[68];
    assign G[83] = in[67] & in2[67];
    assign P[83] = in[67] ^ in2[67];
    assign G[84] = in[66] & in2[66];
    assign P[84] = in[66] ^ in2[66];
    assign G[85] = in[65] & in2[65];
    assign P[85] = in[65] ^ in2[65];
    assign G[86] = in[64] & in2[64];
    assign P[86] = in[64] ^ in2[64];
    assign G[87] = in[63] & in2[63];
    assign P[87] = in[63] ^ in2[63];
    assign G[88] = in[62] & in2[62];
    assign P[88] = in[62] ^ in2[62];
    assign G[89] = in[61] & in2[61];
    assign P[89] = in[61] ^ in2[61];
    assign G[90] = in[60] & in2[60];
    assign P[90] = in[60] ^ in2[60];
    assign G[91] = in[59] & in2[59];
    assign P[91] = in[59] ^ in2[59];
    assign G[92] = in[58] & in2[58];
    assign P[92] = in[58] ^ in2[58];
    assign G[93] = in[57] & in2[57];
    assign P[93] = in[57] ^ in2[57];
    assign G[94] = in[56] & in2[56];
    assign P[94] = in[56] ^ in2[56];
    assign G[95] = in[55] & in2[55];
    assign P[95] = in[55] ^ in2[55];
    assign G[96] = in[54] & in2[54];
    assign P[96] = in[54] ^ in2[54];
    assign G[97] = in[53] & in2[53];
    assign P[97] = in[53] ^ in2[53];
    assign G[98] = in[52] & in2[52];
    assign P[98] = in[52] ^ in2[52];
    assign G[99] = in[51] & in2[51];
    assign P[99] = in[51] ^ in2[51];
    assign G[100] = in[50] & in2[50];
    assign P[100] = in[50] ^ in2[50];
    assign G[101] = in[49] & in2[49];
    assign P[101] = in[49] ^ in2[49];
    assign G[102] = in[48] & in2[48];
    assign P[102] = in[48] ^ in2[48];
    assign G[103] = in[47] & in2[47];
    assign P[103] = in[47] ^ in2[47];
    assign G[104] = in[46] & in2[46];
    assign P[104] = in[46] ^ in2[46];
    assign G[105] = in[45] & in2[45];
    assign P[105] = in[45] ^ in2[45];
    assign G[106] = in[44] & in2[44];
    assign P[106] = in[44] ^ in2[44];
    assign G[107] = in[43] & in2[43];
    assign P[107] = in[43] ^ in2[43];
    assign G[108] = in[42] & in2[42];
    assign P[108] = in[42] ^ in2[42];
    assign G[109] = in[41] & in2[41];
    assign P[109] = in[41] ^ in2[41];
    assign G[110] = in[40] & in2[40];
    assign P[110] = in[40] ^ in2[40];
    assign G[111] = in[39] & in2[39];
    assign P[111] = in[39] ^ in2[39];
    assign G[112] = in[38] & in2[38];
    assign P[112] = in[38] ^ in2[38];
    assign G[113] = in[37] & in2[37];
    assign P[113] = in[37] ^ in2[37];
    assign G[114] = in[36] & in2[36];
    assign P[114] = in[36] ^ in2[36];
    assign G[115] = in[35] & in2[35];
    assign P[115] = in[35] ^ in2[35];
    assign G[116] = in[34] & in2[34];
    assign P[116] = in[34] ^ in2[34];
    assign G[117] = in[33] & in2[33];
    assign P[117] = in[33] ^ in2[33];
    assign G[118] = in[32] & in2[32];
    assign P[118] = in[32] ^ in2[32];
    assign G[119] = in[31] & in2[31];
    assign P[119] = in[31] ^ in2[31];
    assign G[120] = in[30] & in2[30];
    assign P[120] = in[30] ^ in2[30];
    assign G[121] = in[29] & in2[29];
    assign P[121] = in[29] ^ in2[29];
    assign G[122] = in[28] & in2[28];
    assign P[122] = in[28] ^ in2[28];
    assign G[123] = in[27] & in2[27];
    assign P[123] = in[27] ^ in2[27];
    assign G[124] = in[26] & in2[26];
    assign P[124] = in[26] ^ in2[26];
    assign G[125] = in[25] & in2[25];
    assign P[125] = in[25] ^ in2[25];
    assign G[126] = in[24] & in2[24];
    assign P[126] = in[24] ^ in2[24];
    assign G[127] = in[23] & in2[23];
    assign P[127] = in[23] ^ in2[23];
    assign G[128] = in[22] & in2[22];
    assign P[128] = in[22] ^ in2[22];
    assign G[129] = in[21] & in2[21];
    assign P[129] = in[21] ^ in2[21];
    assign G[130] = in[20] & in2[20];
    assign P[130] = in[20] ^ in2[20];
    assign G[131] = in[19] & in2[19];
    assign P[131] = in[19] ^ in2[19];
    assign G[132] = in[18] & in2[18];
    assign P[132] = in[18] ^ in2[18];
    assign G[133] = in[17] & in2[17];
    assign P[133] = in[17] ^ in2[17];
    assign G[134] = in[16] & in2[16];
    assign P[134] = in[16] ^ in2[16];
    assign G[135] = in[15] & in2[15];
    assign P[135] = in[15] ^ in2[15];
    assign G[136] = in[14] & in2[14];
    assign P[136] = in[14] ^ in2[14];
    assign G[137] = in[13] & in2[13];
    assign P[137] = in[13] ^ in2[13];
    assign G[138] = in[12] & in2[12];
    assign P[138] = in[12] ^ in2[12];
    assign G[139] = in[11] & in2[11];
    assign P[139] = in[11] ^ in2[11];
    assign G[140] = in[10] & in2[10];
    assign P[140] = in[10] ^ in2[10];
    assign G[141] = in[9] & in2[9];
    assign P[141] = in[9] ^ in2[9];
    assign G[142] = in[8] & in2[8];
    assign P[142] = in[8] ^ in2[8];
    assign G[143] = in[7] & in2[7];
    assign P[143] = in[7] ^ in2[7];
    assign G[144] = in[6] & in2[6];
    assign P[144] = in[6] ^ in2[6];
    assign G[145] = in[5] & in2[5];
    assign P[145] = in[5] ^ in2[5];
    assign G[146] = in[4] & in2[4];
    assign P[146] = in[4] ^ in2[4];
    assign G[147] = in[3] & in2[3];
    assign P[147] = in[3] ^ in2[3];
    assign G[148] = in[2] & in2[2];
    assign P[148] = in[2] ^ in2[2];
    assign G[149] = in[1] & in2[1];
    assign P[149] = in[1] ^ in2[1];
    assign G[150] = in[0] & in2[0];
    assign P[150] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign C[150] = G[149] | (P[149] & C[149]);
    assign cout = G[150] | (P[150] & C[150]);
    assign sum = P ^ C;
endmodule

module CLA150(output [149:0] sum, output cout, input [149:0] in1, input [149:0] in2;

    wire[149:0] G;
    wire[149:0] C;
    wire[149:0] P;

    assign G[0] = in[149] & in2[149];
    assign P[0] = in[149] ^ in2[149];
    assign G[1] = in[148] & in2[148];
    assign P[1] = in[148] ^ in2[148];
    assign G[2] = in[147] & in2[147];
    assign P[2] = in[147] ^ in2[147];
    assign G[3] = in[146] & in2[146];
    assign P[3] = in[146] ^ in2[146];
    assign G[4] = in[145] & in2[145];
    assign P[4] = in[145] ^ in2[145];
    assign G[5] = in[144] & in2[144];
    assign P[5] = in[144] ^ in2[144];
    assign G[6] = in[143] & in2[143];
    assign P[6] = in[143] ^ in2[143];
    assign G[7] = in[142] & in2[142];
    assign P[7] = in[142] ^ in2[142];
    assign G[8] = in[141] & in2[141];
    assign P[8] = in[141] ^ in2[141];
    assign G[9] = in[140] & in2[140];
    assign P[9] = in[140] ^ in2[140];
    assign G[10] = in[139] & in2[139];
    assign P[10] = in[139] ^ in2[139];
    assign G[11] = in[138] & in2[138];
    assign P[11] = in[138] ^ in2[138];
    assign G[12] = in[137] & in2[137];
    assign P[12] = in[137] ^ in2[137];
    assign G[13] = in[136] & in2[136];
    assign P[13] = in[136] ^ in2[136];
    assign G[14] = in[135] & in2[135];
    assign P[14] = in[135] ^ in2[135];
    assign G[15] = in[134] & in2[134];
    assign P[15] = in[134] ^ in2[134];
    assign G[16] = in[133] & in2[133];
    assign P[16] = in[133] ^ in2[133];
    assign G[17] = in[132] & in2[132];
    assign P[17] = in[132] ^ in2[132];
    assign G[18] = in[131] & in2[131];
    assign P[18] = in[131] ^ in2[131];
    assign G[19] = in[130] & in2[130];
    assign P[19] = in[130] ^ in2[130];
    assign G[20] = in[129] & in2[129];
    assign P[20] = in[129] ^ in2[129];
    assign G[21] = in[128] & in2[128];
    assign P[21] = in[128] ^ in2[128];
    assign G[22] = in[127] & in2[127];
    assign P[22] = in[127] ^ in2[127];
    assign G[23] = in[126] & in2[126];
    assign P[23] = in[126] ^ in2[126];
    assign G[24] = in[125] & in2[125];
    assign P[24] = in[125] ^ in2[125];
    assign G[25] = in[124] & in2[124];
    assign P[25] = in[124] ^ in2[124];
    assign G[26] = in[123] & in2[123];
    assign P[26] = in[123] ^ in2[123];
    assign G[27] = in[122] & in2[122];
    assign P[27] = in[122] ^ in2[122];
    assign G[28] = in[121] & in2[121];
    assign P[28] = in[121] ^ in2[121];
    assign G[29] = in[120] & in2[120];
    assign P[29] = in[120] ^ in2[120];
    assign G[30] = in[119] & in2[119];
    assign P[30] = in[119] ^ in2[119];
    assign G[31] = in[118] & in2[118];
    assign P[31] = in[118] ^ in2[118];
    assign G[32] = in[117] & in2[117];
    assign P[32] = in[117] ^ in2[117];
    assign G[33] = in[116] & in2[116];
    assign P[33] = in[116] ^ in2[116];
    assign G[34] = in[115] & in2[115];
    assign P[34] = in[115] ^ in2[115];
    assign G[35] = in[114] & in2[114];
    assign P[35] = in[114] ^ in2[114];
    assign G[36] = in[113] & in2[113];
    assign P[36] = in[113] ^ in2[113];
    assign G[37] = in[112] & in2[112];
    assign P[37] = in[112] ^ in2[112];
    assign G[38] = in[111] & in2[111];
    assign P[38] = in[111] ^ in2[111];
    assign G[39] = in[110] & in2[110];
    assign P[39] = in[110] ^ in2[110];
    assign G[40] = in[109] & in2[109];
    assign P[40] = in[109] ^ in2[109];
    assign G[41] = in[108] & in2[108];
    assign P[41] = in[108] ^ in2[108];
    assign G[42] = in[107] & in2[107];
    assign P[42] = in[107] ^ in2[107];
    assign G[43] = in[106] & in2[106];
    assign P[43] = in[106] ^ in2[106];
    assign G[44] = in[105] & in2[105];
    assign P[44] = in[105] ^ in2[105];
    assign G[45] = in[104] & in2[104];
    assign P[45] = in[104] ^ in2[104];
    assign G[46] = in[103] & in2[103];
    assign P[46] = in[103] ^ in2[103];
    assign G[47] = in[102] & in2[102];
    assign P[47] = in[102] ^ in2[102];
    assign G[48] = in[101] & in2[101];
    assign P[48] = in[101] ^ in2[101];
    assign G[49] = in[100] & in2[100];
    assign P[49] = in[100] ^ in2[100];
    assign G[50] = in[99] & in2[99];
    assign P[50] = in[99] ^ in2[99];
    assign G[51] = in[98] & in2[98];
    assign P[51] = in[98] ^ in2[98];
    assign G[52] = in[97] & in2[97];
    assign P[52] = in[97] ^ in2[97];
    assign G[53] = in[96] & in2[96];
    assign P[53] = in[96] ^ in2[96];
    assign G[54] = in[95] & in2[95];
    assign P[54] = in[95] ^ in2[95];
    assign G[55] = in[94] & in2[94];
    assign P[55] = in[94] ^ in2[94];
    assign G[56] = in[93] & in2[93];
    assign P[56] = in[93] ^ in2[93];
    assign G[57] = in[92] & in2[92];
    assign P[57] = in[92] ^ in2[92];
    assign G[58] = in[91] & in2[91];
    assign P[58] = in[91] ^ in2[91];
    assign G[59] = in[90] & in2[90];
    assign P[59] = in[90] ^ in2[90];
    assign G[60] = in[89] & in2[89];
    assign P[60] = in[89] ^ in2[89];
    assign G[61] = in[88] & in2[88];
    assign P[61] = in[88] ^ in2[88];
    assign G[62] = in[87] & in2[87];
    assign P[62] = in[87] ^ in2[87];
    assign G[63] = in[86] & in2[86];
    assign P[63] = in[86] ^ in2[86];
    assign G[64] = in[85] & in2[85];
    assign P[64] = in[85] ^ in2[85];
    assign G[65] = in[84] & in2[84];
    assign P[65] = in[84] ^ in2[84];
    assign G[66] = in[83] & in2[83];
    assign P[66] = in[83] ^ in2[83];
    assign G[67] = in[82] & in2[82];
    assign P[67] = in[82] ^ in2[82];
    assign G[68] = in[81] & in2[81];
    assign P[68] = in[81] ^ in2[81];
    assign G[69] = in[80] & in2[80];
    assign P[69] = in[80] ^ in2[80];
    assign G[70] = in[79] & in2[79];
    assign P[70] = in[79] ^ in2[79];
    assign G[71] = in[78] & in2[78];
    assign P[71] = in[78] ^ in2[78];
    assign G[72] = in[77] & in2[77];
    assign P[72] = in[77] ^ in2[77];
    assign G[73] = in[76] & in2[76];
    assign P[73] = in[76] ^ in2[76];
    assign G[74] = in[75] & in2[75];
    assign P[74] = in[75] ^ in2[75];
    assign G[75] = in[74] & in2[74];
    assign P[75] = in[74] ^ in2[74];
    assign G[76] = in[73] & in2[73];
    assign P[76] = in[73] ^ in2[73];
    assign G[77] = in[72] & in2[72];
    assign P[77] = in[72] ^ in2[72];
    assign G[78] = in[71] & in2[71];
    assign P[78] = in[71] ^ in2[71];
    assign G[79] = in[70] & in2[70];
    assign P[79] = in[70] ^ in2[70];
    assign G[80] = in[69] & in2[69];
    assign P[80] = in[69] ^ in2[69];
    assign G[81] = in[68] & in2[68];
    assign P[81] = in[68] ^ in2[68];
    assign G[82] = in[67] & in2[67];
    assign P[82] = in[67] ^ in2[67];
    assign G[83] = in[66] & in2[66];
    assign P[83] = in[66] ^ in2[66];
    assign G[84] = in[65] & in2[65];
    assign P[84] = in[65] ^ in2[65];
    assign G[85] = in[64] & in2[64];
    assign P[85] = in[64] ^ in2[64];
    assign G[86] = in[63] & in2[63];
    assign P[86] = in[63] ^ in2[63];
    assign G[87] = in[62] & in2[62];
    assign P[87] = in[62] ^ in2[62];
    assign G[88] = in[61] & in2[61];
    assign P[88] = in[61] ^ in2[61];
    assign G[89] = in[60] & in2[60];
    assign P[89] = in[60] ^ in2[60];
    assign G[90] = in[59] & in2[59];
    assign P[90] = in[59] ^ in2[59];
    assign G[91] = in[58] & in2[58];
    assign P[91] = in[58] ^ in2[58];
    assign G[92] = in[57] & in2[57];
    assign P[92] = in[57] ^ in2[57];
    assign G[93] = in[56] & in2[56];
    assign P[93] = in[56] ^ in2[56];
    assign G[94] = in[55] & in2[55];
    assign P[94] = in[55] ^ in2[55];
    assign G[95] = in[54] & in2[54];
    assign P[95] = in[54] ^ in2[54];
    assign G[96] = in[53] & in2[53];
    assign P[96] = in[53] ^ in2[53];
    assign G[97] = in[52] & in2[52];
    assign P[97] = in[52] ^ in2[52];
    assign G[98] = in[51] & in2[51];
    assign P[98] = in[51] ^ in2[51];
    assign G[99] = in[50] & in2[50];
    assign P[99] = in[50] ^ in2[50];
    assign G[100] = in[49] & in2[49];
    assign P[100] = in[49] ^ in2[49];
    assign G[101] = in[48] & in2[48];
    assign P[101] = in[48] ^ in2[48];
    assign G[102] = in[47] & in2[47];
    assign P[102] = in[47] ^ in2[47];
    assign G[103] = in[46] & in2[46];
    assign P[103] = in[46] ^ in2[46];
    assign G[104] = in[45] & in2[45];
    assign P[104] = in[45] ^ in2[45];
    assign G[105] = in[44] & in2[44];
    assign P[105] = in[44] ^ in2[44];
    assign G[106] = in[43] & in2[43];
    assign P[106] = in[43] ^ in2[43];
    assign G[107] = in[42] & in2[42];
    assign P[107] = in[42] ^ in2[42];
    assign G[108] = in[41] & in2[41];
    assign P[108] = in[41] ^ in2[41];
    assign G[109] = in[40] & in2[40];
    assign P[109] = in[40] ^ in2[40];
    assign G[110] = in[39] & in2[39];
    assign P[110] = in[39] ^ in2[39];
    assign G[111] = in[38] & in2[38];
    assign P[111] = in[38] ^ in2[38];
    assign G[112] = in[37] & in2[37];
    assign P[112] = in[37] ^ in2[37];
    assign G[113] = in[36] & in2[36];
    assign P[113] = in[36] ^ in2[36];
    assign G[114] = in[35] & in2[35];
    assign P[114] = in[35] ^ in2[35];
    assign G[115] = in[34] & in2[34];
    assign P[115] = in[34] ^ in2[34];
    assign G[116] = in[33] & in2[33];
    assign P[116] = in[33] ^ in2[33];
    assign G[117] = in[32] & in2[32];
    assign P[117] = in[32] ^ in2[32];
    assign G[118] = in[31] & in2[31];
    assign P[118] = in[31] ^ in2[31];
    assign G[119] = in[30] & in2[30];
    assign P[119] = in[30] ^ in2[30];
    assign G[120] = in[29] & in2[29];
    assign P[120] = in[29] ^ in2[29];
    assign G[121] = in[28] & in2[28];
    assign P[121] = in[28] ^ in2[28];
    assign G[122] = in[27] & in2[27];
    assign P[122] = in[27] ^ in2[27];
    assign G[123] = in[26] & in2[26];
    assign P[123] = in[26] ^ in2[26];
    assign G[124] = in[25] & in2[25];
    assign P[124] = in[25] ^ in2[25];
    assign G[125] = in[24] & in2[24];
    assign P[125] = in[24] ^ in2[24];
    assign G[126] = in[23] & in2[23];
    assign P[126] = in[23] ^ in2[23];
    assign G[127] = in[22] & in2[22];
    assign P[127] = in[22] ^ in2[22];
    assign G[128] = in[21] & in2[21];
    assign P[128] = in[21] ^ in2[21];
    assign G[129] = in[20] & in2[20];
    assign P[129] = in[20] ^ in2[20];
    assign G[130] = in[19] & in2[19];
    assign P[130] = in[19] ^ in2[19];
    assign G[131] = in[18] & in2[18];
    assign P[131] = in[18] ^ in2[18];
    assign G[132] = in[17] & in2[17];
    assign P[132] = in[17] ^ in2[17];
    assign G[133] = in[16] & in2[16];
    assign P[133] = in[16] ^ in2[16];
    assign G[134] = in[15] & in2[15];
    assign P[134] = in[15] ^ in2[15];
    assign G[135] = in[14] & in2[14];
    assign P[135] = in[14] ^ in2[14];
    assign G[136] = in[13] & in2[13];
    assign P[136] = in[13] ^ in2[13];
    assign G[137] = in[12] & in2[12];
    assign P[137] = in[12] ^ in2[12];
    assign G[138] = in[11] & in2[11];
    assign P[138] = in[11] ^ in2[11];
    assign G[139] = in[10] & in2[10];
    assign P[139] = in[10] ^ in2[10];
    assign G[140] = in[9] & in2[9];
    assign P[140] = in[9] ^ in2[9];
    assign G[141] = in[8] & in2[8];
    assign P[141] = in[8] ^ in2[8];
    assign G[142] = in[7] & in2[7];
    assign P[142] = in[7] ^ in2[7];
    assign G[143] = in[6] & in2[6];
    assign P[143] = in[6] ^ in2[6];
    assign G[144] = in[5] & in2[5];
    assign P[144] = in[5] ^ in2[5];
    assign G[145] = in[4] & in2[4];
    assign P[145] = in[4] ^ in2[4];
    assign G[146] = in[3] & in2[3];
    assign P[146] = in[3] ^ in2[3];
    assign G[147] = in[2] & in2[2];
    assign P[147] = in[2] ^ in2[2];
    assign G[148] = in[1] & in2[1];
    assign P[148] = in[1] ^ in2[1];
    assign G[149] = in[0] & in2[0];
    assign P[149] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign C[149] = G[148] | (P[148] & C[148]);
    assign cout = G[149] | (P[149] & C[149]);
    assign sum = P ^ C;
endmodule

module CLA149(output [148:0] sum, output cout, input [148:0] in1, input [148:0] in2;

    wire[148:0] G;
    wire[148:0] C;
    wire[148:0] P;

    assign G[0] = in[148] & in2[148];
    assign P[0] = in[148] ^ in2[148];
    assign G[1] = in[147] & in2[147];
    assign P[1] = in[147] ^ in2[147];
    assign G[2] = in[146] & in2[146];
    assign P[2] = in[146] ^ in2[146];
    assign G[3] = in[145] & in2[145];
    assign P[3] = in[145] ^ in2[145];
    assign G[4] = in[144] & in2[144];
    assign P[4] = in[144] ^ in2[144];
    assign G[5] = in[143] & in2[143];
    assign P[5] = in[143] ^ in2[143];
    assign G[6] = in[142] & in2[142];
    assign P[6] = in[142] ^ in2[142];
    assign G[7] = in[141] & in2[141];
    assign P[7] = in[141] ^ in2[141];
    assign G[8] = in[140] & in2[140];
    assign P[8] = in[140] ^ in2[140];
    assign G[9] = in[139] & in2[139];
    assign P[9] = in[139] ^ in2[139];
    assign G[10] = in[138] & in2[138];
    assign P[10] = in[138] ^ in2[138];
    assign G[11] = in[137] & in2[137];
    assign P[11] = in[137] ^ in2[137];
    assign G[12] = in[136] & in2[136];
    assign P[12] = in[136] ^ in2[136];
    assign G[13] = in[135] & in2[135];
    assign P[13] = in[135] ^ in2[135];
    assign G[14] = in[134] & in2[134];
    assign P[14] = in[134] ^ in2[134];
    assign G[15] = in[133] & in2[133];
    assign P[15] = in[133] ^ in2[133];
    assign G[16] = in[132] & in2[132];
    assign P[16] = in[132] ^ in2[132];
    assign G[17] = in[131] & in2[131];
    assign P[17] = in[131] ^ in2[131];
    assign G[18] = in[130] & in2[130];
    assign P[18] = in[130] ^ in2[130];
    assign G[19] = in[129] & in2[129];
    assign P[19] = in[129] ^ in2[129];
    assign G[20] = in[128] & in2[128];
    assign P[20] = in[128] ^ in2[128];
    assign G[21] = in[127] & in2[127];
    assign P[21] = in[127] ^ in2[127];
    assign G[22] = in[126] & in2[126];
    assign P[22] = in[126] ^ in2[126];
    assign G[23] = in[125] & in2[125];
    assign P[23] = in[125] ^ in2[125];
    assign G[24] = in[124] & in2[124];
    assign P[24] = in[124] ^ in2[124];
    assign G[25] = in[123] & in2[123];
    assign P[25] = in[123] ^ in2[123];
    assign G[26] = in[122] & in2[122];
    assign P[26] = in[122] ^ in2[122];
    assign G[27] = in[121] & in2[121];
    assign P[27] = in[121] ^ in2[121];
    assign G[28] = in[120] & in2[120];
    assign P[28] = in[120] ^ in2[120];
    assign G[29] = in[119] & in2[119];
    assign P[29] = in[119] ^ in2[119];
    assign G[30] = in[118] & in2[118];
    assign P[30] = in[118] ^ in2[118];
    assign G[31] = in[117] & in2[117];
    assign P[31] = in[117] ^ in2[117];
    assign G[32] = in[116] & in2[116];
    assign P[32] = in[116] ^ in2[116];
    assign G[33] = in[115] & in2[115];
    assign P[33] = in[115] ^ in2[115];
    assign G[34] = in[114] & in2[114];
    assign P[34] = in[114] ^ in2[114];
    assign G[35] = in[113] & in2[113];
    assign P[35] = in[113] ^ in2[113];
    assign G[36] = in[112] & in2[112];
    assign P[36] = in[112] ^ in2[112];
    assign G[37] = in[111] & in2[111];
    assign P[37] = in[111] ^ in2[111];
    assign G[38] = in[110] & in2[110];
    assign P[38] = in[110] ^ in2[110];
    assign G[39] = in[109] & in2[109];
    assign P[39] = in[109] ^ in2[109];
    assign G[40] = in[108] & in2[108];
    assign P[40] = in[108] ^ in2[108];
    assign G[41] = in[107] & in2[107];
    assign P[41] = in[107] ^ in2[107];
    assign G[42] = in[106] & in2[106];
    assign P[42] = in[106] ^ in2[106];
    assign G[43] = in[105] & in2[105];
    assign P[43] = in[105] ^ in2[105];
    assign G[44] = in[104] & in2[104];
    assign P[44] = in[104] ^ in2[104];
    assign G[45] = in[103] & in2[103];
    assign P[45] = in[103] ^ in2[103];
    assign G[46] = in[102] & in2[102];
    assign P[46] = in[102] ^ in2[102];
    assign G[47] = in[101] & in2[101];
    assign P[47] = in[101] ^ in2[101];
    assign G[48] = in[100] & in2[100];
    assign P[48] = in[100] ^ in2[100];
    assign G[49] = in[99] & in2[99];
    assign P[49] = in[99] ^ in2[99];
    assign G[50] = in[98] & in2[98];
    assign P[50] = in[98] ^ in2[98];
    assign G[51] = in[97] & in2[97];
    assign P[51] = in[97] ^ in2[97];
    assign G[52] = in[96] & in2[96];
    assign P[52] = in[96] ^ in2[96];
    assign G[53] = in[95] & in2[95];
    assign P[53] = in[95] ^ in2[95];
    assign G[54] = in[94] & in2[94];
    assign P[54] = in[94] ^ in2[94];
    assign G[55] = in[93] & in2[93];
    assign P[55] = in[93] ^ in2[93];
    assign G[56] = in[92] & in2[92];
    assign P[56] = in[92] ^ in2[92];
    assign G[57] = in[91] & in2[91];
    assign P[57] = in[91] ^ in2[91];
    assign G[58] = in[90] & in2[90];
    assign P[58] = in[90] ^ in2[90];
    assign G[59] = in[89] & in2[89];
    assign P[59] = in[89] ^ in2[89];
    assign G[60] = in[88] & in2[88];
    assign P[60] = in[88] ^ in2[88];
    assign G[61] = in[87] & in2[87];
    assign P[61] = in[87] ^ in2[87];
    assign G[62] = in[86] & in2[86];
    assign P[62] = in[86] ^ in2[86];
    assign G[63] = in[85] & in2[85];
    assign P[63] = in[85] ^ in2[85];
    assign G[64] = in[84] & in2[84];
    assign P[64] = in[84] ^ in2[84];
    assign G[65] = in[83] & in2[83];
    assign P[65] = in[83] ^ in2[83];
    assign G[66] = in[82] & in2[82];
    assign P[66] = in[82] ^ in2[82];
    assign G[67] = in[81] & in2[81];
    assign P[67] = in[81] ^ in2[81];
    assign G[68] = in[80] & in2[80];
    assign P[68] = in[80] ^ in2[80];
    assign G[69] = in[79] & in2[79];
    assign P[69] = in[79] ^ in2[79];
    assign G[70] = in[78] & in2[78];
    assign P[70] = in[78] ^ in2[78];
    assign G[71] = in[77] & in2[77];
    assign P[71] = in[77] ^ in2[77];
    assign G[72] = in[76] & in2[76];
    assign P[72] = in[76] ^ in2[76];
    assign G[73] = in[75] & in2[75];
    assign P[73] = in[75] ^ in2[75];
    assign G[74] = in[74] & in2[74];
    assign P[74] = in[74] ^ in2[74];
    assign G[75] = in[73] & in2[73];
    assign P[75] = in[73] ^ in2[73];
    assign G[76] = in[72] & in2[72];
    assign P[76] = in[72] ^ in2[72];
    assign G[77] = in[71] & in2[71];
    assign P[77] = in[71] ^ in2[71];
    assign G[78] = in[70] & in2[70];
    assign P[78] = in[70] ^ in2[70];
    assign G[79] = in[69] & in2[69];
    assign P[79] = in[69] ^ in2[69];
    assign G[80] = in[68] & in2[68];
    assign P[80] = in[68] ^ in2[68];
    assign G[81] = in[67] & in2[67];
    assign P[81] = in[67] ^ in2[67];
    assign G[82] = in[66] & in2[66];
    assign P[82] = in[66] ^ in2[66];
    assign G[83] = in[65] & in2[65];
    assign P[83] = in[65] ^ in2[65];
    assign G[84] = in[64] & in2[64];
    assign P[84] = in[64] ^ in2[64];
    assign G[85] = in[63] & in2[63];
    assign P[85] = in[63] ^ in2[63];
    assign G[86] = in[62] & in2[62];
    assign P[86] = in[62] ^ in2[62];
    assign G[87] = in[61] & in2[61];
    assign P[87] = in[61] ^ in2[61];
    assign G[88] = in[60] & in2[60];
    assign P[88] = in[60] ^ in2[60];
    assign G[89] = in[59] & in2[59];
    assign P[89] = in[59] ^ in2[59];
    assign G[90] = in[58] & in2[58];
    assign P[90] = in[58] ^ in2[58];
    assign G[91] = in[57] & in2[57];
    assign P[91] = in[57] ^ in2[57];
    assign G[92] = in[56] & in2[56];
    assign P[92] = in[56] ^ in2[56];
    assign G[93] = in[55] & in2[55];
    assign P[93] = in[55] ^ in2[55];
    assign G[94] = in[54] & in2[54];
    assign P[94] = in[54] ^ in2[54];
    assign G[95] = in[53] & in2[53];
    assign P[95] = in[53] ^ in2[53];
    assign G[96] = in[52] & in2[52];
    assign P[96] = in[52] ^ in2[52];
    assign G[97] = in[51] & in2[51];
    assign P[97] = in[51] ^ in2[51];
    assign G[98] = in[50] & in2[50];
    assign P[98] = in[50] ^ in2[50];
    assign G[99] = in[49] & in2[49];
    assign P[99] = in[49] ^ in2[49];
    assign G[100] = in[48] & in2[48];
    assign P[100] = in[48] ^ in2[48];
    assign G[101] = in[47] & in2[47];
    assign P[101] = in[47] ^ in2[47];
    assign G[102] = in[46] & in2[46];
    assign P[102] = in[46] ^ in2[46];
    assign G[103] = in[45] & in2[45];
    assign P[103] = in[45] ^ in2[45];
    assign G[104] = in[44] & in2[44];
    assign P[104] = in[44] ^ in2[44];
    assign G[105] = in[43] & in2[43];
    assign P[105] = in[43] ^ in2[43];
    assign G[106] = in[42] & in2[42];
    assign P[106] = in[42] ^ in2[42];
    assign G[107] = in[41] & in2[41];
    assign P[107] = in[41] ^ in2[41];
    assign G[108] = in[40] & in2[40];
    assign P[108] = in[40] ^ in2[40];
    assign G[109] = in[39] & in2[39];
    assign P[109] = in[39] ^ in2[39];
    assign G[110] = in[38] & in2[38];
    assign P[110] = in[38] ^ in2[38];
    assign G[111] = in[37] & in2[37];
    assign P[111] = in[37] ^ in2[37];
    assign G[112] = in[36] & in2[36];
    assign P[112] = in[36] ^ in2[36];
    assign G[113] = in[35] & in2[35];
    assign P[113] = in[35] ^ in2[35];
    assign G[114] = in[34] & in2[34];
    assign P[114] = in[34] ^ in2[34];
    assign G[115] = in[33] & in2[33];
    assign P[115] = in[33] ^ in2[33];
    assign G[116] = in[32] & in2[32];
    assign P[116] = in[32] ^ in2[32];
    assign G[117] = in[31] & in2[31];
    assign P[117] = in[31] ^ in2[31];
    assign G[118] = in[30] & in2[30];
    assign P[118] = in[30] ^ in2[30];
    assign G[119] = in[29] & in2[29];
    assign P[119] = in[29] ^ in2[29];
    assign G[120] = in[28] & in2[28];
    assign P[120] = in[28] ^ in2[28];
    assign G[121] = in[27] & in2[27];
    assign P[121] = in[27] ^ in2[27];
    assign G[122] = in[26] & in2[26];
    assign P[122] = in[26] ^ in2[26];
    assign G[123] = in[25] & in2[25];
    assign P[123] = in[25] ^ in2[25];
    assign G[124] = in[24] & in2[24];
    assign P[124] = in[24] ^ in2[24];
    assign G[125] = in[23] & in2[23];
    assign P[125] = in[23] ^ in2[23];
    assign G[126] = in[22] & in2[22];
    assign P[126] = in[22] ^ in2[22];
    assign G[127] = in[21] & in2[21];
    assign P[127] = in[21] ^ in2[21];
    assign G[128] = in[20] & in2[20];
    assign P[128] = in[20] ^ in2[20];
    assign G[129] = in[19] & in2[19];
    assign P[129] = in[19] ^ in2[19];
    assign G[130] = in[18] & in2[18];
    assign P[130] = in[18] ^ in2[18];
    assign G[131] = in[17] & in2[17];
    assign P[131] = in[17] ^ in2[17];
    assign G[132] = in[16] & in2[16];
    assign P[132] = in[16] ^ in2[16];
    assign G[133] = in[15] & in2[15];
    assign P[133] = in[15] ^ in2[15];
    assign G[134] = in[14] & in2[14];
    assign P[134] = in[14] ^ in2[14];
    assign G[135] = in[13] & in2[13];
    assign P[135] = in[13] ^ in2[13];
    assign G[136] = in[12] & in2[12];
    assign P[136] = in[12] ^ in2[12];
    assign G[137] = in[11] & in2[11];
    assign P[137] = in[11] ^ in2[11];
    assign G[138] = in[10] & in2[10];
    assign P[138] = in[10] ^ in2[10];
    assign G[139] = in[9] & in2[9];
    assign P[139] = in[9] ^ in2[9];
    assign G[140] = in[8] & in2[8];
    assign P[140] = in[8] ^ in2[8];
    assign G[141] = in[7] & in2[7];
    assign P[141] = in[7] ^ in2[7];
    assign G[142] = in[6] & in2[6];
    assign P[142] = in[6] ^ in2[6];
    assign G[143] = in[5] & in2[5];
    assign P[143] = in[5] ^ in2[5];
    assign G[144] = in[4] & in2[4];
    assign P[144] = in[4] ^ in2[4];
    assign G[145] = in[3] & in2[3];
    assign P[145] = in[3] ^ in2[3];
    assign G[146] = in[2] & in2[2];
    assign P[146] = in[2] ^ in2[2];
    assign G[147] = in[1] & in2[1];
    assign P[147] = in[1] ^ in2[1];
    assign G[148] = in[0] & in2[0];
    assign P[148] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign C[148] = G[147] | (P[147] & C[147]);
    assign cout = G[148] | (P[148] & C[148]);
    assign sum = P ^ C;
endmodule

module CLA148(output [147:0] sum, output cout, input [147:0] in1, input [147:0] in2;

    wire[147:0] G;
    wire[147:0] C;
    wire[147:0] P;

    assign G[0] = in[147] & in2[147];
    assign P[0] = in[147] ^ in2[147];
    assign G[1] = in[146] & in2[146];
    assign P[1] = in[146] ^ in2[146];
    assign G[2] = in[145] & in2[145];
    assign P[2] = in[145] ^ in2[145];
    assign G[3] = in[144] & in2[144];
    assign P[3] = in[144] ^ in2[144];
    assign G[4] = in[143] & in2[143];
    assign P[4] = in[143] ^ in2[143];
    assign G[5] = in[142] & in2[142];
    assign P[5] = in[142] ^ in2[142];
    assign G[6] = in[141] & in2[141];
    assign P[6] = in[141] ^ in2[141];
    assign G[7] = in[140] & in2[140];
    assign P[7] = in[140] ^ in2[140];
    assign G[8] = in[139] & in2[139];
    assign P[8] = in[139] ^ in2[139];
    assign G[9] = in[138] & in2[138];
    assign P[9] = in[138] ^ in2[138];
    assign G[10] = in[137] & in2[137];
    assign P[10] = in[137] ^ in2[137];
    assign G[11] = in[136] & in2[136];
    assign P[11] = in[136] ^ in2[136];
    assign G[12] = in[135] & in2[135];
    assign P[12] = in[135] ^ in2[135];
    assign G[13] = in[134] & in2[134];
    assign P[13] = in[134] ^ in2[134];
    assign G[14] = in[133] & in2[133];
    assign P[14] = in[133] ^ in2[133];
    assign G[15] = in[132] & in2[132];
    assign P[15] = in[132] ^ in2[132];
    assign G[16] = in[131] & in2[131];
    assign P[16] = in[131] ^ in2[131];
    assign G[17] = in[130] & in2[130];
    assign P[17] = in[130] ^ in2[130];
    assign G[18] = in[129] & in2[129];
    assign P[18] = in[129] ^ in2[129];
    assign G[19] = in[128] & in2[128];
    assign P[19] = in[128] ^ in2[128];
    assign G[20] = in[127] & in2[127];
    assign P[20] = in[127] ^ in2[127];
    assign G[21] = in[126] & in2[126];
    assign P[21] = in[126] ^ in2[126];
    assign G[22] = in[125] & in2[125];
    assign P[22] = in[125] ^ in2[125];
    assign G[23] = in[124] & in2[124];
    assign P[23] = in[124] ^ in2[124];
    assign G[24] = in[123] & in2[123];
    assign P[24] = in[123] ^ in2[123];
    assign G[25] = in[122] & in2[122];
    assign P[25] = in[122] ^ in2[122];
    assign G[26] = in[121] & in2[121];
    assign P[26] = in[121] ^ in2[121];
    assign G[27] = in[120] & in2[120];
    assign P[27] = in[120] ^ in2[120];
    assign G[28] = in[119] & in2[119];
    assign P[28] = in[119] ^ in2[119];
    assign G[29] = in[118] & in2[118];
    assign P[29] = in[118] ^ in2[118];
    assign G[30] = in[117] & in2[117];
    assign P[30] = in[117] ^ in2[117];
    assign G[31] = in[116] & in2[116];
    assign P[31] = in[116] ^ in2[116];
    assign G[32] = in[115] & in2[115];
    assign P[32] = in[115] ^ in2[115];
    assign G[33] = in[114] & in2[114];
    assign P[33] = in[114] ^ in2[114];
    assign G[34] = in[113] & in2[113];
    assign P[34] = in[113] ^ in2[113];
    assign G[35] = in[112] & in2[112];
    assign P[35] = in[112] ^ in2[112];
    assign G[36] = in[111] & in2[111];
    assign P[36] = in[111] ^ in2[111];
    assign G[37] = in[110] & in2[110];
    assign P[37] = in[110] ^ in2[110];
    assign G[38] = in[109] & in2[109];
    assign P[38] = in[109] ^ in2[109];
    assign G[39] = in[108] & in2[108];
    assign P[39] = in[108] ^ in2[108];
    assign G[40] = in[107] & in2[107];
    assign P[40] = in[107] ^ in2[107];
    assign G[41] = in[106] & in2[106];
    assign P[41] = in[106] ^ in2[106];
    assign G[42] = in[105] & in2[105];
    assign P[42] = in[105] ^ in2[105];
    assign G[43] = in[104] & in2[104];
    assign P[43] = in[104] ^ in2[104];
    assign G[44] = in[103] & in2[103];
    assign P[44] = in[103] ^ in2[103];
    assign G[45] = in[102] & in2[102];
    assign P[45] = in[102] ^ in2[102];
    assign G[46] = in[101] & in2[101];
    assign P[46] = in[101] ^ in2[101];
    assign G[47] = in[100] & in2[100];
    assign P[47] = in[100] ^ in2[100];
    assign G[48] = in[99] & in2[99];
    assign P[48] = in[99] ^ in2[99];
    assign G[49] = in[98] & in2[98];
    assign P[49] = in[98] ^ in2[98];
    assign G[50] = in[97] & in2[97];
    assign P[50] = in[97] ^ in2[97];
    assign G[51] = in[96] & in2[96];
    assign P[51] = in[96] ^ in2[96];
    assign G[52] = in[95] & in2[95];
    assign P[52] = in[95] ^ in2[95];
    assign G[53] = in[94] & in2[94];
    assign P[53] = in[94] ^ in2[94];
    assign G[54] = in[93] & in2[93];
    assign P[54] = in[93] ^ in2[93];
    assign G[55] = in[92] & in2[92];
    assign P[55] = in[92] ^ in2[92];
    assign G[56] = in[91] & in2[91];
    assign P[56] = in[91] ^ in2[91];
    assign G[57] = in[90] & in2[90];
    assign P[57] = in[90] ^ in2[90];
    assign G[58] = in[89] & in2[89];
    assign P[58] = in[89] ^ in2[89];
    assign G[59] = in[88] & in2[88];
    assign P[59] = in[88] ^ in2[88];
    assign G[60] = in[87] & in2[87];
    assign P[60] = in[87] ^ in2[87];
    assign G[61] = in[86] & in2[86];
    assign P[61] = in[86] ^ in2[86];
    assign G[62] = in[85] & in2[85];
    assign P[62] = in[85] ^ in2[85];
    assign G[63] = in[84] & in2[84];
    assign P[63] = in[84] ^ in2[84];
    assign G[64] = in[83] & in2[83];
    assign P[64] = in[83] ^ in2[83];
    assign G[65] = in[82] & in2[82];
    assign P[65] = in[82] ^ in2[82];
    assign G[66] = in[81] & in2[81];
    assign P[66] = in[81] ^ in2[81];
    assign G[67] = in[80] & in2[80];
    assign P[67] = in[80] ^ in2[80];
    assign G[68] = in[79] & in2[79];
    assign P[68] = in[79] ^ in2[79];
    assign G[69] = in[78] & in2[78];
    assign P[69] = in[78] ^ in2[78];
    assign G[70] = in[77] & in2[77];
    assign P[70] = in[77] ^ in2[77];
    assign G[71] = in[76] & in2[76];
    assign P[71] = in[76] ^ in2[76];
    assign G[72] = in[75] & in2[75];
    assign P[72] = in[75] ^ in2[75];
    assign G[73] = in[74] & in2[74];
    assign P[73] = in[74] ^ in2[74];
    assign G[74] = in[73] & in2[73];
    assign P[74] = in[73] ^ in2[73];
    assign G[75] = in[72] & in2[72];
    assign P[75] = in[72] ^ in2[72];
    assign G[76] = in[71] & in2[71];
    assign P[76] = in[71] ^ in2[71];
    assign G[77] = in[70] & in2[70];
    assign P[77] = in[70] ^ in2[70];
    assign G[78] = in[69] & in2[69];
    assign P[78] = in[69] ^ in2[69];
    assign G[79] = in[68] & in2[68];
    assign P[79] = in[68] ^ in2[68];
    assign G[80] = in[67] & in2[67];
    assign P[80] = in[67] ^ in2[67];
    assign G[81] = in[66] & in2[66];
    assign P[81] = in[66] ^ in2[66];
    assign G[82] = in[65] & in2[65];
    assign P[82] = in[65] ^ in2[65];
    assign G[83] = in[64] & in2[64];
    assign P[83] = in[64] ^ in2[64];
    assign G[84] = in[63] & in2[63];
    assign P[84] = in[63] ^ in2[63];
    assign G[85] = in[62] & in2[62];
    assign P[85] = in[62] ^ in2[62];
    assign G[86] = in[61] & in2[61];
    assign P[86] = in[61] ^ in2[61];
    assign G[87] = in[60] & in2[60];
    assign P[87] = in[60] ^ in2[60];
    assign G[88] = in[59] & in2[59];
    assign P[88] = in[59] ^ in2[59];
    assign G[89] = in[58] & in2[58];
    assign P[89] = in[58] ^ in2[58];
    assign G[90] = in[57] & in2[57];
    assign P[90] = in[57] ^ in2[57];
    assign G[91] = in[56] & in2[56];
    assign P[91] = in[56] ^ in2[56];
    assign G[92] = in[55] & in2[55];
    assign P[92] = in[55] ^ in2[55];
    assign G[93] = in[54] & in2[54];
    assign P[93] = in[54] ^ in2[54];
    assign G[94] = in[53] & in2[53];
    assign P[94] = in[53] ^ in2[53];
    assign G[95] = in[52] & in2[52];
    assign P[95] = in[52] ^ in2[52];
    assign G[96] = in[51] & in2[51];
    assign P[96] = in[51] ^ in2[51];
    assign G[97] = in[50] & in2[50];
    assign P[97] = in[50] ^ in2[50];
    assign G[98] = in[49] & in2[49];
    assign P[98] = in[49] ^ in2[49];
    assign G[99] = in[48] & in2[48];
    assign P[99] = in[48] ^ in2[48];
    assign G[100] = in[47] & in2[47];
    assign P[100] = in[47] ^ in2[47];
    assign G[101] = in[46] & in2[46];
    assign P[101] = in[46] ^ in2[46];
    assign G[102] = in[45] & in2[45];
    assign P[102] = in[45] ^ in2[45];
    assign G[103] = in[44] & in2[44];
    assign P[103] = in[44] ^ in2[44];
    assign G[104] = in[43] & in2[43];
    assign P[104] = in[43] ^ in2[43];
    assign G[105] = in[42] & in2[42];
    assign P[105] = in[42] ^ in2[42];
    assign G[106] = in[41] & in2[41];
    assign P[106] = in[41] ^ in2[41];
    assign G[107] = in[40] & in2[40];
    assign P[107] = in[40] ^ in2[40];
    assign G[108] = in[39] & in2[39];
    assign P[108] = in[39] ^ in2[39];
    assign G[109] = in[38] & in2[38];
    assign P[109] = in[38] ^ in2[38];
    assign G[110] = in[37] & in2[37];
    assign P[110] = in[37] ^ in2[37];
    assign G[111] = in[36] & in2[36];
    assign P[111] = in[36] ^ in2[36];
    assign G[112] = in[35] & in2[35];
    assign P[112] = in[35] ^ in2[35];
    assign G[113] = in[34] & in2[34];
    assign P[113] = in[34] ^ in2[34];
    assign G[114] = in[33] & in2[33];
    assign P[114] = in[33] ^ in2[33];
    assign G[115] = in[32] & in2[32];
    assign P[115] = in[32] ^ in2[32];
    assign G[116] = in[31] & in2[31];
    assign P[116] = in[31] ^ in2[31];
    assign G[117] = in[30] & in2[30];
    assign P[117] = in[30] ^ in2[30];
    assign G[118] = in[29] & in2[29];
    assign P[118] = in[29] ^ in2[29];
    assign G[119] = in[28] & in2[28];
    assign P[119] = in[28] ^ in2[28];
    assign G[120] = in[27] & in2[27];
    assign P[120] = in[27] ^ in2[27];
    assign G[121] = in[26] & in2[26];
    assign P[121] = in[26] ^ in2[26];
    assign G[122] = in[25] & in2[25];
    assign P[122] = in[25] ^ in2[25];
    assign G[123] = in[24] & in2[24];
    assign P[123] = in[24] ^ in2[24];
    assign G[124] = in[23] & in2[23];
    assign P[124] = in[23] ^ in2[23];
    assign G[125] = in[22] & in2[22];
    assign P[125] = in[22] ^ in2[22];
    assign G[126] = in[21] & in2[21];
    assign P[126] = in[21] ^ in2[21];
    assign G[127] = in[20] & in2[20];
    assign P[127] = in[20] ^ in2[20];
    assign G[128] = in[19] & in2[19];
    assign P[128] = in[19] ^ in2[19];
    assign G[129] = in[18] & in2[18];
    assign P[129] = in[18] ^ in2[18];
    assign G[130] = in[17] & in2[17];
    assign P[130] = in[17] ^ in2[17];
    assign G[131] = in[16] & in2[16];
    assign P[131] = in[16] ^ in2[16];
    assign G[132] = in[15] & in2[15];
    assign P[132] = in[15] ^ in2[15];
    assign G[133] = in[14] & in2[14];
    assign P[133] = in[14] ^ in2[14];
    assign G[134] = in[13] & in2[13];
    assign P[134] = in[13] ^ in2[13];
    assign G[135] = in[12] & in2[12];
    assign P[135] = in[12] ^ in2[12];
    assign G[136] = in[11] & in2[11];
    assign P[136] = in[11] ^ in2[11];
    assign G[137] = in[10] & in2[10];
    assign P[137] = in[10] ^ in2[10];
    assign G[138] = in[9] & in2[9];
    assign P[138] = in[9] ^ in2[9];
    assign G[139] = in[8] & in2[8];
    assign P[139] = in[8] ^ in2[8];
    assign G[140] = in[7] & in2[7];
    assign P[140] = in[7] ^ in2[7];
    assign G[141] = in[6] & in2[6];
    assign P[141] = in[6] ^ in2[6];
    assign G[142] = in[5] & in2[5];
    assign P[142] = in[5] ^ in2[5];
    assign G[143] = in[4] & in2[4];
    assign P[143] = in[4] ^ in2[4];
    assign G[144] = in[3] & in2[3];
    assign P[144] = in[3] ^ in2[3];
    assign G[145] = in[2] & in2[2];
    assign P[145] = in[2] ^ in2[2];
    assign G[146] = in[1] & in2[1];
    assign P[146] = in[1] ^ in2[1];
    assign G[147] = in[0] & in2[0];
    assign P[147] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign C[147] = G[146] | (P[146] & C[146]);
    assign cout = G[147] | (P[147] & C[147]);
    assign sum = P ^ C;
endmodule

module CLA147(output [146:0] sum, output cout, input [146:0] in1, input [146:0] in2;

    wire[146:0] G;
    wire[146:0] C;
    wire[146:0] P;

    assign G[0] = in[146] & in2[146];
    assign P[0] = in[146] ^ in2[146];
    assign G[1] = in[145] & in2[145];
    assign P[1] = in[145] ^ in2[145];
    assign G[2] = in[144] & in2[144];
    assign P[2] = in[144] ^ in2[144];
    assign G[3] = in[143] & in2[143];
    assign P[3] = in[143] ^ in2[143];
    assign G[4] = in[142] & in2[142];
    assign P[4] = in[142] ^ in2[142];
    assign G[5] = in[141] & in2[141];
    assign P[5] = in[141] ^ in2[141];
    assign G[6] = in[140] & in2[140];
    assign P[6] = in[140] ^ in2[140];
    assign G[7] = in[139] & in2[139];
    assign P[7] = in[139] ^ in2[139];
    assign G[8] = in[138] & in2[138];
    assign P[8] = in[138] ^ in2[138];
    assign G[9] = in[137] & in2[137];
    assign P[9] = in[137] ^ in2[137];
    assign G[10] = in[136] & in2[136];
    assign P[10] = in[136] ^ in2[136];
    assign G[11] = in[135] & in2[135];
    assign P[11] = in[135] ^ in2[135];
    assign G[12] = in[134] & in2[134];
    assign P[12] = in[134] ^ in2[134];
    assign G[13] = in[133] & in2[133];
    assign P[13] = in[133] ^ in2[133];
    assign G[14] = in[132] & in2[132];
    assign P[14] = in[132] ^ in2[132];
    assign G[15] = in[131] & in2[131];
    assign P[15] = in[131] ^ in2[131];
    assign G[16] = in[130] & in2[130];
    assign P[16] = in[130] ^ in2[130];
    assign G[17] = in[129] & in2[129];
    assign P[17] = in[129] ^ in2[129];
    assign G[18] = in[128] & in2[128];
    assign P[18] = in[128] ^ in2[128];
    assign G[19] = in[127] & in2[127];
    assign P[19] = in[127] ^ in2[127];
    assign G[20] = in[126] & in2[126];
    assign P[20] = in[126] ^ in2[126];
    assign G[21] = in[125] & in2[125];
    assign P[21] = in[125] ^ in2[125];
    assign G[22] = in[124] & in2[124];
    assign P[22] = in[124] ^ in2[124];
    assign G[23] = in[123] & in2[123];
    assign P[23] = in[123] ^ in2[123];
    assign G[24] = in[122] & in2[122];
    assign P[24] = in[122] ^ in2[122];
    assign G[25] = in[121] & in2[121];
    assign P[25] = in[121] ^ in2[121];
    assign G[26] = in[120] & in2[120];
    assign P[26] = in[120] ^ in2[120];
    assign G[27] = in[119] & in2[119];
    assign P[27] = in[119] ^ in2[119];
    assign G[28] = in[118] & in2[118];
    assign P[28] = in[118] ^ in2[118];
    assign G[29] = in[117] & in2[117];
    assign P[29] = in[117] ^ in2[117];
    assign G[30] = in[116] & in2[116];
    assign P[30] = in[116] ^ in2[116];
    assign G[31] = in[115] & in2[115];
    assign P[31] = in[115] ^ in2[115];
    assign G[32] = in[114] & in2[114];
    assign P[32] = in[114] ^ in2[114];
    assign G[33] = in[113] & in2[113];
    assign P[33] = in[113] ^ in2[113];
    assign G[34] = in[112] & in2[112];
    assign P[34] = in[112] ^ in2[112];
    assign G[35] = in[111] & in2[111];
    assign P[35] = in[111] ^ in2[111];
    assign G[36] = in[110] & in2[110];
    assign P[36] = in[110] ^ in2[110];
    assign G[37] = in[109] & in2[109];
    assign P[37] = in[109] ^ in2[109];
    assign G[38] = in[108] & in2[108];
    assign P[38] = in[108] ^ in2[108];
    assign G[39] = in[107] & in2[107];
    assign P[39] = in[107] ^ in2[107];
    assign G[40] = in[106] & in2[106];
    assign P[40] = in[106] ^ in2[106];
    assign G[41] = in[105] & in2[105];
    assign P[41] = in[105] ^ in2[105];
    assign G[42] = in[104] & in2[104];
    assign P[42] = in[104] ^ in2[104];
    assign G[43] = in[103] & in2[103];
    assign P[43] = in[103] ^ in2[103];
    assign G[44] = in[102] & in2[102];
    assign P[44] = in[102] ^ in2[102];
    assign G[45] = in[101] & in2[101];
    assign P[45] = in[101] ^ in2[101];
    assign G[46] = in[100] & in2[100];
    assign P[46] = in[100] ^ in2[100];
    assign G[47] = in[99] & in2[99];
    assign P[47] = in[99] ^ in2[99];
    assign G[48] = in[98] & in2[98];
    assign P[48] = in[98] ^ in2[98];
    assign G[49] = in[97] & in2[97];
    assign P[49] = in[97] ^ in2[97];
    assign G[50] = in[96] & in2[96];
    assign P[50] = in[96] ^ in2[96];
    assign G[51] = in[95] & in2[95];
    assign P[51] = in[95] ^ in2[95];
    assign G[52] = in[94] & in2[94];
    assign P[52] = in[94] ^ in2[94];
    assign G[53] = in[93] & in2[93];
    assign P[53] = in[93] ^ in2[93];
    assign G[54] = in[92] & in2[92];
    assign P[54] = in[92] ^ in2[92];
    assign G[55] = in[91] & in2[91];
    assign P[55] = in[91] ^ in2[91];
    assign G[56] = in[90] & in2[90];
    assign P[56] = in[90] ^ in2[90];
    assign G[57] = in[89] & in2[89];
    assign P[57] = in[89] ^ in2[89];
    assign G[58] = in[88] & in2[88];
    assign P[58] = in[88] ^ in2[88];
    assign G[59] = in[87] & in2[87];
    assign P[59] = in[87] ^ in2[87];
    assign G[60] = in[86] & in2[86];
    assign P[60] = in[86] ^ in2[86];
    assign G[61] = in[85] & in2[85];
    assign P[61] = in[85] ^ in2[85];
    assign G[62] = in[84] & in2[84];
    assign P[62] = in[84] ^ in2[84];
    assign G[63] = in[83] & in2[83];
    assign P[63] = in[83] ^ in2[83];
    assign G[64] = in[82] & in2[82];
    assign P[64] = in[82] ^ in2[82];
    assign G[65] = in[81] & in2[81];
    assign P[65] = in[81] ^ in2[81];
    assign G[66] = in[80] & in2[80];
    assign P[66] = in[80] ^ in2[80];
    assign G[67] = in[79] & in2[79];
    assign P[67] = in[79] ^ in2[79];
    assign G[68] = in[78] & in2[78];
    assign P[68] = in[78] ^ in2[78];
    assign G[69] = in[77] & in2[77];
    assign P[69] = in[77] ^ in2[77];
    assign G[70] = in[76] & in2[76];
    assign P[70] = in[76] ^ in2[76];
    assign G[71] = in[75] & in2[75];
    assign P[71] = in[75] ^ in2[75];
    assign G[72] = in[74] & in2[74];
    assign P[72] = in[74] ^ in2[74];
    assign G[73] = in[73] & in2[73];
    assign P[73] = in[73] ^ in2[73];
    assign G[74] = in[72] & in2[72];
    assign P[74] = in[72] ^ in2[72];
    assign G[75] = in[71] & in2[71];
    assign P[75] = in[71] ^ in2[71];
    assign G[76] = in[70] & in2[70];
    assign P[76] = in[70] ^ in2[70];
    assign G[77] = in[69] & in2[69];
    assign P[77] = in[69] ^ in2[69];
    assign G[78] = in[68] & in2[68];
    assign P[78] = in[68] ^ in2[68];
    assign G[79] = in[67] & in2[67];
    assign P[79] = in[67] ^ in2[67];
    assign G[80] = in[66] & in2[66];
    assign P[80] = in[66] ^ in2[66];
    assign G[81] = in[65] & in2[65];
    assign P[81] = in[65] ^ in2[65];
    assign G[82] = in[64] & in2[64];
    assign P[82] = in[64] ^ in2[64];
    assign G[83] = in[63] & in2[63];
    assign P[83] = in[63] ^ in2[63];
    assign G[84] = in[62] & in2[62];
    assign P[84] = in[62] ^ in2[62];
    assign G[85] = in[61] & in2[61];
    assign P[85] = in[61] ^ in2[61];
    assign G[86] = in[60] & in2[60];
    assign P[86] = in[60] ^ in2[60];
    assign G[87] = in[59] & in2[59];
    assign P[87] = in[59] ^ in2[59];
    assign G[88] = in[58] & in2[58];
    assign P[88] = in[58] ^ in2[58];
    assign G[89] = in[57] & in2[57];
    assign P[89] = in[57] ^ in2[57];
    assign G[90] = in[56] & in2[56];
    assign P[90] = in[56] ^ in2[56];
    assign G[91] = in[55] & in2[55];
    assign P[91] = in[55] ^ in2[55];
    assign G[92] = in[54] & in2[54];
    assign P[92] = in[54] ^ in2[54];
    assign G[93] = in[53] & in2[53];
    assign P[93] = in[53] ^ in2[53];
    assign G[94] = in[52] & in2[52];
    assign P[94] = in[52] ^ in2[52];
    assign G[95] = in[51] & in2[51];
    assign P[95] = in[51] ^ in2[51];
    assign G[96] = in[50] & in2[50];
    assign P[96] = in[50] ^ in2[50];
    assign G[97] = in[49] & in2[49];
    assign P[97] = in[49] ^ in2[49];
    assign G[98] = in[48] & in2[48];
    assign P[98] = in[48] ^ in2[48];
    assign G[99] = in[47] & in2[47];
    assign P[99] = in[47] ^ in2[47];
    assign G[100] = in[46] & in2[46];
    assign P[100] = in[46] ^ in2[46];
    assign G[101] = in[45] & in2[45];
    assign P[101] = in[45] ^ in2[45];
    assign G[102] = in[44] & in2[44];
    assign P[102] = in[44] ^ in2[44];
    assign G[103] = in[43] & in2[43];
    assign P[103] = in[43] ^ in2[43];
    assign G[104] = in[42] & in2[42];
    assign P[104] = in[42] ^ in2[42];
    assign G[105] = in[41] & in2[41];
    assign P[105] = in[41] ^ in2[41];
    assign G[106] = in[40] & in2[40];
    assign P[106] = in[40] ^ in2[40];
    assign G[107] = in[39] & in2[39];
    assign P[107] = in[39] ^ in2[39];
    assign G[108] = in[38] & in2[38];
    assign P[108] = in[38] ^ in2[38];
    assign G[109] = in[37] & in2[37];
    assign P[109] = in[37] ^ in2[37];
    assign G[110] = in[36] & in2[36];
    assign P[110] = in[36] ^ in2[36];
    assign G[111] = in[35] & in2[35];
    assign P[111] = in[35] ^ in2[35];
    assign G[112] = in[34] & in2[34];
    assign P[112] = in[34] ^ in2[34];
    assign G[113] = in[33] & in2[33];
    assign P[113] = in[33] ^ in2[33];
    assign G[114] = in[32] & in2[32];
    assign P[114] = in[32] ^ in2[32];
    assign G[115] = in[31] & in2[31];
    assign P[115] = in[31] ^ in2[31];
    assign G[116] = in[30] & in2[30];
    assign P[116] = in[30] ^ in2[30];
    assign G[117] = in[29] & in2[29];
    assign P[117] = in[29] ^ in2[29];
    assign G[118] = in[28] & in2[28];
    assign P[118] = in[28] ^ in2[28];
    assign G[119] = in[27] & in2[27];
    assign P[119] = in[27] ^ in2[27];
    assign G[120] = in[26] & in2[26];
    assign P[120] = in[26] ^ in2[26];
    assign G[121] = in[25] & in2[25];
    assign P[121] = in[25] ^ in2[25];
    assign G[122] = in[24] & in2[24];
    assign P[122] = in[24] ^ in2[24];
    assign G[123] = in[23] & in2[23];
    assign P[123] = in[23] ^ in2[23];
    assign G[124] = in[22] & in2[22];
    assign P[124] = in[22] ^ in2[22];
    assign G[125] = in[21] & in2[21];
    assign P[125] = in[21] ^ in2[21];
    assign G[126] = in[20] & in2[20];
    assign P[126] = in[20] ^ in2[20];
    assign G[127] = in[19] & in2[19];
    assign P[127] = in[19] ^ in2[19];
    assign G[128] = in[18] & in2[18];
    assign P[128] = in[18] ^ in2[18];
    assign G[129] = in[17] & in2[17];
    assign P[129] = in[17] ^ in2[17];
    assign G[130] = in[16] & in2[16];
    assign P[130] = in[16] ^ in2[16];
    assign G[131] = in[15] & in2[15];
    assign P[131] = in[15] ^ in2[15];
    assign G[132] = in[14] & in2[14];
    assign P[132] = in[14] ^ in2[14];
    assign G[133] = in[13] & in2[13];
    assign P[133] = in[13] ^ in2[13];
    assign G[134] = in[12] & in2[12];
    assign P[134] = in[12] ^ in2[12];
    assign G[135] = in[11] & in2[11];
    assign P[135] = in[11] ^ in2[11];
    assign G[136] = in[10] & in2[10];
    assign P[136] = in[10] ^ in2[10];
    assign G[137] = in[9] & in2[9];
    assign P[137] = in[9] ^ in2[9];
    assign G[138] = in[8] & in2[8];
    assign P[138] = in[8] ^ in2[8];
    assign G[139] = in[7] & in2[7];
    assign P[139] = in[7] ^ in2[7];
    assign G[140] = in[6] & in2[6];
    assign P[140] = in[6] ^ in2[6];
    assign G[141] = in[5] & in2[5];
    assign P[141] = in[5] ^ in2[5];
    assign G[142] = in[4] & in2[4];
    assign P[142] = in[4] ^ in2[4];
    assign G[143] = in[3] & in2[3];
    assign P[143] = in[3] ^ in2[3];
    assign G[144] = in[2] & in2[2];
    assign P[144] = in[2] ^ in2[2];
    assign G[145] = in[1] & in2[1];
    assign P[145] = in[1] ^ in2[1];
    assign G[146] = in[0] & in2[0];
    assign P[146] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign C[146] = G[145] | (P[145] & C[145]);
    assign cout = G[146] | (P[146] & C[146]);
    assign sum = P ^ C;
endmodule

module CLA146(output [145:0] sum, output cout, input [145:0] in1, input [145:0] in2;

    wire[145:0] G;
    wire[145:0] C;
    wire[145:0] P;

    assign G[0] = in[145] & in2[145];
    assign P[0] = in[145] ^ in2[145];
    assign G[1] = in[144] & in2[144];
    assign P[1] = in[144] ^ in2[144];
    assign G[2] = in[143] & in2[143];
    assign P[2] = in[143] ^ in2[143];
    assign G[3] = in[142] & in2[142];
    assign P[3] = in[142] ^ in2[142];
    assign G[4] = in[141] & in2[141];
    assign P[4] = in[141] ^ in2[141];
    assign G[5] = in[140] & in2[140];
    assign P[5] = in[140] ^ in2[140];
    assign G[6] = in[139] & in2[139];
    assign P[6] = in[139] ^ in2[139];
    assign G[7] = in[138] & in2[138];
    assign P[7] = in[138] ^ in2[138];
    assign G[8] = in[137] & in2[137];
    assign P[8] = in[137] ^ in2[137];
    assign G[9] = in[136] & in2[136];
    assign P[9] = in[136] ^ in2[136];
    assign G[10] = in[135] & in2[135];
    assign P[10] = in[135] ^ in2[135];
    assign G[11] = in[134] & in2[134];
    assign P[11] = in[134] ^ in2[134];
    assign G[12] = in[133] & in2[133];
    assign P[12] = in[133] ^ in2[133];
    assign G[13] = in[132] & in2[132];
    assign P[13] = in[132] ^ in2[132];
    assign G[14] = in[131] & in2[131];
    assign P[14] = in[131] ^ in2[131];
    assign G[15] = in[130] & in2[130];
    assign P[15] = in[130] ^ in2[130];
    assign G[16] = in[129] & in2[129];
    assign P[16] = in[129] ^ in2[129];
    assign G[17] = in[128] & in2[128];
    assign P[17] = in[128] ^ in2[128];
    assign G[18] = in[127] & in2[127];
    assign P[18] = in[127] ^ in2[127];
    assign G[19] = in[126] & in2[126];
    assign P[19] = in[126] ^ in2[126];
    assign G[20] = in[125] & in2[125];
    assign P[20] = in[125] ^ in2[125];
    assign G[21] = in[124] & in2[124];
    assign P[21] = in[124] ^ in2[124];
    assign G[22] = in[123] & in2[123];
    assign P[22] = in[123] ^ in2[123];
    assign G[23] = in[122] & in2[122];
    assign P[23] = in[122] ^ in2[122];
    assign G[24] = in[121] & in2[121];
    assign P[24] = in[121] ^ in2[121];
    assign G[25] = in[120] & in2[120];
    assign P[25] = in[120] ^ in2[120];
    assign G[26] = in[119] & in2[119];
    assign P[26] = in[119] ^ in2[119];
    assign G[27] = in[118] & in2[118];
    assign P[27] = in[118] ^ in2[118];
    assign G[28] = in[117] & in2[117];
    assign P[28] = in[117] ^ in2[117];
    assign G[29] = in[116] & in2[116];
    assign P[29] = in[116] ^ in2[116];
    assign G[30] = in[115] & in2[115];
    assign P[30] = in[115] ^ in2[115];
    assign G[31] = in[114] & in2[114];
    assign P[31] = in[114] ^ in2[114];
    assign G[32] = in[113] & in2[113];
    assign P[32] = in[113] ^ in2[113];
    assign G[33] = in[112] & in2[112];
    assign P[33] = in[112] ^ in2[112];
    assign G[34] = in[111] & in2[111];
    assign P[34] = in[111] ^ in2[111];
    assign G[35] = in[110] & in2[110];
    assign P[35] = in[110] ^ in2[110];
    assign G[36] = in[109] & in2[109];
    assign P[36] = in[109] ^ in2[109];
    assign G[37] = in[108] & in2[108];
    assign P[37] = in[108] ^ in2[108];
    assign G[38] = in[107] & in2[107];
    assign P[38] = in[107] ^ in2[107];
    assign G[39] = in[106] & in2[106];
    assign P[39] = in[106] ^ in2[106];
    assign G[40] = in[105] & in2[105];
    assign P[40] = in[105] ^ in2[105];
    assign G[41] = in[104] & in2[104];
    assign P[41] = in[104] ^ in2[104];
    assign G[42] = in[103] & in2[103];
    assign P[42] = in[103] ^ in2[103];
    assign G[43] = in[102] & in2[102];
    assign P[43] = in[102] ^ in2[102];
    assign G[44] = in[101] & in2[101];
    assign P[44] = in[101] ^ in2[101];
    assign G[45] = in[100] & in2[100];
    assign P[45] = in[100] ^ in2[100];
    assign G[46] = in[99] & in2[99];
    assign P[46] = in[99] ^ in2[99];
    assign G[47] = in[98] & in2[98];
    assign P[47] = in[98] ^ in2[98];
    assign G[48] = in[97] & in2[97];
    assign P[48] = in[97] ^ in2[97];
    assign G[49] = in[96] & in2[96];
    assign P[49] = in[96] ^ in2[96];
    assign G[50] = in[95] & in2[95];
    assign P[50] = in[95] ^ in2[95];
    assign G[51] = in[94] & in2[94];
    assign P[51] = in[94] ^ in2[94];
    assign G[52] = in[93] & in2[93];
    assign P[52] = in[93] ^ in2[93];
    assign G[53] = in[92] & in2[92];
    assign P[53] = in[92] ^ in2[92];
    assign G[54] = in[91] & in2[91];
    assign P[54] = in[91] ^ in2[91];
    assign G[55] = in[90] & in2[90];
    assign P[55] = in[90] ^ in2[90];
    assign G[56] = in[89] & in2[89];
    assign P[56] = in[89] ^ in2[89];
    assign G[57] = in[88] & in2[88];
    assign P[57] = in[88] ^ in2[88];
    assign G[58] = in[87] & in2[87];
    assign P[58] = in[87] ^ in2[87];
    assign G[59] = in[86] & in2[86];
    assign P[59] = in[86] ^ in2[86];
    assign G[60] = in[85] & in2[85];
    assign P[60] = in[85] ^ in2[85];
    assign G[61] = in[84] & in2[84];
    assign P[61] = in[84] ^ in2[84];
    assign G[62] = in[83] & in2[83];
    assign P[62] = in[83] ^ in2[83];
    assign G[63] = in[82] & in2[82];
    assign P[63] = in[82] ^ in2[82];
    assign G[64] = in[81] & in2[81];
    assign P[64] = in[81] ^ in2[81];
    assign G[65] = in[80] & in2[80];
    assign P[65] = in[80] ^ in2[80];
    assign G[66] = in[79] & in2[79];
    assign P[66] = in[79] ^ in2[79];
    assign G[67] = in[78] & in2[78];
    assign P[67] = in[78] ^ in2[78];
    assign G[68] = in[77] & in2[77];
    assign P[68] = in[77] ^ in2[77];
    assign G[69] = in[76] & in2[76];
    assign P[69] = in[76] ^ in2[76];
    assign G[70] = in[75] & in2[75];
    assign P[70] = in[75] ^ in2[75];
    assign G[71] = in[74] & in2[74];
    assign P[71] = in[74] ^ in2[74];
    assign G[72] = in[73] & in2[73];
    assign P[72] = in[73] ^ in2[73];
    assign G[73] = in[72] & in2[72];
    assign P[73] = in[72] ^ in2[72];
    assign G[74] = in[71] & in2[71];
    assign P[74] = in[71] ^ in2[71];
    assign G[75] = in[70] & in2[70];
    assign P[75] = in[70] ^ in2[70];
    assign G[76] = in[69] & in2[69];
    assign P[76] = in[69] ^ in2[69];
    assign G[77] = in[68] & in2[68];
    assign P[77] = in[68] ^ in2[68];
    assign G[78] = in[67] & in2[67];
    assign P[78] = in[67] ^ in2[67];
    assign G[79] = in[66] & in2[66];
    assign P[79] = in[66] ^ in2[66];
    assign G[80] = in[65] & in2[65];
    assign P[80] = in[65] ^ in2[65];
    assign G[81] = in[64] & in2[64];
    assign P[81] = in[64] ^ in2[64];
    assign G[82] = in[63] & in2[63];
    assign P[82] = in[63] ^ in2[63];
    assign G[83] = in[62] & in2[62];
    assign P[83] = in[62] ^ in2[62];
    assign G[84] = in[61] & in2[61];
    assign P[84] = in[61] ^ in2[61];
    assign G[85] = in[60] & in2[60];
    assign P[85] = in[60] ^ in2[60];
    assign G[86] = in[59] & in2[59];
    assign P[86] = in[59] ^ in2[59];
    assign G[87] = in[58] & in2[58];
    assign P[87] = in[58] ^ in2[58];
    assign G[88] = in[57] & in2[57];
    assign P[88] = in[57] ^ in2[57];
    assign G[89] = in[56] & in2[56];
    assign P[89] = in[56] ^ in2[56];
    assign G[90] = in[55] & in2[55];
    assign P[90] = in[55] ^ in2[55];
    assign G[91] = in[54] & in2[54];
    assign P[91] = in[54] ^ in2[54];
    assign G[92] = in[53] & in2[53];
    assign P[92] = in[53] ^ in2[53];
    assign G[93] = in[52] & in2[52];
    assign P[93] = in[52] ^ in2[52];
    assign G[94] = in[51] & in2[51];
    assign P[94] = in[51] ^ in2[51];
    assign G[95] = in[50] & in2[50];
    assign P[95] = in[50] ^ in2[50];
    assign G[96] = in[49] & in2[49];
    assign P[96] = in[49] ^ in2[49];
    assign G[97] = in[48] & in2[48];
    assign P[97] = in[48] ^ in2[48];
    assign G[98] = in[47] & in2[47];
    assign P[98] = in[47] ^ in2[47];
    assign G[99] = in[46] & in2[46];
    assign P[99] = in[46] ^ in2[46];
    assign G[100] = in[45] & in2[45];
    assign P[100] = in[45] ^ in2[45];
    assign G[101] = in[44] & in2[44];
    assign P[101] = in[44] ^ in2[44];
    assign G[102] = in[43] & in2[43];
    assign P[102] = in[43] ^ in2[43];
    assign G[103] = in[42] & in2[42];
    assign P[103] = in[42] ^ in2[42];
    assign G[104] = in[41] & in2[41];
    assign P[104] = in[41] ^ in2[41];
    assign G[105] = in[40] & in2[40];
    assign P[105] = in[40] ^ in2[40];
    assign G[106] = in[39] & in2[39];
    assign P[106] = in[39] ^ in2[39];
    assign G[107] = in[38] & in2[38];
    assign P[107] = in[38] ^ in2[38];
    assign G[108] = in[37] & in2[37];
    assign P[108] = in[37] ^ in2[37];
    assign G[109] = in[36] & in2[36];
    assign P[109] = in[36] ^ in2[36];
    assign G[110] = in[35] & in2[35];
    assign P[110] = in[35] ^ in2[35];
    assign G[111] = in[34] & in2[34];
    assign P[111] = in[34] ^ in2[34];
    assign G[112] = in[33] & in2[33];
    assign P[112] = in[33] ^ in2[33];
    assign G[113] = in[32] & in2[32];
    assign P[113] = in[32] ^ in2[32];
    assign G[114] = in[31] & in2[31];
    assign P[114] = in[31] ^ in2[31];
    assign G[115] = in[30] & in2[30];
    assign P[115] = in[30] ^ in2[30];
    assign G[116] = in[29] & in2[29];
    assign P[116] = in[29] ^ in2[29];
    assign G[117] = in[28] & in2[28];
    assign P[117] = in[28] ^ in2[28];
    assign G[118] = in[27] & in2[27];
    assign P[118] = in[27] ^ in2[27];
    assign G[119] = in[26] & in2[26];
    assign P[119] = in[26] ^ in2[26];
    assign G[120] = in[25] & in2[25];
    assign P[120] = in[25] ^ in2[25];
    assign G[121] = in[24] & in2[24];
    assign P[121] = in[24] ^ in2[24];
    assign G[122] = in[23] & in2[23];
    assign P[122] = in[23] ^ in2[23];
    assign G[123] = in[22] & in2[22];
    assign P[123] = in[22] ^ in2[22];
    assign G[124] = in[21] & in2[21];
    assign P[124] = in[21] ^ in2[21];
    assign G[125] = in[20] & in2[20];
    assign P[125] = in[20] ^ in2[20];
    assign G[126] = in[19] & in2[19];
    assign P[126] = in[19] ^ in2[19];
    assign G[127] = in[18] & in2[18];
    assign P[127] = in[18] ^ in2[18];
    assign G[128] = in[17] & in2[17];
    assign P[128] = in[17] ^ in2[17];
    assign G[129] = in[16] & in2[16];
    assign P[129] = in[16] ^ in2[16];
    assign G[130] = in[15] & in2[15];
    assign P[130] = in[15] ^ in2[15];
    assign G[131] = in[14] & in2[14];
    assign P[131] = in[14] ^ in2[14];
    assign G[132] = in[13] & in2[13];
    assign P[132] = in[13] ^ in2[13];
    assign G[133] = in[12] & in2[12];
    assign P[133] = in[12] ^ in2[12];
    assign G[134] = in[11] & in2[11];
    assign P[134] = in[11] ^ in2[11];
    assign G[135] = in[10] & in2[10];
    assign P[135] = in[10] ^ in2[10];
    assign G[136] = in[9] & in2[9];
    assign P[136] = in[9] ^ in2[9];
    assign G[137] = in[8] & in2[8];
    assign P[137] = in[8] ^ in2[8];
    assign G[138] = in[7] & in2[7];
    assign P[138] = in[7] ^ in2[7];
    assign G[139] = in[6] & in2[6];
    assign P[139] = in[6] ^ in2[6];
    assign G[140] = in[5] & in2[5];
    assign P[140] = in[5] ^ in2[5];
    assign G[141] = in[4] & in2[4];
    assign P[141] = in[4] ^ in2[4];
    assign G[142] = in[3] & in2[3];
    assign P[142] = in[3] ^ in2[3];
    assign G[143] = in[2] & in2[2];
    assign P[143] = in[2] ^ in2[2];
    assign G[144] = in[1] & in2[1];
    assign P[144] = in[1] ^ in2[1];
    assign G[145] = in[0] & in2[0];
    assign P[145] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign C[145] = G[144] | (P[144] & C[144]);
    assign cout = G[145] | (P[145] & C[145]);
    assign sum = P ^ C;
endmodule

module CLA145(output [144:0] sum, output cout, input [144:0] in1, input [144:0] in2;

    wire[144:0] G;
    wire[144:0] C;
    wire[144:0] P;

    assign G[0] = in[144] & in2[144];
    assign P[0] = in[144] ^ in2[144];
    assign G[1] = in[143] & in2[143];
    assign P[1] = in[143] ^ in2[143];
    assign G[2] = in[142] & in2[142];
    assign P[2] = in[142] ^ in2[142];
    assign G[3] = in[141] & in2[141];
    assign P[3] = in[141] ^ in2[141];
    assign G[4] = in[140] & in2[140];
    assign P[4] = in[140] ^ in2[140];
    assign G[5] = in[139] & in2[139];
    assign P[5] = in[139] ^ in2[139];
    assign G[6] = in[138] & in2[138];
    assign P[6] = in[138] ^ in2[138];
    assign G[7] = in[137] & in2[137];
    assign P[7] = in[137] ^ in2[137];
    assign G[8] = in[136] & in2[136];
    assign P[8] = in[136] ^ in2[136];
    assign G[9] = in[135] & in2[135];
    assign P[9] = in[135] ^ in2[135];
    assign G[10] = in[134] & in2[134];
    assign P[10] = in[134] ^ in2[134];
    assign G[11] = in[133] & in2[133];
    assign P[11] = in[133] ^ in2[133];
    assign G[12] = in[132] & in2[132];
    assign P[12] = in[132] ^ in2[132];
    assign G[13] = in[131] & in2[131];
    assign P[13] = in[131] ^ in2[131];
    assign G[14] = in[130] & in2[130];
    assign P[14] = in[130] ^ in2[130];
    assign G[15] = in[129] & in2[129];
    assign P[15] = in[129] ^ in2[129];
    assign G[16] = in[128] & in2[128];
    assign P[16] = in[128] ^ in2[128];
    assign G[17] = in[127] & in2[127];
    assign P[17] = in[127] ^ in2[127];
    assign G[18] = in[126] & in2[126];
    assign P[18] = in[126] ^ in2[126];
    assign G[19] = in[125] & in2[125];
    assign P[19] = in[125] ^ in2[125];
    assign G[20] = in[124] & in2[124];
    assign P[20] = in[124] ^ in2[124];
    assign G[21] = in[123] & in2[123];
    assign P[21] = in[123] ^ in2[123];
    assign G[22] = in[122] & in2[122];
    assign P[22] = in[122] ^ in2[122];
    assign G[23] = in[121] & in2[121];
    assign P[23] = in[121] ^ in2[121];
    assign G[24] = in[120] & in2[120];
    assign P[24] = in[120] ^ in2[120];
    assign G[25] = in[119] & in2[119];
    assign P[25] = in[119] ^ in2[119];
    assign G[26] = in[118] & in2[118];
    assign P[26] = in[118] ^ in2[118];
    assign G[27] = in[117] & in2[117];
    assign P[27] = in[117] ^ in2[117];
    assign G[28] = in[116] & in2[116];
    assign P[28] = in[116] ^ in2[116];
    assign G[29] = in[115] & in2[115];
    assign P[29] = in[115] ^ in2[115];
    assign G[30] = in[114] & in2[114];
    assign P[30] = in[114] ^ in2[114];
    assign G[31] = in[113] & in2[113];
    assign P[31] = in[113] ^ in2[113];
    assign G[32] = in[112] & in2[112];
    assign P[32] = in[112] ^ in2[112];
    assign G[33] = in[111] & in2[111];
    assign P[33] = in[111] ^ in2[111];
    assign G[34] = in[110] & in2[110];
    assign P[34] = in[110] ^ in2[110];
    assign G[35] = in[109] & in2[109];
    assign P[35] = in[109] ^ in2[109];
    assign G[36] = in[108] & in2[108];
    assign P[36] = in[108] ^ in2[108];
    assign G[37] = in[107] & in2[107];
    assign P[37] = in[107] ^ in2[107];
    assign G[38] = in[106] & in2[106];
    assign P[38] = in[106] ^ in2[106];
    assign G[39] = in[105] & in2[105];
    assign P[39] = in[105] ^ in2[105];
    assign G[40] = in[104] & in2[104];
    assign P[40] = in[104] ^ in2[104];
    assign G[41] = in[103] & in2[103];
    assign P[41] = in[103] ^ in2[103];
    assign G[42] = in[102] & in2[102];
    assign P[42] = in[102] ^ in2[102];
    assign G[43] = in[101] & in2[101];
    assign P[43] = in[101] ^ in2[101];
    assign G[44] = in[100] & in2[100];
    assign P[44] = in[100] ^ in2[100];
    assign G[45] = in[99] & in2[99];
    assign P[45] = in[99] ^ in2[99];
    assign G[46] = in[98] & in2[98];
    assign P[46] = in[98] ^ in2[98];
    assign G[47] = in[97] & in2[97];
    assign P[47] = in[97] ^ in2[97];
    assign G[48] = in[96] & in2[96];
    assign P[48] = in[96] ^ in2[96];
    assign G[49] = in[95] & in2[95];
    assign P[49] = in[95] ^ in2[95];
    assign G[50] = in[94] & in2[94];
    assign P[50] = in[94] ^ in2[94];
    assign G[51] = in[93] & in2[93];
    assign P[51] = in[93] ^ in2[93];
    assign G[52] = in[92] & in2[92];
    assign P[52] = in[92] ^ in2[92];
    assign G[53] = in[91] & in2[91];
    assign P[53] = in[91] ^ in2[91];
    assign G[54] = in[90] & in2[90];
    assign P[54] = in[90] ^ in2[90];
    assign G[55] = in[89] & in2[89];
    assign P[55] = in[89] ^ in2[89];
    assign G[56] = in[88] & in2[88];
    assign P[56] = in[88] ^ in2[88];
    assign G[57] = in[87] & in2[87];
    assign P[57] = in[87] ^ in2[87];
    assign G[58] = in[86] & in2[86];
    assign P[58] = in[86] ^ in2[86];
    assign G[59] = in[85] & in2[85];
    assign P[59] = in[85] ^ in2[85];
    assign G[60] = in[84] & in2[84];
    assign P[60] = in[84] ^ in2[84];
    assign G[61] = in[83] & in2[83];
    assign P[61] = in[83] ^ in2[83];
    assign G[62] = in[82] & in2[82];
    assign P[62] = in[82] ^ in2[82];
    assign G[63] = in[81] & in2[81];
    assign P[63] = in[81] ^ in2[81];
    assign G[64] = in[80] & in2[80];
    assign P[64] = in[80] ^ in2[80];
    assign G[65] = in[79] & in2[79];
    assign P[65] = in[79] ^ in2[79];
    assign G[66] = in[78] & in2[78];
    assign P[66] = in[78] ^ in2[78];
    assign G[67] = in[77] & in2[77];
    assign P[67] = in[77] ^ in2[77];
    assign G[68] = in[76] & in2[76];
    assign P[68] = in[76] ^ in2[76];
    assign G[69] = in[75] & in2[75];
    assign P[69] = in[75] ^ in2[75];
    assign G[70] = in[74] & in2[74];
    assign P[70] = in[74] ^ in2[74];
    assign G[71] = in[73] & in2[73];
    assign P[71] = in[73] ^ in2[73];
    assign G[72] = in[72] & in2[72];
    assign P[72] = in[72] ^ in2[72];
    assign G[73] = in[71] & in2[71];
    assign P[73] = in[71] ^ in2[71];
    assign G[74] = in[70] & in2[70];
    assign P[74] = in[70] ^ in2[70];
    assign G[75] = in[69] & in2[69];
    assign P[75] = in[69] ^ in2[69];
    assign G[76] = in[68] & in2[68];
    assign P[76] = in[68] ^ in2[68];
    assign G[77] = in[67] & in2[67];
    assign P[77] = in[67] ^ in2[67];
    assign G[78] = in[66] & in2[66];
    assign P[78] = in[66] ^ in2[66];
    assign G[79] = in[65] & in2[65];
    assign P[79] = in[65] ^ in2[65];
    assign G[80] = in[64] & in2[64];
    assign P[80] = in[64] ^ in2[64];
    assign G[81] = in[63] & in2[63];
    assign P[81] = in[63] ^ in2[63];
    assign G[82] = in[62] & in2[62];
    assign P[82] = in[62] ^ in2[62];
    assign G[83] = in[61] & in2[61];
    assign P[83] = in[61] ^ in2[61];
    assign G[84] = in[60] & in2[60];
    assign P[84] = in[60] ^ in2[60];
    assign G[85] = in[59] & in2[59];
    assign P[85] = in[59] ^ in2[59];
    assign G[86] = in[58] & in2[58];
    assign P[86] = in[58] ^ in2[58];
    assign G[87] = in[57] & in2[57];
    assign P[87] = in[57] ^ in2[57];
    assign G[88] = in[56] & in2[56];
    assign P[88] = in[56] ^ in2[56];
    assign G[89] = in[55] & in2[55];
    assign P[89] = in[55] ^ in2[55];
    assign G[90] = in[54] & in2[54];
    assign P[90] = in[54] ^ in2[54];
    assign G[91] = in[53] & in2[53];
    assign P[91] = in[53] ^ in2[53];
    assign G[92] = in[52] & in2[52];
    assign P[92] = in[52] ^ in2[52];
    assign G[93] = in[51] & in2[51];
    assign P[93] = in[51] ^ in2[51];
    assign G[94] = in[50] & in2[50];
    assign P[94] = in[50] ^ in2[50];
    assign G[95] = in[49] & in2[49];
    assign P[95] = in[49] ^ in2[49];
    assign G[96] = in[48] & in2[48];
    assign P[96] = in[48] ^ in2[48];
    assign G[97] = in[47] & in2[47];
    assign P[97] = in[47] ^ in2[47];
    assign G[98] = in[46] & in2[46];
    assign P[98] = in[46] ^ in2[46];
    assign G[99] = in[45] & in2[45];
    assign P[99] = in[45] ^ in2[45];
    assign G[100] = in[44] & in2[44];
    assign P[100] = in[44] ^ in2[44];
    assign G[101] = in[43] & in2[43];
    assign P[101] = in[43] ^ in2[43];
    assign G[102] = in[42] & in2[42];
    assign P[102] = in[42] ^ in2[42];
    assign G[103] = in[41] & in2[41];
    assign P[103] = in[41] ^ in2[41];
    assign G[104] = in[40] & in2[40];
    assign P[104] = in[40] ^ in2[40];
    assign G[105] = in[39] & in2[39];
    assign P[105] = in[39] ^ in2[39];
    assign G[106] = in[38] & in2[38];
    assign P[106] = in[38] ^ in2[38];
    assign G[107] = in[37] & in2[37];
    assign P[107] = in[37] ^ in2[37];
    assign G[108] = in[36] & in2[36];
    assign P[108] = in[36] ^ in2[36];
    assign G[109] = in[35] & in2[35];
    assign P[109] = in[35] ^ in2[35];
    assign G[110] = in[34] & in2[34];
    assign P[110] = in[34] ^ in2[34];
    assign G[111] = in[33] & in2[33];
    assign P[111] = in[33] ^ in2[33];
    assign G[112] = in[32] & in2[32];
    assign P[112] = in[32] ^ in2[32];
    assign G[113] = in[31] & in2[31];
    assign P[113] = in[31] ^ in2[31];
    assign G[114] = in[30] & in2[30];
    assign P[114] = in[30] ^ in2[30];
    assign G[115] = in[29] & in2[29];
    assign P[115] = in[29] ^ in2[29];
    assign G[116] = in[28] & in2[28];
    assign P[116] = in[28] ^ in2[28];
    assign G[117] = in[27] & in2[27];
    assign P[117] = in[27] ^ in2[27];
    assign G[118] = in[26] & in2[26];
    assign P[118] = in[26] ^ in2[26];
    assign G[119] = in[25] & in2[25];
    assign P[119] = in[25] ^ in2[25];
    assign G[120] = in[24] & in2[24];
    assign P[120] = in[24] ^ in2[24];
    assign G[121] = in[23] & in2[23];
    assign P[121] = in[23] ^ in2[23];
    assign G[122] = in[22] & in2[22];
    assign P[122] = in[22] ^ in2[22];
    assign G[123] = in[21] & in2[21];
    assign P[123] = in[21] ^ in2[21];
    assign G[124] = in[20] & in2[20];
    assign P[124] = in[20] ^ in2[20];
    assign G[125] = in[19] & in2[19];
    assign P[125] = in[19] ^ in2[19];
    assign G[126] = in[18] & in2[18];
    assign P[126] = in[18] ^ in2[18];
    assign G[127] = in[17] & in2[17];
    assign P[127] = in[17] ^ in2[17];
    assign G[128] = in[16] & in2[16];
    assign P[128] = in[16] ^ in2[16];
    assign G[129] = in[15] & in2[15];
    assign P[129] = in[15] ^ in2[15];
    assign G[130] = in[14] & in2[14];
    assign P[130] = in[14] ^ in2[14];
    assign G[131] = in[13] & in2[13];
    assign P[131] = in[13] ^ in2[13];
    assign G[132] = in[12] & in2[12];
    assign P[132] = in[12] ^ in2[12];
    assign G[133] = in[11] & in2[11];
    assign P[133] = in[11] ^ in2[11];
    assign G[134] = in[10] & in2[10];
    assign P[134] = in[10] ^ in2[10];
    assign G[135] = in[9] & in2[9];
    assign P[135] = in[9] ^ in2[9];
    assign G[136] = in[8] & in2[8];
    assign P[136] = in[8] ^ in2[8];
    assign G[137] = in[7] & in2[7];
    assign P[137] = in[7] ^ in2[7];
    assign G[138] = in[6] & in2[6];
    assign P[138] = in[6] ^ in2[6];
    assign G[139] = in[5] & in2[5];
    assign P[139] = in[5] ^ in2[5];
    assign G[140] = in[4] & in2[4];
    assign P[140] = in[4] ^ in2[4];
    assign G[141] = in[3] & in2[3];
    assign P[141] = in[3] ^ in2[3];
    assign G[142] = in[2] & in2[2];
    assign P[142] = in[2] ^ in2[2];
    assign G[143] = in[1] & in2[1];
    assign P[143] = in[1] ^ in2[1];
    assign G[144] = in[0] & in2[0];
    assign P[144] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign C[144] = G[143] | (P[143] & C[143]);
    assign cout = G[144] | (P[144] & C[144]);
    assign sum = P ^ C;
endmodule

module CLA144(output [143:0] sum, output cout, input [143:0] in1, input [143:0] in2;

    wire[143:0] G;
    wire[143:0] C;
    wire[143:0] P;

    assign G[0] = in[143] & in2[143];
    assign P[0] = in[143] ^ in2[143];
    assign G[1] = in[142] & in2[142];
    assign P[1] = in[142] ^ in2[142];
    assign G[2] = in[141] & in2[141];
    assign P[2] = in[141] ^ in2[141];
    assign G[3] = in[140] & in2[140];
    assign P[3] = in[140] ^ in2[140];
    assign G[4] = in[139] & in2[139];
    assign P[4] = in[139] ^ in2[139];
    assign G[5] = in[138] & in2[138];
    assign P[5] = in[138] ^ in2[138];
    assign G[6] = in[137] & in2[137];
    assign P[6] = in[137] ^ in2[137];
    assign G[7] = in[136] & in2[136];
    assign P[7] = in[136] ^ in2[136];
    assign G[8] = in[135] & in2[135];
    assign P[8] = in[135] ^ in2[135];
    assign G[9] = in[134] & in2[134];
    assign P[9] = in[134] ^ in2[134];
    assign G[10] = in[133] & in2[133];
    assign P[10] = in[133] ^ in2[133];
    assign G[11] = in[132] & in2[132];
    assign P[11] = in[132] ^ in2[132];
    assign G[12] = in[131] & in2[131];
    assign P[12] = in[131] ^ in2[131];
    assign G[13] = in[130] & in2[130];
    assign P[13] = in[130] ^ in2[130];
    assign G[14] = in[129] & in2[129];
    assign P[14] = in[129] ^ in2[129];
    assign G[15] = in[128] & in2[128];
    assign P[15] = in[128] ^ in2[128];
    assign G[16] = in[127] & in2[127];
    assign P[16] = in[127] ^ in2[127];
    assign G[17] = in[126] & in2[126];
    assign P[17] = in[126] ^ in2[126];
    assign G[18] = in[125] & in2[125];
    assign P[18] = in[125] ^ in2[125];
    assign G[19] = in[124] & in2[124];
    assign P[19] = in[124] ^ in2[124];
    assign G[20] = in[123] & in2[123];
    assign P[20] = in[123] ^ in2[123];
    assign G[21] = in[122] & in2[122];
    assign P[21] = in[122] ^ in2[122];
    assign G[22] = in[121] & in2[121];
    assign P[22] = in[121] ^ in2[121];
    assign G[23] = in[120] & in2[120];
    assign P[23] = in[120] ^ in2[120];
    assign G[24] = in[119] & in2[119];
    assign P[24] = in[119] ^ in2[119];
    assign G[25] = in[118] & in2[118];
    assign P[25] = in[118] ^ in2[118];
    assign G[26] = in[117] & in2[117];
    assign P[26] = in[117] ^ in2[117];
    assign G[27] = in[116] & in2[116];
    assign P[27] = in[116] ^ in2[116];
    assign G[28] = in[115] & in2[115];
    assign P[28] = in[115] ^ in2[115];
    assign G[29] = in[114] & in2[114];
    assign P[29] = in[114] ^ in2[114];
    assign G[30] = in[113] & in2[113];
    assign P[30] = in[113] ^ in2[113];
    assign G[31] = in[112] & in2[112];
    assign P[31] = in[112] ^ in2[112];
    assign G[32] = in[111] & in2[111];
    assign P[32] = in[111] ^ in2[111];
    assign G[33] = in[110] & in2[110];
    assign P[33] = in[110] ^ in2[110];
    assign G[34] = in[109] & in2[109];
    assign P[34] = in[109] ^ in2[109];
    assign G[35] = in[108] & in2[108];
    assign P[35] = in[108] ^ in2[108];
    assign G[36] = in[107] & in2[107];
    assign P[36] = in[107] ^ in2[107];
    assign G[37] = in[106] & in2[106];
    assign P[37] = in[106] ^ in2[106];
    assign G[38] = in[105] & in2[105];
    assign P[38] = in[105] ^ in2[105];
    assign G[39] = in[104] & in2[104];
    assign P[39] = in[104] ^ in2[104];
    assign G[40] = in[103] & in2[103];
    assign P[40] = in[103] ^ in2[103];
    assign G[41] = in[102] & in2[102];
    assign P[41] = in[102] ^ in2[102];
    assign G[42] = in[101] & in2[101];
    assign P[42] = in[101] ^ in2[101];
    assign G[43] = in[100] & in2[100];
    assign P[43] = in[100] ^ in2[100];
    assign G[44] = in[99] & in2[99];
    assign P[44] = in[99] ^ in2[99];
    assign G[45] = in[98] & in2[98];
    assign P[45] = in[98] ^ in2[98];
    assign G[46] = in[97] & in2[97];
    assign P[46] = in[97] ^ in2[97];
    assign G[47] = in[96] & in2[96];
    assign P[47] = in[96] ^ in2[96];
    assign G[48] = in[95] & in2[95];
    assign P[48] = in[95] ^ in2[95];
    assign G[49] = in[94] & in2[94];
    assign P[49] = in[94] ^ in2[94];
    assign G[50] = in[93] & in2[93];
    assign P[50] = in[93] ^ in2[93];
    assign G[51] = in[92] & in2[92];
    assign P[51] = in[92] ^ in2[92];
    assign G[52] = in[91] & in2[91];
    assign P[52] = in[91] ^ in2[91];
    assign G[53] = in[90] & in2[90];
    assign P[53] = in[90] ^ in2[90];
    assign G[54] = in[89] & in2[89];
    assign P[54] = in[89] ^ in2[89];
    assign G[55] = in[88] & in2[88];
    assign P[55] = in[88] ^ in2[88];
    assign G[56] = in[87] & in2[87];
    assign P[56] = in[87] ^ in2[87];
    assign G[57] = in[86] & in2[86];
    assign P[57] = in[86] ^ in2[86];
    assign G[58] = in[85] & in2[85];
    assign P[58] = in[85] ^ in2[85];
    assign G[59] = in[84] & in2[84];
    assign P[59] = in[84] ^ in2[84];
    assign G[60] = in[83] & in2[83];
    assign P[60] = in[83] ^ in2[83];
    assign G[61] = in[82] & in2[82];
    assign P[61] = in[82] ^ in2[82];
    assign G[62] = in[81] & in2[81];
    assign P[62] = in[81] ^ in2[81];
    assign G[63] = in[80] & in2[80];
    assign P[63] = in[80] ^ in2[80];
    assign G[64] = in[79] & in2[79];
    assign P[64] = in[79] ^ in2[79];
    assign G[65] = in[78] & in2[78];
    assign P[65] = in[78] ^ in2[78];
    assign G[66] = in[77] & in2[77];
    assign P[66] = in[77] ^ in2[77];
    assign G[67] = in[76] & in2[76];
    assign P[67] = in[76] ^ in2[76];
    assign G[68] = in[75] & in2[75];
    assign P[68] = in[75] ^ in2[75];
    assign G[69] = in[74] & in2[74];
    assign P[69] = in[74] ^ in2[74];
    assign G[70] = in[73] & in2[73];
    assign P[70] = in[73] ^ in2[73];
    assign G[71] = in[72] & in2[72];
    assign P[71] = in[72] ^ in2[72];
    assign G[72] = in[71] & in2[71];
    assign P[72] = in[71] ^ in2[71];
    assign G[73] = in[70] & in2[70];
    assign P[73] = in[70] ^ in2[70];
    assign G[74] = in[69] & in2[69];
    assign P[74] = in[69] ^ in2[69];
    assign G[75] = in[68] & in2[68];
    assign P[75] = in[68] ^ in2[68];
    assign G[76] = in[67] & in2[67];
    assign P[76] = in[67] ^ in2[67];
    assign G[77] = in[66] & in2[66];
    assign P[77] = in[66] ^ in2[66];
    assign G[78] = in[65] & in2[65];
    assign P[78] = in[65] ^ in2[65];
    assign G[79] = in[64] & in2[64];
    assign P[79] = in[64] ^ in2[64];
    assign G[80] = in[63] & in2[63];
    assign P[80] = in[63] ^ in2[63];
    assign G[81] = in[62] & in2[62];
    assign P[81] = in[62] ^ in2[62];
    assign G[82] = in[61] & in2[61];
    assign P[82] = in[61] ^ in2[61];
    assign G[83] = in[60] & in2[60];
    assign P[83] = in[60] ^ in2[60];
    assign G[84] = in[59] & in2[59];
    assign P[84] = in[59] ^ in2[59];
    assign G[85] = in[58] & in2[58];
    assign P[85] = in[58] ^ in2[58];
    assign G[86] = in[57] & in2[57];
    assign P[86] = in[57] ^ in2[57];
    assign G[87] = in[56] & in2[56];
    assign P[87] = in[56] ^ in2[56];
    assign G[88] = in[55] & in2[55];
    assign P[88] = in[55] ^ in2[55];
    assign G[89] = in[54] & in2[54];
    assign P[89] = in[54] ^ in2[54];
    assign G[90] = in[53] & in2[53];
    assign P[90] = in[53] ^ in2[53];
    assign G[91] = in[52] & in2[52];
    assign P[91] = in[52] ^ in2[52];
    assign G[92] = in[51] & in2[51];
    assign P[92] = in[51] ^ in2[51];
    assign G[93] = in[50] & in2[50];
    assign P[93] = in[50] ^ in2[50];
    assign G[94] = in[49] & in2[49];
    assign P[94] = in[49] ^ in2[49];
    assign G[95] = in[48] & in2[48];
    assign P[95] = in[48] ^ in2[48];
    assign G[96] = in[47] & in2[47];
    assign P[96] = in[47] ^ in2[47];
    assign G[97] = in[46] & in2[46];
    assign P[97] = in[46] ^ in2[46];
    assign G[98] = in[45] & in2[45];
    assign P[98] = in[45] ^ in2[45];
    assign G[99] = in[44] & in2[44];
    assign P[99] = in[44] ^ in2[44];
    assign G[100] = in[43] & in2[43];
    assign P[100] = in[43] ^ in2[43];
    assign G[101] = in[42] & in2[42];
    assign P[101] = in[42] ^ in2[42];
    assign G[102] = in[41] & in2[41];
    assign P[102] = in[41] ^ in2[41];
    assign G[103] = in[40] & in2[40];
    assign P[103] = in[40] ^ in2[40];
    assign G[104] = in[39] & in2[39];
    assign P[104] = in[39] ^ in2[39];
    assign G[105] = in[38] & in2[38];
    assign P[105] = in[38] ^ in2[38];
    assign G[106] = in[37] & in2[37];
    assign P[106] = in[37] ^ in2[37];
    assign G[107] = in[36] & in2[36];
    assign P[107] = in[36] ^ in2[36];
    assign G[108] = in[35] & in2[35];
    assign P[108] = in[35] ^ in2[35];
    assign G[109] = in[34] & in2[34];
    assign P[109] = in[34] ^ in2[34];
    assign G[110] = in[33] & in2[33];
    assign P[110] = in[33] ^ in2[33];
    assign G[111] = in[32] & in2[32];
    assign P[111] = in[32] ^ in2[32];
    assign G[112] = in[31] & in2[31];
    assign P[112] = in[31] ^ in2[31];
    assign G[113] = in[30] & in2[30];
    assign P[113] = in[30] ^ in2[30];
    assign G[114] = in[29] & in2[29];
    assign P[114] = in[29] ^ in2[29];
    assign G[115] = in[28] & in2[28];
    assign P[115] = in[28] ^ in2[28];
    assign G[116] = in[27] & in2[27];
    assign P[116] = in[27] ^ in2[27];
    assign G[117] = in[26] & in2[26];
    assign P[117] = in[26] ^ in2[26];
    assign G[118] = in[25] & in2[25];
    assign P[118] = in[25] ^ in2[25];
    assign G[119] = in[24] & in2[24];
    assign P[119] = in[24] ^ in2[24];
    assign G[120] = in[23] & in2[23];
    assign P[120] = in[23] ^ in2[23];
    assign G[121] = in[22] & in2[22];
    assign P[121] = in[22] ^ in2[22];
    assign G[122] = in[21] & in2[21];
    assign P[122] = in[21] ^ in2[21];
    assign G[123] = in[20] & in2[20];
    assign P[123] = in[20] ^ in2[20];
    assign G[124] = in[19] & in2[19];
    assign P[124] = in[19] ^ in2[19];
    assign G[125] = in[18] & in2[18];
    assign P[125] = in[18] ^ in2[18];
    assign G[126] = in[17] & in2[17];
    assign P[126] = in[17] ^ in2[17];
    assign G[127] = in[16] & in2[16];
    assign P[127] = in[16] ^ in2[16];
    assign G[128] = in[15] & in2[15];
    assign P[128] = in[15] ^ in2[15];
    assign G[129] = in[14] & in2[14];
    assign P[129] = in[14] ^ in2[14];
    assign G[130] = in[13] & in2[13];
    assign P[130] = in[13] ^ in2[13];
    assign G[131] = in[12] & in2[12];
    assign P[131] = in[12] ^ in2[12];
    assign G[132] = in[11] & in2[11];
    assign P[132] = in[11] ^ in2[11];
    assign G[133] = in[10] & in2[10];
    assign P[133] = in[10] ^ in2[10];
    assign G[134] = in[9] & in2[9];
    assign P[134] = in[9] ^ in2[9];
    assign G[135] = in[8] & in2[8];
    assign P[135] = in[8] ^ in2[8];
    assign G[136] = in[7] & in2[7];
    assign P[136] = in[7] ^ in2[7];
    assign G[137] = in[6] & in2[6];
    assign P[137] = in[6] ^ in2[6];
    assign G[138] = in[5] & in2[5];
    assign P[138] = in[5] ^ in2[5];
    assign G[139] = in[4] & in2[4];
    assign P[139] = in[4] ^ in2[4];
    assign G[140] = in[3] & in2[3];
    assign P[140] = in[3] ^ in2[3];
    assign G[141] = in[2] & in2[2];
    assign P[141] = in[2] ^ in2[2];
    assign G[142] = in[1] & in2[1];
    assign P[142] = in[1] ^ in2[1];
    assign G[143] = in[0] & in2[0];
    assign P[143] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign C[143] = G[142] | (P[142] & C[142]);
    assign cout = G[143] | (P[143] & C[143]);
    assign sum = P ^ C;
endmodule

module CLA143(output [142:0] sum, output cout, input [142:0] in1, input [142:0] in2;

    wire[142:0] G;
    wire[142:0] C;
    wire[142:0] P;

    assign G[0] = in[142] & in2[142];
    assign P[0] = in[142] ^ in2[142];
    assign G[1] = in[141] & in2[141];
    assign P[1] = in[141] ^ in2[141];
    assign G[2] = in[140] & in2[140];
    assign P[2] = in[140] ^ in2[140];
    assign G[3] = in[139] & in2[139];
    assign P[3] = in[139] ^ in2[139];
    assign G[4] = in[138] & in2[138];
    assign P[4] = in[138] ^ in2[138];
    assign G[5] = in[137] & in2[137];
    assign P[5] = in[137] ^ in2[137];
    assign G[6] = in[136] & in2[136];
    assign P[6] = in[136] ^ in2[136];
    assign G[7] = in[135] & in2[135];
    assign P[7] = in[135] ^ in2[135];
    assign G[8] = in[134] & in2[134];
    assign P[8] = in[134] ^ in2[134];
    assign G[9] = in[133] & in2[133];
    assign P[9] = in[133] ^ in2[133];
    assign G[10] = in[132] & in2[132];
    assign P[10] = in[132] ^ in2[132];
    assign G[11] = in[131] & in2[131];
    assign P[11] = in[131] ^ in2[131];
    assign G[12] = in[130] & in2[130];
    assign P[12] = in[130] ^ in2[130];
    assign G[13] = in[129] & in2[129];
    assign P[13] = in[129] ^ in2[129];
    assign G[14] = in[128] & in2[128];
    assign P[14] = in[128] ^ in2[128];
    assign G[15] = in[127] & in2[127];
    assign P[15] = in[127] ^ in2[127];
    assign G[16] = in[126] & in2[126];
    assign P[16] = in[126] ^ in2[126];
    assign G[17] = in[125] & in2[125];
    assign P[17] = in[125] ^ in2[125];
    assign G[18] = in[124] & in2[124];
    assign P[18] = in[124] ^ in2[124];
    assign G[19] = in[123] & in2[123];
    assign P[19] = in[123] ^ in2[123];
    assign G[20] = in[122] & in2[122];
    assign P[20] = in[122] ^ in2[122];
    assign G[21] = in[121] & in2[121];
    assign P[21] = in[121] ^ in2[121];
    assign G[22] = in[120] & in2[120];
    assign P[22] = in[120] ^ in2[120];
    assign G[23] = in[119] & in2[119];
    assign P[23] = in[119] ^ in2[119];
    assign G[24] = in[118] & in2[118];
    assign P[24] = in[118] ^ in2[118];
    assign G[25] = in[117] & in2[117];
    assign P[25] = in[117] ^ in2[117];
    assign G[26] = in[116] & in2[116];
    assign P[26] = in[116] ^ in2[116];
    assign G[27] = in[115] & in2[115];
    assign P[27] = in[115] ^ in2[115];
    assign G[28] = in[114] & in2[114];
    assign P[28] = in[114] ^ in2[114];
    assign G[29] = in[113] & in2[113];
    assign P[29] = in[113] ^ in2[113];
    assign G[30] = in[112] & in2[112];
    assign P[30] = in[112] ^ in2[112];
    assign G[31] = in[111] & in2[111];
    assign P[31] = in[111] ^ in2[111];
    assign G[32] = in[110] & in2[110];
    assign P[32] = in[110] ^ in2[110];
    assign G[33] = in[109] & in2[109];
    assign P[33] = in[109] ^ in2[109];
    assign G[34] = in[108] & in2[108];
    assign P[34] = in[108] ^ in2[108];
    assign G[35] = in[107] & in2[107];
    assign P[35] = in[107] ^ in2[107];
    assign G[36] = in[106] & in2[106];
    assign P[36] = in[106] ^ in2[106];
    assign G[37] = in[105] & in2[105];
    assign P[37] = in[105] ^ in2[105];
    assign G[38] = in[104] & in2[104];
    assign P[38] = in[104] ^ in2[104];
    assign G[39] = in[103] & in2[103];
    assign P[39] = in[103] ^ in2[103];
    assign G[40] = in[102] & in2[102];
    assign P[40] = in[102] ^ in2[102];
    assign G[41] = in[101] & in2[101];
    assign P[41] = in[101] ^ in2[101];
    assign G[42] = in[100] & in2[100];
    assign P[42] = in[100] ^ in2[100];
    assign G[43] = in[99] & in2[99];
    assign P[43] = in[99] ^ in2[99];
    assign G[44] = in[98] & in2[98];
    assign P[44] = in[98] ^ in2[98];
    assign G[45] = in[97] & in2[97];
    assign P[45] = in[97] ^ in2[97];
    assign G[46] = in[96] & in2[96];
    assign P[46] = in[96] ^ in2[96];
    assign G[47] = in[95] & in2[95];
    assign P[47] = in[95] ^ in2[95];
    assign G[48] = in[94] & in2[94];
    assign P[48] = in[94] ^ in2[94];
    assign G[49] = in[93] & in2[93];
    assign P[49] = in[93] ^ in2[93];
    assign G[50] = in[92] & in2[92];
    assign P[50] = in[92] ^ in2[92];
    assign G[51] = in[91] & in2[91];
    assign P[51] = in[91] ^ in2[91];
    assign G[52] = in[90] & in2[90];
    assign P[52] = in[90] ^ in2[90];
    assign G[53] = in[89] & in2[89];
    assign P[53] = in[89] ^ in2[89];
    assign G[54] = in[88] & in2[88];
    assign P[54] = in[88] ^ in2[88];
    assign G[55] = in[87] & in2[87];
    assign P[55] = in[87] ^ in2[87];
    assign G[56] = in[86] & in2[86];
    assign P[56] = in[86] ^ in2[86];
    assign G[57] = in[85] & in2[85];
    assign P[57] = in[85] ^ in2[85];
    assign G[58] = in[84] & in2[84];
    assign P[58] = in[84] ^ in2[84];
    assign G[59] = in[83] & in2[83];
    assign P[59] = in[83] ^ in2[83];
    assign G[60] = in[82] & in2[82];
    assign P[60] = in[82] ^ in2[82];
    assign G[61] = in[81] & in2[81];
    assign P[61] = in[81] ^ in2[81];
    assign G[62] = in[80] & in2[80];
    assign P[62] = in[80] ^ in2[80];
    assign G[63] = in[79] & in2[79];
    assign P[63] = in[79] ^ in2[79];
    assign G[64] = in[78] & in2[78];
    assign P[64] = in[78] ^ in2[78];
    assign G[65] = in[77] & in2[77];
    assign P[65] = in[77] ^ in2[77];
    assign G[66] = in[76] & in2[76];
    assign P[66] = in[76] ^ in2[76];
    assign G[67] = in[75] & in2[75];
    assign P[67] = in[75] ^ in2[75];
    assign G[68] = in[74] & in2[74];
    assign P[68] = in[74] ^ in2[74];
    assign G[69] = in[73] & in2[73];
    assign P[69] = in[73] ^ in2[73];
    assign G[70] = in[72] & in2[72];
    assign P[70] = in[72] ^ in2[72];
    assign G[71] = in[71] & in2[71];
    assign P[71] = in[71] ^ in2[71];
    assign G[72] = in[70] & in2[70];
    assign P[72] = in[70] ^ in2[70];
    assign G[73] = in[69] & in2[69];
    assign P[73] = in[69] ^ in2[69];
    assign G[74] = in[68] & in2[68];
    assign P[74] = in[68] ^ in2[68];
    assign G[75] = in[67] & in2[67];
    assign P[75] = in[67] ^ in2[67];
    assign G[76] = in[66] & in2[66];
    assign P[76] = in[66] ^ in2[66];
    assign G[77] = in[65] & in2[65];
    assign P[77] = in[65] ^ in2[65];
    assign G[78] = in[64] & in2[64];
    assign P[78] = in[64] ^ in2[64];
    assign G[79] = in[63] & in2[63];
    assign P[79] = in[63] ^ in2[63];
    assign G[80] = in[62] & in2[62];
    assign P[80] = in[62] ^ in2[62];
    assign G[81] = in[61] & in2[61];
    assign P[81] = in[61] ^ in2[61];
    assign G[82] = in[60] & in2[60];
    assign P[82] = in[60] ^ in2[60];
    assign G[83] = in[59] & in2[59];
    assign P[83] = in[59] ^ in2[59];
    assign G[84] = in[58] & in2[58];
    assign P[84] = in[58] ^ in2[58];
    assign G[85] = in[57] & in2[57];
    assign P[85] = in[57] ^ in2[57];
    assign G[86] = in[56] & in2[56];
    assign P[86] = in[56] ^ in2[56];
    assign G[87] = in[55] & in2[55];
    assign P[87] = in[55] ^ in2[55];
    assign G[88] = in[54] & in2[54];
    assign P[88] = in[54] ^ in2[54];
    assign G[89] = in[53] & in2[53];
    assign P[89] = in[53] ^ in2[53];
    assign G[90] = in[52] & in2[52];
    assign P[90] = in[52] ^ in2[52];
    assign G[91] = in[51] & in2[51];
    assign P[91] = in[51] ^ in2[51];
    assign G[92] = in[50] & in2[50];
    assign P[92] = in[50] ^ in2[50];
    assign G[93] = in[49] & in2[49];
    assign P[93] = in[49] ^ in2[49];
    assign G[94] = in[48] & in2[48];
    assign P[94] = in[48] ^ in2[48];
    assign G[95] = in[47] & in2[47];
    assign P[95] = in[47] ^ in2[47];
    assign G[96] = in[46] & in2[46];
    assign P[96] = in[46] ^ in2[46];
    assign G[97] = in[45] & in2[45];
    assign P[97] = in[45] ^ in2[45];
    assign G[98] = in[44] & in2[44];
    assign P[98] = in[44] ^ in2[44];
    assign G[99] = in[43] & in2[43];
    assign P[99] = in[43] ^ in2[43];
    assign G[100] = in[42] & in2[42];
    assign P[100] = in[42] ^ in2[42];
    assign G[101] = in[41] & in2[41];
    assign P[101] = in[41] ^ in2[41];
    assign G[102] = in[40] & in2[40];
    assign P[102] = in[40] ^ in2[40];
    assign G[103] = in[39] & in2[39];
    assign P[103] = in[39] ^ in2[39];
    assign G[104] = in[38] & in2[38];
    assign P[104] = in[38] ^ in2[38];
    assign G[105] = in[37] & in2[37];
    assign P[105] = in[37] ^ in2[37];
    assign G[106] = in[36] & in2[36];
    assign P[106] = in[36] ^ in2[36];
    assign G[107] = in[35] & in2[35];
    assign P[107] = in[35] ^ in2[35];
    assign G[108] = in[34] & in2[34];
    assign P[108] = in[34] ^ in2[34];
    assign G[109] = in[33] & in2[33];
    assign P[109] = in[33] ^ in2[33];
    assign G[110] = in[32] & in2[32];
    assign P[110] = in[32] ^ in2[32];
    assign G[111] = in[31] & in2[31];
    assign P[111] = in[31] ^ in2[31];
    assign G[112] = in[30] & in2[30];
    assign P[112] = in[30] ^ in2[30];
    assign G[113] = in[29] & in2[29];
    assign P[113] = in[29] ^ in2[29];
    assign G[114] = in[28] & in2[28];
    assign P[114] = in[28] ^ in2[28];
    assign G[115] = in[27] & in2[27];
    assign P[115] = in[27] ^ in2[27];
    assign G[116] = in[26] & in2[26];
    assign P[116] = in[26] ^ in2[26];
    assign G[117] = in[25] & in2[25];
    assign P[117] = in[25] ^ in2[25];
    assign G[118] = in[24] & in2[24];
    assign P[118] = in[24] ^ in2[24];
    assign G[119] = in[23] & in2[23];
    assign P[119] = in[23] ^ in2[23];
    assign G[120] = in[22] & in2[22];
    assign P[120] = in[22] ^ in2[22];
    assign G[121] = in[21] & in2[21];
    assign P[121] = in[21] ^ in2[21];
    assign G[122] = in[20] & in2[20];
    assign P[122] = in[20] ^ in2[20];
    assign G[123] = in[19] & in2[19];
    assign P[123] = in[19] ^ in2[19];
    assign G[124] = in[18] & in2[18];
    assign P[124] = in[18] ^ in2[18];
    assign G[125] = in[17] & in2[17];
    assign P[125] = in[17] ^ in2[17];
    assign G[126] = in[16] & in2[16];
    assign P[126] = in[16] ^ in2[16];
    assign G[127] = in[15] & in2[15];
    assign P[127] = in[15] ^ in2[15];
    assign G[128] = in[14] & in2[14];
    assign P[128] = in[14] ^ in2[14];
    assign G[129] = in[13] & in2[13];
    assign P[129] = in[13] ^ in2[13];
    assign G[130] = in[12] & in2[12];
    assign P[130] = in[12] ^ in2[12];
    assign G[131] = in[11] & in2[11];
    assign P[131] = in[11] ^ in2[11];
    assign G[132] = in[10] & in2[10];
    assign P[132] = in[10] ^ in2[10];
    assign G[133] = in[9] & in2[9];
    assign P[133] = in[9] ^ in2[9];
    assign G[134] = in[8] & in2[8];
    assign P[134] = in[8] ^ in2[8];
    assign G[135] = in[7] & in2[7];
    assign P[135] = in[7] ^ in2[7];
    assign G[136] = in[6] & in2[6];
    assign P[136] = in[6] ^ in2[6];
    assign G[137] = in[5] & in2[5];
    assign P[137] = in[5] ^ in2[5];
    assign G[138] = in[4] & in2[4];
    assign P[138] = in[4] ^ in2[4];
    assign G[139] = in[3] & in2[3];
    assign P[139] = in[3] ^ in2[3];
    assign G[140] = in[2] & in2[2];
    assign P[140] = in[2] ^ in2[2];
    assign G[141] = in[1] & in2[1];
    assign P[141] = in[1] ^ in2[1];
    assign G[142] = in[0] & in2[0];
    assign P[142] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign C[142] = G[141] | (P[141] & C[141]);
    assign cout = G[142] | (P[142] & C[142]);
    assign sum = P ^ C;
endmodule

module CLA142(output [141:0] sum, output cout, input [141:0] in1, input [141:0] in2;

    wire[141:0] G;
    wire[141:0] C;
    wire[141:0] P;

    assign G[0] = in[141] & in2[141];
    assign P[0] = in[141] ^ in2[141];
    assign G[1] = in[140] & in2[140];
    assign P[1] = in[140] ^ in2[140];
    assign G[2] = in[139] & in2[139];
    assign P[2] = in[139] ^ in2[139];
    assign G[3] = in[138] & in2[138];
    assign P[3] = in[138] ^ in2[138];
    assign G[4] = in[137] & in2[137];
    assign P[4] = in[137] ^ in2[137];
    assign G[5] = in[136] & in2[136];
    assign P[5] = in[136] ^ in2[136];
    assign G[6] = in[135] & in2[135];
    assign P[6] = in[135] ^ in2[135];
    assign G[7] = in[134] & in2[134];
    assign P[7] = in[134] ^ in2[134];
    assign G[8] = in[133] & in2[133];
    assign P[8] = in[133] ^ in2[133];
    assign G[9] = in[132] & in2[132];
    assign P[9] = in[132] ^ in2[132];
    assign G[10] = in[131] & in2[131];
    assign P[10] = in[131] ^ in2[131];
    assign G[11] = in[130] & in2[130];
    assign P[11] = in[130] ^ in2[130];
    assign G[12] = in[129] & in2[129];
    assign P[12] = in[129] ^ in2[129];
    assign G[13] = in[128] & in2[128];
    assign P[13] = in[128] ^ in2[128];
    assign G[14] = in[127] & in2[127];
    assign P[14] = in[127] ^ in2[127];
    assign G[15] = in[126] & in2[126];
    assign P[15] = in[126] ^ in2[126];
    assign G[16] = in[125] & in2[125];
    assign P[16] = in[125] ^ in2[125];
    assign G[17] = in[124] & in2[124];
    assign P[17] = in[124] ^ in2[124];
    assign G[18] = in[123] & in2[123];
    assign P[18] = in[123] ^ in2[123];
    assign G[19] = in[122] & in2[122];
    assign P[19] = in[122] ^ in2[122];
    assign G[20] = in[121] & in2[121];
    assign P[20] = in[121] ^ in2[121];
    assign G[21] = in[120] & in2[120];
    assign P[21] = in[120] ^ in2[120];
    assign G[22] = in[119] & in2[119];
    assign P[22] = in[119] ^ in2[119];
    assign G[23] = in[118] & in2[118];
    assign P[23] = in[118] ^ in2[118];
    assign G[24] = in[117] & in2[117];
    assign P[24] = in[117] ^ in2[117];
    assign G[25] = in[116] & in2[116];
    assign P[25] = in[116] ^ in2[116];
    assign G[26] = in[115] & in2[115];
    assign P[26] = in[115] ^ in2[115];
    assign G[27] = in[114] & in2[114];
    assign P[27] = in[114] ^ in2[114];
    assign G[28] = in[113] & in2[113];
    assign P[28] = in[113] ^ in2[113];
    assign G[29] = in[112] & in2[112];
    assign P[29] = in[112] ^ in2[112];
    assign G[30] = in[111] & in2[111];
    assign P[30] = in[111] ^ in2[111];
    assign G[31] = in[110] & in2[110];
    assign P[31] = in[110] ^ in2[110];
    assign G[32] = in[109] & in2[109];
    assign P[32] = in[109] ^ in2[109];
    assign G[33] = in[108] & in2[108];
    assign P[33] = in[108] ^ in2[108];
    assign G[34] = in[107] & in2[107];
    assign P[34] = in[107] ^ in2[107];
    assign G[35] = in[106] & in2[106];
    assign P[35] = in[106] ^ in2[106];
    assign G[36] = in[105] & in2[105];
    assign P[36] = in[105] ^ in2[105];
    assign G[37] = in[104] & in2[104];
    assign P[37] = in[104] ^ in2[104];
    assign G[38] = in[103] & in2[103];
    assign P[38] = in[103] ^ in2[103];
    assign G[39] = in[102] & in2[102];
    assign P[39] = in[102] ^ in2[102];
    assign G[40] = in[101] & in2[101];
    assign P[40] = in[101] ^ in2[101];
    assign G[41] = in[100] & in2[100];
    assign P[41] = in[100] ^ in2[100];
    assign G[42] = in[99] & in2[99];
    assign P[42] = in[99] ^ in2[99];
    assign G[43] = in[98] & in2[98];
    assign P[43] = in[98] ^ in2[98];
    assign G[44] = in[97] & in2[97];
    assign P[44] = in[97] ^ in2[97];
    assign G[45] = in[96] & in2[96];
    assign P[45] = in[96] ^ in2[96];
    assign G[46] = in[95] & in2[95];
    assign P[46] = in[95] ^ in2[95];
    assign G[47] = in[94] & in2[94];
    assign P[47] = in[94] ^ in2[94];
    assign G[48] = in[93] & in2[93];
    assign P[48] = in[93] ^ in2[93];
    assign G[49] = in[92] & in2[92];
    assign P[49] = in[92] ^ in2[92];
    assign G[50] = in[91] & in2[91];
    assign P[50] = in[91] ^ in2[91];
    assign G[51] = in[90] & in2[90];
    assign P[51] = in[90] ^ in2[90];
    assign G[52] = in[89] & in2[89];
    assign P[52] = in[89] ^ in2[89];
    assign G[53] = in[88] & in2[88];
    assign P[53] = in[88] ^ in2[88];
    assign G[54] = in[87] & in2[87];
    assign P[54] = in[87] ^ in2[87];
    assign G[55] = in[86] & in2[86];
    assign P[55] = in[86] ^ in2[86];
    assign G[56] = in[85] & in2[85];
    assign P[56] = in[85] ^ in2[85];
    assign G[57] = in[84] & in2[84];
    assign P[57] = in[84] ^ in2[84];
    assign G[58] = in[83] & in2[83];
    assign P[58] = in[83] ^ in2[83];
    assign G[59] = in[82] & in2[82];
    assign P[59] = in[82] ^ in2[82];
    assign G[60] = in[81] & in2[81];
    assign P[60] = in[81] ^ in2[81];
    assign G[61] = in[80] & in2[80];
    assign P[61] = in[80] ^ in2[80];
    assign G[62] = in[79] & in2[79];
    assign P[62] = in[79] ^ in2[79];
    assign G[63] = in[78] & in2[78];
    assign P[63] = in[78] ^ in2[78];
    assign G[64] = in[77] & in2[77];
    assign P[64] = in[77] ^ in2[77];
    assign G[65] = in[76] & in2[76];
    assign P[65] = in[76] ^ in2[76];
    assign G[66] = in[75] & in2[75];
    assign P[66] = in[75] ^ in2[75];
    assign G[67] = in[74] & in2[74];
    assign P[67] = in[74] ^ in2[74];
    assign G[68] = in[73] & in2[73];
    assign P[68] = in[73] ^ in2[73];
    assign G[69] = in[72] & in2[72];
    assign P[69] = in[72] ^ in2[72];
    assign G[70] = in[71] & in2[71];
    assign P[70] = in[71] ^ in2[71];
    assign G[71] = in[70] & in2[70];
    assign P[71] = in[70] ^ in2[70];
    assign G[72] = in[69] & in2[69];
    assign P[72] = in[69] ^ in2[69];
    assign G[73] = in[68] & in2[68];
    assign P[73] = in[68] ^ in2[68];
    assign G[74] = in[67] & in2[67];
    assign P[74] = in[67] ^ in2[67];
    assign G[75] = in[66] & in2[66];
    assign P[75] = in[66] ^ in2[66];
    assign G[76] = in[65] & in2[65];
    assign P[76] = in[65] ^ in2[65];
    assign G[77] = in[64] & in2[64];
    assign P[77] = in[64] ^ in2[64];
    assign G[78] = in[63] & in2[63];
    assign P[78] = in[63] ^ in2[63];
    assign G[79] = in[62] & in2[62];
    assign P[79] = in[62] ^ in2[62];
    assign G[80] = in[61] & in2[61];
    assign P[80] = in[61] ^ in2[61];
    assign G[81] = in[60] & in2[60];
    assign P[81] = in[60] ^ in2[60];
    assign G[82] = in[59] & in2[59];
    assign P[82] = in[59] ^ in2[59];
    assign G[83] = in[58] & in2[58];
    assign P[83] = in[58] ^ in2[58];
    assign G[84] = in[57] & in2[57];
    assign P[84] = in[57] ^ in2[57];
    assign G[85] = in[56] & in2[56];
    assign P[85] = in[56] ^ in2[56];
    assign G[86] = in[55] & in2[55];
    assign P[86] = in[55] ^ in2[55];
    assign G[87] = in[54] & in2[54];
    assign P[87] = in[54] ^ in2[54];
    assign G[88] = in[53] & in2[53];
    assign P[88] = in[53] ^ in2[53];
    assign G[89] = in[52] & in2[52];
    assign P[89] = in[52] ^ in2[52];
    assign G[90] = in[51] & in2[51];
    assign P[90] = in[51] ^ in2[51];
    assign G[91] = in[50] & in2[50];
    assign P[91] = in[50] ^ in2[50];
    assign G[92] = in[49] & in2[49];
    assign P[92] = in[49] ^ in2[49];
    assign G[93] = in[48] & in2[48];
    assign P[93] = in[48] ^ in2[48];
    assign G[94] = in[47] & in2[47];
    assign P[94] = in[47] ^ in2[47];
    assign G[95] = in[46] & in2[46];
    assign P[95] = in[46] ^ in2[46];
    assign G[96] = in[45] & in2[45];
    assign P[96] = in[45] ^ in2[45];
    assign G[97] = in[44] & in2[44];
    assign P[97] = in[44] ^ in2[44];
    assign G[98] = in[43] & in2[43];
    assign P[98] = in[43] ^ in2[43];
    assign G[99] = in[42] & in2[42];
    assign P[99] = in[42] ^ in2[42];
    assign G[100] = in[41] & in2[41];
    assign P[100] = in[41] ^ in2[41];
    assign G[101] = in[40] & in2[40];
    assign P[101] = in[40] ^ in2[40];
    assign G[102] = in[39] & in2[39];
    assign P[102] = in[39] ^ in2[39];
    assign G[103] = in[38] & in2[38];
    assign P[103] = in[38] ^ in2[38];
    assign G[104] = in[37] & in2[37];
    assign P[104] = in[37] ^ in2[37];
    assign G[105] = in[36] & in2[36];
    assign P[105] = in[36] ^ in2[36];
    assign G[106] = in[35] & in2[35];
    assign P[106] = in[35] ^ in2[35];
    assign G[107] = in[34] & in2[34];
    assign P[107] = in[34] ^ in2[34];
    assign G[108] = in[33] & in2[33];
    assign P[108] = in[33] ^ in2[33];
    assign G[109] = in[32] & in2[32];
    assign P[109] = in[32] ^ in2[32];
    assign G[110] = in[31] & in2[31];
    assign P[110] = in[31] ^ in2[31];
    assign G[111] = in[30] & in2[30];
    assign P[111] = in[30] ^ in2[30];
    assign G[112] = in[29] & in2[29];
    assign P[112] = in[29] ^ in2[29];
    assign G[113] = in[28] & in2[28];
    assign P[113] = in[28] ^ in2[28];
    assign G[114] = in[27] & in2[27];
    assign P[114] = in[27] ^ in2[27];
    assign G[115] = in[26] & in2[26];
    assign P[115] = in[26] ^ in2[26];
    assign G[116] = in[25] & in2[25];
    assign P[116] = in[25] ^ in2[25];
    assign G[117] = in[24] & in2[24];
    assign P[117] = in[24] ^ in2[24];
    assign G[118] = in[23] & in2[23];
    assign P[118] = in[23] ^ in2[23];
    assign G[119] = in[22] & in2[22];
    assign P[119] = in[22] ^ in2[22];
    assign G[120] = in[21] & in2[21];
    assign P[120] = in[21] ^ in2[21];
    assign G[121] = in[20] & in2[20];
    assign P[121] = in[20] ^ in2[20];
    assign G[122] = in[19] & in2[19];
    assign P[122] = in[19] ^ in2[19];
    assign G[123] = in[18] & in2[18];
    assign P[123] = in[18] ^ in2[18];
    assign G[124] = in[17] & in2[17];
    assign P[124] = in[17] ^ in2[17];
    assign G[125] = in[16] & in2[16];
    assign P[125] = in[16] ^ in2[16];
    assign G[126] = in[15] & in2[15];
    assign P[126] = in[15] ^ in2[15];
    assign G[127] = in[14] & in2[14];
    assign P[127] = in[14] ^ in2[14];
    assign G[128] = in[13] & in2[13];
    assign P[128] = in[13] ^ in2[13];
    assign G[129] = in[12] & in2[12];
    assign P[129] = in[12] ^ in2[12];
    assign G[130] = in[11] & in2[11];
    assign P[130] = in[11] ^ in2[11];
    assign G[131] = in[10] & in2[10];
    assign P[131] = in[10] ^ in2[10];
    assign G[132] = in[9] & in2[9];
    assign P[132] = in[9] ^ in2[9];
    assign G[133] = in[8] & in2[8];
    assign P[133] = in[8] ^ in2[8];
    assign G[134] = in[7] & in2[7];
    assign P[134] = in[7] ^ in2[7];
    assign G[135] = in[6] & in2[6];
    assign P[135] = in[6] ^ in2[6];
    assign G[136] = in[5] & in2[5];
    assign P[136] = in[5] ^ in2[5];
    assign G[137] = in[4] & in2[4];
    assign P[137] = in[4] ^ in2[4];
    assign G[138] = in[3] & in2[3];
    assign P[138] = in[3] ^ in2[3];
    assign G[139] = in[2] & in2[2];
    assign P[139] = in[2] ^ in2[2];
    assign G[140] = in[1] & in2[1];
    assign P[140] = in[1] ^ in2[1];
    assign G[141] = in[0] & in2[0];
    assign P[141] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign C[141] = G[140] | (P[140] & C[140]);
    assign cout = G[141] | (P[141] & C[141]);
    assign sum = P ^ C;
endmodule

module CLA141(output [140:0] sum, output cout, input [140:0] in1, input [140:0] in2;

    wire[140:0] G;
    wire[140:0] C;
    wire[140:0] P;

    assign G[0] = in[140] & in2[140];
    assign P[0] = in[140] ^ in2[140];
    assign G[1] = in[139] & in2[139];
    assign P[1] = in[139] ^ in2[139];
    assign G[2] = in[138] & in2[138];
    assign P[2] = in[138] ^ in2[138];
    assign G[3] = in[137] & in2[137];
    assign P[3] = in[137] ^ in2[137];
    assign G[4] = in[136] & in2[136];
    assign P[4] = in[136] ^ in2[136];
    assign G[5] = in[135] & in2[135];
    assign P[5] = in[135] ^ in2[135];
    assign G[6] = in[134] & in2[134];
    assign P[6] = in[134] ^ in2[134];
    assign G[7] = in[133] & in2[133];
    assign P[7] = in[133] ^ in2[133];
    assign G[8] = in[132] & in2[132];
    assign P[8] = in[132] ^ in2[132];
    assign G[9] = in[131] & in2[131];
    assign P[9] = in[131] ^ in2[131];
    assign G[10] = in[130] & in2[130];
    assign P[10] = in[130] ^ in2[130];
    assign G[11] = in[129] & in2[129];
    assign P[11] = in[129] ^ in2[129];
    assign G[12] = in[128] & in2[128];
    assign P[12] = in[128] ^ in2[128];
    assign G[13] = in[127] & in2[127];
    assign P[13] = in[127] ^ in2[127];
    assign G[14] = in[126] & in2[126];
    assign P[14] = in[126] ^ in2[126];
    assign G[15] = in[125] & in2[125];
    assign P[15] = in[125] ^ in2[125];
    assign G[16] = in[124] & in2[124];
    assign P[16] = in[124] ^ in2[124];
    assign G[17] = in[123] & in2[123];
    assign P[17] = in[123] ^ in2[123];
    assign G[18] = in[122] & in2[122];
    assign P[18] = in[122] ^ in2[122];
    assign G[19] = in[121] & in2[121];
    assign P[19] = in[121] ^ in2[121];
    assign G[20] = in[120] & in2[120];
    assign P[20] = in[120] ^ in2[120];
    assign G[21] = in[119] & in2[119];
    assign P[21] = in[119] ^ in2[119];
    assign G[22] = in[118] & in2[118];
    assign P[22] = in[118] ^ in2[118];
    assign G[23] = in[117] & in2[117];
    assign P[23] = in[117] ^ in2[117];
    assign G[24] = in[116] & in2[116];
    assign P[24] = in[116] ^ in2[116];
    assign G[25] = in[115] & in2[115];
    assign P[25] = in[115] ^ in2[115];
    assign G[26] = in[114] & in2[114];
    assign P[26] = in[114] ^ in2[114];
    assign G[27] = in[113] & in2[113];
    assign P[27] = in[113] ^ in2[113];
    assign G[28] = in[112] & in2[112];
    assign P[28] = in[112] ^ in2[112];
    assign G[29] = in[111] & in2[111];
    assign P[29] = in[111] ^ in2[111];
    assign G[30] = in[110] & in2[110];
    assign P[30] = in[110] ^ in2[110];
    assign G[31] = in[109] & in2[109];
    assign P[31] = in[109] ^ in2[109];
    assign G[32] = in[108] & in2[108];
    assign P[32] = in[108] ^ in2[108];
    assign G[33] = in[107] & in2[107];
    assign P[33] = in[107] ^ in2[107];
    assign G[34] = in[106] & in2[106];
    assign P[34] = in[106] ^ in2[106];
    assign G[35] = in[105] & in2[105];
    assign P[35] = in[105] ^ in2[105];
    assign G[36] = in[104] & in2[104];
    assign P[36] = in[104] ^ in2[104];
    assign G[37] = in[103] & in2[103];
    assign P[37] = in[103] ^ in2[103];
    assign G[38] = in[102] & in2[102];
    assign P[38] = in[102] ^ in2[102];
    assign G[39] = in[101] & in2[101];
    assign P[39] = in[101] ^ in2[101];
    assign G[40] = in[100] & in2[100];
    assign P[40] = in[100] ^ in2[100];
    assign G[41] = in[99] & in2[99];
    assign P[41] = in[99] ^ in2[99];
    assign G[42] = in[98] & in2[98];
    assign P[42] = in[98] ^ in2[98];
    assign G[43] = in[97] & in2[97];
    assign P[43] = in[97] ^ in2[97];
    assign G[44] = in[96] & in2[96];
    assign P[44] = in[96] ^ in2[96];
    assign G[45] = in[95] & in2[95];
    assign P[45] = in[95] ^ in2[95];
    assign G[46] = in[94] & in2[94];
    assign P[46] = in[94] ^ in2[94];
    assign G[47] = in[93] & in2[93];
    assign P[47] = in[93] ^ in2[93];
    assign G[48] = in[92] & in2[92];
    assign P[48] = in[92] ^ in2[92];
    assign G[49] = in[91] & in2[91];
    assign P[49] = in[91] ^ in2[91];
    assign G[50] = in[90] & in2[90];
    assign P[50] = in[90] ^ in2[90];
    assign G[51] = in[89] & in2[89];
    assign P[51] = in[89] ^ in2[89];
    assign G[52] = in[88] & in2[88];
    assign P[52] = in[88] ^ in2[88];
    assign G[53] = in[87] & in2[87];
    assign P[53] = in[87] ^ in2[87];
    assign G[54] = in[86] & in2[86];
    assign P[54] = in[86] ^ in2[86];
    assign G[55] = in[85] & in2[85];
    assign P[55] = in[85] ^ in2[85];
    assign G[56] = in[84] & in2[84];
    assign P[56] = in[84] ^ in2[84];
    assign G[57] = in[83] & in2[83];
    assign P[57] = in[83] ^ in2[83];
    assign G[58] = in[82] & in2[82];
    assign P[58] = in[82] ^ in2[82];
    assign G[59] = in[81] & in2[81];
    assign P[59] = in[81] ^ in2[81];
    assign G[60] = in[80] & in2[80];
    assign P[60] = in[80] ^ in2[80];
    assign G[61] = in[79] & in2[79];
    assign P[61] = in[79] ^ in2[79];
    assign G[62] = in[78] & in2[78];
    assign P[62] = in[78] ^ in2[78];
    assign G[63] = in[77] & in2[77];
    assign P[63] = in[77] ^ in2[77];
    assign G[64] = in[76] & in2[76];
    assign P[64] = in[76] ^ in2[76];
    assign G[65] = in[75] & in2[75];
    assign P[65] = in[75] ^ in2[75];
    assign G[66] = in[74] & in2[74];
    assign P[66] = in[74] ^ in2[74];
    assign G[67] = in[73] & in2[73];
    assign P[67] = in[73] ^ in2[73];
    assign G[68] = in[72] & in2[72];
    assign P[68] = in[72] ^ in2[72];
    assign G[69] = in[71] & in2[71];
    assign P[69] = in[71] ^ in2[71];
    assign G[70] = in[70] & in2[70];
    assign P[70] = in[70] ^ in2[70];
    assign G[71] = in[69] & in2[69];
    assign P[71] = in[69] ^ in2[69];
    assign G[72] = in[68] & in2[68];
    assign P[72] = in[68] ^ in2[68];
    assign G[73] = in[67] & in2[67];
    assign P[73] = in[67] ^ in2[67];
    assign G[74] = in[66] & in2[66];
    assign P[74] = in[66] ^ in2[66];
    assign G[75] = in[65] & in2[65];
    assign P[75] = in[65] ^ in2[65];
    assign G[76] = in[64] & in2[64];
    assign P[76] = in[64] ^ in2[64];
    assign G[77] = in[63] & in2[63];
    assign P[77] = in[63] ^ in2[63];
    assign G[78] = in[62] & in2[62];
    assign P[78] = in[62] ^ in2[62];
    assign G[79] = in[61] & in2[61];
    assign P[79] = in[61] ^ in2[61];
    assign G[80] = in[60] & in2[60];
    assign P[80] = in[60] ^ in2[60];
    assign G[81] = in[59] & in2[59];
    assign P[81] = in[59] ^ in2[59];
    assign G[82] = in[58] & in2[58];
    assign P[82] = in[58] ^ in2[58];
    assign G[83] = in[57] & in2[57];
    assign P[83] = in[57] ^ in2[57];
    assign G[84] = in[56] & in2[56];
    assign P[84] = in[56] ^ in2[56];
    assign G[85] = in[55] & in2[55];
    assign P[85] = in[55] ^ in2[55];
    assign G[86] = in[54] & in2[54];
    assign P[86] = in[54] ^ in2[54];
    assign G[87] = in[53] & in2[53];
    assign P[87] = in[53] ^ in2[53];
    assign G[88] = in[52] & in2[52];
    assign P[88] = in[52] ^ in2[52];
    assign G[89] = in[51] & in2[51];
    assign P[89] = in[51] ^ in2[51];
    assign G[90] = in[50] & in2[50];
    assign P[90] = in[50] ^ in2[50];
    assign G[91] = in[49] & in2[49];
    assign P[91] = in[49] ^ in2[49];
    assign G[92] = in[48] & in2[48];
    assign P[92] = in[48] ^ in2[48];
    assign G[93] = in[47] & in2[47];
    assign P[93] = in[47] ^ in2[47];
    assign G[94] = in[46] & in2[46];
    assign P[94] = in[46] ^ in2[46];
    assign G[95] = in[45] & in2[45];
    assign P[95] = in[45] ^ in2[45];
    assign G[96] = in[44] & in2[44];
    assign P[96] = in[44] ^ in2[44];
    assign G[97] = in[43] & in2[43];
    assign P[97] = in[43] ^ in2[43];
    assign G[98] = in[42] & in2[42];
    assign P[98] = in[42] ^ in2[42];
    assign G[99] = in[41] & in2[41];
    assign P[99] = in[41] ^ in2[41];
    assign G[100] = in[40] & in2[40];
    assign P[100] = in[40] ^ in2[40];
    assign G[101] = in[39] & in2[39];
    assign P[101] = in[39] ^ in2[39];
    assign G[102] = in[38] & in2[38];
    assign P[102] = in[38] ^ in2[38];
    assign G[103] = in[37] & in2[37];
    assign P[103] = in[37] ^ in2[37];
    assign G[104] = in[36] & in2[36];
    assign P[104] = in[36] ^ in2[36];
    assign G[105] = in[35] & in2[35];
    assign P[105] = in[35] ^ in2[35];
    assign G[106] = in[34] & in2[34];
    assign P[106] = in[34] ^ in2[34];
    assign G[107] = in[33] & in2[33];
    assign P[107] = in[33] ^ in2[33];
    assign G[108] = in[32] & in2[32];
    assign P[108] = in[32] ^ in2[32];
    assign G[109] = in[31] & in2[31];
    assign P[109] = in[31] ^ in2[31];
    assign G[110] = in[30] & in2[30];
    assign P[110] = in[30] ^ in2[30];
    assign G[111] = in[29] & in2[29];
    assign P[111] = in[29] ^ in2[29];
    assign G[112] = in[28] & in2[28];
    assign P[112] = in[28] ^ in2[28];
    assign G[113] = in[27] & in2[27];
    assign P[113] = in[27] ^ in2[27];
    assign G[114] = in[26] & in2[26];
    assign P[114] = in[26] ^ in2[26];
    assign G[115] = in[25] & in2[25];
    assign P[115] = in[25] ^ in2[25];
    assign G[116] = in[24] & in2[24];
    assign P[116] = in[24] ^ in2[24];
    assign G[117] = in[23] & in2[23];
    assign P[117] = in[23] ^ in2[23];
    assign G[118] = in[22] & in2[22];
    assign P[118] = in[22] ^ in2[22];
    assign G[119] = in[21] & in2[21];
    assign P[119] = in[21] ^ in2[21];
    assign G[120] = in[20] & in2[20];
    assign P[120] = in[20] ^ in2[20];
    assign G[121] = in[19] & in2[19];
    assign P[121] = in[19] ^ in2[19];
    assign G[122] = in[18] & in2[18];
    assign P[122] = in[18] ^ in2[18];
    assign G[123] = in[17] & in2[17];
    assign P[123] = in[17] ^ in2[17];
    assign G[124] = in[16] & in2[16];
    assign P[124] = in[16] ^ in2[16];
    assign G[125] = in[15] & in2[15];
    assign P[125] = in[15] ^ in2[15];
    assign G[126] = in[14] & in2[14];
    assign P[126] = in[14] ^ in2[14];
    assign G[127] = in[13] & in2[13];
    assign P[127] = in[13] ^ in2[13];
    assign G[128] = in[12] & in2[12];
    assign P[128] = in[12] ^ in2[12];
    assign G[129] = in[11] & in2[11];
    assign P[129] = in[11] ^ in2[11];
    assign G[130] = in[10] & in2[10];
    assign P[130] = in[10] ^ in2[10];
    assign G[131] = in[9] & in2[9];
    assign P[131] = in[9] ^ in2[9];
    assign G[132] = in[8] & in2[8];
    assign P[132] = in[8] ^ in2[8];
    assign G[133] = in[7] & in2[7];
    assign P[133] = in[7] ^ in2[7];
    assign G[134] = in[6] & in2[6];
    assign P[134] = in[6] ^ in2[6];
    assign G[135] = in[5] & in2[5];
    assign P[135] = in[5] ^ in2[5];
    assign G[136] = in[4] & in2[4];
    assign P[136] = in[4] ^ in2[4];
    assign G[137] = in[3] & in2[3];
    assign P[137] = in[3] ^ in2[3];
    assign G[138] = in[2] & in2[2];
    assign P[138] = in[2] ^ in2[2];
    assign G[139] = in[1] & in2[1];
    assign P[139] = in[1] ^ in2[1];
    assign G[140] = in[0] & in2[0];
    assign P[140] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign C[140] = G[139] | (P[139] & C[139]);
    assign cout = G[140] | (P[140] & C[140]);
    assign sum = P ^ C;
endmodule

module CLA140(output [139:0] sum, output cout, input [139:0] in1, input [139:0] in2;

    wire[139:0] G;
    wire[139:0] C;
    wire[139:0] P;

    assign G[0] = in[139] & in2[139];
    assign P[0] = in[139] ^ in2[139];
    assign G[1] = in[138] & in2[138];
    assign P[1] = in[138] ^ in2[138];
    assign G[2] = in[137] & in2[137];
    assign P[2] = in[137] ^ in2[137];
    assign G[3] = in[136] & in2[136];
    assign P[3] = in[136] ^ in2[136];
    assign G[4] = in[135] & in2[135];
    assign P[4] = in[135] ^ in2[135];
    assign G[5] = in[134] & in2[134];
    assign P[5] = in[134] ^ in2[134];
    assign G[6] = in[133] & in2[133];
    assign P[6] = in[133] ^ in2[133];
    assign G[7] = in[132] & in2[132];
    assign P[7] = in[132] ^ in2[132];
    assign G[8] = in[131] & in2[131];
    assign P[8] = in[131] ^ in2[131];
    assign G[9] = in[130] & in2[130];
    assign P[9] = in[130] ^ in2[130];
    assign G[10] = in[129] & in2[129];
    assign P[10] = in[129] ^ in2[129];
    assign G[11] = in[128] & in2[128];
    assign P[11] = in[128] ^ in2[128];
    assign G[12] = in[127] & in2[127];
    assign P[12] = in[127] ^ in2[127];
    assign G[13] = in[126] & in2[126];
    assign P[13] = in[126] ^ in2[126];
    assign G[14] = in[125] & in2[125];
    assign P[14] = in[125] ^ in2[125];
    assign G[15] = in[124] & in2[124];
    assign P[15] = in[124] ^ in2[124];
    assign G[16] = in[123] & in2[123];
    assign P[16] = in[123] ^ in2[123];
    assign G[17] = in[122] & in2[122];
    assign P[17] = in[122] ^ in2[122];
    assign G[18] = in[121] & in2[121];
    assign P[18] = in[121] ^ in2[121];
    assign G[19] = in[120] & in2[120];
    assign P[19] = in[120] ^ in2[120];
    assign G[20] = in[119] & in2[119];
    assign P[20] = in[119] ^ in2[119];
    assign G[21] = in[118] & in2[118];
    assign P[21] = in[118] ^ in2[118];
    assign G[22] = in[117] & in2[117];
    assign P[22] = in[117] ^ in2[117];
    assign G[23] = in[116] & in2[116];
    assign P[23] = in[116] ^ in2[116];
    assign G[24] = in[115] & in2[115];
    assign P[24] = in[115] ^ in2[115];
    assign G[25] = in[114] & in2[114];
    assign P[25] = in[114] ^ in2[114];
    assign G[26] = in[113] & in2[113];
    assign P[26] = in[113] ^ in2[113];
    assign G[27] = in[112] & in2[112];
    assign P[27] = in[112] ^ in2[112];
    assign G[28] = in[111] & in2[111];
    assign P[28] = in[111] ^ in2[111];
    assign G[29] = in[110] & in2[110];
    assign P[29] = in[110] ^ in2[110];
    assign G[30] = in[109] & in2[109];
    assign P[30] = in[109] ^ in2[109];
    assign G[31] = in[108] & in2[108];
    assign P[31] = in[108] ^ in2[108];
    assign G[32] = in[107] & in2[107];
    assign P[32] = in[107] ^ in2[107];
    assign G[33] = in[106] & in2[106];
    assign P[33] = in[106] ^ in2[106];
    assign G[34] = in[105] & in2[105];
    assign P[34] = in[105] ^ in2[105];
    assign G[35] = in[104] & in2[104];
    assign P[35] = in[104] ^ in2[104];
    assign G[36] = in[103] & in2[103];
    assign P[36] = in[103] ^ in2[103];
    assign G[37] = in[102] & in2[102];
    assign P[37] = in[102] ^ in2[102];
    assign G[38] = in[101] & in2[101];
    assign P[38] = in[101] ^ in2[101];
    assign G[39] = in[100] & in2[100];
    assign P[39] = in[100] ^ in2[100];
    assign G[40] = in[99] & in2[99];
    assign P[40] = in[99] ^ in2[99];
    assign G[41] = in[98] & in2[98];
    assign P[41] = in[98] ^ in2[98];
    assign G[42] = in[97] & in2[97];
    assign P[42] = in[97] ^ in2[97];
    assign G[43] = in[96] & in2[96];
    assign P[43] = in[96] ^ in2[96];
    assign G[44] = in[95] & in2[95];
    assign P[44] = in[95] ^ in2[95];
    assign G[45] = in[94] & in2[94];
    assign P[45] = in[94] ^ in2[94];
    assign G[46] = in[93] & in2[93];
    assign P[46] = in[93] ^ in2[93];
    assign G[47] = in[92] & in2[92];
    assign P[47] = in[92] ^ in2[92];
    assign G[48] = in[91] & in2[91];
    assign P[48] = in[91] ^ in2[91];
    assign G[49] = in[90] & in2[90];
    assign P[49] = in[90] ^ in2[90];
    assign G[50] = in[89] & in2[89];
    assign P[50] = in[89] ^ in2[89];
    assign G[51] = in[88] & in2[88];
    assign P[51] = in[88] ^ in2[88];
    assign G[52] = in[87] & in2[87];
    assign P[52] = in[87] ^ in2[87];
    assign G[53] = in[86] & in2[86];
    assign P[53] = in[86] ^ in2[86];
    assign G[54] = in[85] & in2[85];
    assign P[54] = in[85] ^ in2[85];
    assign G[55] = in[84] & in2[84];
    assign P[55] = in[84] ^ in2[84];
    assign G[56] = in[83] & in2[83];
    assign P[56] = in[83] ^ in2[83];
    assign G[57] = in[82] & in2[82];
    assign P[57] = in[82] ^ in2[82];
    assign G[58] = in[81] & in2[81];
    assign P[58] = in[81] ^ in2[81];
    assign G[59] = in[80] & in2[80];
    assign P[59] = in[80] ^ in2[80];
    assign G[60] = in[79] & in2[79];
    assign P[60] = in[79] ^ in2[79];
    assign G[61] = in[78] & in2[78];
    assign P[61] = in[78] ^ in2[78];
    assign G[62] = in[77] & in2[77];
    assign P[62] = in[77] ^ in2[77];
    assign G[63] = in[76] & in2[76];
    assign P[63] = in[76] ^ in2[76];
    assign G[64] = in[75] & in2[75];
    assign P[64] = in[75] ^ in2[75];
    assign G[65] = in[74] & in2[74];
    assign P[65] = in[74] ^ in2[74];
    assign G[66] = in[73] & in2[73];
    assign P[66] = in[73] ^ in2[73];
    assign G[67] = in[72] & in2[72];
    assign P[67] = in[72] ^ in2[72];
    assign G[68] = in[71] & in2[71];
    assign P[68] = in[71] ^ in2[71];
    assign G[69] = in[70] & in2[70];
    assign P[69] = in[70] ^ in2[70];
    assign G[70] = in[69] & in2[69];
    assign P[70] = in[69] ^ in2[69];
    assign G[71] = in[68] & in2[68];
    assign P[71] = in[68] ^ in2[68];
    assign G[72] = in[67] & in2[67];
    assign P[72] = in[67] ^ in2[67];
    assign G[73] = in[66] & in2[66];
    assign P[73] = in[66] ^ in2[66];
    assign G[74] = in[65] & in2[65];
    assign P[74] = in[65] ^ in2[65];
    assign G[75] = in[64] & in2[64];
    assign P[75] = in[64] ^ in2[64];
    assign G[76] = in[63] & in2[63];
    assign P[76] = in[63] ^ in2[63];
    assign G[77] = in[62] & in2[62];
    assign P[77] = in[62] ^ in2[62];
    assign G[78] = in[61] & in2[61];
    assign P[78] = in[61] ^ in2[61];
    assign G[79] = in[60] & in2[60];
    assign P[79] = in[60] ^ in2[60];
    assign G[80] = in[59] & in2[59];
    assign P[80] = in[59] ^ in2[59];
    assign G[81] = in[58] & in2[58];
    assign P[81] = in[58] ^ in2[58];
    assign G[82] = in[57] & in2[57];
    assign P[82] = in[57] ^ in2[57];
    assign G[83] = in[56] & in2[56];
    assign P[83] = in[56] ^ in2[56];
    assign G[84] = in[55] & in2[55];
    assign P[84] = in[55] ^ in2[55];
    assign G[85] = in[54] & in2[54];
    assign P[85] = in[54] ^ in2[54];
    assign G[86] = in[53] & in2[53];
    assign P[86] = in[53] ^ in2[53];
    assign G[87] = in[52] & in2[52];
    assign P[87] = in[52] ^ in2[52];
    assign G[88] = in[51] & in2[51];
    assign P[88] = in[51] ^ in2[51];
    assign G[89] = in[50] & in2[50];
    assign P[89] = in[50] ^ in2[50];
    assign G[90] = in[49] & in2[49];
    assign P[90] = in[49] ^ in2[49];
    assign G[91] = in[48] & in2[48];
    assign P[91] = in[48] ^ in2[48];
    assign G[92] = in[47] & in2[47];
    assign P[92] = in[47] ^ in2[47];
    assign G[93] = in[46] & in2[46];
    assign P[93] = in[46] ^ in2[46];
    assign G[94] = in[45] & in2[45];
    assign P[94] = in[45] ^ in2[45];
    assign G[95] = in[44] & in2[44];
    assign P[95] = in[44] ^ in2[44];
    assign G[96] = in[43] & in2[43];
    assign P[96] = in[43] ^ in2[43];
    assign G[97] = in[42] & in2[42];
    assign P[97] = in[42] ^ in2[42];
    assign G[98] = in[41] & in2[41];
    assign P[98] = in[41] ^ in2[41];
    assign G[99] = in[40] & in2[40];
    assign P[99] = in[40] ^ in2[40];
    assign G[100] = in[39] & in2[39];
    assign P[100] = in[39] ^ in2[39];
    assign G[101] = in[38] & in2[38];
    assign P[101] = in[38] ^ in2[38];
    assign G[102] = in[37] & in2[37];
    assign P[102] = in[37] ^ in2[37];
    assign G[103] = in[36] & in2[36];
    assign P[103] = in[36] ^ in2[36];
    assign G[104] = in[35] & in2[35];
    assign P[104] = in[35] ^ in2[35];
    assign G[105] = in[34] & in2[34];
    assign P[105] = in[34] ^ in2[34];
    assign G[106] = in[33] & in2[33];
    assign P[106] = in[33] ^ in2[33];
    assign G[107] = in[32] & in2[32];
    assign P[107] = in[32] ^ in2[32];
    assign G[108] = in[31] & in2[31];
    assign P[108] = in[31] ^ in2[31];
    assign G[109] = in[30] & in2[30];
    assign P[109] = in[30] ^ in2[30];
    assign G[110] = in[29] & in2[29];
    assign P[110] = in[29] ^ in2[29];
    assign G[111] = in[28] & in2[28];
    assign P[111] = in[28] ^ in2[28];
    assign G[112] = in[27] & in2[27];
    assign P[112] = in[27] ^ in2[27];
    assign G[113] = in[26] & in2[26];
    assign P[113] = in[26] ^ in2[26];
    assign G[114] = in[25] & in2[25];
    assign P[114] = in[25] ^ in2[25];
    assign G[115] = in[24] & in2[24];
    assign P[115] = in[24] ^ in2[24];
    assign G[116] = in[23] & in2[23];
    assign P[116] = in[23] ^ in2[23];
    assign G[117] = in[22] & in2[22];
    assign P[117] = in[22] ^ in2[22];
    assign G[118] = in[21] & in2[21];
    assign P[118] = in[21] ^ in2[21];
    assign G[119] = in[20] & in2[20];
    assign P[119] = in[20] ^ in2[20];
    assign G[120] = in[19] & in2[19];
    assign P[120] = in[19] ^ in2[19];
    assign G[121] = in[18] & in2[18];
    assign P[121] = in[18] ^ in2[18];
    assign G[122] = in[17] & in2[17];
    assign P[122] = in[17] ^ in2[17];
    assign G[123] = in[16] & in2[16];
    assign P[123] = in[16] ^ in2[16];
    assign G[124] = in[15] & in2[15];
    assign P[124] = in[15] ^ in2[15];
    assign G[125] = in[14] & in2[14];
    assign P[125] = in[14] ^ in2[14];
    assign G[126] = in[13] & in2[13];
    assign P[126] = in[13] ^ in2[13];
    assign G[127] = in[12] & in2[12];
    assign P[127] = in[12] ^ in2[12];
    assign G[128] = in[11] & in2[11];
    assign P[128] = in[11] ^ in2[11];
    assign G[129] = in[10] & in2[10];
    assign P[129] = in[10] ^ in2[10];
    assign G[130] = in[9] & in2[9];
    assign P[130] = in[9] ^ in2[9];
    assign G[131] = in[8] & in2[8];
    assign P[131] = in[8] ^ in2[8];
    assign G[132] = in[7] & in2[7];
    assign P[132] = in[7] ^ in2[7];
    assign G[133] = in[6] & in2[6];
    assign P[133] = in[6] ^ in2[6];
    assign G[134] = in[5] & in2[5];
    assign P[134] = in[5] ^ in2[5];
    assign G[135] = in[4] & in2[4];
    assign P[135] = in[4] ^ in2[4];
    assign G[136] = in[3] & in2[3];
    assign P[136] = in[3] ^ in2[3];
    assign G[137] = in[2] & in2[2];
    assign P[137] = in[2] ^ in2[2];
    assign G[138] = in[1] & in2[1];
    assign P[138] = in[1] ^ in2[1];
    assign G[139] = in[0] & in2[0];
    assign P[139] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign C[139] = G[138] | (P[138] & C[138]);
    assign cout = G[139] | (P[139] & C[139]);
    assign sum = P ^ C;
endmodule

module CLA139(output [138:0] sum, output cout, input [138:0] in1, input [138:0] in2;

    wire[138:0] G;
    wire[138:0] C;
    wire[138:0] P;

    assign G[0] = in[138] & in2[138];
    assign P[0] = in[138] ^ in2[138];
    assign G[1] = in[137] & in2[137];
    assign P[1] = in[137] ^ in2[137];
    assign G[2] = in[136] & in2[136];
    assign P[2] = in[136] ^ in2[136];
    assign G[3] = in[135] & in2[135];
    assign P[3] = in[135] ^ in2[135];
    assign G[4] = in[134] & in2[134];
    assign P[4] = in[134] ^ in2[134];
    assign G[5] = in[133] & in2[133];
    assign P[5] = in[133] ^ in2[133];
    assign G[6] = in[132] & in2[132];
    assign P[6] = in[132] ^ in2[132];
    assign G[7] = in[131] & in2[131];
    assign P[7] = in[131] ^ in2[131];
    assign G[8] = in[130] & in2[130];
    assign P[8] = in[130] ^ in2[130];
    assign G[9] = in[129] & in2[129];
    assign P[9] = in[129] ^ in2[129];
    assign G[10] = in[128] & in2[128];
    assign P[10] = in[128] ^ in2[128];
    assign G[11] = in[127] & in2[127];
    assign P[11] = in[127] ^ in2[127];
    assign G[12] = in[126] & in2[126];
    assign P[12] = in[126] ^ in2[126];
    assign G[13] = in[125] & in2[125];
    assign P[13] = in[125] ^ in2[125];
    assign G[14] = in[124] & in2[124];
    assign P[14] = in[124] ^ in2[124];
    assign G[15] = in[123] & in2[123];
    assign P[15] = in[123] ^ in2[123];
    assign G[16] = in[122] & in2[122];
    assign P[16] = in[122] ^ in2[122];
    assign G[17] = in[121] & in2[121];
    assign P[17] = in[121] ^ in2[121];
    assign G[18] = in[120] & in2[120];
    assign P[18] = in[120] ^ in2[120];
    assign G[19] = in[119] & in2[119];
    assign P[19] = in[119] ^ in2[119];
    assign G[20] = in[118] & in2[118];
    assign P[20] = in[118] ^ in2[118];
    assign G[21] = in[117] & in2[117];
    assign P[21] = in[117] ^ in2[117];
    assign G[22] = in[116] & in2[116];
    assign P[22] = in[116] ^ in2[116];
    assign G[23] = in[115] & in2[115];
    assign P[23] = in[115] ^ in2[115];
    assign G[24] = in[114] & in2[114];
    assign P[24] = in[114] ^ in2[114];
    assign G[25] = in[113] & in2[113];
    assign P[25] = in[113] ^ in2[113];
    assign G[26] = in[112] & in2[112];
    assign P[26] = in[112] ^ in2[112];
    assign G[27] = in[111] & in2[111];
    assign P[27] = in[111] ^ in2[111];
    assign G[28] = in[110] & in2[110];
    assign P[28] = in[110] ^ in2[110];
    assign G[29] = in[109] & in2[109];
    assign P[29] = in[109] ^ in2[109];
    assign G[30] = in[108] & in2[108];
    assign P[30] = in[108] ^ in2[108];
    assign G[31] = in[107] & in2[107];
    assign P[31] = in[107] ^ in2[107];
    assign G[32] = in[106] & in2[106];
    assign P[32] = in[106] ^ in2[106];
    assign G[33] = in[105] & in2[105];
    assign P[33] = in[105] ^ in2[105];
    assign G[34] = in[104] & in2[104];
    assign P[34] = in[104] ^ in2[104];
    assign G[35] = in[103] & in2[103];
    assign P[35] = in[103] ^ in2[103];
    assign G[36] = in[102] & in2[102];
    assign P[36] = in[102] ^ in2[102];
    assign G[37] = in[101] & in2[101];
    assign P[37] = in[101] ^ in2[101];
    assign G[38] = in[100] & in2[100];
    assign P[38] = in[100] ^ in2[100];
    assign G[39] = in[99] & in2[99];
    assign P[39] = in[99] ^ in2[99];
    assign G[40] = in[98] & in2[98];
    assign P[40] = in[98] ^ in2[98];
    assign G[41] = in[97] & in2[97];
    assign P[41] = in[97] ^ in2[97];
    assign G[42] = in[96] & in2[96];
    assign P[42] = in[96] ^ in2[96];
    assign G[43] = in[95] & in2[95];
    assign P[43] = in[95] ^ in2[95];
    assign G[44] = in[94] & in2[94];
    assign P[44] = in[94] ^ in2[94];
    assign G[45] = in[93] & in2[93];
    assign P[45] = in[93] ^ in2[93];
    assign G[46] = in[92] & in2[92];
    assign P[46] = in[92] ^ in2[92];
    assign G[47] = in[91] & in2[91];
    assign P[47] = in[91] ^ in2[91];
    assign G[48] = in[90] & in2[90];
    assign P[48] = in[90] ^ in2[90];
    assign G[49] = in[89] & in2[89];
    assign P[49] = in[89] ^ in2[89];
    assign G[50] = in[88] & in2[88];
    assign P[50] = in[88] ^ in2[88];
    assign G[51] = in[87] & in2[87];
    assign P[51] = in[87] ^ in2[87];
    assign G[52] = in[86] & in2[86];
    assign P[52] = in[86] ^ in2[86];
    assign G[53] = in[85] & in2[85];
    assign P[53] = in[85] ^ in2[85];
    assign G[54] = in[84] & in2[84];
    assign P[54] = in[84] ^ in2[84];
    assign G[55] = in[83] & in2[83];
    assign P[55] = in[83] ^ in2[83];
    assign G[56] = in[82] & in2[82];
    assign P[56] = in[82] ^ in2[82];
    assign G[57] = in[81] & in2[81];
    assign P[57] = in[81] ^ in2[81];
    assign G[58] = in[80] & in2[80];
    assign P[58] = in[80] ^ in2[80];
    assign G[59] = in[79] & in2[79];
    assign P[59] = in[79] ^ in2[79];
    assign G[60] = in[78] & in2[78];
    assign P[60] = in[78] ^ in2[78];
    assign G[61] = in[77] & in2[77];
    assign P[61] = in[77] ^ in2[77];
    assign G[62] = in[76] & in2[76];
    assign P[62] = in[76] ^ in2[76];
    assign G[63] = in[75] & in2[75];
    assign P[63] = in[75] ^ in2[75];
    assign G[64] = in[74] & in2[74];
    assign P[64] = in[74] ^ in2[74];
    assign G[65] = in[73] & in2[73];
    assign P[65] = in[73] ^ in2[73];
    assign G[66] = in[72] & in2[72];
    assign P[66] = in[72] ^ in2[72];
    assign G[67] = in[71] & in2[71];
    assign P[67] = in[71] ^ in2[71];
    assign G[68] = in[70] & in2[70];
    assign P[68] = in[70] ^ in2[70];
    assign G[69] = in[69] & in2[69];
    assign P[69] = in[69] ^ in2[69];
    assign G[70] = in[68] & in2[68];
    assign P[70] = in[68] ^ in2[68];
    assign G[71] = in[67] & in2[67];
    assign P[71] = in[67] ^ in2[67];
    assign G[72] = in[66] & in2[66];
    assign P[72] = in[66] ^ in2[66];
    assign G[73] = in[65] & in2[65];
    assign P[73] = in[65] ^ in2[65];
    assign G[74] = in[64] & in2[64];
    assign P[74] = in[64] ^ in2[64];
    assign G[75] = in[63] & in2[63];
    assign P[75] = in[63] ^ in2[63];
    assign G[76] = in[62] & in2[62];
    assign P[76] = in[62] ^ in2[62];
    assign G[77] = in[61] & in2[61];
    assign P[77] = in[61] ^ in2[61];
    assign G[78] = in[60] & in2[60];
    assign P[78] = in[60] ^ in2[60];
    assign G[79] = in[59] & in2[59];
    assign P[79] = in[59] ^ in2[59];
    assign G[80] = in[58] & in2[58];
    assign P[80] = in[58] ^ in2[58];
    assign G[81] = in[57] & in2[57];
    assign P[81] = in[57] ^ in2[57];
    assign G[82] = in[56] & in2[56];
    assign P[82] = in[56] ^ in2[56];
    assign G[83] = in[55] & in2[55];
    assign P[83] = in[55] ^ in2[55];
    assign G[84] = in[54] & in2[54];
    assign P[84] = in[54] ^ in2[54];
    assign G[85] = in[53] & in2[53];
    assign P[85] = in[53] ^ in2[53];
    assign G[86] = in[52] & in2[52];
    assign P[86] = in[52] ^ in2[52];
    assign G[87] = in[51] & in2[51];
    assign P[87] = in[51] ^ in2[51];
    assign G[88] = in[50] & in2[50];
    assign P[88] = in[50] ^ in2[50];
    assign G[89] = in[49] & in2[49];
    assign P[89] = in[49] ^ in2[49];
    assign G[90] = in[48] & in2[48];
    assign P[90] = in[48] ^ in2[48];
    assign G[91] = in[47] & in2[47];
    assign P[91] = in[47] ^ in2[47];
    assign G[92] = in[46] & in2[46];
    assign P[92] = in[46] ^ in2[46];
    assign G[93] = in[45] & in2[45];
    assign P[93] = in[45] ^ in2[45];
    assign G[94] = in[44] & in2[44];
    assign P[94] = in[44] ^ in2[44];
    assign G[95] = in[43] & in2[43];
    assign P[95] = in[43] ^ in2[43];
    assign G[96] = in[42] & in2[42];
    assign P[96] = in[42] ^ in2[42];
    assign G[97] = in[41] & in2[41];
    assign P[97] = in[41] ^ in2[41];
    assign G[98] = in[40] & in2[40];
    assign P[98] = in[40] ^ in2[40];
    assign G[99] = in[39] & in2[39];
    assign P[99] = in[39] ^ in2[39];
    assign G[100] = in[38] & in2[38];
    assign P[100] = in[38] ^ in2[38];
    assign G[101] = in[37] & in2[37];
    assign P[101] = in[37] ^ in2[37];
    assign G[102] = in[36] & in2[36];
    assign P[102] = in[36] ^ in2[36];
    assign G[103] = in[35] & in2[35];
    assign P[103] = in[35] ^ in2[35];
    assign G[104] = in[34] & in2[34];
    assign P[104] = in[34] ^ in2[34];
    assign G[105] = in[33] & in2[33];
    assign P[105] = in[33] ^ in2[33];
    assign G[106] = in[32] & in2[32];
    assign P[106] = in[32] ^ in2[32];
    assign G[107] = in[31] & in2[31];
    assign P[107] = in[31] ^ in2[31];
    assign G[108] = in[30] & in2[30];
    assign P[108] = in[30] ^ in2[30];
    assign G[109] = in[29] & in2[29];
    assign P[109] = in[29] ^ in2[29];
    assign G[110] = in[28] & in2[28];
    assign P[110] = in[28] ^ in2[28];
    assign G[111] = in[27] & in2[27];
    assign P[111] = in[27] ^ in2[27];
    assign G[112] = in[26] & in2[26];
    assign P[112] = in[26] ^ in2[26];
    assign G[113] = in[25] & in2[25];
    assign P[113] = in[25] ^ in2[25];
    assign G[114] = in[24] & in2[24];
    assign P[114] = in[24] ^ in2[24];
    assign G[115] = in[23] & in2[23];
    assign P[115] = in[23] ^ in2[23];
    assign G[116] = in[22] & in2[22];
    assign P[116] = in[22] ^ in2[22];
    assign G[117] = in[21] & in2[21];
    assign P[117] = in[21] ^ in2[21];
    assign G[118] = in[20] & in2[20];
    assign P[118] = in[20] ^ in2[20];
    assign G[119] = in[19] & in2[19];
    assign P[119] = in[19] ^ in2[19];
    assign G[120] = in[18] & in2[18];
    assign P[120] = in[18] ^ in2[18];
    assign G[121] = in[17] & in2[17];
    assign P[121] = in[17] ^ in2[17];
    assign G[122] = in[16] & in2[16];
    assign P[122] = in[16] ^ in2[16];
    assign G[123] = in[15] & in2[15];
    assign P[123] = in[15] ^ in2[15];
    assign G[124] = in[14] & in2[14];
    assign P[124] = in[14] ^ in2[14];
    assign G[125] = in[13] & in2[13];
    assign P[125] = in[13] ^ in2[13];
    assign G[126] = in[12] & in2[12];
    assign P[126] = in[12] ^ in2[12];
    assign G[127] = in[11] & in2[11];
    assign P[127] = in[11] ^ in2[11];
    assign G[128] = in[10] & in2[10];
    assign P[128] = in[10] ^ in2[10];
    assign G[129] = in[9] & in2[9];
    assign P[129] = in[9] ^ in2[9];
    assign G[130] = in[8] & in2[8];
    assign P[130] = in[8] ^ in2[8];
    assign G[131] = in[7] & in2[7];
    assign P[131] = in[7] ^ in2[7];
    assign G[132] = in[6] & in2[6];
    assign P[132] = in[6] ^ in2[6];
    assign G[133] = in[5] & in2[5];
    assign P[133] = in[5] ^ in2[5];
    assign G[134] = in[4] & in2[4];
    assign P[134] = in[4] ^ in2[4];
    assign G[135] = in[3] & in2[3];
    assign P[135] = in[3] ^ in2[3];
    assign G[136] = in[2] & in2[2];
    assign P[136] = in[2] ^ in2[2];
    assign G[137] = in[1] & in2[1];
    assign P[137] = in[1] ^ in2[1];
    assign G[138] = in[0] & in2[0];
    assign P[138] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign C[138] = G[137] | (P[137] & C[137]);
    assign cout = G[138] | (P[138] & C[138]);
    assign sum = P ^ C;
endmodule

module CLA138(output [137:0] sum, output cout, input [137:0] in1, input [137:0] in2;

    wire[137:0] G;
    wire[137:0] C;
    wire[137:0] P;

    assign G[0] = in[137] & in2[137];
    assign P[0] = in[137] ^ in2[137];
    assign G[1] = in[136] & in2[136];
    assign P[1] = in[136] ^ in2[136];
    assign G[2] = in[135] & in2[135];
    assign P[2] = in[135] ^ in2[135];
    assign G[3] = in[134] & in2[134];
    assign P[3] = in[134] ^ in2[134];
    assign G[4] = in[133] & in2[133];
    assign P[4] = in[133] ^ in2[133];
    assign G[5] = in[132] & in2[132];
    assign P[5] = in[132] ^ in2[132];
    assign G[6] = in[131] & in2[131];
    assign P[6] = in[131] ^ in2[131];
    assign G[7] = in[130] & in2[130];
    assign P[7] = in[130] ^ in2[130];
    assign G[8] = in[129] & in2[129];
    assign P[8] = in[129] ^ in2[129];
    assign G[9] = in[128] & in2[128];
    assign P[9] = in[128] ^ in2[128];
    assign G[10] = in[127] & in2[127];
    assign P[10] = in[127] ^ in2[127];
    assign G[11] = in[126] & in2[126];
    assign P[11] = in[126] ^ in2[126];
    assign G[12] = in[125] & in2[125];
    assign P[12] = in[125] ^ in2[125];
    assign G[13] = in[124] & in2[124];
    assign P[13] = in[124] ^ in2[124];
    assign G[14] = in[123] & in2[123];
    assign P[14] = in[123] ^ in2[123];
    assign G[15] = in[122] & in2[122];
    assign P[15] = in[122] ^ in2[122];
    assign G[16] = in[121] & in2[121];
    assign P[16] = in[121] ^ in2[121];
    assign G[17] = in[120] & in2[120];
    assign P[17] = in[120] ^ in2[120];
    assign G[18] = in[119] & in2[119];
    assign P[18] = in[119] ^ in2[119];
    assign G[19] = in[118] & in2[118];
    assign P[19] = in[118] ^ in2[118];
    assign G[20] = in[117] & in2[117];
    assign P[20] = in[117] ^ in2[117];
    assign G[21] = in[116] & in2[116];
    assign P[21] = in[116] ^ in2[116];
    assign G[22] = in[115] & in2[115];
    assign P[22] = in[115] ^ in2[115];
    assign G[23] = in[114] & in2[114];
    assign P[23] = in[114] ^ in2[114];
    assign G[24] = in[113] & in2[113];
    assign P[24] = in[113] ^ in2[113];
    assign G[25] = in[112] & in2[112];
    assign P[25] = in[112] ^ in2[112];
    assign G[26] = in[111] & in2[111];
    assign P[26] = in[111] ^ in2[111];
    assign G[27] = in[110] & in2[110];
    assign P[27] = in[110] ^ in2[110];
    assign G[28] = in[109] & in2[109];
    assign P[28] = in[109] ^ in2[109];
    assign G[29] = in[108] & in2[108];
    assign P[29] = in[108] ^ in2[108];
    assign G[30] = in[107] & in2[107];
    assign P[30] = in[107] ^ in2[107];
    assign G[31] = in[106] & in2[106];
    assign P[31] = in[106] ^ in2[106];
    assign G[32] = in[105] & in2[105];
    assign P[32] = in[105] ^ in2[105];
    assign G[33] = in[104] & in2[104];
    assign P[33] = in[104] ^ in2[104];
    assign G[34] = in[103] & in2[103];
    assign P[34] = in[103] ^ in2[103];
    assign G[35] = in[102] & in2[102];
    assign P[35] = in[102] ^ in2[102];
    assign G[36] = in[101] & in2[101];
    assign P[36] = in[101] ^ in2[101];
    assign G[37] = in[100] & in2[100];
    assign P[37] = in[100] ^ in2[100];
    assign G[38] = in[99] & in2[99];
    assign P[38] = in[99] ^ in2[99];
    assign G[39] = in[98] & in2[98];
    assign P[39] = in[98] ^ in2[98];
    assign G[40] = in[97] & in2[97];
    assign P[40] = in[97] ^ in2[97];
    assign G[41] = in[96] & in2[96];
    assign P[41] = in[96] ^ in2[96];
    assign G[42] = in[95] & in2[95];
    assign P[42] = in[95] ^ in2[95];
    assign G[43] = in[94] & in2[94];
    assign P[43] = in[94] ^ in2[94];
    assign G[44] = in[93] & in2[93];
    assign P[44] = in[93] ^ in2[93];
    assign G[45] = in[92] & in2[92];
    assign P[45] = in[92] ^ in2[92];
    assign G[46] = in[91] & in2[91];
    assign P[46] = in[91] ^ in2[91];
    assign G[47] = in[90] & in2[90];
    assign P[47] = in[90] ^ in2[90];
    assign G[48] = in[89] & in2[89];
    assign P[48] = in[89] ^ in2[89];
    assign G[49] = in[88] & in2[88];
    assign P[49] = in[88] ^ in2[88];
    assign G[50] = in[87] & in2[87];
    assign P[50] = in[87] ^ in2[87];
    assign G[51] = in[86] & in2[86];
    assign P[51] = in[86] ^ in2[86];
    assign G[52] = in[85] & in2[85];
    assign P[52] = in[85] ^ in2[85];
    assign G[53] = in[84] & in2[84];
    assign P[53] = in[84] ^ in2[84];
    assign G[54] = in[83] & in2[83];
    assign P[54] = in[83] ^ in2[83];
    assign G[55] = in[82] & in2[82];
    assign P[55] = in[82] ^ in2[82];
    assign G[56] = in[81] & in2[81];
    assign P[56] = in[81] ^ in2[81];
    assign G[57] = in[80] & in2[80];
    assign P[57] = in[80] ^ in2[80];
    assign G[58] = in[79] & in2[79];
    assign P[58] = in[79] ^ in2[79];
    assign G[59] = in[78] & in2[78];
    assign P[59] = in[78] ^ in2[78];
    assign G[60] = in[77] & in2[77];
    assign P[60] = in[77] ^ in2[77];
    assign G[61] = in[76] & in2[76];
    assign P[61] = in[76] ^ in2[76];
    assign G[62] = in[75] & in2[75];
    assign P[62] = in[75] ^ in2[75];
    assign G[63] = in[74] & in2[74];
    assign P[63] = in[74] ^ in2[74];
    assign G[64] = in[73] & in2[73];
    assign P[64] = in[73] ^ in2[73];
    assign G[65] = in[72] & in2[72];
    assign P[65] = in[72] ^ in2[72];
    assign G[66] = in[71] & in2[71];
    assign P[66] = in[71] ^ in2[71];
    assign G[67] = in[70] & in2[70];
    assign P[67] = in[70] ^ in2[70];
    assign G[68] = in[69] & in2[69];
    assign P[68] = in[69] ^ in2[69];
    assign G[69] = in[68] & in2[68];
    assign P[69] = in[68] ^ in2[68];
    assign G[70] = in[67] & in2[67];
    assign P[70] = in[67] ^ in2[67];
    assign G[71] = in[66] & in2[66];
    assign P[71] = in[66] ^ in2[66];
    assign G[72] = in[65] & in2[65];
    assign P[72] = in[65] ^ in2[65];
    assign G[73] = in[64] & in2[64];
    assign P[73] = in[64] ^ in2[64];
    assign G[74] = in[63] & in2[63];
    assign P[74] = in[63] ^ in2[63];
    assign G[75] = in[62] & in2[62];
    assign P[75] = in[62] ^ in2[62];
    assign G[76] = in[61] & in2[61];
    assign P[76] = in[61] ^ in2[61];
    assign G[77] = in[60] & in2[60];
    assign P[77] = in[60] ^ in2[60];
    assign G[78] = in[59] & in2[59];
    assign P[78] = in[59] ^ in2[59];
    assign G[79] = in[58] & in2[58];
    assign P[79] = in[58] ^ in2[58];
    assign G[80] = in[57] & in2[57];
    assign P[80] = in[57] ^ in2[57];
    assign G[81] = in[56] & in2[56];
    assign P[81] = in[56] ^ in2[56];
    assign G[82] = in[55] & in2[55];
    assign P[82] = in[55] ^ in2[55];
    assign G[83] = in[54] & in2[54];
    assign P[83] = in[54] ^ in2[54];
    assign G[84] = in[53] & in2[53];
    assign P[84] = in[53] ^ in2[53];
    assign G[85] = in[52] & in2[52];
    assign P[85] = in[52] ^ in2[52];
    assign G[86] = in[51] & in2[51];
    assign P[86] = in[51] ^ in2[51];
    assign G[87] = in[50] & in2[50];
    assign P[87] = in[50] ^ in2[50];
    assign G[88] = in[49] & in2[49];
    assign P[88] = in[49] ^ in2[49];
    assign G[89] = in[48] & in2[48];
    assign P[89] = in[48] ^ in2[48];
    assign G[90] = in[47] & in2[47];
    assign P[90] = in[47] ^ in2[47];
    assign G[91] = in[46] & in2[46];
    assign P[91] = in[46] ^ in2[46];
    assign G[92] = in[45] & in2[45];
    assign P[92] = in[45] ^ in2[45];
    assign G[93] = in[44] & in2[44];
    assign P[93] = in[44] ^ in2[44];
    assign G[94] = in[43] & in2[43];
    assign P[94] = in[43] ^ in2[43];
    assign G[95] = in[42] & in2[42];
    assign P[95] = in[42] ^ in2[42];
    assign G[96] = in[41] & in2[41];
    assign P[96] = in[41] ^ in2[41];
    assign G[97] = in[40] & in2[40];
    assign P[97] = in[40] ^ in2[40];
    assign G[98] = in[39] & in2[39];
    assign P[98] = in[39] ^ in2[39];
    assign G[99] = in[38] & in2[38];
    assign P[99] = in[38] ^ in2[38];
    assign G[100] = in[37] & in2[37];
    assign P[100] = in[37] ^ in2[37];
    assign G[101] = in[36] & in2[36];
    assign P[101] = in[36] ^ in2[36];
    assign G[102] = in[35] & in2[35];
    assign P[102] = in[35] ^ in2[35];
    assign G[103] = in[34] & in2[34];
    assign P[103] = in[34] ^ in2[34];
    assign G[104] = in[33] & in2[33];
    assign P[104] = in[33] ^ in2[33];
    assign G[105] = in[32] & in2[32];
    assign P[105] = in[32] ^ in2[32];
    assign G[106] = in[31] & in2[31];
    assign P[106] = in[31] ^ in2[31];
    assign G[107] = in[30] & in2[30];
    assign P[107] = in[30] ^ in2[30];
    assign G[108] = in[29] & in2[29];
    assign P[108] = in[29] ^ in2[29];
    assign G[109] = in[28] & in2[28];
    assign P[109] = in[28] ^ in2[28];
    assign G[110] = in[27] & in2[27];
    assign P[110] = in[27] ^ in2[27];
    assign G[111] = in[26] & in2[26];
    assign P[111] = in[26] ^ in2[26];
    assign G[112] = in[25] & in2[25];
    assign P[112] = in[25] ^ in2[25];
    assign G[113] = in[24] & in2[24];
    assign P[113] = in[24] ^ in2[24];
    assign G[114] = in[23] & in2[23];
    assign P[114] = in[23] ^ in2[23];
    assign G[115] = in[22] & in2[22];
    assign P[115] = in[22] ^ in2[22];
    assign G[116] = in[21] & in2[21];
    assign P[116] = in[21] ^ in2[21];
    assign G[117] = in[20] & in2[20];
    assign P[117] = in[20] ^ in2[20];
    assign G[118] = in[19] & in2[19];
    assign P[118] = in[19] ^ in2[19];
    assign G[119] = in[18] & in2[18];
    assign P[119] = in[18] ^ in2[18];
    assign G[120] = in[17] & in2[17];
    assign P[120] = in[17] ^ in2[17];
    assign G[121] = in[16] & in2[16];
    assign P[121] = in[16] ^ in2[16];
    assign G[122] = in[15] & in2[15];
    assign P[122] = in[15] ^ in2[15];
    assign G[123] = in[14] & in2[14];
    assign P[123] = in[14] ^ in2[14];
    assign G[124] = in[13] & in2[13];
    assign P[124] = in[13] ^ in2[13];
    assign G[125] = in[12] & in2[12];
    assign P[125] = in[12] ^ in2[12];
    assign G[126] = in[11] & in2[11];
    assign P[126] = in[11] ^ in2[11];
    assign G[127] = in[10] & in2[10];
    assign P[127] = in[10] ^ in2[10];
    assign G[128] = in[9] & in2[9];
    assign P[128] = in[9] ^ in2[9];
    assign G[129] = in[8] & in2[8];
    assign P[129] = in[8] ^ in2[8];
    assign G[130] = in[7] & in2[7];
    assign P[130] = in[7] ^ in2[7];
    assign G[131] = in[6] & in2[6];
    assign P[131] = in[6] ^ in2[6];
    assign G[132] = in[5] & in2[5];
    assign P[132] = in[5] ^ in2[5];
    assign G[133] = in[4] & in2[4];
    assign P[133] = in[4] ^ in2[4];
    assign G[134] = in[3] & in2[3];
    assign P[134] = in[3] ^ in2[3];
    assign G[135] = in[2] & in2[2];
    assign P[135] = in[2] ^ in2[2];
    assign G[136] = in[1] & in2[1];
    assign P[136] = in[1] ^ in2[1];
    assign G[137] = in[0] & in2[0];
    assign P[137] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign C[137] = G[136] | (P[136] & C[136]);
    assign cout = G[137] | (P[137] & C[137]);
    assign sum = P ^ C;
endmodule

module CLA137(output [136:0] sum, output cout, input [136:0] in1, input [136:0] in2;

    wire[136:0] G;
    wire[136:0] C;
    wire[136:0] P;

    assign G[0] = in[136] & in2[136];
    assign P[0] = in[136] ^ in2[136];
    assign G[1] = in[135] & in2[135];
    assign P[1] = in[135] ^ in2[135];
    assign G[2] = in[134] & in2[134];
    assign P[2] = in[134] ^ in2[134];
    assign G[3] = in[133] & in2[133];
    assign P[3] = in[133] ^ in2[133];
    assign G[4] = in[132] & in2[132];
    assign P[4] = in[132] ^ in2[132];
    assign G[5] = in[131] & in2[131];
    assign P[5] = in[131] ^ in2[131];
    assign G[6] = in[130] & in2[130];
    assign P[6] = in[130] ^ in2[130];
    assign G[7] = in[129] & in2[129];
    assign P[7] = in[129] ^ in2[129];
    assign G[8] = in[128] & in2[128];
    assign P[8] = in[128] ^ in2[128];
    assign G[9] = in[127] & in2[127];
    assign P[9] = in[127] ^ in2[127];
    assign G[10] = in[126] & in2[126];
    assign P[10] = in[126] ^ in2[126];
    assign G[11] = in[125] & in2[125];
    assign P[11] = in[125] ^ in2[125];
    assign G[12] = in[124] & in2[124];
    assign P[12] = in[124] ^ in2[124];
    assign G[13] = in[123] & in2[123];
    assign P[13] = in[123] ^ in2[123];
    assign G[14] = in[122] & in2[122];
    assign P[14] = in[122] ^ in2[122];
    assign G[15] = in[121] & in2[121];
    assign P[15] = in[121] ^ in2[121];
    assign G[16] = in[120] & in2[120];
    assign P[16] = in[120] ^ in2[120];
    assign G[17] = in[119] & in2[119];
    assign P[17] = in[119] ^ in2[119];
    assign G[18] = in[118] & in2[118];
    assign P[18] = in[118] ^ in2[118];
    assign G[19] = in[117] & in2[117];
    assign P[19] = in[117] ^ in2[117];
    assign G[20] = in[116] & in2[116];
    assign P[20] = in[116] ^ in2[116];
    assign G[21] = in[115] & in2[115];
    assign P[21] = in[115] ^ in2[115];
    assign G[22] = in[114] & in2[114];
    assign P[22] = in[114] ^ in2[114];
    assign G[23] = in[113] & in2[113];
    assign P[23] = in[113] ^ in2[113];
    assign G[24] = in[112] & in2[112];
    assign P[24] = in[112] ^ in2[112];
    assign G[25] = in[111] & in2[111];
    assign P[25] = in[111] ^ in2[111];
    assign G[26] = in[110] & in2[110];
    assign P[26] = in[110] ^ in2[110];
    assign G[27] = in[109] & in2[109];
    assign P[27] = in[109] ^ in2[109];
    assign G[28] = in[108] & in2[108];
    assign P[28] = in[108] ^ in2[108];
    assign G[29] = in[107] & in2[107];
    assign P[29] = in[107] ^ in2[107];
    assign G[30] = in[106] & in2[106];
    assign P[30] = in[106] ^ in2[106];
    assign G[31] = in[105] & in2[105];
    assign P[31] = in[105] ^ in2[105];
    assign G[32] = in[104] & in2[104];
    assign P[32] = in[104] ^ in2[104];
    assign G[33] = in[103] & in2[103];
    assign P[33] = in[103] ^ in2[103];
    assign G[34] = in[102] & in2[102];
    assign P[34] = in[102] ^ in2[102];
    assign G[35] = in[101] & in2[101];
    assign P[35] = in[101] ^ in2[101];
    assign G[36] = in[100] & in2[100];
    assign P[36] = in[100] ^ in2[100];
    assign G[37] = in[99] & in2[99];
    assign P[37] = in[99] ^ in2[99];
    assign G[38] = in[98] & in2[98];
    assign P[38] = in[98] ^ in2[98];
    assign G[39] = in[97] & in2[97];
    assign P[39] = in[97] ^ in2[97];
    assign G[40] = in[96] & in2[96];
    assign P[40] = in[96] ^ in2[96];
    assign G[41] = in[95] & in2[95];
    assign P[41] = in[95] ^ in2[95];
    assign G[42] = in[94] & in2[94];
    assign P[42] = in[94] ^ in2[94];
    assign G[43] = in[93] & in2[93];
    assign P[43] = in[93] ^ in2[93];
    assign G[44] = in[92] & in2[92];
    assign P[44] = in[92] ^ in2[92];
    assign G[45] = in[91] & in2[91];
    assign P[45] = in[91] ^ in2[91];
    assign G[46] = in[90] & in2[90];
    assign P[46] = in[90] ^ in2[90];
    assign G[47] = in[89] & in2[89];
    assign P[47] = in[89] ^ in2[89];
    assign G[48] = in[88] & in2[88];
    assign P[48] = in[88] ^ in2[88];
    assign G[49] = in[87] & in2[87];
    assign P[49] = in[87] ^ in2[87];
    assign G[50] = in[86] & in2[86];
    assign P[50] = in[86] ^ in2[86];
    assign G[51] = in[85] & in2[85];
    assign P[51] = in[85] ^ in2[85];
    assign G[52] = in[84] & in2[84];
    assign P[52] = in[84] ^ in2[84];
    assign G[53] = in[83] & in2[83];
    assign P[53] = in[83] ^ in2[83];
    assign G[54] = in[82] & in2[82];
    assign P[54] = in[82] ^ in2[82];
    assign G[55] = in[81] & in2[81];
    assign P[55] = in[81] ^ in2[81];
    assign G[56] = in[80] & in2[80];
    assign P[56] = in[80] ^ in2[80];
    assign G[57] = in[79] & in2[79];
    assign P[57] = in[79] ^ in2[79];
    assign G[58] = in[78] & in2[78];
    assign P[58] = in[78] ^ in2[78];
    assign G[59] = in[77] & in2[77];
    assign P[59] = in[77] ^ in2[77];
    assign G[60] = in[76] & in2[76];
    assign P[60] = in[76] ^ in2[76];
    assign G[61] = in[75] & in2[75];
    assign P[61] = in[75] ^ in2[75];
    assign G[62] = in[74] & in2[74];
    assign P[62] = in[74] ^ in2[74];
    assign G[63] = in[73] & in2[73];
    assign P[63] = in[73] ^ in2[73];
    assign G[64] = in[72] & in2[72];
    assign P[64] = in[72] ^ in2[72];
    assign G[65] = in[71] & in2[71];
    assign P[65] = in[71] ^ in2[71];
    assign G[66] = in[70] & in2[70];
    assign P[66] = in[70] ^ in2[70];
    assign G[67] = in[69] & in2[69];
    assign P[67] = in[69] ^ in2[69];
    assign G[68] = in[68] & in2[68];
    assign P[68] = in[68] ^ in2[68];
    assign G[69] = in[67] & in2[67];
    assign P[69] = in[67] ^ in2[67];
    assign G[70] = in[66] & in2[66];
    assign P[70] = in[66] ^ in2[66];
    assign G[71] = in[65] & in2[65];
    assign P[71] = in[65] ^ in2[65];
    assign G[72] = in[64] & in2[64];
    assign P[72] = in[64] ^ in2[64];
    assign G[73] = in[63] & in2[63];
    assign P[73] = in[63] ^ in2[63];
    assign G[74] = in[62] & in2[62];
    assign P[74] = in[62] ^ in2[62];
    assign G[75] = in[61] & in2[61];
    assign P[75] = in[61] ^ in2[61];
    assign G[76] = in[60] & in2[60];
    assign P[76] = in[60] ^ in2[60];
    assign G[77] = in[59] & in2[59];
    assign P[77] = in[59] ^ in2[59];
    assign G[78] = in[58] & in2[58];
    assign P[78] = in[58] ^ in2[58];
    assign G[79] = in[57] & in2[57];
    assign P[79] = in[57] ^ in2[57];
    assign G[80] = in[56] & in2[56];
    assign P[80] = in[56] ^ in2[56];
    assign G[81] = in[55] & in2[55];
    assign P[81] = in[55] ^ in2[55];
    assign G[82] = in[54] & in2[54];
    assign P[82] = in[54] ^ in2[54];
    assign G[83] = in[53] & in2[53];
    assign P[83] = in[53] ^ in2[53];
    assign G[84] = in[52] & in2[52];
    assign P[84] = in[52] ^ in2[52];
    assign G[85] = in[51] & in2[51];
    assign P[85] = in[51] ^ in2[51];
    assign G[86] = in[50] & in2[50];
    assign P[86] = in[50] ^ in2[50];
    assign G[87] = in[49] & in2[49];
    assign P[87] = in[49] ^ in2[49];
    assign G[88] = in[48] & in2[48];
    assign P[88] = in[48] ^ in2[48];
    assign G[89] = in[47] & in2[47];
    assign P[89] = in[47] ^ in2[47];
    assign G[90] = in[46] & in2[46];
    assign P[90] = in[46] ^ in2[46];
    assign G[91] = in[45] & in2[45];
    assign P[91] = in[45] ^ in2[45];
    assign G[92] = in[44] & in2[44];
    assign P[92] = in[44] ^ in2[44];
    assign G[93] = in[43] & in2[43];
    assign P[93] = in[43] ^ in2[43];
    assign G[94] = in[42] & in2[42];
    assign P[94] = in[42] ^ in2[42];
    assign G[95] = in[41] & in2[41];
    assign P[95] = in[41] ^ in2[41];
    assign G[96] = in[40] & in2[40];
    assign P[96] = in[40] ^ in2[40];
    assign G[97] = in[39] & in2[39];
    assign P[97] = in[39] ^ in2[39];
    assign G[98] = in[38] & in2[38];
    assign P[98] = in[38] ^ in2[38];
    assign G[99] = in[37] & in2[37];
    assign P[99] = in[37] ^ in2[37];
    assign G[100] = in[36] & in2[36];
    assign P[100] = in[36] ^ in2[36];
    assign G[101] = in[35] & in2[35];
    assign P[101] = in[35] ^ in2[35];
    assign G[102] = in[34] & in2[34];
    assign P[102] = in[34] ^ in2[34];
    assign G[103] = in[33] & in2[33];
    assign P[103] = in[33] ^ in2[33];
    assign G[104] = in[32] & in2[32];
    assign P[104] = in[32] ^ in2[32];
    assign G[105] = in[31] & in2[31];
    assign P[105] = in[31] ^ in2[31];
    assign G[106] = in[30] & in2[30];
    assign P[106] = in[30] ^ in2[30];
    assign G[107] = in[29] & in2[29];
    assign P[107] = in[29] ^ in2[29];
    assign G[108] = in[28] & in2[28];
    assign P[108] = in[28] ^ in2[28];
    assign G[109] = in[27] & in2[27];
    assign P[109] = in[27] ^ in2[27];
    assign G[110] = in[26] & in2[26];
    assign P[110] = in[26] ^ in2[26];
    assign G[111] = in[25] & in2[25];
    assign P[111] = in[25] ^ in2[25];
    assign G[112] = in[24] & in2[24];
    assign P[112] = in[24] ^ in2[24];
    assign G[113] = in[23] & in2[23];
    assign P[113] = in[23] ^ in2[23];
    assign G[114] = in[22] & in2[22];
    assign P[114] = in[22] ^ in2[22];
    assign G[115] = in[21] & in2[21];
    assign P[115] = in[21] ^ in2[21];
    assign G[116] = in[20] & in2[20];
    assign P[116] = in[20] ^ in2[20];
    assign G[117] = in[19] & in2[19];
    assign P[117] = in[19] ^ in2[19];
    assign G[118] = in[18] & in2[18];
    assign P[118] = in[18] ^ in2[18];
    assign G[119] = in[17] & in2[17];
    assign P[119] = in[17] ^ in2[17];
    assign G[120] = in[16] & in2[16];
    assign P[120] = in[16] ^ in2[16];
    assign G[121] = in[15] & in2[15];
    assign P[121] = in[15] ^ in2[15];
    assign G[122] = in[14] & in2[14];
    assign P[122] = in[14] ^ in2[14];
    assign G[123] = in[13] & in2[13];
    assign P[123] = in[13] ^ in2[13];
    assign G[124] = in[12] & in2[12];
    assign P[124] = in[12] ^ in2[12];
    assign G[125] = in[11] & in2[11];
    assign P[125] = in[11] ^ in2[11];
    assign G[126] = in[10] & in2[10];
    assign P[126] = in[10] ^ in2[10];
    assign G[127] = in[9] & in2[9];
    assign P[127] = in[9] ^ in2[9];
    assign G[128] = in[8] & in2[8];
    assign P[128] = in[8] ^ in2[8];
    assign G[129] = in[7] & in2[7];
    assign P[129] = in[7] ^ in2[7];
    assign G[130] = in[6] & in2[6];
    assign P[130] = in[6] ^ in2[6];
    assign G[131] = in[5] & in2[5];
    assign P[131] = in[5] ^ in2[5];
    assign G[132] = in[4] & in2[4];
    assign P[132] = in[4] ^ in2[4];
    assign G[133] = in[3] & in2[3];
    assign P[133] = in[3] ^ in2[3];
    assign G[134] = in[2] & in2[2];
    assign P[134] = in[2] ^ in2[2];
    assign G[135] = in[1] & in2[1];
    assign P[135] = in[1] ^ in2[1];
    assign G[136] = in[0] & in2[0];
    assign P[136] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign C[136] = G[135] | (P[135] & C[135]);
    assign cout = G[136] | (P[136] & C[136]);
    assign sum = P ^ C;
endmodule

module CLA136(output [135:0] sum, output cout, input [135:0] in1, input [135:0] in2;

    wire[135:0] G;
    wire[135:0] C;
    wire[135:0] P;

    assign G[0] = in[135] & in2[135];
    assign P[0] = in[135] ^ in2[135];
    assign G[1] = in[134] & in2[134];
    assign P[1] = in[134] ^ in2[134];
    assign G[2] = in[133] & in2[133];
    assign P[2] = in[133] ^ in2[133];
    assign G[3] = in[132] & in2[132];
    assign P[3] = in[132] ^ in2[132];
    assign G[4] = in[131] & in2[131];
    assign P[4] = in[131] ^ in2[131];
    assign G[5] = in[130] & in2[130];
    assign P[5] = in[130] ^ in2[130];
    assign G[6] = in[129] & in2[129];
    assign P[6] = in[129] ^ in2[129];
    assign G[7] = in[128] & in2[128];
    assign P[7] = in[128] ^ in2[128];
    assign G[8] = in[127] & in2[127];
    assign P[8] = in[127] ^ in2[127];
    assign G[9] = in[126] & in2[126];
    assign P[9] = in[126] ^ in2[126];
    assign G[10] = in[125] & in2[125];
    assign P[10] = in[125] ^ in2[125];
    assign G[11] = in[124] & in2[124];
    assign P[11] = in[124] ^ in2[124];
    assign G[12] = in[123] & in2[123];
    assign P[12] = in[123] ^ in2[123];
    assign G[13] = in[122] & in2[122];
    assign P[13] = in[122] ^ in2[122];
    assign G[14] = in[121] & in2[121];
    assign P[14] = in[121] ^ in2[121];
    assign G[15] = in[120] & in2[120];
    assign P[15] = in[120] ^ in2[120];
    assign G[16] = in[119] & in2[119];
    assign P[16] = in[119] ^ in2[119];
    assign G[17] = in[118] & in2[118];
    assign P[17] = in[118] ^ in2[118];
    assign G[18] = in[117] & in2[117];
    assign P[18] = in[117] ^ in2[117];
    assign G[19] = in[116] & in2[116];
    assign P[19] = in[116] ^ in2[116];
    assign G[20] = in[115] & in2[115];
    assign P[20] = in[115] ^ in2[115];
    assign G[21] = in[114] & in2[114];
    assign P[21] = in[114] ^ in2[114];
    assign G[22] = in[113] & in2[113];
    assign P[22] = in[113] ^ in2[113];
    assign G[23] = in[112] & in2[112];
    assign P[23] = in[112] ^ in2[112];
    assign G[24] = in[111] & in2[111];
    assign P[24] = in[111] ^ in2[111];
    assign G[25] = in[110] & in2[110];
    assign P[25] = in[110] ^ in2[110];
    assign G[26] = in[109] & in2[109];
    assign P[26] = in[109] ^ in2[109];
    assign G[27] = in[108] & in2[108];
    assign P[27] = in[108] ^ in2[108];
    assign G[28] = in[107] & in2[107];
    assign P[28] = in[107] ^ in2[107];
    assign G[29] = in[106] & in2[106];
    assign P[29] = in[106] ^ in2[106];
    assign G[30] = in[105] & in2[105];
    assign P[30] = in[105] ^ in2[105];
    assign G[31] = in[104] & in2[104];
    assign P[31] = in[104] ^ in2[104];
    assign G[32] = in[103] & in2[103];
    assign P[32] = in[103] ^ in2[103];
    assign G[33] = in[102] & in2[102];
    assign P[33] = in[102] ^ in2[102];
    assign G[34] = in[101] & in2[101];
    assign P[34] = in[101] ^ in2[101];
    assign G[35] = in[100] & in2[100];
    assign P[35] = in[100] ^ in2[100];
    assign G[36] = in[99] & in2[99];
    assign P[36] = in[99] ^ in2[99];
    assign G[37] = in[98] & in2[98];
    assign P[37] = in[98] ^ in2[98];
    assign G[38] = in[97] & in2[97];
    assign P[38] = in[97] ^ in2[97];
    assign G[39] = in[96] & in2[96];
    assign P[39] = in[96] ^ in2[96];
    assign G[40] = in[95] & in2[95];
    assign P[40] = in[95] ^ in2[95];
    assign G[41] = in[94] & in2[94];
    assign P[41] = in[94] ^ in2[94];
    assign G[42] = in[93] & in2[93];
    assign P[42] = in[93] ^ in2[93];
    assign G[43] = in[92] & in2[92];
    assign P[43] = in[92] ^ in2[92];
    assign G[44] = in[91] & in2[91];
    assign P[44] = in[91] ^ in2[91];
    assign G[45] = in[90] & in2[90];
    assign P[45] = in[90] ^ in2[90];
    assign G[46] = in[89] & in2[89];
    assign P[46] = in[89] ^ in2[89];
    assign G[47] = in[88] & in2[88];
    assign P[47] = in[88] ^ in2[88];
    assign G[48] = in[87] & in2[87];
    assign P[48] = in[87] ^ in2[87];
    assign G[49] = in[86] & in2[86];
    assign P[49] = in[86] ^ in2[86];
    assign G[50] = in[85] & in2[85];
    assign P[50] = in[85] ^ in2[85];
    assign G[51] = in[84] & in2[84];
    assign P[51] = in[84] ^ in2[84];
    assign G[52] = in[83] & in2[83];
    assign P[52] = in[83] ^ in2[83];
    assign G[53] = in[82] & in2[82];
    assign P[53] = in[82] ^ in2[82];
    assign G[54] = in[81] & in2[81];
    assign P[54] = in[81] ^ in2[81];
    assign G[55] = in[80] & in2[80];
    assign P[55] = in[80] ^ in2[80];
    assign G[56] = in[79] & in2[79];
    assign P[56] = in[79] ^ in2[79];
    assign G[57] = in[78] & in2[78];
    assign P[57] = in[78] ^ in2[78];
    assign G[58] = in[77] & in2[77];
    assign P[58] = in[77] ^ in2[77];
    assign G[59] = in[76] & in2[76];
    assign P[59] = in[76] ^ in2[76];
    assign G[60] = in[75] & in2[75];
    assign P[60] = in[75] ^ in2[75];
    assign G[61] = in[74] & in2[74];
    assign P[61] = in[74] ^ in2[74];
    assign G[62] = in[73] & in2[73];
    assign P[62] = in[73] ^ in2[73];
    assign G[63] = in[72] & in2[72];
    assign P[63] = in[72] ^ in2[72];
    assign G[64] = in[71] & in2[71];
    assign P[64] = in[71] ^ in2[71];
    assign G[65] = in[70] & in2[70];
    assign P[65] = in[70] ^ in2[70];
    assign G[66] = in[69] & in2[69];
    assign P[66] = in[69] ^ in2[69];
    assign G[67] = in[68] & in2[68];
    assign P[67] = in[68] ^ in2[68];
    assign G[68] = in[67] & in2[67];
    assign P[68] = in[67] ^ in2[67];
    assign G[69] = in[66] & in2[66];
    assign P[69] = in[66] ^ in2[66];
    assign G[70] = in[65] & in2[65];
    assign P[70] = in[65] ^ in2[65];
    assign G[71] = in[64] & in2[64];
    assign P[71] = in[64] ^ in2[64];
    assign G[72] = in[63] & in2[63];
    assign P[72] = in[63] ^ in2[63];
    assign G[73] = in[62] & in2[62];
    assign P[73] = in[62] ^ in2[62];
    assign G[74] = in[61] & in2[61];
    assign P[74] = in[61] ^ in2[61];
    assign G[75] = in[60] & in2[60];
    assign P[75] = in[60] ^ in2[60];
    assign G[76] = in[59] & in2[59];
    assign P[76] = in[59] ^ in2[59];
    assign G[77] = in[58] & in2[58];
    assign P[77] = in[58] ^ in2[58];
    assign G[78] = in[57] & in2[57];
    assign P[78] = in[57] ^ in2[57];
    assign G[79] = in[56] & in2[56];
    assign P[79] = in[56] ^ in2[56];
    assign G[80] = in[55] & in2[55];
    assign P[80] = in[55] ^ in2[55];
    assign G[81] = in[54] & in2[54];
    assign P[81] = in[54] ^ in2[54];
    assign G[82] = in[53] & in2[53];
    assign P[82] = in[53] ^ in2[53];
    assign G[83] = in[52] & in2[52];
    assign P[83] = in[52] ^ in2[52];
    assign G[84] = in[51] & in2[51];
    assign P[84] = in[51] ^ in2[51];
    assign G[85] = in[50] & in2[50];
    assign P[85] = in[50] ^ in2[50];
    assign G[86] = in[49] & in2[49];
    assign P[86] = in[49] ^ in2[49];
    assign G[87] = in[48] & in2[48];
    assign P[87] = in[48] ^ in2[48];
    assign G[88] = in[47] & in2[47];
    assign P[88] = in[47] ^ in2[47];
    assign G[89] = in[46] & in2[46];
    assign P[89] = in[46] ^ in2[46];
    assign G[90] = in[45] & in2[45];
    assign P[90] = in[45] ^ in2[45];
    assign G[91] = in[44] & in2[44];
    assign P[91] = in[44] ^ in2[44];
    assign G[92] = in[43] & in2[43];
    assign P[92] = in[43] ^ in2[43];
    assign G[93] = in[42] & in2[42];
    assign P[93] = in[42] ^ in2[42];
    assign G[94] = in[41] & in2[41];
    assign P[94] = in[41] ^ in2[41];
    assign G[95] = in[40] & in2[40];
    assign P[95] = in[40] ^ in2[40];
    assign G[96] = in[39] & in2[39];
    assign P[96] = in[39] ^ in2[39];
    assign G[97] = in[38] & in2[38];
    assign P[97] = in[38] ^ in2[38];
    assign G[98] = in[37] & in2[37];
    assign P[98] = in[37] ^ in2[37];
    assign G[99] = in[36] & in2[36];
    assign P[99] = in[36] ^ in2[36];
    assign G[100] = in[35] & in2[35];
    assign P[100] = in[35] ^ in2[35];
    assign G[101] = in[34] & in2[34];
    assign P[101] = in[34] ^ in2[34];
    assign G[102] = in[33] & in2[33];
    assign P[102] = in[33] ^ in2[33];
    assign G[103] = in[32] & in2[32];
    assign P[103] = in[32] ^ in2[32];
    assign G[104] = in[31] & in2[31];
    assign P[104] = in[31] ^ in2[31];
    assign G[105] = in[30] & in2[30];
    assign P[105] = in[30] ^ in2[30];
    assign G[106] = in[29] & in2[29];
    assign P[106] = in[29] ^ in2[29];
    assign G[107] = in[28] & in2[28];
    assign P[107] = in[28] ^ in2[28];
    assign G[108] = in[27] & in2[27];
    assign P[108] = in[27] ^ in2[27];
    assign G[109] = in[26] & in2[26];
    assign P[109] = in[26] ^ in2[26];
    assign G[110] = in[25] & in2[25];
    assign P[110] = in[25] ^ in2[25];
    assign G[111] = in[24] & in2[24];
    assign P[111] = in[24] ^ in2[24];
    assign G[112] = in[23] & in2[23];
    assign P[112] = in[23] ^ in2[23];
    assign G[113] = in[22] & in2[22];
    assign P[113] = in[22] ^ in2[22];
    assign G[114] = in[21] & in2[21];
    assign P[114] = in[21] ^ in2[21];
    assign G[115] = in[20] & in2[20];
    assign P[115] = in[20] ^ in2[20];
    assign G[116] = in[19] & in2[19];
    assign P[116] = in[19] ^ in2[19];
    assign G[117] = in[18] & in2[18];
    assign P[117] = in[18] ^ in2[18];
    assign G[118] = in[17] & in2[17];
    assign P[118] = in[17] ^ in2[17];
    assign G[119] = in[16] & in2[16];
    assign P[119] = in[16] ^ in2[16];
    assign G[120] = in[15] & in2[15];
    assign P[120] = in[15] ^ in2[15];
    assign G[121] = in[14] & in2[14];
    assign P[121] = in[14] ^ in2[14];
    assign G[122] = in[13] & in2[13];
    assign P[122] = in[13] ^ in2[13];
    assign G[123] = in[12] & in2[12];
    assign P[123] = in[12] ^ in2[12];
    assign G[124] = in[11] & in2[11];
    assign P[124] = in[11] ^ in2[11];
    assign G[125] = in[10] & in2[10];
    assign P[125] = in[10] ^ in2[10];
    assign G[126] = in[9] & in2[9];
    assign P[126] = in[9] ^ in2[9];
    assign G[127] = in[8] & in2[8];
    assign P[127] = in[8] ^ in2[8];
    assign G[128] = in[7] & in2[7];
    assign P[128] = in[7] ^ in2[7];
    assign G[129] = in[6] & in2[6];
    assign P[129] = in[6] ^ in2[6];
    assign G[130] = in[5] & in2[5];
    assign P[130] = in[5] ^ in2[5];
    assign G[131] = in[4] & in2[4];
    assign P[131] = in[4] ^ in2[4];
    assign G[132] = in[3] & in2[3];
    assign P[132] = in[3] ^ in2[3];
    assign G[133] = in[2] & in2[2];
    assign P[133] = in[2] ^ in2[2];
    assign G[134] = in[1] & in2[1];
    assign P[134] = in[1] ^ in2[1];
    assign G[135] = in[0] & in2[0];
    assign P[135] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign C[135] = G[134] | (P[134] & C[134]);
    assign cout = G[135] | (P[135] & C[135]);
    assign sum = P ^ C;
endmodule

module CLA135(output [134:0] sum, output cout, input [134:0] in1, input [134:0] in2;

    wire[134:0] G;
    wire[134:0] C;
    wire[134:0] P;

    assign G[0] = in[134] & in2[134];
    assign P[0] = in[134] ^ in2[134];
    assign G[1] = in[133] & in2[133];
    assign P[1] = in[133] ^ in2[133];
    assign G[2] = in[132] & in2[132];
    assign P[2] = in[132] ^ in2[132];
    assign G[3] = in[131] & in2[131];
    assign P[3] = in[131] ^ in2[131];
    assign G[4] = in[130] & in2[130];
    assign P[4] = in[130] ^ in2[130];
    assign G[5] = in[129] & in2[129];
    assign P[5] = in[129] ^ in2[129];
    assign G[6] = in[128] & in2[128];
    assign P[6] = in[128] ^ in2[128];
    assign G[7] = in[127] & in2[127];
    assign P[7] = in[127] ^ in2[127];
    assign G[8] = in[126] & in2[126];
    assign P[8] = in[126] ^ in2[126];
    assign G[9] = in[125] & in2[125];
    assign P[9] = in[125] ^ in2[125];
    assign G[10] = in[124] & in2[124];
    assign P[10] = in[124] ^ in2[124];
    assign G[11] = in[123] & in2[123];
    assign P[11] = in[123] ^ in2[123];
    assign G[12] = in[122] & in2[122];
    assign P[12] = in[122] ^ in2[122];
    assign G[13] = in[121] & in2[121];
    assign P[13] = in[121] ^ in2[121];
    assign G[14] = in[120] & in2[120];
    assign P[14] = in[120] ^ in2[120];
    assign G[15] = in[119] & in2[119];
    assign P[15] = in[119] ^ in2[119];
    assign G[16] = in[118] & in2[118];
    assign P[16] = in[118] ^ in2[118];
    assign G[17] = in[117] & in2[117];
    assign P[17] = in[117] ^ in2[117];
    assign G[18] = in[116] & in2[116];
    assign P[18] = in[116] ^ in2[116];
    assign G[19] = in[115] & in2[115];
    assign P[19] = in[115] ^ in2[115];
    assign G[20] = in[114] & in2[114];
    assign P[20] = in[114] ^ in2[114];
    assign G[21] = in[113] & in2[113];
    assign P[21] = in[113] ^ in2[113];
    assign G[22] = in[112] & in2[112];
    assign P[22] = in[112] ^ in2[112];
    assign G[23] = in[111] & in2[111];
    assign P[23] = in[111] ^ in2[111];
    assign G[24] = in[110] & in2[110];
    assign P[24] = in[110] ^ in2[110];
    assign G[25] = in[109] & in2[109];
    assign P[25] = in[109] ^ in2[109];
    assign G[26] = in[108] & in2[108];
    assign P[26] = in[108] ^ in2[108];
    assign G[27] = in[107] & in2[107];
    assign P[27] = in[107] ^ in2[107];
    assign G[28] = in[106] & in2[106];
    assign P[28] = in[106] ^ in2[106];
    assign G[29] = in[105] & in2[105];
    assign P[29] = in[105] ^ in2[105];
    assign G[30] = in[104] & in2[104];
    assign P[30] = in[104] ^ in2[104];
    assign G[31] = in[103] & in2[103];
    assign P[31] = in[103] ^ in2[103];
    assign G[32] = in[102] & in2[102];
    assign P[32] = in[102] ^ in2[102];
    assign G[33] = in[101] & in2[101];
    assign P[33] = in[101] ^ in2[101];
    assign G[34] = in[100] & in2[100];
    assign P[34] = in[100] ^ in2[100];
    assign G[35] = in[99] & in2[99];
    assign P[35] = in[99] ^ in2[99];
    assign G[36] = in[98] & in2[98];
    assign P[36] = in[98] ^ in2[98];
    assign G[37] = in[97] & in2[97];
    assign P[37] = in[97] ^ in2[97];
    assign G[38] = in[96] & in2[96];
    assign P[38] = in[96] ^ in2[96];
    assign G[39] = in[95] & in2[95];
    assign P[39] = in[95] ^ in2[95];
    assign G[40] = in[94] & in2[94];
    assign P[40] = in[94] ^ in2[94];
    assign G[41] = in[93] & in2[93];
    assign P[41] = in[93] ^ in2[93];
    assign G[42] = in[92] & in2[92];
    assign P[42] = in[92] ^ in2[92];
    assign G[43] = in[91] & in2[91];
    assign P[43] = in[91] ^ in2[91];
    assign G[44] = in[90] & in2[90];
    assign P[44] = in[90] ^ in2[90];
    assign G[45] = in[89] & in2[89];
    assign P[45] = in[89] ^ in2[89];
    assign G[46] = in[88] & in2[88];
    assign P[46] = in[88] ^ in2[88];
    assign G[47] = in[87] & in2[87];
    assign P[47] = in[87] ^ in2[87];
    assign G[48] = in[86] & in2[86];
    assign P[48] = in[86] ^ in2[86];
    assign G[49] = in[85] & in2[85];
    assign P[49] = in[85] ^ in2[85];
    assign G[50] = in[84] & in2[84];
    assign P[50] = in[84] ^ in2[84];
    assign G[51] = in[83] & in2[83];
    assign P[51] = in[83] ^ in2[83];
    assign G[52] = in[82] & in2[82];
    assign P[52] = in[82] ^ in2[82];
    assign G[53] = in[81] & in2[81];
    assign P[53] = in[81] ^ in2[81];
    assign G[54] = in[80] & in2[80];
    assign P[54] = in[80] ^ in2[80];
    assign G[55] = in[79] & in2[79];
    assign P[55] = in[79] ^ in2[79];
    assign G[56] = in[78] & in2[78];
    assign P[56] = in[78] ^ in2[78];
    assign G[57] = in[77] & in2[77];
    assign P[57] = in[77] ^ in2[77];
    assign G[58] = in[76] & in2[76];
    assign P[58] = in[76] ^ in2[76];
    assign G[59] = in[75] & in2[75];
    assign P[59] = in[75] ^ in2[75];
    assign G[60] = in[74] & in2[74];
    assign P[60] = in[74] ^ in2[74];
    assign G[61] = in[73] & in2[73];
    assign P[61] = in[73] ^ in2[73];
    assign G[62] = in[72] & in2[72];
    assign P[62] = in[72] ^ in2[72];
    assign G[63] = in[71] & in2[71];
    assign P[63] = in[71] ^ in2[71];
    assign G[64] = in[70] & in2[70];
    assign P[64] = in[70] ^ in2[70];
    assign G[65] = in[69] & in2[69];
    assign P[65] = in[69] ^ in2[69];
    assign G[66] = in[68] & in2[68];
    assign P[66] = in[68] ^ in2[68];
    assign G[67] = in[67] & in2[67];
    assign P[67] = in[67] ^ in2[67];
    assign G[68] = in[66] & in2[66];
    assign P[68] = in[66] ^ in2[66];
    assign G[69] = in[65] & in2[65];
    assign P[69] = in[65] ^ in2[65];
    assign G[70] = in[64] & in2[64];
    assign P[70] = in[64] ^ in2[64];
    assign G[71] = in[63] & in2[63];
    assign P[71] = in[63] ^ in2[63];
    assign G[72] = in[62] & in2[62];
    assign P[72] = in[62] ^ in2[62];
    assign G[73] = in[61] & in2[61];
    assign P[73] = in[61] ^ in2[61];
    assign G[74] = in[60] & in2[60];
    assign P[74] = in[60] ^ in2[60];
    assign G[75] = in[59] & in2[59];
    assign P[75] = in[59] ^ in2[59];
    assign G[76] = in[58] & in2[58];
    assign P[76] = in[58] ^ in2[58];
    assign G[77] = in[57] & in2[57];
    assign P[77] = in[57] ^ in2[57];
    assign G[78] = in[56] & in2[56];
    assign P[78] = in[56] ^ in2[56];
    assign G[79] = in[55] & in2[55];
    assign P[79] = in[55] ^ in2[55];
    assign G[80] = in[54] & in2[54];
    assign P[80] = in[54] ^ in2[54];
    assign G[81] = in[53] & in2[53];
    assign P[81] = in[53] ^ in2[53];
    assign G[82] = in[52] & in2[52];
    assign P[82] = in[52] ^ in2[52];
    assign G[83] = in[51] & in2[51];
    assign P[83] = in[51] ^ in2[51];
    assign G[84] = in[50] & in2[50];
    assign P[84] = in[50] ^ in2[50];
    assign G[85] = in[49] & in2[49];
    assign P[85] = in[49] ^ in2[49];
    assign G[86] = in[48] & in2[48];
    assign P[86] = in[48] ^ in2[48];
    assign G[87] = in[47] & in2[47];
    assign P[87] = in[47] ^ in2[47];
    assign G[88] = in[46] & in2[46];
    assign P[88] = in[46] ^ in2[46];
    assign G[89] = in[45] & in2[45];
    assign P[89] = in[45] ^ in2[45];
    assign G[90] = in[44] & in2[44];
    assign P[90] = in[44] ^ in2[44];
    assign G[91] = in[43] & in2[43];
    assign P[91] = in[43] ^ in2[43];
    assign G[92] = in[42] & in2[42];
    assign P[92] = in[42] ^ in2[42];
    assign G[93] = in[41] & in2[41];
    assign P[93] = in[41] ^ in2[41];
    assign G[94] = in[40] & in2[40];
    assign P[94] = in[40] ^ in2[40];
    assign G[95] = in[39] & in2[39];
    assign P[95] = in[39] ^ in2[39];
    assign G[96] = in[38] & in2[38];
    assign P[96] = in[38] ^ in2[38];
    assign G[97] = in[37] & in2[37];
    assign P[97] = in[37] ^ in2[37];
    assign G[98] = in[36] & in2[36];
    assign P[98] = in[36] ^ in2[36];
    assign G[99] = in[35] & in2[35];
    assign P[99] = in[35] ^ in2[35];
    assign G[100] = in[34] & in2[34];
    assign P[100] = in[34] ^ in2[34];
    assign G[101] = in[33] & in2[33];
    assign P[101] = in[33] ^ in2[33];
    assign G[102] = in[32] & in2[32];
    assign P[102] = in[32] ^ in2[32];
    assign G[103] = in[31] & in2[31];
    assign P[103] = in[31] ^ in2[31];
    assign G[104] = in[30] & in2[30];
    assign P[104] = in[30] ^ in2[30];
    assign G[105] = in[29] & in2[29];
    assign P[105] = in[29] ^ in2[29];
    assign G[106] = in[28] & in2[28];
    assign P[106] = in[28] ^ in2[28];
    assign G[107] = in[27] & in2[27];
    assign P[107] = in[27] ^ in2[27];
    assign G[108] = in[26] & in2[26];
    assign P[108] = in[26] ^ in2[26];
    assign G[109] = in[25] & in2[25];
    assign P[109] = in[25] ^ in2[25];
    assign G[110] = in[24] & in2[24];
    assign P[110] = in[24] ^ in2[24];
    assign G[111] = in[23] & in2[23];
    assign P[111] = in[23] ^ in2[23];
    assign G[112] = in[22] & in2[22];
    assign P[112] = in[22] ^ in2[22];
    assign G[113] = in[21] & in2[21];
    assign P[113] = in[21] ^ in2[21];
    assign G[114] = in[20] & in2[20];
    assign P[114] = in[20] ^ in2[20];
    assign G[115] = in[19] & in2[19];
    assign P[115] = in[19] ^ in2[19];
    assign G[116] = in[18] & in2[18];
    assign P[116] = in[18] ^ in2[18];
    assign G[117] = in[17] & in2[17];
    assign P[117] = in[17] ^ in2[17];
    assign G[118] = in[16] & in2[16];
    assign P[118] = in[16] ^ in2[16];
    assign G[119] = in[15] & in2[15];
    assign P[119] = in[15] ^ in2[15];
    assign G[120] = in[14] & in2[14];
    assign P[120] = in[14] ^ in2[14];
    assign G[121] = in[13] & in2[13];
    assign P[121] = in[13] ^ in2[13];
    assign G[122] = in[12] & in2[12];
    assign P[122] = in[12] ^ in2[12];
    assign G[123] = in[11] & in2[11];
    assign P[123] = in[11] ^ in2[11];
    assign G[124] = in[10] & in2[10];
    assign P[124] = in[10] ^ in2[10];
    assign G[125] = in[9] & in2[9];
    assign P[125] = in[9] ^ in2[9];
    assign G[126] = in[8] & in2[8];
    assign P[126] = in[8] ^ in2[8];
    assign G[127] = in[7] & in2[7];
    assign P[127] = in[7] ^ in2[7];
    assign G[128] = in[6] & in2[6];
    assign P[128] = in[6] ^ in2[6];
    assign G[129] = in[5] & in2[5];
    assign P[129] = in[5] ^ in2[5];
    assign G[130] = in[4] & in2[4];
    assign P[130] = in[4] ^ in2[4];
    assign G[131] = in[3] & in2[3];
    assign P[131] = in[3] ^ in2[3];
    assign G[132] = in[2] & in2[2];
    assign P[132] = in[2] ^ in2[2];
    assign G[133] = in[1] & in2[1];
    assign P[133] = in[1] ^ in2[1];
    assign G[134] = in[0] & in2[0];
    assign P[134] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign C[134] = G[133] | (P[133] & C[133]);
    assign cout = G[134] | (P[134] & C[134]);
    assign sum = P ^ C;
endmodule

module CLA134(output [133:0] sum, output cout, input [133:0] in1, input [133:0] in2;

    wire[133:0] G;
    wire[133:0] C;
    wire[133:0] P;

    assign G[0] = in[133] & in2[133];
    assign P[0] = in[133] ^ in2[133];
    assign G[1] = in[132] & in2[132];
    assign P[1] = in[132] ^ in2[132];
    assign G[2] = in[131] & in2[131];
    assign P[2] = in[131] ^ in2[131];
    assign G[3] = in[130] & in2[130];
    assign P[3] = in[130] ^ in2[130];
    assign G[4] = in[129] & in2[129];
    assign P[4] = in[129] ^ in2[129];
    assign G[5] = in[128] & in2[128];
    assign P[5] = in[128] ^ in2[128];
    assign G[6] = in[127] & in2[127];
    assign P[6] = in[127] ^ in2[127];
    assign G[7] = in[126] & in2[126];
    assign P[7] = in[126] ^ in2[126];
    assign G[8] = in[125] & in2[125];
    assign P[8] = in[125] ^ in2[125];
    assign G[9] = in[124] & in2[124];
    assign P[9] = in[124] ^ in2[124];
    assign G[10] = in[123] & in2[123];
    assign P[10] = in[123] ^ in2[123];
    assign G[11] = in[122] & in2[122];
    assign P[11] = in[122] ^ in2[122];
    assign G[12] = in[121] & in2[121];
    assign P[12] = in[121] ^ in2[121];
    assign G[13] = in[120] & in2[120];
    assign P[13] = in[120] ^ in2[120];
    assign G[14] = in[119] & in2[119];
    assign P[14] = in[119] ^ in2[119];
    assign G[15] = in[118] & in2[118];
    assign P[15] = in[118] ^ in2[118];
    assign G[16] = in[117] & in2[117];
    assign P[16] = in[117] ^ in2[117];
    assign G[17] = in[116] & in2[116];
    assign P[17] = in[116] ^ in2[116];
    assign G[18] = in[115] & in2[115];
    assign P[18] = in[115] ^ in2[115];
    assign G[19] = in[114] & in2[114];
    assign P[19] = in[114] ^ in2[114];
    assign G[20] = in[113] & in2[113];
    assign P[20] = in[113] ^ in2[113];
    assign G[21] = in[112] & in2[112];
    assign P[21] = in[112] ^ in2[112];
    assign G[22] = in[111] & in2[111];
    assign P[22] = in[111] ^ in2[111];
    assign G[23] = in[110] & in2[110];
    assign P[23] = in[110] ^ in2[110];
    assign G[24] = in[109] & in2[109];
    assign P[24] = in[109] ^ in2[109];
    assign G[25] = in[108] & in2[108];
    assign P[25] = in[108] ^ in2[108];
    assign G[26] = in[107] & in2[107];
    assign P[26] = in[107] ^ in2[107];
    assign G[27] = in[106] & in2[106];
    assign P[27] = in[106] ^ in2[106];
    assign G[28] = in[105] & in2[105];
    assign P[28] = in[105] ^ in2[105];
    assign G[29] = in[104] & in2[104];
    assign P[29] = in[104] ^ in2[104];
    assign G[30] = in[103] & in2[103];
    assign P[30] = in[103] ^ in2[103];
    assign G[31] = in[102] & in2[102];
    assign P[31] = in[102] ^ in2[102];
    assign G[32] = in[101] & in2[101];
    assign P[32] = in[101] ^ in2[101];
    assign G[33] = in[100] & in2[100];
    assign P[33] = in[100] ^ in2[100];
    assign G[34] = in[99] & in2[99];
    assign P[34] = in[99] ^ in2[99];
    assign G[35] = in[98] & in2[98];
    assign P[35] = in[98] ^ in2[98];
    assign G[36] = in[97] & in2[97];
    assign P[36] = in[97] ^ in2[97];
    assign G[37] = in[96] & in2[96];
    assign P[37] = in[96] ^ in2[96];
    assign G[38] = in[95] & in2[95];
    assign P[38] = in[95] ^ in2[95];
    assign G[39] = in[94] & in2[94];
    assign P[39] = in[94] ^ in2[94];
    assign G[40] = in[93] & in2[93];
    assign P[40] = in[93] ^ in2[93];
    assign G[41] = in[92] & in2[92];
    assign P[41] = in[92] ^ in2[92];
    assign G[42] = in[91] & in2[91];
    assign P[42] = in[91] ^ in2[91];
    assign G[43] = in[90] & in2[90];
    assign P[43] = in[90] ^ in2[90];
    assign G[44] = in[89] & in2[89];
    assign P[44] = in[89] ^ in2[89];
    assign G[45] = in[88] & in2[88];
    assign P[45] = in[88] ^ in2[88];
    assign G[46] = in[87] & in2[87];
    assign P[46] = in[87] ^ in2[87];
    assign G[47] = in[86] & in2[86];
    assign P[47] = in[86] ^ in2[86];
    assign G[48] = in[85] & in2[85];
    assign P[48] = in[85] ^ in2[85];
    assign G[49] = in[84] & in2[84];
    assign P[49] = in[84] ^ in2[84];
    assign G[50] = in[83] & in2[83];
    assign P[50] = in[83] ^ in2[83];
    assign G[51] = in[82] & in2[82];
    assign P[51] = in[82] ^ in2[82];
    assign G[52] = in[81] & in2[81];
    assign P[52] = in[81] ^ in2[81];
    assign G[53] = in[80] & in2[80];
    assign P[53] = in[80] ^ in2[80];
    assign G[54] = in[79] & in2[79];
    assign P[54] = in[79] ^ in2[79];
    assign G[55] = in[78] & in2[78];
    assign P[55] = in[78] ^ in2[78];
    assign G[56] = in[77] & in2[77];
    assign P[56] = in[77] ^ in2[77];
    assign G[57] = in[76] & in2[76];
    assign P[57] = in[76] ^ in2[76];
    assign G[58] = in[75] & in2[75];
    assign P[58] = in[75] ^ in2[75];
    assign G[59] = in[74] & in2[74];
    assign P[59] = in[74] ^ in2[74];
    assign G[60] = in[73] & in2[73];
    assign P[60] = in[73] ^ in2[73];
    assign G[61] = in[72] & in2[72];
    assign P[61] = in[72] ^ in2[72];
    assign G[62] = in[71] & in2[71];
    assign P[62] = in[71] ^ in2[71];
    assign G[63] = in[70] & in2[70];
    assign P[63] = in[70] ^ in2[70];
    assign G[64] = in[69] & in2[69];
    assign P[64] = in[69] ^ in2[69];
    assign G[65] = in[68] & in2[68];
    assign P[65] = in[68] ^ in2[68];
    assign G[66] = in[67] & in2[67];
    assign P[66] = in[67] ^ in2[67];
    assign G[67] = in[66] & in2[66];
    assign P[67] = in[66] ^ in2[66];
    assign G[68] = in[65] & in2[65];
    assign P[68] = in[65] ^ in2[65];
    assign G[69] = in[64] & in2[64];
    assign P[69] = in[64] ^ in2[64];
    assign G[70] = in[63] & in2[63];
    assign P[70] = in[63] ^ in2[63];
    assign G[71] = in[62] & in2[62];
    assign P[71] = in[62] ^ in2[62];
    assign G[72] = in[61] & in2[61];
    assign P[72] = in[61] ^ in2[61];
    assign G[73] = in[60] & in2[60];
    assign P[73] = in[60] ^ in2[60];
    assign G[74] = in[59] & in2[59];
    assign P[74] = in[59] ^ in2[59];
    assign G[75] = in[58] & in2[58];
    assign P[75] = in[58] ^ in2[58];
    assign G[76] = in[57] & in2[57];
    assign P[76] = in[57] ^ in2[57];
    assign G[77] = in[56] & in2[56];
    assign P[77] = in[56] ^ in2[56];
    assign G[78] = in[55] & in2[55];
    assign P[78] = in[55] ^ in2[55];
    assign G[79] = in[54] & in2[54];
    assign P[79] = in[54] ^ in2[54];
    assign G[80] = in[53] & in2[53];
    assign P[80] = in[53] ^ in2[53];
    assign G[81] = in[52] & in2[52];
    assign P[81] = in[52] ^ in2[52];
    assign G[82] = in[51] & in2[51];
    assign P[82] = in[51] ^ in2[51];
    assign G[83] = in[50] & in2[50];
    assign P[83] = in[50] ^ in2[50];
    assign G[84] = in[49] & in2[49];
    assign P[84] = in[49] ^ in2[49];
    assign G[85] = in[48] & in2[48];
    assign P[85] = in[48] ^ in2[48];
    assign G[86] = in[47] & in2[47];
    assign P[86] = in[47] ^ in2[47];
    assign G[87] = in[46] & in2[46];
    assign P[87] = in[46] ^ in2[46];
    assign G[88] = in[45] & in2[45];
    assign P[88] = in[45] ^ in2[45];
    assign G[89] = in[44] & in2[44];
    assign P[89] = in[44] ^ in2[44];
    assign G[90] = in[43] & in2[43];
    assign P[90] = in[43] ^ in2[43];
    assign G[91] = in[42] & in2[42];
    assign P[91] = in[42] ^ in2[42];
    assign G[92] = in[41] & in2[41];
    assign P[92] = in[41] ^ in2[41];
    assign G[93] = in[40] & in2[40];
    assign P[93] = in[40] ^ in2[40];
    assign G[94] = in[39] & in2[39];
    assign P[94] = in[39] ^ in2[39];
    assign G[95] = in[38] & in2[38];
    assign P[95] = in[38] ^ in2[38];
    assign G[96] = in[37] & in2[37];
    assign P[96] = in[37] ^ in2[37];
    assign G[97] = in[36] & in2[36];
    assign P[97] = in[36] ^ in2[36];
    assign G[98] = in[35] & in2[35];
    assign P[98] = in[35] ^ in2[35];
    assign G[99] = in[34] & in2[34];
    assign P[99] = in[34] ^ in2[34];
    assign G[100] = in[33] & in2[33];
    assign P[100] = in[33] ^ in2[33];
    assign G[101] = in[32] & in2[32];
    assign P[101] = in[32] ^ in2[32];
    assign G[102] = in[31] & in2[31];
    assign P[102] = in[31] ^ in2[31];
    assign G[103] = in[30] & in2[30];
    assign P[103] = in[30] ^ in2[30];
    assign G[104] = in[29] & in2[29];
    assign P[104] = in[29] ^ in2[29];
    assign G[105] = in[28] & in2[28];
    assign P[105] = in[28] ^ in2[28];
    assign G[106] = in[27] & in2[27];
    assign P[106] = in[27] ^ in2[27];
    assign G[107] = in[26] & in2[26];
    assign P[107] = in[26] ^ in2[26];
    assign G[108] = in[25] & in2[25];
    assign P[108] = in[25] ^ in2[25];
    assign G[109] = in[24] & in2[24];
    assign P[109] = in[24] ^ in2[24];
    assign G[110] = in[23] & in2[23];
    assign P[110] = in[23] ^ in2[23];
    assign G[111] = in[22] & in2[22];
    assign P[111] = in[22] ^ in2[22];
    assign G[112] = in[21] & in2[21];
    assign P[112] = in[21] ^ in2[21];
    assign G[113] = in[20] & in2[20];
    assign P[113] = in[20] ^ in2[20];
    assign G[114] = in[19] & in2[19];
    assign P[114] = in[19] ^ in2[19];
    assign G[115] = in[18] & in2[18];
    assign P[115] = in[18] ^ in2[18];
    assign G[116] = in[17] & in2[17];
    assign P[116] = in[17] ^ in2[17];
    assign G[117] = in[16] & in2[16];
    assign P[117] = in[16] ^ in2[16];
    assign G[118] = in[15] & in2[15];
    assign P[118] = in[15] ^ in2[15];
    assign G[119] = in[14] & in2[14];
    assign P[119] = in[14] ^ in2[14];
    assign G[120] = in[13] & in2[13];
    assign P[120] = in[13] ^ in2[13];
    assign G[121] = in[12] & in2[12];
    assign P[121] = in[12] ^ in2[12];
    assign G[122] = in[11] & in2[11];
    assign P[122] = in[11] ^ in2[11];
    assign G[123] = in[10] & in2[10];
    assign P[123] = in[10] ^ in2[10];
    assign G[124] = in[9] & in2[9];
    assign P[124] = in[9] ^ in2[9];
    assign G[125] = in[8] & in2[8];
    assign P[125] = in[8] ^ in2[8];
    assign G[126] = in[7] & in2[7];
    assign P[126] = in[7] ^ in2[7];
    assign G[127] = in[6] & in2[6];
    assign P[127] = in[6] ^ in2[6];
    assign G[128] = in[5] & in2[5];
    assign P[128] = in[5] ^ in2[5];
    assign G[129] = in[4] & in2[4];
    assign P[129] = in[4] ^ in2[4];
    assign G[130] = in[3] & in2[3];
    assign P[130] = in[3] ^ in2[3];
    assign G[131] = in[2] & in2[2];
    assign P[131] = in[2] ^ in2[2];
    assign G[132] = in[1] & in2[1];
    assign P[132] = in[1] ^ in2[1];
    assign G[133] = in[0] & in2[0];
    assign P[133] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign C[133] = G[132] | (P[132] & C[132]);
    assign cout = G[133] | (P[133] & C[133]);
    assign sum = P ^ C;
endmodule

module CLA133(output [132:0] sum, output cout, input [132:0] in1, input [132:0] in2;

    wire[132:0] G;
    wire[132:0] C;
    wire[132:0] P;

    assign G[0] = in[132] & in2[132];
    assign P[0] = in[132] ^ in2[132];
    assign G[1] = in[131] & in2[131];
    assign P[1] = in[131] ^ in2[131];
    assign G[2] = in[130] & in2[130];
    assign P[2] = in[130] ^ in2[130];
    assign G[3] = in[129] & in2[129];
    assign P[3] = in[129] ^ in2[129];
    assign G[4] = in[128] & in2[128];
    assign P[4] = in[128] ^ in2[128];
    assign G[5] = in[127] & in2[127];
    assign P[5] = in[127] ^ in2[127];
    assign G[6] = in[126] & in2[126];
    assign P[6] = in[126] ^ in2[126];
    assign G[7] = in[125] & in2[125];
    assign P[7] = in[125] ^ in2[125];
    assign G[8] = in[124] & in2[124];
    assign P[8] = in[124] ^ in2[124];
    assign G[9] = in[123] & in2[123];
    assign P[9] = in[123] ^ in2[123];
    assign G[10] = in[122] & in2[122];
    assign P[10] = in[122] ^ in2[122];
    assign G[11] = in[121] & in2[121];
    assign P[11] = in[121] ^ in2[121];
    assign G[12] = in[120] & in2[120];
    assign P[12] = in[120] ^ in2[120];
    assign G[13] = in[119] & in2[119];
    assign P[13] = in[119] ^ in2[119];
    assign G[14] = in[118] & in2[118];
    assign P[14] = in[118] ^ in2[118];
    assign G[15] = in[117] & in2[117];
    assign P[15] = in[117] ^ in2[117];
    assign G[16] = in[116] & in2[116];
    assign P[16] = in[116] ^ in2[116];
    assign G[17] = in[115] & in2[115];
    assign P[17] = in[115] ^ in2[115];
    assign G[18] = in[114] & in2[114];
    assign P[18] = in[114] ^ in2[114];
    assign G[19] = in[113] & in2[113];
    assign P[19] = in[113] ^ in2[113];
    assign G[20] = in[112] & in2[112];
    assign P[20] = in[112] ^ in2[112];
    assign G[21] = in[111] & in2[111];
    assign P[21] = in[111] ^ in2[111];
    assign G[22] = in[110] & in2[110];
    assign P[22] = in[110] ^ in2[110];
    assign G[23] = in[109] & in2[109];
    assign P[23] = in[109] ^ in2[109];
    assign G[24] = in[108] & in2[108];
    assign P[24] = in[108] ^ in2[108];
    assign G[25] = in[107] & in2[107];
    assign P[25] = in[107] ^ in2[107];
    assign G[26] = in[106] & in2[106];
    assign P[26] = in[106] ^ in2[106];
    assign G[27] = in[105] & in2[105];
    assign P[27] = in[105] ^ in2[105];
    assign G[28] = in[104] & in2[104];
    assign P[28] = in[104] ^ in2[104];
    assign G[29] = in[103] & in2[103];
    assign P[29] = in[103] ^ in2[103];
    assign G[30] = in[102] & in2[102];
    assign P[30] = in[102] ^ in2[102];
    assign G[31] = in[101] & in2[101];
    assign P[31] = in[101] ^ in2[101];
    assign G[32] = in[100] & in2[100];
    assign P[32] = in[100] ^ in2[100];
    assign G[33] = in[99] & in2[99];
    assign P[33] = in[99] ^ in2[99];
    assign G[34] = in[98] & in2[98];
    assign P[34] = in[98] ^ in2[98];
    assign G[35] = in[97] & in2[97];
    assign P[35] = in[97] ^ in2[97];
    assign G[36] = in[96] & in2[96];
    assign P[36] = in[96] ^ in2[96];
    assign G[37] = in[95] & in2[95];
    assign P[37] = in[95] ^ in2[95];
    assign G[38] = in[94] & in2[94];
    assign P[38] = in[94] ^ in2[94];
    assign G[39] = in[93] & in2[93];
    assign P[39] = in[93] ^ in2[93];
    assign G[40] = in[92] & in2[92];
    assign P[40] = in[92] ^ in2[92];
    assign G[41] = in[91] & in2[91];
    assign P[41] = in[91] ^ in2[91];
    assign G[42] = in[90] & in2[90];
    assign P[42] = in[90] ^ in2[90];
    assign G[43] = in[89] & in2[89];
    assign P[43] = in[89] ^ in2[89];
    assign G[44] = in[88] & in2[88];
    assign P[44] = in[88] ^ in2[88];
    assign G[45] = in[87] & in2[87];
    assign P[45] = in[87] ^ in2[87];
    assign G[46] = in[86] & in2[86];
    assign P[46] = in[86] ^ in2[86];
    assign G[47] = in[85] & in2[85];
    assign P[47] = in[85] ^ in2[85];
    assign G[48] = in[84] & in2[84];
    assign P[48] = in[84] ^ in2[84];
    assign G[49] = in[83] & in2[83];
    assign P[49] = in[83] ^ in2[83];
    assign G[50] = in[82] & in2[82];
    assign P[50] = in[82] ^ in2[82];
    assign G[51] = in[81] & in2[81];
    assign P[51] = in[81] ^ in2[81];
    assign G[52] = in[80] & in2[80];
    assign P[52] = in[80] ^ in2[80];
    assign G[53] = in[79] & in2[79];
    assign P[53] = in[79] ^ in2[79];
    assign G[54] = in[78] & in2[78];
    assign P[54] = in[78] ^ in2[78];
    assign G[55] = in[77] & in2[77];
    assign P[55] = in[77] ^ in2[77];
    assign G[56] = in[76] & in2[76];
    assign P[56] = in[76] ^ in2[76];
    assign G[57] = in[75] & in2[75];
    assign P[57] = in[75] ^ in2[75];
    assign G[58] = in[74] & in2[74];
    assign P[58] = in[74] ^ in2[74];
    assign G[59] = in[73] & in2[73];
    assign P[59] = in[73] ^ in2[73];
    assign G[60] = in[72] & in2[72];
    assign P[60] = in[72] ^ in2[72];
    assign G[61] = in[71] & in2[71];
    assign P[61] = in[71] ^ in2[71];
    assign G[62] = in[70] & in2[70];
    assign P[62] = in[70] ^ in2[70];
    assign G[63] = in[69] & in2[69];
    assign P[63] = in[69] ^ in2[69];
    assign G[64] = in[68] & in2[68];
    assign P[64] = in[68] ^ in2[68];
    assign G[65] = in[67] & in2[67];
    assign P[65] = in[67] ^ in2[67];
    assign G[66] = in[66] & in2[66];
    assign P[66] = in[66] ^ in2[66];
    assign G[67] = in[65] & in2[65];
    assign P[67] = in[65] ^ in2[65];
    assign G[68] = in[64] & in2[64];
    assign P[68] = in[64] ^ in2[64];
    assign G[69] = in[63] & in2[63];
    assign P[69] = in[63] ^ in2[63];
    assign G[70] = in[62] & in2[62];
    assign P[70] = in[62] ^ in2[62];
    assign G[71] = in[61] & in2[61];
    assign P[71] = in[61] ^ in2[61];
    assign G[72] = in[60] & in2[60];
    assign P[72] = in[60] ^ in2[60];
    assign G[73] = in[59] & in2[59];
    assign P[73] = in[59] ^ in2[59];
    assign G[74] = in[58] & in2[58];
    assign P[74] = in[58] ^ in2[58];
    assign G[75] = in[57] & in2[57];
    assign P[75] = in[57] ^ in2[57];
    assign G[76] = in[56] & in2[56];
    assign P[76] = in[56] ^ in2[56];
    assign G[77] = in[55] & in2[55];
    assign P[77] = in[55] ^ in2[55];
    assign G[78] = in[54] & in2[54];
    assign P[78] = in[54] ^ in2[54];
    assign G[79] = in[53] & in2[53];
    assign P[79] = in[53] ^ in2[53];
    assign G[80] = in[52] & in2[52];
    assign P[80] = in[52] ^ in2[52];
    assign G[81] = in[51] & in2[51];
    assign P[81] = in[51] ^ in2[51];
    assign G[82] = in[50] & in2[50];
    assign P[82] = in[50] ^ in2[50];
    assign G[83] = in[49] & in2[49];
    assign P[83] = in[49] ^ in2[49];
    assign G[84] = in[48] & in2[48];
    assign P[84] = in[48] ^ in2[48];
    assign G[85] = in[47] & in2[47];
    assign P[85] = in[47] ^ in2[47];
    assign G[86] = in[46] & in2[46];
    assign P[86] = in[46] ^ in2[46];
    assign G[87] = in[45] & in2[45];
    assign P[87] = in[45] ^ in2[45];
    assign G[88] = in[44] & in2[44];
    assign P[88] = in[44] ^ in2[44];
    assign G[89] = in[43] & in2[43];
    assign P[89] = in[43] ^ in2[43];
    assign G[90] = in[42] & in2[42];
    assign P[90] = in[42] ^ in2[42];
    assign G[91] = in[41] & in2[41];
    assign P[91] = in[41] ^ in2[41];
    assign G[92] = in[40] & in2[40];
    assign P[92] = in[40] ^ in2[40];
    assign G[93] = in[39] & in2[39];
    assign P[93] = in[39] ^ in2[39];
    assign G[94] = in[38] & in2[38];
    assign P[94] = in[38] ^ in2[38];
    assign G[95] = in[37] & in2[37];
    assign P[95] = in[37] ^ in2[37];
    assign G[96] = in[36] & in2[36];
    assign P[96] = in[36] ^ in2[36];
    assign G[97] = in[35] & in2[35];
    assign P[97] = in[35] ^ in2[35];
    assign G[98] = in[34] & in2[34];
    assign P[98] = in[34] ^ in2[34];
    assign G[99] = in[33] & in2[33];
    assign P[99] = in[33] ^ in2[33];
    assign G[100] = in[32] & in2[32];
    assign P[100] = in[32] ^ in2[32];
    assign G[101] = in[31] & in2[31];
    assign P[101] = in[31] ^ in2[31];
    assign G[102] = in[30] & in2[30];
    assign P[102] = in[30] ^ in2[30];
    assign G[103] = in[29] & in2[29];
    assign P[103] = in[29] ^ in2[29];
    assign G[104] = in[28] & in2[28];
    assign P[104] = in[28] ^ in2[28];
    assign G[105] = in[27] & in2[27];
    assign P[105] = in[27] ^ in2[27];
    assign G[106] = in[26] & in2[26];
    assign P[106] = in[26] ^ in2[26];
    assign G[107] = in[25] & in2[25];
    assign P[107] = in[25] ^ in2[25];
    assign G[108] = in[24] & in2[24];
    assign P[108] = in[24] ^ in2[24];
    assign G[109] = in[23] & in2[23];
    assign P[109] = in[23] ^ in2[23];
    assign G[110] = in[22] & in2[22];
    assign P[110] = in[22] ^ in2[22];
    assign G[111] = in[21] & in2[21];
    assign P[111] = in[21] ^ in2[21];
    assign G[112] = in[20] & in2[20];
    assign P[112] = in[20] ^ in2[20];
    assign G[113] = in[19] & in2[19];
    assign P[113] = in[19] ^ in2[19];
    assign G[114] = in[18] & in2[18];
    assign P[114] = in[18] ^ in2[18];
    assign G[115] = in[17] & in2[17];
    assign P[115] = in[17] ^ in2[17];
    assign G[116] = in[16] & in2[16];
    assign P[116] = in[16] ^ in2[16];
    assign G[117] = in[15] & in2[15];
    assign P[117] = in[15] ^ in2[15];
    assign G[118] = in[14] & in2[14];
    assign P[118] = in[14] ^ in2[14];
    assign G[119] = in[13] & in2[13];
    assign P[119] = in[13] ^ in2[13];
    assign G[120] = in[12] & in2[12];
    assign P[120] = in[12] ^ in2[12];
    assign G[121] = in[11] & in2[11];
    assign P[121] = in[11] ^ in2[11];
    assign G[122] = in[10] & in2[10];
    assign P[122] = in[10] ^ in2[10];
    assign G[123] = in[9] & in2[9];
    assign P[123] = in[9] ^ in2[9];
    assign G[124] = in[8] & in2[8];
    assign P[124] = in[8] ^ in2[8];
    assign G[125] = in[7] & in2[7];
    assign P[125] = in[7] ^ in2[7];
    assign G[126] = in[6] & in2[6];
    assign P[126] = in[6] ^ in2[6];
    assign G[127] = in[5] & in2[5];
    assign P[127] = in[5] ^ in2[5];
    assign G[128] = in[4] & in2[4];
    assign P[128] = in[4] ^ in2[4];
    assign G[129] = in[3] & in2[3];
    assign P[129] = in[3] ^ in2[3];
    assign G[130] = in[2] & in2[2];
    assign P[130] = in[2] ^ in2[2];
    assign G[131] = in[1] & in2[1];
    assign P[131] = in[1] ^ in2[1];
    assign G[132] = in[0] & in2[0];
    assign P[132] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign C[132] = G[131] | (P[131] & C[131]);
    assign cout = G[132] | (P[132] & C[132]);
    assign sum = P ^ C;
endmodule

module CLA132(output [131:0] sum, output cout, input [131:0] in1, input [131:0] in2;

    wire[131:0] G;
    wire[131:0] C;
    wire[131:0] P;

    assign G[0] = in[131] & in2[131];
    assign P[0] = in[131] ^ in2[131];
    assign G[1] = in[130] & in2[130];
    assign P[1] = in[130] ^ in2[130];
    assign G[2] = in[129] & in2[129];
    assign P[2] = in[129] ^ in2[129];
    assign G[3] = in[128] & in2[128];
    assign P[3] = in[128] ^ in2[128];
    assign G[4] = in[127] & in2[127];
    assign P[4] = in[127] ^ in2[127];
    assign G[5] = in[126] & in2[126];
    assign P[5] = in[126] ^ in2[126];
    assign G[6] = in[125] & in2[125];
    assign P[6] = in[125] ^ in2[125];
    assign G[7] = in[124] & in2[124];
    assign P[7] = in[124] ^ in2[124];
    assign G[8] = in[123] & in2[123];
    assign P[8] = in[123] ^ in2[123];
    assign G[9] = in[122] & in2[122];
    assign P[9] = in[122] ^ in2[122];
    assign G[10] = in[121] & in2[121];
    assign P[10] = in[121] ^ in2[121];
    assign G[11] = in[120] & in2[120];
    assign P[11] = in[120] ^ in2[120];
    assign G[12] = in[119] & in2[119];
    assign P[12] = in[119] ^ in2[119];
    assign G[13] = in[118] & in2[118];
    assign P[13] = in[118] ^ in2[118];
    assign G[14] = in[117] & in2[117];
    assign P[14] = in[117] ^ in2[117];
    assign G[15] = in[116] & in2[116];
    assign P[15] = in[116] ^ in2[116];
    assign G[16] = in[115] & in2[115];
    assign P[16] = in[115] ^ in2[115];
    assign G[17] = in[114] & in2[114];
    assign P[17] = in[114] ^ in2[114];
    assign G[18] = in[113] & in2[113];
    assign P[18] = in[113] ^ in2[113];
    assign G[19] = in[112] & in2[112];
    assign P[19] = in[112] ^ in2[112];
    assign G[20] = in[111] & in2[111];
    assign P[20] = in[111] ^ in2[111];
    assign G[21] = in[110] & in2[110];
    assign P[21] = in[110] ^ in2[110];
    assign G[22] = in[109] & in2[109];
    assign P[22] = in[109] ^ in2[109];
    assign G[23] = in[108] & in2[108];
    assign P[23] = in[108] ^ in2[108];
    assign G[24] = in[107] & in2[107];
    assign P[24] = in[107] ^ in2[107];
    assign G[25] = in[106] & in2[106];
    assign P[25] = in[106] ^ in2[106];
    assign G[26] = in[105] & in2[105];
    assign P[26] = in[105] ^ in2[105];
    assign G[27] = in[104] & in2[104];
    assign P[27] = in[104] ^ in2[104];
    assign G[28] = in[103] & in2[103];
    assign P[28] = in[103] ^ in2[103];
    assign G[29] = in[102] & in2[102];
    assign P[29] = in[102] ^ in2[102];
    assign G[30] = in[101] & in2[101];
    assign P[30] = in[101] ^ in2[101];
    assign G[31] = in[100] & in2[100];
    assign P[31] = in[100] ^ in2[100];
    assign G[32] = in[99] & in2[99];
    assign P[32] = in[99] ^ in2[99];
    assign G[33] = in[98] & in2[98];
    assign P[33] = in[98] ^ in2[98];
    assign G[34] = in[97] & in2[97];
    assign P[34] = in[97] ^ in2[97];
    assign G[35] = in[96] & in2[96];
    assign P[35] = in[96] ^ in2[96];
    assign G[36] = in[95] & in2[95];
    assign P[36] = in[95] ^ in2[95];
    assign G[37] = in[94] & in2[94];
    assign P[37] = in[94] ^ in2[94];
    assign G[38] = in[93] & in2[93];
    assign P[38] = in[93] ^ in2[93];
    assign G[39] = in[92] & in2[92];
    assign P[39] = in[92] ^ in2[92];
    assign G[40] = in[91] & in2[91];
    assign P[40] = in[91] ^ in2[91];
    assign G[41] = in[90] & in2[90];
    assign P[41] = in[90] ^ in2[90];
    assign G[42] = in[89] & in2[89];
    assign P[42] = in[89] ^ in2[89];
    assign G[43] = in[88] & in2[88];
    assign P[43] = in[88] ^ in2[88];
    assign G[44] = in[87] & in2[87];
    assign P[44] = in[87] ^ in2[87];
    assign G[45] = in[86] & in2[86];
    assign P[45] = in[86] ^ in2[86];
    assign G[46] = in[85] & in2[85];
    assign P[46] = in[85] ^ in2[85];
    assign G[47] = in[84] & in2[84];
    assign P[47] = in[84] ^ in2[84];
    assign G[48] = in[83] & in2[83];
    assign P[48] = in[83] ^ in2[83];
    assign G[49] = in[82] & in2[82];
    assign P[49] = in[82] ^ in2[82];
    assign G[50] = in[81] & in2[81];
    assign P[50] = in[81] ^ in2[81];
    assign G[51] = in[80] & in2[80];
    assign P[51] = in[80] ^ in2[80];
    assign G[52] = in[79] & in2[79];
    assign P[52] = in[79] ^ in2[79];
    assign G[53] = in[78] & in2[78];
    assign P[53] = in[78] ^ in2[78];
    assign G[54] = in[77] & in2[77];
    assign P[54] = in[77] ^ in2[77];
    assign G[55] = in[76] & in2[76];
    assign P[55] = in[76] ^ in2[76];
    assign G[56] = in[75] & in2[75];
    assign P[56] = in[75] ^ in2[75];
    assign G[57] = in[74] & in2[74];
    assign P[57] = in[74] ^ in2[74];
    assign G[58] = in[73] & in2[73];
    assign P[58] = in[73] ^ in2[73];
    assign G[59] = in[72] & in2[72];
    assign P[59] = in[72] ^ in2[72];
    assign G[60] = in[71] & in2[71];
    assign P[60] = in[71] ^ in2[71];
    assign G[61] = in[70] & in2[70];
    assign P[61] = in[70] ^ in2[70];
    assign G[62] = in[69] & in2[69];
    assign P[62] = in[69] ^ in2[69];
    assign G[63] = in[68] & in2[68];
    assign P[63] = in[68] ^ in2[68];
    assign G[64] = in[67] & in2[67];
    assign P[64] = in[67] ^ in2[67];
    assign G[65] = in[66] & in2[66];
    assign P[65] = in[66] ^ in2[66];
    assign G[66] = in[65] & in2[65];
    assign P[66] = in[65] ^ in2[65];
    assign G[67] = in[64] & in2[64];
    assign P[67] = in[64] ^ in2[64];
    assign G[68] = in[63] & in2[63];
    assign P[68] = in[63] ^ in2[63];
    assign G[69] = in[62] & in2[62];
    assign P[69] = in[62] ^ in2[62];
    assign G[70] = in[61] & in2[61];
    assign P[70] = in[61] ^ in2[61];
    assign G[71] = in[60] & in2[60];
    assign P[71] = in[60] ^ in2[60];
    assign G[72] = in[59] & in2[59];
    assign P[72] = in[59] ^ in2[59];
    assign G[73] = in[58] & in2[58];
    assign P[73] = in[58] ^ in2[58];
    assign G[74] = in[57] & in2[57];
    assign P[74] = in[57] ^ in2[57];
    assign G[75] = in[56] & in2[56];
    assign P[75] = in[56] ^ in2[56];
    assign G[76] = in[55] & in2[55];
    assign P[76] = in[55] ^ in2[55];
    assign G[77] = in[54] & in2[54];
    assign P[77] = in[54] ^ in2[54];
    assign G[78] = in[53] & in2[53];
    assign P[78] = in[53] ^ in2[53];
    assign G[79] = in[52] & in2[52];
    assign P[79] = in[52] ^ in2[52];
    assign G[80] = in[51] & in2[51];
    assign P[80] = in[51] ^ in2[51];
    assign G[81] = in[50] & in2[50];
    assign P[81] = in[50] ^ in2[50];
    assign G[82] = in[49] & in2[49];
    assign P[82] = in[49] ^ in2[49];
    assign G[83] = in[48] & in2[48];
    assign P[83] = in[48] ^ in2[48];
    assign G[84] = in[47] & in2[47];
    assign P[84] = in[47] ^ in2[47];
    assign G[85] = in[46] & in2[46];
    assign P[85] = in[46] ^ in2[46];
    assign G[86] = in[45] & in2[45];
    assign P[86] = in[45] ^ in2[45];
    assign G[87] = in[44] & in2[44];
    assign P[87] = in[44] ^ in2[44];
    assign G[88] = in[43] & in2[43];
    assign P[88] = in[43] ^ in2[43];
    assign G[89] = in[42] & in2[42];
    assign P[89] = in[42] ^ in2[42];
    assign G[90] = in[41] & in2[41];
    assign P[90] = in[41] ^ in2[41];
    assign G[91] = in[40] & in2[40];
    assign P[91] = in[40] ^ in2[40];
    assign G[92] = in[39] & in2[39];
    assign P[92] = in[39] ^ in2[39];
    assign G[93] = in[38] & in2[38];
    assign P[93] = in[38] ^ in2[38];
    assign G[94] = in[37] & in2[37];
    assign P[94] = in[37] ^ in2[37];
    assign G[95] = in[36] & in2[36];
    assign P[95] = in[36] ^ in2[36];
    assign G[96] = in[35] & in2[35];
    assign P[96] = in[35] ^ in2[35];
    assign G[97] = in[34] & in2[34];
    assign P[97] = in[34] ^ in2[34];
    assign G[98] = in[33] & in2[33];
    assign P[98] = in[33] ^ in2[33];
    assign G[99] = in[32] & in2[32];
    assign P[99] = in[32] ^ in2[32];
    assign G[100] = in[31] & in2[31];
    assign P[100] = in[31] ^ in2[31];
    assign G[101] = in[30] & in2[30];
    assign P[101] = in[30] ^ in2[30];
    assign G[102] = in[29] & in2[29];
    assign P[102] = in[29] ^ in2[29];
    assign G[103] = in[28] & in2[28];
    assign P[103] = in[28] ^ in2[28];
    assign G[104] = in[27] & in2[27];
    assign P[104] = in[27] ^ in2[27];
    assign G[105] = in[26] & in2[26];
    assign P[105] = in[26] ^ in2[26];
    assign G[106] = in[25] & in2[25];
    assign P[106] = in[25] ^ in2[25];
    assign G[107] = in[24] & in2[24];
    assign P[107] = in[24] ^ in2[24];
    assign G[108] = in[23] & in2[23];
    assign P[108] = in[23] ^ in2[23];
    assign G[109] = in[22] & in2[22];
    assign P[109] = in[22] ^ in2[22];
    assign G[110] = in[21] & in2[21];
    assign P[110] = in[21] ^ in2[21];
    assign G[111] = in[20] & in2[20];
    assign P[111] = in[20] ^ in2[20];
    assign G[112] = in[19] & in2[19];
    assign P[112] = in[19] ^ in2[19];
    assign G[113] = in[18] & in2[18];
    assign P[113] = in[18] ^ in2[18];
    assign G[114] = in[17] & in2[17];
    assign P[114] = in[17] ^ in2[17];
    assign G[115] = in[16] & in2[16];
    assign P[115] = in[16] ^ in2[16];
    assign G[116] = in[15] & in2[15];
    assign P[116] = in[15] ^ in2[15];
    assign G[117] = in[14] & in2[14];
    assign P[117] = in[14] ^ in2[14];
    assign G[118] = in[13] & in2[13];
    assign P[118] = in[13] ^ in2[13];
    assign G[119] = in[12] & in2[12];
    assign P[119] = in[12] ^ in2[12];
    assign G[120] = in[11] & in2[11];
    assign P[120] = in[11] ^ in2[11];
    assign G[121] = in[10] & in2[10];
    assign P[121] = in[10] ^ in2[10];
    assign G[122] = in[9] & in2[9];
    assign P[122] = in[9] ^ in2[9];
    assign G[123] = in[8] & in2[8];
    assign P[123] = in[8] ^ in2[8];
    assign G[124] = in[7] & in2[7];
    assign P[124] = in[7] ^ in2[7];
    assign G[125] = in[6] & in2[6];
    assign P[125] = in[6] ^ in2[6];
    assign G[126] = in[5] & in2[5];
    assign P[126] = in[5] ^ in2[5];
    assign G[127] = in[4] & in2[4];
    assign P[127] = in[4] ^ in2[4];
    assign G[128] = in[3] & in2[3];
    assign P[128] = in[3] ^ in2[3];
    assign G[129] = in[2] & in2[2];
    assign P[129] = in[2] ^ in2[2];
    assign G[130] = in[1] & in2[1];
    assign P[130] = in[1] ^ in2[1];
    assign G[131] = in[0] & in2[0];
    assign P[131] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign C[131] = G[130] | (P[130] & C[130]);
    assign cout = G[131] | (P[131] & C[131]);
    assign sum = P ^ C;
endmodule

module CLA131(output [130:0] sum, output cout, input [130:0] in1, input [130:0] in2;

    wire[130:0] G;
    wire[130:0] C;
    wire[130:0] P;

    assign G[0] = in[130] & in2[130];
    assign P[0] = in[130] ^ in2[130];
    assign G[1] = in[129] & in2[129];
    assign P[1] = in[129] ^ in2[129];
    assign G[2] = in[128] & in2[128];
    assign P[2] = in[128] ^ in2[128];
    assign G[3] = in[127] & in2[127];
    assign P[3] = in[127] ^ in2[127];
    assign G[4] = in[126] & in2[126];
    assign P[4] = in[126] ^ in2[126];
    assign G[5] = in[125] & in2[125];
    assign P[5] = in[125] ^ in2[125];
    assign G[6] = in[124] & in2[124];
    assign P[6] = in[124] ^ in2[124];
    assign G[7] = in[123] & in2[123];
    assign P[7] = in[123] ^ in2[123];
    assign G[8] = in[122] & in2[122];
    assign P[8] = in[122] ^ in2[122];
    assign G[9] = in[121] & in2[121];
    assign P[9] = in[121] ^ in2[121];
    assign G[10] = in[120] & in2[120];
    assign P[10] = in[120] ^ in2[120];
    assign G[11] = in[119] & in2[119];
    assign P[11] = in[119] ^ in2[119];
    assign G[12] = in[118] & in2[118];
    assign P[12] = in[118] ^ in2[118];
    assign G[13] = in[117] & in2[117];
    assign P[13] = in[117] ^ in2[117];
    assign G[14] = in[116] & in2[116];
    assign P[14] = in[116] ^ in2[116];
    assign G[15] = in[115] & in2[115];
    assign P[15] = in[115] ^ in2[115];
    assign G[16] = in[114] & in2[114];
    assign P[16] = in[114] ^ in2[114];
    assign G[17] = in[113] & in2[113];
    assign P[17] = in[113] ^ in2[113];
    assign G[18] = in[112] & in2[112];
    assign P[18] = in[112] ^ in2[112];
    assign G[19] = in[111] & in2[111];
    assign P[19] = in[111] ^ in2[111];
    assign G[20] = in[110] & in2[110];
    assign P[20] = in[110] ^ in2[110];
    assign G[21] = in[109] & in2[109];
    assign P[21] = in[109] ^ in2[109];
    assign G[22] = in[108] & in2[108];
    assign P[22] = in[108] ^ in2[108];
    assign G[23] = in[107] & in2[107];
    assign P[23] = in[107] ^ in2[107];
    assign G[24] = in[106] & in2[106];
    assign P[24] = in[106] ^ in2[106];
    assign G[25] = in[105] & in2[105];
    assign P[25] = in[105] ^ in2[105];
    assign G[26] = in[104] & in2[104];
    assign P[26] = in[104] ^ in2[104];
    assign G[27] = in[103] & in2[103];
    assign P[27] = in[103] ^ in2[103];
    assign G[28] = in[102] & in2[102];
    assign P[28] = in[102] ^ in2[102];
    assign G[29] = in[101] & in2[101];
    assign P[29] = in[101] ^ in2[101];
    assign G[30] = in[100] & in2[100];
    assign P[30] = in[100] ^ in2[100];
    assign G[31] = in[99] & in2[99];
    assign P[31] = in[99] ^ in2[99];
    assign G[32] = in[98] & in2[98];
    assign P[32] = in[98] ^ in2[98];
    assign G[33] = in[97] & in2[97];
    assign P[33] = in[97] ^ in2[97];
    assign G[34] = in[96] & in2[96];
    assign P[34] = in[96] ^ in2[96];
    assign G[35] = in[95] & in2[95];
    assign P[35] = in[95] ^ in2[95];
    assign G[36] = in[94] & in2[94];
    assign P[36] = in[94] ^ in2[94];
    assign G[37] = in[93] & in2[93];
    assign P[37] = in[93] ^ in2[93];
    assign G[38] = in[92] & in2[92];
    assign P[38] = in[92] ^ in2[92];
    assign G[39] = in[91] & in2[91];
    assign P[39] = in[91] ^ in2[91];
    assign G[40] = in[90] & in2[90];
    assign P[40] = in[90] ^ in2[90];
    assign G[41] = in[89] & in2[89];
    assign P[41] = in[89] ^ in2[89];
    assign G[42] = in[88] & in2[88];
    assign P[42] = in[88] ^ in2[88];
    assign G[43] = in[87] & in2[87];
    assign P[43] = in[87] ^ in2[87];
    assign G[44] = in[86] & in2[86];
    assign P[44] = in[86] ^ in2[86];
    assign G[45] = in[85] & in2[85];
    assign P[45] = in[85] ^ in2[85];
    assign G[46] = in[84] & in2[84];
    assign P[46] = in[84] ^ in2[84];
    assign G[47] = in[83] & in2[83];
    assign P[47] = in[83] ^ in2[83];
    assign G[48] = in[82] & in2[82];
    assign P[48] = in[82] ^ in2[82];
    assign G[49] = in[81] & in2[81];
    assign P[49] = in[81] ^ in2[81];
    assign G[50] = in[80] & in2[80];
    assign P[50] = in[80] ^ in2[80];
    assign G[51] = in[79] & in2[79];
    assign P[51] = in[79] ^ in2[79];
    assign G[52] = in[78] & in2[78];
    assign P[52] = in[78] ^ in2[78];
    assign G[53] = in[77] & in2[77];
    assign P[53] = in[77] ^ in2[77];
    assign G[54] = in[76] & in2[76];
    assign P[54] = in[76] ^ in2[76];
    assign G[55] = in[75] & in2[75];
    assign P[55] = in[75] ^ in2[75];
    assign G[56] = in[74] & in2[74];
    assign P[56] = in[74] ^ in2[74];
    assign G[57] = in[73] & in2[73];
    assign P[57] = in[73] ^ in2[73];
    assign G[58] = in[72] & in2[72];
    assign P[58] = in[72] ^ in2[72];
    assign G[59] = in[71] & in2[71];
    assign P[59] = in[71] ^ in2[71];
    assign G[60] = in[70] & in2[70];
    assign P[60] = in[70] ^ in2[70];
    assign G[61] = in[69] & in2[69];
    assign P[61] = in[69] ^ in2[69];
    assign G[62] = in[68] & in2[68];
    assign P[62] = in[68] ^ in2[68];
    assign G[63] = in[67] & in2[67];
    assign P[63] = in[67] ^ in2[67];
    assign G[64] = in[66] & in2[66];
    assign P[64] = in[66] ^ in2[66];
    assign G[65] = in[65] & in2[65];
    assign P[65] = in[65] ^ in2[65];
    assign G[66] = in[64] & in2[64];
    assign P[66] = in[64] ^ in2[64];
    assign G[67] = in[63] & in2[63];
    assign P[67] = in[63] ^ in2[63];
    assign G[68] = in[62] & in2[62];
    assign P[68] = in[62] ^ in2[62];
    assign G[69] = in[61] & in2[61];
    assign P[69] = in[61] ^ in2[61];
    assign G[70] = in[60] & in2[60];
    assign P[70] = in[60] ^ in2[60];
    assign G[71] = in[59] & in2[59];
    assign P[71] = in[59] ^ in2[59];
    assign G[72] = in[58] & in2[58];
    assign P[72] = in[58] ^ in2[58];
    assign G[73] = in[57] & in2[57];
    assign P[73] = in[57] ^ in2[57];
    assign G[74] = in[56] & in2[56];
    assign P[74] = in[56] ^ in2[56];
    assign G[75] = in[55] & in2[55];
    assign P[75] = in[55] ^ in2[55];
    assign G[76] = in[54] & in2[54];
    assign P[76] = in[54] ^ in2[54];
    assign G[77] = in[53] & in2[53];
    assign P[77] = in[53] ^ in2[53];
    assign G[78] = in[52] & in2[52];
    assign P[78] = in[52] ^ in2[52];
    assign G[79] = in[51] & in2[51];
    assign P[79] = in[51] ^ in2[51];
    assign G[80] = in[50] & in2[50];
    assign P[80] = in[50] ^ in2[50];
    assign G[81] = in[49] & in2[49];
    assign P[81] = in[49] ^ in2[49];
    assign G[82] = in[48] & in2[48];
    assign P[82] = in[48] ^ in2[48];
    assign G[83] = in[47] & in2[47];
    assign P[83] = in[47] ^ in2[47];
    assign G[84] = in[46] & in2[46];
    assign P[84] = in[46] ^ in2[46];
    assign G[85] = in[45] & in2[45];
    assign P[85] = in[45] ^ in2[45];
    assign G[86] = in[44] & in2[44];
    assign P[86] = in[44] ^ in2[44];
    assign G[87] = in[43] & in2[43];
    assign P[87] = in[43] ^ in2[43];
    assign G[88] = in[42] & in2[42];
    assign P[88] = in[42] ^ in2[42];
    assign G[89] = in[41] & in2[41];
    assign P[89] = in[41] ^ in2[41];
    assign G[90] = in[40] & in2[40];
    assign P[90] = in[40] ^ in2[40];
    assign G[91] = in[39] & in2[39];
    assign P[91] = in[39] ^ in2[39];
    assign G[92] = in[38] & in2[38];
    assign P[92] = in[38] ^ in2[38];
    assign G[93] = in[37] & in2[37];
    assign P[93] = in[37] ^ in2[37];
    assign G[94] = in[36] & in2[36];
    assign P[94] = in[36] ^ in2[36];
    assign G[95] = in[35] & in2[35];
    assign P[95] = in[35] ^ in2[35];
    assign G[96] = in[34] & in2[34];
    assign P[96] = in[34] ^ in2[34];
    assign G[97] = in[33] & in2[33];
    assign P[97] = in[33] ^ in2[33];
    assign G[98] = in[32] & in2[32];
    assign P[98] = in[32] ^ in2[32];
    assign G[99] = in[31] & in2[31];
    assign P[99] = in[31] ^ in2[31];
    assign G[100] = in[30] & in2[30];
    assign P[100] = in[30] ^ in2[30];
    assign G[101] = in[29] & in2[29];
    assign P[101] = in[29] ^ in2[29];
    assign G[102] = in[28] & in2[28];
    assign P[102] = in[28] ^ in2[28];
    assign G[103] = in[27] & in2[27];
    assign P[103] = in[27] ^ in2[27];
    assign G[104] = in[26] & in2[26];
    assign P[104] = in[26] ^ in2[26];
    assign G[105] = in[25] & in2[25];
    assign P[105] = in[25] ^ in2[25];
    assign G[106] = in[24] & in2[24];
    assign P[106] = in[24] ^ in2[24];
    assign G[107] = in[23] & in2[23];
    assign P[107] = in[23] ^ in2[23];
    assign G[108] = in[22] & in2[22];
    assign P[108] = in[22] ^ in2[22];
    assign G[109] = in[21] & in2[21];
    assign P[109] = in[21] ^ in2[21];
    assign G[110] = in[20] & in2[20];
    assign P[110] = in[20] ^ in2[20];
    assign G[111] = in[19] & in2[19];
    assign P[111] = in[19] ^ in2[19];
    assign G[112] = in[18] & in2[18];
    assign P[112] = in[18] ^ in2[18];
    assign G[113] = in[17] & in2[17];
    assign P[113] = in[17] ^ in2[17];
    assign G[114] = in[16] & in2[16];
    assign P[114] = in[16] ^ in2[16];
    assign G[115] = in[15] & in2[15];
    assign P[115] = in[15] ^ in2[15];
    assign G[116] = in[14] & in2[14];
    assign P[116] = in[14] ^ in2[14];
    assign G[117] = in[13] & in2[13];
    assign P[117] = in[13] ^ in2[13];
    assign G[118] = in[12] & in2[12];
    assign P[118] = in[12] ^ in2[12];
    assign G[119] = in[11] & in2[11];
    assign P[119] = in[11] ^ in2[11];
    assign G[120] = in[10] & in2[10];
    assign P[120] = in[10] ^ in2[10];
    assign G[121] = in[9] & in2[9];
    assign P[121] = in[9] ^ in2[9];
    assign G[122] = in[8] & in2[8];
    assign P[122] = in[8] ^ in2[8];
    assign G[123] = in[7] & in2[7];
    assign P[123] = in[7] ^ in2[7];
    assign G[124] = in[6] & in2[6];
    assign P[124] = in[6] ^ in2[6];
    assign G[125] = in[5] & in2[5];
    assign P[125] = in[5] ^ in2[5];
    assign G[126] = in[4] & in2[4];
    assign P[126] = in[4] ^ in2[4];
    assign G[127] = in[3] & in2[3];
    assign P[127] = in[3] ^ in2[3];
    assign G[128] = in[2] & in2[2];
    assign P[128] = in[2] ^ in2[2];
    assign G[129] = in[1] & in2[1];
    assign P[129] = in[1] ^ in2[1];
    assign G[130] = in[0] & in2[0];
    assign P[130] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign C[130] = G[129] | (P[129] & C[129]);
    assign cout = G[130] | (P[130] & C[130]);
    assign sum = P ^ C;
endmodule

module CLA130(output [129:0] sum, output cout, input [129:0] in1, input [129:0] in2;

    wire[129:0] G;
    wire[129:0] C;
    wire[129:0] P;

    assign G[0] = in[129] & in2[129];
    assign P[0] = in[129] ^ in2[129];
    assign G[1] = in[128] & in2[128];
    assign P[1] = in[128] ^ in2[128];
    assign G[2] = in[127] & in2[127];
    assign P[2] = in[127] ^ in2[127];
    assign G[3] = in[126] & in2[126];
    assign P[3] = in[126] ^ in2[126];
    assign G[4] = in[125] & in2[125];
    assign P[4] = in[125] ^ in2[125];
    assign G[5] = in[124] & in2[124];
    assign P[5] = in[124] ^ in2[124];
    assign G[6] = in[123] & in2[123];
    assign P[6] = in[123] ^ in2[123];
    assign G[7] = in[122] & in2[122];
    assign P[7] = in[122] ^ in2[122];
    assign G[8] = in[121] & in2[121];
    assign P[8] = in[121] ^ in2[121];
    assign G[9] = in[120] & in2[120];
    assign P[9] = in[120] ^ in2[120];
    assign G[10] = in[119] & in2[119];
    assign P[10] = in[119] ^ in2[119];
    assign G[11] = in[118] & in2[118];
    assign P[11] = in[118] ^ in2[118];
    assign G[12] = in[117] & in2[117];
    assign P[12] = in[117] ^ in2[117];
    assign G[13] = in[116] & in2[116];
    assign P[13] = in[116] ^ in2[116];
    assign G[14] = in[115] & in2[115];
    assign P[14] = in[115] ^ in2[115];
    assign G[15] = in[114] & in2[114];
    assign P[15] = in[114] ^ in2[114];
    assign G[16] = in[113] & in2[113];
    assign P[16] = in[113] ^ in2[113];
    assign G[17] = in[112] & in2[112];
    assign P[17] = in[112] ^ in2[112];
    assign G[18] = in[111] & in2[111];
    assign P[18] = in[111] ^ in2[111];
    assign G[19] = in[110] & in2[110];
    assign P[19] = in[110] ^ in2[110];
    assign G[20] = in[109] & in2[109];
    assign P[20] = in[109] ^ in2[109];
    assign G[21] = in[108] & in2[108];
    assign P[21] = in[108] ^ in2[108];
    assign G[22] = in[107] & in2[107];
    assign P[22] = in[107] ^ in2[107];
    assign G[23] = in[106] & in2[106];
    assign P[23] = in[106] ^ in2[106];
    assign G[24] = in[105] & in2[105];
    assign P[24] = in[105] ^ in2[105];
    assign G[25] = in[104] & in2[104];
    assign P[25] = in[104] ^ in2[104];
    assign G[26] = in[103] & in2[103];
    assign P[26] = in[103] ^ in2[103];
    assign G[27] = in[102] & in2[102];
    assign P[27] = in[102] ^ in2[102];
    assign G[28] = in[101] & in2[101];
    assign P[28] = in[101] ^ in2[101];
    assign G[29] = in[100] & in2[100];
    assign P[29] = in[100] ^ in2[100];
    assign G[30] = in[99] & in2[99];
    assign P[30] = in[99] ^ in2[99];
    assign G[31] = in[98] & in2[98];
    assign P[31] = in[98] ^ in2[98];
    assign G[32] = in[97] & in2[97];
    assign P[32] = in[97] ^ in2[97];
    assign G[33] = in[96] & in2[96];
    assign P[33] = in[96] ^ in2[96];
    assign G[34] = in[95] & in2[95];
    assign P[34] = in[95] ^ in2[95];
    assign G[35] = in[94] & in2[94];
    assign P[35] = in[94] ^ in2[94];
    assign G[36] = in[93] & in2[93];
    assign P[36] = in[93] ^ in2[93];
    assign G[37] = in[92] & in2[92];
    assign P[37] = in[92] ^ in2[92];
    assign G[38] = in[91] & in2[91];
    assign P[38] = in[91] ^ in2[91];
    assign G[39] = in[90] & in2[90];
    assign P[39] = in[90] ^ in2[90];
    assign G[40] = in[89] & in2[89];
    assign P[40] = in[89] ^ in2[89];
    assign G[41] = in[88] & in2[88];
    assign P[41] = in[88] ^ in2[88];
    assign G[42] = in[87] & in2[87];
    assign P[42] = in[87] ^ in2[87];
    assign G[43] = in[86] & in2[86];
    assign P[43] = in[86] ^ in2[86];
    assign G[44] = in[85] & in2[85];
    assign P[44] = in[85] ^ in2[85];
    assign G[45] = in[84] & in2[84];
    assign P[45] = in[84] ^ in2[84];
    assign G[46] = in[83] & in2[83];
    assign P[46] = in[83] ^ in2[83];
    assign G[47] = in[82] & in2[82];
    assign P[47] = in[82] ^ in2[82];
    assign G[48] = in[81] & in2[81];
    assign P[48] = in[81] ^ in2[81];
    assign G[49] = in[80] & in2[80];
    assign P[49] = in[80] ^ in2[80];
    assign G[50] = in[79] & in2[79];
    assign P[50] = in[79] ^ in2[79];
    assign G[51] = in[78] & in2[78];
    assign P[51] = in[78] ^ in2[78];
    assign G[52] = in[77] & in2[77];
    assign P[52] = in[77] ^ in2[77];
    assign G[53] = in[76] & in2[76];
    assign P[53] = in[76] ^ in2[76];
    assign G[54] = in[75] & in2[75];
    assign P[54] = in[75] ^ in2[75];
    assign G[55] = in[74] & in2[74];
    assign P[55] = in[74] ^ in2[74];
    assign G[56] = in[73] & in2[73];
    assign P[56] = in[73] ^ in2[73];
    assign G[57] = in[72] & in2[72];
    assign P[57] = in[72] ^ in2[72];
    assign G[58] = in[71] & in2[71];
    assign P[58] = in[71] ^ in2[71];
    assign G[59] = in[70] & in2[70];
    assign P[59] = in[70] ^ in2[70];
    assign G[60] = in[69] & in2[69];
    assign P[60] = in[69] ^ in2[69];
    assign G[61] = in[68] & in2[68];
    assign P[61] = in[68] ^ in2[68];
    assign G[62] = in[67] & in2[67];
    assign P[62] = in[67] ^ in2[67];
    assign G[63] = in[66] & in2[66];
    assign P[63] = in[66] ^ in2[66];
    assign G[64] = in[65] & in2[65];
    assign P[64] = in[65] ^ in2[65];
    assign G[65] = in[64] & in2[64];
    assign P[65] = in[64] ^ in2[64];
    assign G[66] = in[63] & in2[63];
    assign P[66] = in[63] ^ in2[63];
    assign G[67] = in[62] & in2[62];
    assign P[67] = in[62] ^ in2[62];
    assign G[68] = in[61] & in2[61];
    assign P[68] = in[61] ^ in2[61];
    assign G[69] = in[60] & in2[60];
    assign P[69] = in[60] ^ in2[60];
    assign G[70] = in[59] & in2[59];
    assign P[70] = in[59] ^ in2[59];
    assign G[71] = in[58] & in2[58];
    assign P[71] = in[58] ^ in2[58];
    assign G[72] = in[57] & in2[57];
    assign P[72] = in[57] ^ in2[57];
    assign G[73] = in[56] & in2[56];
    assign P[73] = in[56] ^ in2[56];
    assign G[74] = in[55] & in2[55];
    assign P[74] = in[55] ^ in2[55];
    assign G[75] = in[54] & in2[54];
    assign P[75] = in[54] ^ in2[54];
    assign G[76] = in[53] & in2[53];
    assign P[76] = in[53] ^ in2[53];
    assign G[77] = in[52] & in2[52];
    assign P[77] = in[52] ^ in2[52];
    assign G[78] = in[51] & in2[51];
    assign P[78] = in[51] ^ in2[51];
    assign G[79] = in[50] & in2[50];
    assign P[79] = in[50] ^ in2[50];
    assign G[80] = in[49] & in2[49];
    assign P[80] = in[49] ^ in2[49];
    assign G[81] = in[48] & in2[48];
    assign P[81] = in[48] ^ in2[48];
    assign G[82] = in[47] & in2[47];
    assign P[82] = in[47] ^ in2[47];
    assign G[83] = in[46] & in2[46];
    assign P[83] = in[46] ^ in2[46];
    assign G[84] = in[45] & in2[45];
    assign P[84] = in[45] ^ in2[45];
    assign G[85] = in[44] & in2[44];
    assign P[85] = in[44] ^ in2[44];
    assign G[86] = in[43] & in2[43];
    assign P[86] = in[43] ^ in2[43];
    assign G[87] = in[42] & in2[42];
    assign P[87] = in[42] ^ in2[42];
    assign G[88] = in[41] & in2[41];
    assign P[88] = in[41] ^ in2[41];
    assign G[89] = in[40] & in2[40];
    assign P[89] = in[40] ^ in2[40];
    assign G[90] = in[39] & in2[39];
    assign P[90] = in[39] ^ in2[39];
    assign G[91] = in[38] & in2[38];
    assign P[91] = in[38] ^ in2[38];
    assign G[92] = in[37] & in2[37];
    assign P[92] = in[37] ^ in2[37];
    assign G[93] = in[36] & in2[36];
    assign P[93] = in[36] ^ in2[36];
    assign G[94] = in[35] & in2[35];
    assign P[94] = in[35] ^ in2[35];
    assign G[95] = in[34] & in2[34];
    assign P[95] = in[34] ^ in2[34];
    assign G[96] = in[33] & in2[33];
    assign P[96] = in[33] ^ in2[33];
    assign G[97] = in[32] & in2[32];
    assign P[97] = in[32] ^ in2[32];
    assign G[98] = in[31] & in2[31];
    assign P[98] = in[31] ^ in2[31];
    assign G[99] = in[30] & in2[30];
    assign P[99] = in[30] ^ in2[30];
    assign G[100] = in[29] & in2[29];
    assign P[100] = in[29] ^ in2[29];
    assign G[101] = in[28] & in2[28];
    assign P[101] = in[28] ^ in2[28];
    assign G[102] = in[27] & in2[27];
    assign P[102] = in[27] ^ in2[27];
    assign G[103] = in[26] & in2[26];
    assign P[103] = in[26] ^ in2[26];
    assign G[104] = in[25] & in2[25];
    assign P[104] = in[25] ^ in2[25];
    assign G[105] = in[24] & in2[24];
    assign P[105] = in[24] ^ in2[24];
    assign G[106] = in[23] & in2[23];
    assign P[106] = in[23] ^ in2[23];
    assign G[107] = in[22] & in2[22];
    assign P[107] = in[22] ^ in2[22];
    assign G[108] = in[21] & in2[21];
    assign P[108] = in[21] ^ in2[21];
    assign G[109] = in[20] & in2[20];
    assign P[109] = in[20] ^ in2[20];
    assign G[110] = in[19] & in2[19];
    assign P[110] = in[19] ^ in2[19];
    assign G[111] = in[18] & in2[18];
    assign P[111] = in[18] ^ in2[18];
    assign G[112] = in[17] & in2[17];
    assign P[112] = in[17] ^ in2[17];
    assign G[113] = in[16] & in2[16];
    assign P[113] = in[16] ^ in2[16];
    assign G[114] = in[15] & in2[15];
    assign P[114] = in[15] ^ in2[15];
    assign G[115] = in[14] & in2[14];
    assign P[115] = in[14] ^ in2[14];
    assign G[116] = in[13] & in2[13];
    assign P[116] = in[13] ^ in2[13];
    assign G[117] = in[12] & in2[12];
    assign P[117] = in[12] ^ in2[12];
    assign G[118] = in[11] & in2[11];
    assign P[118] = in[11] ^ in2[11];
    assign G[119] = in[10] & in2[10];
    assign P[119] = in[10] ^ in2[10];
    assign G[120] = in[9] & in2[9];
    assign P[120] = in[9] ^ in2[9];
    assign G[121] = in[8] & in2[8];
    assign P[121] = in[8] ^ in2[8];
    assign G[122] = in[7] & in2[7];
    assign P[122] = in[7] ^ in2[7];
    assign G[123] = in[6] & in2[6];
    assign P[123] = in[6] ^ in2[6];
    assign G[124] = in[5] & in2[5];
    assign P[124] = in[5] ^ in2[5];
    assign G[125] = in[4] & in2[4];
    assign P[125] = in[4] ^ in2[4];
    assign G[126] = in[3] & in2[3];
    assign P[126] = in[3] ^ in2[3];
    assign G[127] = in[2] & in2[2];
    assign P[127] = in[2] ^ in2[2];
    assign G[128] = in[1] & in2[1];
    assign P[128] = in[1] ^ in2[1];
    assign G[129] = in[0] & in2[0];
    assign P[129] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign C[129] = G[128] | (P[128] & C[128]);
    assign cout = G[129] | (P[129] & C[129]);
    assign sum = P ^ C;
endmodule

module CLA129(output [128:0] sum, output cout, input [128:0] in1, input [128:0] in2;

    wire[128:0] G;
    wire[128:0] C;
    wire[128:0] P;

    assign G[0] = in[128] & in2[128];
    assign P[0] = in[128] ^ in2[128];
    assign G[1] = in[127] & in2[127];
    assign P[1] = in[127] ^ in2[127];
    assign G[2] = in[126] & in2[126];
    assign P[2] = in[126] ^ in2[126];
    assign G[3] = in[125] & in2[125];
    assign P[3] = in[125] ^ in2[125];
    assign G[4] = in[124] & in2[124];
    assign P[4] = in[124] ^ in2[124];
    assign G[5] = in[123] & in2[123];
    assign P[5] = in[123] ^ in2[123];
    assign G[6] = in[122] & in2[122];
    assign P[6] = in[122] ^ in2[122];
    assign G[7] = in[121] & in2[121];
    assign P[7] = in[121] ^ in2[121];
    assign G[8] = in[120] & in2[120];
    assign P[8] = in[120] ^ in2[120];
    assign G[9] = in[119] & in2[119];
    assign P[9] = in[119] ^ in2[119];
    assign G[10] = in[118] & in2[118];
    assign P[10] = in[118] ^ in2[118];
    assign G[11] = in[117] & in2[117];
    assign P[11] = in[117] ^ in2[117];
    assign G[12] = in[116] & in2[116];
    assign P[12] = in[116] ^ in2[116];
    assign G[13] = in[115] & in2[115];
    assign P[13] = in[115] ^ in2[115];
    assign G[14] = in[114] & in2[114];
    assign P[14] = in[114] ^ in2[114];
    assign G[15] = in[113] & in2[113];
    assign P[15] = in[113] ^ in2[113];
    assign G[16] = in[112] & in2[112];
    assign P[16] = in[112] ^ in2[112];
    assign G[17] = in[111] & in2[111];
    assign P[17] = in[111] ^ in2[111];
    assign G[18] = in[110] & in2[110];
    assign P[18] = in[110] ^ in2[110];
    assign G[19] = in[109] & in2[109];
    assign P[19] = in[109] ^ in2[109];
    assign G[20] = in[108] & in2[108];
    assign P[20] = in[108] ^ in2[108];
    assign G[21] = in[107] & in2[107];
    assign P[21] = in[107] ^ in2[107];
    assign G[22] = in[106] & in2[106];
    assign P[22] = in[106] ^ in2[106];
    assign G[23] = in[105] & in2[105];
    assign P[23] = in[105] ^ in2[105];
    assign G[24] = in[104] & in2[104];
    assign P[24] = in[104] ^ in2[104];
    assign G[25] = in[103] & in2[103];
    assign P[25] = in[103] ^ in2[103];
    assign G[26] = in[102] & in2[102];
    assign P[26] = in[102] ^ in2[102];
    assign G[27] = in[101] & in2[101];
    assign P[27] = in[101] ^ in2[101];
    assign G[28] = in[100] & in2[100];
    assign P[28] = in[100] ^ in2[100];
    assign G[29] = in[99] & in2[99];
    assign P[29] = in[99] ^ in2[99];
    assign G[30] = in[98] & in2[98];
    assign P[30] = in[98] ^ in2[98];
    assign G[31] = in[97] & in2[97];
    assign P[31] = in[97] ^ in2[97];
    assign G[32] = in[96] & in2[96];
    assign P[32] = in[96] ^ in2[96];
    assign G[33] = in[95] & in2[95];
    assign P[33] = in[95] ^ in2[95];
    assign G[34] = in[94] & in2[94];
    assign P[34] = in[94] ^ in2[94];
    assign G[35] = in[93] & in2[93];
    assign P[35] = in[93] ^ in2[93];
    assign G[36] = in[92] & in2[92];
    assign P[36] = in[92] ^ in2[92];
    assign G[37] = in[91] & in2[91];
    assign P[37] = in[91] ^ in2[91];
    assign G[38] = in[90] & in2[90];
    assign P[38] = in[90] ^ in2[90];
    assign G[39] = in[89] & in2[89];
    assign P[39] = in[89] ^ in2[89];
    assign G[40] = in[88] & in2[88];
    assign P[40] = in[88] ^ in2[88];
    assign G[41] = in[87] & in2[87];
    assign P[41] = in[87] ^ in2[87];
    assign G[42] = in[86] & in2[86];
    assign P[42] = in[86] ^ in2[86];
    assign G[43] = in[85] & in2[85];
    assign P[43] = in[85] ^ in2[85];
    assign G[44] = in[84] & in2[84];
    assign P[44] = in[84] ^ in2[84];
    assign G[45] = in[83] & in2[83];
    assign P[45] = in[83] ^ in2[83];
    assign G[46] = in[82] & in2[82];
    assign P[46] = in[82] ^ in2[82];
    assign G[47] = in[81] & in2[81];
    assign P[47] = in[81] ^ in2[81];
    assign G[48] = in[80] & in2[80];
    assign P[48] = in[80] ^ in2[80];
    assign G[49] = in[79] & in2[79];
    assign P[49] = in[79] ^ in2[79];
    assign G[50] = in[78] & in2[78];
    assign P[50] = in[78] ^ in2[78];
    assign G[51] = in[77] & in2[77];
    assign P[51] = in[77] ^ in2[77];
    assign G[52] = in[76] & in2[76];
    assign P[52] = in[76] ^ in2[76];
    assign G[53] = in[75] & in2[75];
    assign P[53] = in[75] ^ in2[75];
    assign G[54] = in[74] & in2[74];
    assign P[54] = in[74] ^ in2[74];
    assign G[55] = in[73] & in2[73];
    assign P[55] = in[73] ^ in2[73];
    assign G[56] = in[72] & in2[72];
    assign P[56] = in[72] ^ in2[72];
    assign G[57] = in[71] & in2[71];
    assign P[57] = in[71] ^ in2[71];
    assign G[58] = in[70] & in2[70];
    assign P[58] = in[70] ^ in2[70];
    assign G[59] = in[69] & in2[69];
    assign P[59] = in[69] ^ in2[69];
    assign G[60] = in[68] & in2[68];
    assign P[60] = in[68] ^ in2[68];
    assign G[61] = in[67] & in2[67];
    assign P[61] = in[67] ^ in2[67];
    assign G[62] = in[66] & in2[66];
    assign P[62] = in[66] ^ in2[66];
    assign G[63] = in[65] & in2[65];
    assign P[63] = in[65] ^ in2[65];
    assign G[64] = in[64] & in2[64];
    assign P[64] = in[64] ^ in2[64];
    assign G[65] = in[63] & in2[63];
    assign P[65] = in[63] ^ in2[63];
    assign G[66] = in[62] & in2[62];
    assign P[66] = in[62] ^ in2[62];
    assign G[67] = in[61] & in2[61];
    assign P[67] = in[61] ^ in2[61];
    assign G[68] = in[60] & in2[60];
    assign P[68] = in[60] ^ in2[60];
    assign G[69] = in[59] & in2[59];
    assign P[69] = in[59] ^ in2[59];
    assign G[70] = in[58] & in2[58];
    assign P[70] = in[58] ^ in2[58];
    assign G[71] = in[57] & in2[57];
    assign P[71] = in[57] ^ in2[57];
    assign G[72] = in[56] & in2[56];
    assign P[72] = in[56] ^ in2[56];
    assign G[73] = in[55] & in2[55];
    assign P[73] = in[55] ^ in2[55];
    assign G[74] = in[54] & in2[54];
    assign P[74] = in[54] ^ in2[54];
    assign G[75] = in[53] & in2[53];
    assign P[75] = in[53] ^ in2[53];
    assign G[76] = in[52] & in2[52];
    assign P[76] = in[52] ^ in2[52];
    assign G[77] = in[51] & in2[51];
    assign P[77] = in[51] ^ in2[51];
    assign G[78] = in[50] & in2[50];
    assign P[78] = in[50] ^ in2[50];
    assign G[79] = in[49] & in2[49];
    assign P[79] = in[49] ^ in2[49];
    assign G[80] = in[48] & in2[48];
    assign P[80] = in[48] ^ in2[48];
    assign G[81] = in[47] & in2[47];
    assign P[81] = in[47] ^ in2[47];
    assign G[82] = in[46] & in2[46];
    assign P[82] = in[46] ^ in2[46];
    assign G[83] = in[45] & in2[45];
    assign P[83] = in[45] ^ in2[45];
    assign G[84] = in[44] & in2[44];
    assign P[84] = in[44] ^ in2[44];
    assign G[85] = in[43] & in2[43];
    assign P[85] = in[43] ^ in2[43];
    assign G[86] = in[42] & in2[42];
    assign P[86] = in[42] ^ in2[42];
    assign G[87] = in[41] & in2[41];
    assign P[87] = in[41] ^ in2[41];
    assign G[88] = in[40] & in2[40];
    assign P[88] = in[40] ^ in2[40];
    assign G[89] = in[39] & in2[39];
    assign P[89] = in[39] ^ in2[39];
    assign G[90] = in[38] & in2[38];
    assign P[90] = in[38] ^ in2[38];
    assign G[91] = in[37] & in2[37];
    assign P[91] = in[37] ^ in2[37];
    assign G[92] = in[36] & in2[36];
    assign P[92] = in[36] ^ in2[36];
    assign G[93] = in[35] & in2[35];
    assign P[93] = in[35] ^ in2[35];
    assign G[94] = in[34] & in2[34];
    assign P[94] = in[34] ^ in2[34];
    assign G[95] = in[33] & in2[33];
    assign P[95] = in[33] ^ in2[33];
    assign G[96] = in[32] & in2[32];
    assign P[96] = in[32] ^ in2[32];
    assign G[97] = in[31] & in2[31];
    assign P[97] = in[31] ^ in2[31];
    assign G[98] = in[30] & in2[30];
    assign P[98] = in[30] ^ in2[30];
    assign G[99] = in[29] & in2[29];
    assign P[99] = in[29] ^ in2[29];
    assign G[100] = in[28] & in2[28];
    assign P[100] = in[28] ^ in2[28];
    assign G[101] = in[27] & in2[27];
    assign P[101] = in[27] ^ in2[27];
    assign G[102] = in[26] & in2[26];
    assign P[102] = in[26] ^ in2[26];
    assign G[103] = in[25] & in2[25];
    assign P[103] = in[25] ^ in2[25];
    assign G[104] = in[24] & in2[24];
    assign P[104] = in[24] ^ in2[24];
    assign G[105] = in[23] & in2[23];
    assign P[105] = in[23] ^ in2[23];
    assign G[106] = in[22] & in2[22];
    assign P[106] = in[22] ^ in2[22];
    assign G[107] = in[21] & in2[21];
    assign P[107] = in[21] ^ in2[21];
    assign G[108] = in[20] & in2[20];
    assign P[108] = in[20] ^ in2[20];
    assign G[109] = in[19] & in2[19];
    assign P[109] = in[19] ^ in2[19];
    assign G[110] = in[18] & in2[18];
    assign P[110] = in[18] ^ in2[18];
    assign G[111] = in[17] & in2[17];
    assign P[111] = in[17] ^ in2[17];
    assign G[112] = in[16] & in2[16];
    assign P[112] = in[16] ^ in2[16];
    assign G[113] = in[15] & in2[15];
    assign P[113] = in[15] ^ in2[15];
    assign G[114] = in[14] & in2[14];
    assign P[114] = in[14] ^ in2[14];
    assign G[115] = in[13] & in2[13];
    assign P[115] = in[13] ^ in2[13];
    assign G[116] = in[12] & in2[12];
    assign P[116] = in[12] ^ in2[12];
    assign G[117] = in[11] & in2[11];
    assign P[117] = in[11] ^ in2[11];
    assign G[118] = in[10] & in2[10];
    assign P[118] = in[10] ^ in2[10];
    assign G[119] = in[9] & in2[9];
    assign P[119] = in[9] ^ in2[9];
    assign G[120] = in[8] & in2[8];
    assign P[120] = in[8] ^ in2[8];
    assign G[121] = in[7] & in2[7];
    assign P[121] = in[7] ^ in2[7];
    assign G[122] = in[6] & in2[6];
    assign P[122] = in[6] ^ in2[6];
    assign G[123] = in[5] & in2[5];
    assign P[123] = in[5] ^ in2[5];
    assign G[124] = in[4] & in2[4];
    assign P[124] = in[4] ^ in2[4];
    assign G[125] = in[3] & in2[3];
    assign P[125] = in[3] ^ in2[3];
    assign G[126] = in[2] & in2[2];
    assign P[126] = in[2] ^ in2[2];
    assign G[127] = in[1] & in2[1];
    assign P[127] = in[1] ^ in2[1];
    assign G[128] = in[0] & in2[0];
    assign P[128] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign C[128] = G[127] | (P[127] & C[127]);
    assign cout = G[128] | (P[128] & C[128]);
    assign sum = P ^ C;
endmodule

module CLA128(output [127:0] sum, output cout, input [127:0] in1, input [127:0] in2;

    wire[127:0] G;
    wire[127:0] C;
    wire[127:0] P;

    assign G[0] = in[127] & in2[127];
    assign P[0] = in[127] ^ in2[127];
    assign G[1] = in[126] & in2[126];
    assign P[1] = in[126] ^ in2[126];
    assign G[2] = in[125] & in2[125];
    assign P[2] = in[125] ^ in2[125];
    assign G[3] = in[124] & in2[124];
    assign P[3] = in[124] ^ in2[124];
    assign G[4] = in[123] & in2[123];
    assign P[4] = in[123] ^ in2[123];
    assign G[5] = in[122] & in2[122];
    assign P[5] = in[122] ^ in2[122];
    assign G[6] = in[121] & in2[121];
    assign P[6] = in[121] ^ in2[121];
    assign G[7] = in[120] & in2[120];
    assign P[7] = in[120] ^ in2[120];
    assign G[8] = in[119] & in2[119];
    assign P[8] = in[119] ^ in2[119];
    assign G[9] = in[118] & in2[118];
    assign P[9] = in[118] ^ in2[118];
    assign G[10] = in[117] & in2[117];
    assign P[10] = in[117] ^ in2[117];
    assign G[11] = in[116] & in2[116];
    assign P[11] = in[116] ^ in2[116];
    assign G[12] = in[115] & in2[115];
    assign P[12] = in[115] ^ in2[115];
    assign G[13] = in[114] & in2[114];
    assign P[13] = in[114] ^ in2[114];
    assign G[14] = in[113] & in2[113];
    assign P[14] = in[113] ^ in2[113];
    assign G[15] = in[112] & in2[112];
    assign P[15] = in[112] ^ in2[112];
    assign G[16] = in[111] & in2[111];
    assign P[16] = in[111] ^ in2[111];
    assign G[17] = in[110] & in2[110];
    assign P[17] = in[110] ^ in2[110];
    assign G[18] = in[109] & in2[109];
    assign P[18] = in[109] ^ in2[109];
    assign G[19] = in[108] & in2[108];
    assign P[19] = in[108] ^ in2[108];
    assign G[20] = in[107] & in2[107];
    assign P[20] = in[107] ^ in2[107];
    assign G[21] = in[106] & in2[106];
    assign P[21] = in[106] ^ in2[106];
    assign G[22] = in[105] & in2[105];
    assign P[22] = in[105] ^ in2[105];
    assign G[23] = in[104] & in2[104];
    assign P[23] = in[104] ^ in2[104];
    assign G[24] = in[103] & in2[103];
    assign P[24] = in[103] ^ in2[103];
    assign G[25] = in[102] & in2[102];
    assign P[25] = in[102] ^ in2[102];
    assign G[26] = in[101] & in2[101];
    assign P[26] = in[101] ^ in2[101];
    assign G[27] = in[100] & in2[100];
    assign P[27] = in[100] ^ in2[100];
    assign G[28] = in[99] & in2[99];
    assign P[28] = in[99] ^ in2[99];
    assign G[29] = in[98] & in2[98];
    assign P[29] = in[98] ^ in2[98];
    assign G[30] = in[97] & in2[97];
    assign P[30] = in[97] ^ in2[97];
    assign G[31] = in[96] & in2[96];
    assign P[31] = in[96] ^ in2[96];
    assign G[32] = in[95] & in2[95];
    assign P[32] = in[95] ^ in2[95];
    assign G[33] = in[94] & in2[94];
    assign P[33] = in[94] ^ in2[94];
    assign G[34] = in[93] & in2[93];
    assign P[34] = in[93] ^ in2[93];
    assign G[35] = in[92] & in2[92];
    assign P[35] = in[92] ^ in2[92];
    assign G[36] = in[91] & in2[91];
    assign P[36] = in[91] ^ in2[91];
    assign G[37] = in[90] & in2[90];
    assign P[37] = in[90] ^ in2[90];
    assign G[38] = in[89] & in2[89];
    assign P[38] = in[89] ^ in2[89];
    assign G[39] = in[88] & in2[88];
    assign P[39] = in[88] ^ in2[88];
    assign G[40] = in[87] & in2[87];
    assign P[40] = in[87] ^ in2[87];
    assign G[41] = in[86] & in2[86];
    assign P[41] = in[86] ^ in2[86];
    assign G[42] = in[85] & in2[85];
    assign P[42] = in[85] ^ in2[85];
    assign G[43] = in[84] & in2[84];
    assign P[43] = in[84] ^ in2[84];
    assign G[44] = in[83] & in2[83];
    assign P[44] = in[83] ^ in2[83];
    assign G[45] = in[82] & in2[82];
    assign P[45] = in[82] ^ in2[82];
    assign G[46] = in[81] & in2[81];
    assign P[46] = in[81] ^ in2[81];
    assign G[47] = in[80] & in2[80];
    assign P[47] = in[80] ^ in2[80];
    assign G[48] = in[79] & in2[79];
    assign P[48] = in[79] ^ in2[79];
    assign G[49] = in[78] & in2[78];
    assign P[49] = in[78] ^ in2[78];
    assign G[50] = in[77] & in2[77];
    assign P[50] = in[77] ^ in2[77];
    assign G[51] = in[76] & in2[76];
    assign P[51] = in[76] ^ in2[76];
    assign G[52] = in[75] & in2[75];
    assign P[52] = in[75] ^ in2[75];
    assign G[53] = in[74] & in2[74];
    assign P[53] = in[74] ^ in2[74];
    assign G[54] = in[73] & in2[73];
    assign P[54] = in[73] ^ in2[73];
    assign G[55] = in[72] & in2[72];
    assign P[55] = in[72] ^ in2[72];
    assign G[56] = in[71] & in2[71];
    assign P[56] = in[71] ^ in2[71];
    assign G[57] = in[70] & in2[70];
    assign P[57] = in[70] ^ in2[70];
    assign G[58] = in[69] & in2[69];
    assign P[58] = in[69] ^ in2[69];
    assign G[59] = in[68] & in2[68];
    assign P[59] = in[68] ^ in2[68];
    assign G[60] = in[67] & in2[67];
    assign P[60] = in[67] ^ in2[67];
    assign G[61] = in[66] & in2[66];
    assign P[61] = in[66] ^ in2[66];
    assign G[62] = in[65] & in2[65];
    assign P[62] = in[65] ^ in2[65];
    assign G[63] = in[64] & in2[64];
    assign P[63] = in[64] ^ in2[64];
    assign G[64] = in[63] & in2[63];
    assign P[64] = in[63] ^ in2[63];
    assign G[65] = in[62] & in2[62];
    assign P[65] = in[62] ^ in2[62];
    assign G[66] = in[61] & in2[61];
    assign P[66] = in[61] ^ in2[61];
    assign G[67] = in[60] & in2[60];
    assign P[67] = in[60] ^ in2[60];
    assign G[68] = in[59] & in2[59];
    assign P[68] = in[59] ^ in2[59];
    assign G[69] = in[58] & in2[58];
    assign P[69] = in[58] ^ in2[58];
    assign G[70] = in[57] & in2[57];
    assign P[70] = in[57] ^ in2[57];
    assign G[71] = in[56] & in2[56];
    assign P[71] = in[56] ^ in2[56];
    assign G[72] = in[55] & in2[55];
    assign P[72] = in[55] ^ in2[55];
    assign G[73] = in[54] & in2[54];
    assign P[73] = in[54] ^ in2[54];
    assign G[74] = in[53] & in2[53];
    assign P[74] = in[53] ^ in2[53];
    assign G[75] = in[52] & in2[52];
    assign P[75] = in[52] ^ in2[52];
    assign G[76] = in[51] & in2[51];
    assign P[76] = in[51] ^ in2[51];
    assign G[77] = in[50] & in2[50];
    assign P[77] = in[50] ^ in2[50];
    assign G[78] = in[49] & in2[49];
    assign P[78] = in[49] ^ in2[49];
    assign G[79] = in[48] & in2[48];
    assign P[79] = in[48] ^ in2[48];
    assign G[80] = in[47] & in2[47];
    assign P[80] = in[47] ^ in2[47];
    assign G[81] = in[46] & in2[46];
    assign P[81] = in[46] ^ in2[46];
    assign G[82] = in[45] & in2[45];
    assign P[82] = in[45] ^ in2[45];
    assign G[83] = in[44] & in2[44];
    assign P[83] = in[44] ^ in2[44];
    assign G[84] = in[43] & in2[43];
    assign P[84] = in[43] ^ in2[43];
    assign G[85] = in[42] & in2[42];
    assign P[85] = in[42] ^ in2[42];
    assign G[86] = in[41] & in2[41];
    assign P[86] = in[41] ^ in2[41];
    assign G[87] = in[40] & in2[40];
    assign P[87] = in[40] ^ in2[40];
    assign G[88] = in[39] & in2[39];
    assign P[88] = in[39] ^ in2[39];
    assign G[89] = in[38] & in2[38];
    assign P[89] = in[38] ^ in2[38];
    assign G[90] = in[37] & in2[37];
    assign P[90] = in[37] ^ in2[37];
    assign G[91] = in[36] & in2[36];
    assign P[91] = in[36] ^ in2[36];
    assign G[92] = in[35] & in2[35];
    assign P[92] = in[35] ^ in2[35];
    assign G[93] = in[34] & in2[34];
    assign P[93] = in[34] ^ in2[34];
    assign G[94] = in[33] & in2[33];
    assign P[94] = in[33] ^ in2[33];
    assign G[95] = in[32] & in2[32];
    assign P[95] = in[32] ^ in2[32];
    assign G[96] = in[31] & in2[31];
    assign P[96] = in[31] ^ in2[31];
    assign G[97] = in[30] & in2[30];
    assign P[97] = in[30] ^ in2[30];
    assign G[98] = in[29] & in2[29];
    assign P[98] = in[29] ^ in2[29];
    assign G[99] = in[28] & in2[28];
    assign P[99] = in[28] ^ in2[28];
    assign G[100] = in[27] & in2[27];
    assign P[100] = in[27] ^ in2[27];
    assign G[101] = in[26] & in2[26];
    assign P[101] = in[26] ^ in2[26];
    assign G[102] = in[25] & in2[25];
    assign P[102] = in[25] ^ in2[25];
    assign G[103] = in[24] & in2[24];
    assign P[103] = in[24] ^ in2[24];
    assign G[104] = in[23] & in2[23];
    assign P[104] = in[23] ^ in2[23];
    assign G[105] = in[22] & in2[22];
    assign P[105] = in[22] ^ in2[22];
    assign G[106] = in[21] & in2[21];
    assign P[106] = in[21] ^ in2[21];
    assign G[107] = in[20] & in2[20];
    assign P[107] = in[20] ^ in2[20];
    assign G[108] = in[19] & in2[19];
    assign P[108] = in[19] ^ in2[19];
    assign G[109] = in[18] & in2[18];
    assign P[109] = in[18] ^ in2[18];
    assign G[110] = in[17] & in2[17];
    assign P[110] = in[17] ^ in2[17];
    assign G[111] = in[16] & in2[16];
    assign P[111] = in[16] ^ in2[16];
    assign G[112] = in[15] & in2[15];
    assign P[112] = in[15] ^ in2[15];
    assign G[113] = in[14] & in2[14];
    assign P[113] = in[14] ^ in2[14];
    assign G[114] = in[13] & in2[13];
    assign P[114] = in[13] ^ in2[13];
    assign G[115] = in[12] & in2[12];
    assign P[115] = in[12] ^ in2[12];
    assign G[116] = in[11] & in2[11];
    assign P[116] = in[11] ^ in2[11];
    assign G[117] = in[10] & in2[10];
    assign P[117] = in[10] ^ in2[10];
    assign G[118] = in[9] & in2[9];
    assign P[118] = in[9] ^ in2[9];
    assign G[119] = in[8] & in2[8];
    assign P[119] = in[8] ^ in2[8];
    assign G[120] = in[7] & in2[7];
    assign P[120] = in[7] ^ in2[7];
    assign G[121] = in[6] & in2[6];
    assign P[121] = in[6] ^ in2[6];
    assign G[122] = in[5] & in2[5];
    assign P[122] = in[5] ^ in2[5];
    assign G[123] = in[4] & in2[4];
    assign P[123] = in[4] ^ in2[4];
    assign G[124] = in[3] & in2[3];
    assign P[124] = in[3] ^ in2[3];
    assign G[125] = in[2] & in2[2];
    assign P[125] = in[2] ^ in2[2];
    assign G[126] = in[1] & in2[1];
    assign P[126] = in[1] ^ in2[1];
    assign G[127] = in[0] & in2[0];
    assign P[127] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign C[127] = G[126] | (P[126] & C[126]);
    assign cout = G[127] | (P[127] & C[127]);
    assign sum = P ^ C;
endmodule

module CLA127(output [126:0] sum, output cout, input [126:0] in1, input [126:0] in2;

    wire[126:0] G;
    wire[126:0] C;
    wire[126:0] P;

    assign G[0] = in[126] & in2[126];
    assign P[0] = in[126] ^ in2[126];
    assign G[1] = in[125] & in2[125];
    assign P[1] = in[125] ^ in2[125];
    assign G[2] = in[124] & in2[124];
    assign P[2] = in[124] ^ in2[124];
    assign G[3] = in[123] & in2[123];
    assign P[3] = in[123] ^ in2[123];
    assign G[4] = in[122] & in2[122];
    assign P[4] = in[122] ^ in2[122];
    assign G[5] = in[121] & in2[121];
    assign P[5] = in[121] ^ in2[121];
    assign G[6] = in[120] & in2[120];
    assign P[6] = in[120] ^ in2[120];
    assign G[7] = in[119] & in2[119];
    assign P[7] = in[119] ^ in2[119];
    assign G[8] = in[118] & in2[118];
    assign P[8] = in[118] ^ in2[118];
    assign G[9] = in[117] & in2[117];
    assign P[9] = in[117] ^ in2[117];
    assign G[10] = in[116] & in2[116];
    assign P[10] = in[116] ^ in2[116];
    assign G[11] = in[115] & in2[115];
    assign P[11] = in[115] ^ in2[115];
    assign G[12] = in[114] & in2[114];
    assign P[12] = in[114] ^ in2[114];
    assign G[13] = in[113] & in2[113];
    assign P[13] = in[113] ^ in2[113];
    assign G[14] = in[112] & in2[112];
    assign P[14] = in[112] ^ in2[112];
    assign G[15] = in[111] & in2[111];
    assign P[15] = in[111] ^ in2[111];
    assign G[16] = in[110] & in2[110];
    assign P[16] = in[110] ^ in2[110];
    assign G[17] = in[109] & in2[109];
    assign P[17] = in[109] ^ in2[109];
    assign G[18] = in[108] & in2[108];
    assign P[18] = in[108] ^ in2[108];
    assign G[19] = in[107] & in2[107];
    assign P[19] = in[107] ^ in2[107];
    assign G[20] = in[106] & in2[106];
    assign P[20] = in[106] ^ in2[106];
    assign G[21] = in[105] & in2[105];
    assign P[21] = in[105] ^ in2[105];
    assign G[22] = in[104] & in2[104];
    assign P[22] = in[104] ^ in2[104];
    assign G[23] = in[103] & in2[103];
    assign P[23] = in[103] ^ in2[103];
    assign G[24] = in[102] & in2[102];
    assign P[24] = in[102] ^ in2[102];
    assign G[25] = in[101] & in2[101];
    assign P[25] = in[101] ^ in2[101];
    assign G[26] = in[100] & in2[100];
    assign P[26] = in[100] ^ in2[100];
    assign G[27] = in[99] & in2[99];
    assign P[27] = in[99] ^ in2[99];
    assign G[28] = in[98] & in2[98];
    assign P[28] = in[98] ^ in2[98];
    assign G[29] = in[97] & in2[97];
    assign P[29] = in[97] ^ in2[97];
    assign G[30] = in[96] & in2[96];
    assign P[30] = in[96] ^ in2[96];
    assign G[31] = in[95] & in2[95];
    assign P[31] = in[95] ^ in2[95];
    assign G[32] = in[94] & in2[94];
    assign P[32] = in[94] ^ in2[94];
    assign G[33] = in[93] & in2[93];
    assign P[33] = in[93] ^ in2[93];
    assign G[34] = in[92] & in2[92];
    assign P[34] = in[92] ^ in2[92];
    assign G[35] = in[91] & in2[91];
    assign P[35] = in[91] ^ in2[91];
    assign G[36] = in[90] & in2[90];
    assign P[36] = in[90] ^ in2[90];
    assign G[37] = in[89] & in2[89];
    assign P[37] = in[89] ^ in2[89];
    assign G[38] = in[88] & in2[88];
    assign P[38] = in[88] ^ in2[88];
    assign G[39] = in[87] & in2[87];
    assign P[39] = in[87] ^ in2[87];
    assign G[40] = in[86] & in2[86];
    assign P[40] = in[86] ^ in2[86];
    assign G[41] = in[85] & in2[85];
    assign P[41] = in[85] ^ in2[85];
    assign G[42] = in[84] & in2[84];
    assign P[42] = in[84] ^ in2[84];
    assign G[43] = in[83] & in2[83];
    assign P[43] = in[83] ^ in2[83];
    assign G[44] = in[82] & in2[82];
    assign P[44] = in[82] ^ in2[82];
    assign G[45] = in[81] & in2[81];
    assign P[45] = in[81] ^ in2[81];
    assign G[46] = in[80] & in2[80];
    assign P[46] = in[80] ^ in2[80];
    assign G[47] = in[79] & in2[79];
    assign P[47] = in[79] ^ in2[79];
    assign G[48] = in[78] & in2[78];
    assign P[48] = in[78] ^ in2[78];
    assign G[49] = in[77] & in2[77];
    assign P[49] = in[77] ^ in2[77];
    assign G[50] = in[76] & in2[76];
    assign P[50] = in[76] ^ in2[76];
    assign G[51] = in[75] & in2[75];
    assign P[51] = in[75] ^ in2[75];
    assign G[52] = in[74] & in2[74];
    assign P[52] = in[74] ^ in2[74];
    assign G[53] = in[73] & in2[73];
    assign P[53] = in[73] ^ in2[73];
    assign G[54] = in[72] & in2[72];
    assign P[54] = in[72] ^ in2[72];
    assign G[55] = in[71] & in2[71];
    assign P[55] = in[71] ^ in2[71];
    assign G[56] = in[70] & in2[70];
    assign P[56] = in[70] ^ in2[70];
    assign G[57] = in[69] & in2[69];
    assign P[57] = in[69] ^ in2[69];
    assign G[58] = in[68] & in2[68];
    assign P[58] = in[68] ^ in2[68];
    assign G[59] = in[67] & in2[67];
    assign P[59] = in[67] ^ in2[67];
    assign G[60] = in[66] & in2[66];
    assign P[60] = in[66] ^ in2[66];
    assign G[61] = in[65] & in2[65];
    assign P[61] = in[65] ^ in2[65];
    assign G[62] = in[64] & in2[64];
    assign P[62] = in[64] ^ in2[64];
    assign G[63] = in[63] & in2[63];
    assign P[63] = in[63] ^ in2[63];
    assign G[64] = in[62] & in2[62];
    assign P[64] = in[62] ^ in2[62];
    assign G[65] = in[61] & in2[61];
    assign P[65] = in[61] ^ in2[61];
    assign G[66] = in[60] & in2[60];
    assign P[66] = in[60] ^ in2[60];
    assign G[67] = in[59] & in2[59];
    assign P[67] = in[59] ^ in2[59];
    assign G[68] = in[58] & in2[58];
    assign P[68] = in[58] ^ in2[58];
    assign G[69] = in[57] & in2[57];
    assign P[69] = in[57] ^ in2[57];
    assign G[70] = in[56] & in2[56];
    assign P[70] = in[56] ^ in2[56];
    assign G[71] = in[55] & in2[55];
    assign P[71] = in[55] ^ in2[55];
    assign G[72] = in[54] & in2[54];
    assign P[72] = in[54] ^ in2[54];
    assign G[73] = in[53] & in2[53];
    assign P[73] = in[53] ^ in2[53];
    assign G[74] = in[52] & in2[52];
    assign P[74] = in[52] ^ in2[52];
    assign G[75] = in[51] & in2[51];
    assign P[75] = in[51] ^ in2[51];
    assign G[76] = in[50] & in2[50];
    assign P[76] = in[50] ^ in2[50];
    assign G[77] = in[49] & in2[49];
    assign P[77] = in[49] ^ in2[49];
    assign G[78] = in[48] & in2[48];
    assign P[78] = in[48] ^ in2[48];
    assign G[79] = in[47] & in2[47];
    assign P[79] = in[47] ^ in2[47];
    assign G[80] = in[46] & in2[46];
    assign P[80] = in[46] ^ in2[46];
    assign G[81] = in[45] & in2[45];
    assign P[81] = in[45] ^ in2[45];
    assign G[82] = in[44] & in2[44];
    assign P[82] = in[44] ^ in2[44];
    assign G[83] = in[43] & in2[43];
    assign P[83] = in[43] ^ in2[43];
    assign G[84] = in[42] & in2[42];
    assign P[84] = in[42] ^ in2[42];
    assign G[85] = in[41] & in2[41];
    assign P[85] = in[41] ^ in2[41];
    assign G[86] = in[40] & in2[40];
    assign P[86] = in[40] ^ in2[40];
    assign G[87] = in[39] & in2[39];
    assign P[87] = in[39] ^ in2[39];
    assign G[88] = in[38] & in2[38];
    assign P[88] = in[38] ^ in2[38];
    assign G[89] = in[37] & in2[37];
    assign P[89] = in[37] ^ in2[37];
    assign G[90] = in[36] & in2[36];
    assign P[90] = in[36] ^ in2[36];
    assign G[91] = in[35] & in2[35];
    assign P[91] = in[35] ^ in2[35];
    assign G[92] = in[34] & in2[34];
    assign P[92] = in[34] ^ in2[34];
    assign G[93] = in[33] & in2[33];
    assign P[93] = in[33] ^ in2[33];
    assign G[94] = in[32] & in2[32];
    assign P[94] = in[32] ^ in2[32];
    assign G[95] = in[31] & in2[31];
    assign P[95] = in[31] ^ in2[31];
    assign G[96] = in[30] & in2[30];
    assign P[96] = in[30] ^ in2[30];
    assign G[97] = in[29] & in2[29];
    assign P[97] = in[29] ^ in2[29];
    assign G[98] = in[28] & in2[28];
    assign P[98] = in[28] ^ in2[28];
    assign G[99] = in[27] & in2[27];
    assign P[99] = in[27] ^ in2[27];
    assign G[100] = in[26] & in2[26];
    assign P[100] = in[26] ^ in2[26];
    assign G[101] = in[25] & in2[25];
    assign P[101] = in[25] ^ in2[25];
    assign G[102] = in[24] & in2[24];
    assign P[102] = in[24] ^ in2[24];
    assign G[103] = in[23] & in2[23];
    assign P[103] = in[23] ^ in2[23];
    assign G[104] = in[22] & in2[22];
    assign P[104] = in[22] ^ in2[22];
    assign G[105] = in[21] & in2[21];
    assign P[105] = in[21] ^ in2[21];
    assign G[106] = in[20] & in2[20];
    assign P[106] = in[20] ^ in2[20];
    assign G[107] = in[19] & in2[19];
    assign P[107] = in[19] ^ in2[19];
    assign G[108] = in[18] & in2[18];
    assign P[108] = in[18] ^ in2[18];
    assign G[109] = in[17] & in2[17];
    assign P[109] = in[17] ^ in2[17];
    assign G[110] = in[16] & in2[16];
    assign P[110] = in[16] ^ in2[16];
    assign G[111] = in[15] & in2[15];
    assign P[111] = in[15] ^ in2[15];
    assign G[112] = in[14] & in2[14];
    assign P[112] = in[14] ^ in2[14];
    assign G[113] = in[13] & in2[13];
    assign P[113] = in[13] ^ in2[13];
    assign G[114] = in[12] & in2[12];
    assign P[114] = in[12] ^ in2[12];
    assign G[115] = in[11] & in2[11];
    assign P[115] = in[11] ^ in2[11];
    assign G[116] = in[10] & in2[10];
    assign P[116] = in[10] ^ in2[10];
    assign G[117] = in[9] & in2[9];
    assign P[117] = in[9] ^ in2[9];
    assign G[118] = in[8] & in2[8];
    assign P[118] = in[8] ^ in2[8];
    assign G[119] = in[7] & in2[7];
    assign P[119] = in[7] ^ in2[7];
    assign G[120] = in[6] & in2[6];
    assign P[120] = in[6] ^ in2[6];
    assign G[121] = in[5] & in2[5];
    assign P[121] = in[5] ^ in2[5];
    assign G[122] = in[4] & in2[4];
    assign P[122] = in[4] ^ in2[4];
    assign G[123] = in[3] & in2[3];
    assign P[123] = in[3] ^ in2[3];
    assign G[124] = in[2] & in2[2];
    assign P[124] = in[2] ^ in2[2];
    assign G[125] = in[1] & in2[1];
    assign P[125] = in[1] ^ in2[1];
    assign G[126] = in[0] & in2[0];
    assign P[126] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign C[126] = G[125] | (P[125] & C[125]);
    assign cout = G[126] | (P[126] & C[126]);
    assign sum = P ^ C;
endmodule

module CLA126(output [125:0] sum, output cout, input [125:0] in1, input [125:0] in2;

    wire[125:0] G;
    wire[125:0] C;
    wire[125:0] P;

    assign G[0] = in[125] & in2[125];
    assign P[0] = in[125] ^ in2[125];
    assign G[1] = in[124] & in2[124];
    assign P[1] = in[124] ^ in2[124];
    assign G[2] = in[123] & in2[123];
    assign P[2] = in[123] ^ in2[123];
    assign G[3] = in[122] & in2[122];
    assign P[3] = in[122] ^ in2[122];
    assign G[4] = in[121] & in2[121];
    assign P[4] = in[121] ^ in2[121];
    assign G[5] = in[120] & in2[120];
    assign P[5] = in[120] ^ in2[120];
    assign G[6] = in[119] & in2[119];
    assign P[6] = in[119] ^ in2[119];
    assign G[7] = in[118] & in2[118];
    assign P[7] = in[118] ^ in2[118];
    assign G[8] = in[117] & in2[117];
    assign P[8] = in[117] ^ in2[117];
    assign G[9] = in[116] & in2[116];
    assign P[9] = in[116] ^ in2[116];
    assign G[10] = in[115] & in2[115];
    assign P[10] = in[115] ^ in2[115];
    assign G[11] = in[114] & in2[114];
    assign P[11] = in[114] ^ in2[114];
    assign G[12] = in[113] & in2[113];
    assign P[12] = in[113] ^ in2[113];
    assign G[13] = in[112] & in2[112];
    assign P[13] = in[112] ^ in2[112];
    assign G[14] = in[111] & in2[111];
    assign P[14] = in[111] ^ in2[111];
    assign G[15] = in[110] & in2[110];
    assign P[15] = in[110] ^ in2[110];
    assign G[16] = in[109] & in2[109];
    assign P[16] = in[109] ^ in2[109];
    assign G[17] = in[108] & in2[108];
    assign P[17] = in[108] ^ in2[108];
    assign G[18] = in[107] & in2[107];
    assign P[18] = in[107] ^ in2[107];
    assign G[19] = in[106] & in2[106];
    assign P[19] = in[106] ^ in2[106];
    assign G[20] = in[105] & in2[105];
    assign P[20] = in[105] ^ in2[105];
    assign G[21] = in[104] & in2[104];
    assign P[21] = in[104] ^ in2[104];
    assign G[22] = in[103] & in2[103];
    assign P[22] = in[103] ^ in2[103];
    assign G[23] = in[102] & in2[102];
    assign P[23] = in[102] ^ in2[102];
    assign G[24] = in[101] & in2[101];
    assign P[24] = in[101] ^ in2[101];
    assign G[25] = in[100] & in2[100];
    assign P[25] = in[100] ^ in2[100];
    assign G[26] = in[99] & in2[99];
    assign P[26] = in[99] ^ in2[99];
    assign G[27] = in[98] & in2[98];
    assign P[27] = in[98] ^ in2[98];
    assign G[28] = in[97] & in2[97];
    assign P[28] = in[97] ^ in2[97];
    assign G[29] = in[96] & in2[96];
    assign P[29] = in[96] ^ in2[96];
    assign G[30] = in[95] & in2[95];
    assign P[30] = in[95] ^ in2[95];
    assign G[31] = in[94] & in2[94];
    assign P[31] = in[94] ^ in2[94];
    assign G[32] = in[93] & in2[93];
    assign P[32] = in[93] ^ in2[93];
    assign G[33] = in[92] & in2[92];
    assign P[33] = in[92] ^ in2[92];
    assign G[34] = in[91] & in2[91];
    assign P[34] = in[91] ^ in2[91];
    assign G[35] = in[90] & in2[90];
    assign P[35] = in[90] ^ in2[90];
    assign G[36] = in[89] & in2[89];
    assign P[36] = in[89] ^ in2[89];
    assign G[37] = in[88] & in2[88];
    assign P[37] = in[88] ^ in2[88];
    assign G[38] = in[87] & in2[87];
    assign P[38] = in[87] ^ in2[87];
    assign G[39] = in[86] & in2[86];
    assign P[39] = in[86] ^ in2[86];
    assign G[40] = in[85] & in2[85];
    assign P[40] = in[85] ^ in2[85];
    assign G[41] = in[84] & in2[84];
    assign P[41] = in[84] ^ in2[84];
    assign G[42] = in[83] & in2[83];
    assign P[42] = in[83] ^ in2[83];
    assign G[43] = in[82] & in2[82];
    assign P[43] = in[82] ^ in2[82];
    assign G[44] = in[81] & in2[81];
    assign P[44] = in[81] ^ in2[81];
    assign G[45] = in[80] & in2[80];
    assign P[45] = in[80] ^ in2[80];
    assign G[46] = in[79] & in2[79];
    assign P[46] = in[79] ^ in2[79];
    assign G[47] = in[78] & in2[78];
    assign P[47] = in[78] ^ in2[78];
    assign G[48] = in[77] & in2[77];
    assign P[48] = in[77] ^ in2[77];
    assign G[49] = in[76] & in2[76];
    assign P[49] = in[76] ^ in2[76];
    assign G[50] = in[75] & in2[75];
    assign P[50] = in[75] ^ in2[75];
    assign G[51] = in[74] & in2[74];
    assign P[51] = in[74] ^ in2[74];
    assign G[52] = in[73] & in2[73];
    assign P[52] = in[73] ^ in2[73];
    assign G[53] = in[72] & in2[72];
    assign P[53] = in[72] ^ in2[72];
    assign G[54] = in[71] & in2[71];
    assign P[54] = in[71] ^ in2[71];
    assign G[55] = in[70] & in2[70];
    assign P[55] = in[70] ^ in2[70];
    assign G[56] = in[69] & in2[69];
    assign P[56] = in[69] ^ in2[69];
    assign G[57] = in[68] & in2[68];
    assign P[57] = in[68] ^ in2[68];
    assign G[58] = in[67] & in2[67];
    assign P[58] = in[67] ^ in2[67];
    assign G[59] = in[66] & in2[66];
    assign P[59] = in[66] ^ in2[66];
    assign G[60] = in[65] & in2[65];
    assign P[60] = in[65] ^ in2[65];
    assign G[61] = in[64] & in2[64];
    assign P[61] = in[64] ^ in2[64];
    assign G[62] = in[63] & in2[63];
    assign P[62] = in[63] ^ in2[63];
    assign G[63] = in[62] & in2[62];
    assign P[63] = in[62] ^ in2[62];
    assign G[64] = in[61] & in2[61];
    assign P[64] = in[61] ^ in2[61];
    assign G[65] = in[60] & in2[60];
    assign P[65] = in[60] ^ in2[60];
    assign G[66] = in[59] & in2[59];
    assign P[66] = in[59] ^ in2[59];
    assign G[67] = in[58] & in2[58];
    assign P[67] = in[58] ^ in2[58];
    assign G[68] = in[57] & in2[57];
    assign P[68] = in[57] ^ in2[57];
    assign G[69] = in[56] & in2[56];
    assign P[69] = in[56] ^ in2[56];
    assign G[70] = in[55] & in2[55];
    assign P[70] = in[55] ^ in2[55];
    assign G[71] = in[54] & in2[54];
    assign P[71] = in[54] ^ in2[54];
    assign G[72] = in[53] & in2[53];
    assign P[72] = in[53] ^ in2[53];
    assign G[73] = in[52] & in2[52];
    assign P[73] = in[52] ^ in2[52];
    assign G[74] = in[51] & in2[51];
    assign P[74] = in[51] ^ in2[51];
    assign G[75] = in[50] & in2[50];
    assign P[75] = in[50] ^ in2[50];
    assign G[76] = in[49] & in2[49];
    assign P[76] = in[49] ^ in2[49];
    assign G[77] = in[48] & in2[48];
    assign P[77] = in[48] ^ in2[48];
    assign G[78] = in[47] & in2[47];
    assign P[78] = in[47] ^ in2[47];
    assign G[79] = in[46] & in2[46];
    assign P[79] = in[46] ^ in2[46];
    assign G[80] = in[45] & in2[45];
    assign P[80] = in[45] ^ in2[45];
    assign G[81] = in[44] & in2[44];
    assign P[81] = in[44] ^ in2[44];
    assign G[82] = in[43] & in2[43];
    assign P[82] = in[43] ^ in2[43];
    assign G[83] = in[42] & in2[42];
    assign P[83] = in[42] ^ in2[42];
    assign G[84] = in[41] & in2[41];
    assign P[84] = in[41] ^ in2[41];
    assign G[85] = in[40] & in2[40];
    assign P[85] = in[40] ^ in2[40];
    assign G[86] = in[39] & in2[39];
    assign P[86] = in[39] ^ in2[39];
    assign G[87] = in[38] & in2[38];
    assign P[87] = in[38] ^ in2[38];
    assign G[88] = in[37] & in2[37];
    assign P[88] = in[37] ^ in2[37];
    assign G[89] = in[36] & in2[36];
    assign P[89] = in[36] ^ in2[36];
    assign G[90] = in[35] & in2[35];
    assign P[90] = in[35] ^ in2[35];
    assign G[91] = in[34] & in2[34];
    assign P[91] = in[34] ^ in2[34];
    assign G[92] = in[33] & in2[33];
    assign P[92] = in[33] ^ in2[33];
    assign G[93] = in[32] & in2[32];
    assign P[93] = in[32] ^ in2[32];
    assign G[94] = in[31] & in2[31];
    assign P[94] = in[31] ^ in2[31];
    assign G[95] = in[30] & in2[30];
    assign P[95] = in[30] ^ in2[30];
    assign G[96] = in[29] & in2[29];
    assign P[96] = in[29] ^ in2[29];
    assign G[97] = in[28] & in2[28];
    assign P[97] = in[28] ^ in2[28];
    assign G[98] = in[27] & in2[27];
    assign P[98] = in[27] ^ in2[27];
    assign G[99] = in[26] & in2[26];
    assign P[99] = in[26] ^ in2[26];
    assign G[100] = in[25] & in2[25];
    assign P[100] = in[25] ^ in2[25];
    assign G[101] = in[24] & in2[24];
    assign P[101] = in[24] ^ in2[24];
    assign G[102] = in[23] & in2[23];
    assign P[102] = in[23] ^ in2[23];
    assign G[103] = in[22] & in2[22];
    assign P[103] = in[22] ^ in2[22];
    assign G[104] = in[21] & in2[21];
    assign P[104] = in[21] ^ in2[21];
    assign G[105] = in[20] & in2[20];
    assign P[105] = in[20] ^ in2[20];
    assign G[106] = in[19] & in2[19];
    assign P[106] = in[19] ^ in2[19];
    assign G[107] = in[18] & in2[18];
    assign P[107] = in[18] ^ in2[18];
    assign G[108] = in[17] & in2[17];
    assign P[108] = in[17] ^ in2[17];
    assign G[109] = in[16] & in2[16];
    assign P[109] = in[16] ^ in2[16];
    assign G[110] = in[15] & in2[15];
    assign P[110] = in[15] ^ in2[15];
    assign G[111] = in[14] & in2[14];
    assign P[111] = in[14] ^ in2[14];
    assign G[112] = in[13] & in2[13];
    assign P[112] = in[13] ^ in2[13];
    assign G[113] = in[12] & in2[12];
    assign P[113] = in[12] ^ in2[12];
    assign G[114] = in[11] & in2[11];
    assign P[114] = in[11] ^ in2[11];
    assign G[115] = in[10] & in2[10];
    assign P[115] = in[10] ^ in2[10];
    assign G[116] = in[9] & in2[9];
    assign P[116] = in[9] ^ in2[9];
    assign G[117] = in[8] & in2[8];
    assign P[117] = in[8] ^ in2[8];
    assign G[118] = in[7] & in2[7];
    assign P[118] = in[7] ^ in2[7];
    assign G[119] = in[6] & in2[6];
    assign P[119] = in[6] ^ in2[6];
    assign G[120] = in[5] & in2[5];
    assign P[120] = in[5] ^ in2[5];
    assign G[121] = in[4] & in2[4];
    assign P[121] = in[4] ^ in2[4];
    assign G[122] = in[3] & in2[3];
    assign P[122] = in[3] ^ in2[3];
    assign G[123] = in[2] & in2[2];
    assign P[123] = in[2] ^ in2[2];
    assign G[124] = in[1] & in2[1];
    assign P[124] = in[1] ^ in2[1];
    assign G[125] = in[0] & in2[0];
    assign P[125] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign C[125] = G[124] | (P[124] & C[124]);
    assign cout = G[125] | (P[125] & C[125]);
    assign sum = P ^ C;
endmodule

module CLA125(output [124:0] sum, output cout, input [124:0] in1, input [124:0] in2;

    wire[124:0] G;
    wire[124:0] C;
    wire[124:0] P;

    assign G[0] = in[124] & in2[124];
    assign P[0] = in[124] ^ in2[124];
    assign G[1] = in[123] & in2[123];
    assign P[1] = in[123] ^ in2[123];
    assign G[2] = in[122] & in2[122];
    assign P[2] = in[122] ^ in2[122];
    assign G[3] = in[121] & in2[121];
    assign P[3] = in[121] ^ in2[121];
    assign G[4] = in[120] & in2[120];
    assign P[4] = in[120] ^ in2[120];
    assign G[5] = in[119] & in2[119];
    assign P[5] = in[119] ^ in2[119];
    assign G[6] = in[118] & in2[118];
    assign P[6] = in[118] ^ in2[118];
    assign G[7] = in[117] & in2[117];
    assign P[7] = in[117] ^ in2[117];
    assign G[8] = in[116] & in2[116];
    assign P[8] = in[116] ^ in2[116];
    assign G[9] = in[115] & in2[115];
    assign P[9] = in[115] ^ in2[115];
    assign G[10] = in[114] & in2[114];
    assign P[10] = in[114] ^ in2[114];
    assign G[11] = in[113] & in2[113];
    assign P[11] = in[113] ^ in2[113];
    assign G[12] = in[112] & in2[112];
    assign P[12] = in[112] ^ in2[112];
    assign G[13] = in[111] & in2[111];
    assign P[13] = in[111] ^ in2[111];
    assign G[14] = in[110] & in2[110];
    assign P[14] = in[110] ^ in2[110];
    assign G[15] = in[109] & in2[109];
    assign P[15] = in[109] ^ in2[109];
    assign G[16] = in[108] & in2[108];
    assign P[16] = in[108] ^ in2[108];
    assign G[17] = in[107] & in2[107];
    assign P[17] = in[107] ^ in2[107];
    assign G[18] = in[106] & in2[106];
    assign P[18] = in[106] ^ in2[106];
    assign G[19] = in[105] & in2[105];
    assign P[19] = in[105] ^ in2[105];
    assign G[20] = in[104] & in2[104];
    assign P[20] = in[104] ^ in2[104];
    assign G[21] = in[103] & in2[103];
    assign P[21] = in[103] ^ in2[103];
    assign G[22] = in[102] & in2[102];
    assign P[22] = in[102] ^ in2[102];
    assign G[23] = in[101] & in2[101];
    assign P[23] = in[101] ^ in2[101];
    assign G[24] = in[100] & in2[100];
    assign P[24] = in[100] ^ in2[100];
    assign G[25] = in[99] & in2[99];
    assign P[25] = in[99] ^ in2[99];
    assign G[26] = in[98] & in2[98];
    assign P[26] = in[98] ^ in2[98];
    assign G[27] = in[97] & in2[97];
    assign P[27] = in[97] ^ in2[97];
    assign G[28] = in[96] & in2[96];
    assign P[28] = in[96] ^ in2[96];
    assign G[29] = in[95] & in2[95];
    assign P[29] = in[95] ^ in2[95];
    assign G[30] = in[94] & in2[94];
    assign P[30] = in[94] ^ in2[94];
    assign G[31] = in[93] & in2[93];
    assign P[31] = in[93] ^ in2[93];
    assign G[32] = in[92] & in2[92];
    assign P[32] = in[92] ^ in2[92];
    assign G[33] = in[91] & in2[91];
    assign P[33] = in[91] ^ in2[91];
    assign G[34] = in[90] & in2[90];
    assign P[34] = in[90] ^ in2[90];
    assign G[35] = in[89] & in2[89];
    assign P[35] = in[89] ^ in2[89];
    assign G[36] = in[88] & in2[88];
    assign P[36] = in[88] ^ in2[88];
    assign G[37] = in[87] & in2[87];
    assign P[37] = in[87] ^ in2[87];
    assign G[38] = in[86] & in2[86];
    assign P[38] = in[86] ^ in2[86];
    assign G[39] = in[85] & in2[85];
    assign P[39] = in[85] ^ in2[85];
    assign G[40] = in[84] & in2[84];
    assign P[40] = in[84] ^ in2[84];
    assign G[41] = in[83] & in2[83];
    assign P[41] = in[83] ^ in2[83];
    assign G[42] = in[82] & in2[82];
    assign P[42] = in[82] ^ in2[82];
    assign G[43] = in[81] & in2[81];
    assign P[43] = in[81] ^ in2[81];
    assign G[44] = in[80] & in2[80];
    assign P[44] = in[80] ^ in2[80];
    assign G[45] = in[79] & in2[79];
    assign P[45] = in[79] ^ in2[79];
    assign G[46] = in[78] & in2[78];
    assign P[46] = in[78] ^ in2[78];
    assign G[47] = in[77] & in2[77];
    assign P[47] = in[77] ^ in2[77];
    assign G[48] = in[76] & in2[76];
    assign P[48] = in[76] ^ in2[76];
    assign G[49] = in[75] & in2[75];
    assign P[49] = in[75] ^ in2[75];
    assign G[50] = in[74] & in2[74];
    assign P[50] = in[74] ^ in2[74];
    assign G[51] = in[73] & in2[73];
    assign P[51] = in[73] ^ in2[73];
    assign G[52] = in[72] & in2[72];
    assign P[52] = in[72] ^ in2[72];
    assign G[53] = in[71] & in2[71];
    assign P[53] = in[71] ^ in2[71];
    assign G[54] = in[70] & in2[70];
    assign P[54] = in[70] ^ in2[70];
    assign G[55] = in[69] & in2[69];
    assign P[55] = in[69] ^ in2[69];
    assign G[56] = in[68] & in2[68];
    assign P[56] = in[68] ^ in2[68];
    assign G[57] = in[67] & in2[67];
    assign P[57] = in[67] ^ in2[67];
    assign G[58] = in[66] & in2[66];
    assign P[58] = in[66] ^ in2[66];
    assign G[59] = in[65] & in2[65];
    assign P[59] = in[65] ^ in2[65];
    assign G[60] = in[64] & in2[64];
    assign P[60] = in[64] ^ in2[64];
    assign G[61] = in[63] & in2[63];
    assign P[61] = in[63] ^ in2[63];
    assign G[62] = in[62] & in2[62];
    assign P[62] = in[62] ^ in2[62];
    assign G[63] = in[61] & in2[61];
    assign P[63] = in[61] ^ in2[61];
    assign G[64] = in[60] & in2[60];
    assign P[64] = in[60] ^ in2[60];
    assign G[65] = in[59] & in2[59];
    assign P[65] = in[59] ^ in2[59];
    assign G[66] = in[58] & in2[58];
    assign P[66] = in[58] ^ in2[58];
    assign G[67] = in[57] & in2[57];
    assign P[67] = in[57] ^ in2[57];
    assign G[68] = in[56] & in2[56];
    assign P[68] = in[56] ^ in2[56];
    assign G[69] = in[55] & in2[55];
    assign P[69] = in[55] ^ in2[55];
    assign G[70] = in[54] & in2[54];
    assign P[70] = in[54] ^ in2[54];
    assign G[71] = in[53] & in2[53];
    assign P[71] = in[53] ^ in2[53];
    assign G[72] = in[52] & in2[52];
    assign P[72] = in[52] ^ in2[52];
    assign G[73] = in[51] & in2[51];
    assign P[73] = in[51] ^ in2[51];
    assign G[74] = in[50] & in2[50];
    assign P[74] = in[50] ^ in2[50];
    assign G[75] = in[49] & in2[49];
    assign P[75] = in[49] ^ in2[49];
    assign G[76] = in[48] & in2[48];
    assign P[76] = in[48] ^ in2[48];
    assign G[77] = in[47] & in2[47];
    assign P[77] = in[47] ^ in2[47];
    assign G[78] = in[46] & in2[46];
    assign P[78] = in[46] ^ in2[46];
    assign G[79] = in[45] & in2[45];
    assign P[79] = in[45] ^ in2[45];
    assign G[80] = in[44] & in2[44];
    assign P[80] = in[44] ^ in2[44];
    assign G[81] = in[43] & in2[43];
    assign P[81] = in[43] ^ in2[43];
    assign G[82] = in[42] & in2[42];
    assign P[82] = in[42] ^ in2[42];
    assign G[83] = in[41] & in2[41];
    assign P[83] = in[41] ^ in2[41];
    assign G[84] = in[40] & in2[40];
    assign P[84] = in[40] ^ in2[40];
    assign G[85] = in[39] & in2[39];
    assign P[85] = in[39] ^ in2[39];
    assign G[86] = in[38] & in2[38];
    assign P[86] = in[38] ^ in2[38];
    assign G[87] = in[37] & in2[37];
    assign P[87] = in[37] ^ in2[37];
    assign G[88] = in[36] & in2[36];
    assign P[88] = in[36] ^ in2[36];
    assign G[89] = in[35] & in2[35];
    assign P[89] = in[35] ^ in2[35];
    assign G[90] = in[34] & in2[34];
    assign P[90] = in[34] ^ in2[34];
    assign G[91] = in[33] & in2[33];
    assign P[91] = in[33] ^ in2[33];
    assign G[92] = in[32] & in2[32];
    assign P[92] = in[32] ^ in2[32];
    assign G[93] = in[31] & in2[31];
    assign P[93] = in[31] ^ in2[31];
    assign G[94] = in[30] & in2[30];
    assign P[94] = in[30] ^ in2[30];
    assign G[95] = in[29] & in2[29];
    assign P[95] = in[29] ^ in2[29];
    assign G[96] = in[28] & in2[28];
    assign P[96] = in[28] ^ in2[28];
    assign G[97] = in[27] & in2[27];
    assign P[97] = in[27] ^ in2[27];
    assign G[98] = in[26] & in2[26];
    assign P[98] = in[26] ^ in2[26];
    assign G[99] = in[25] & in2[25];
    assign P[99] = in[25] ^ in2[25];
    assign G[100] = in[24] & in2[24];
    assign P[100] = in[24] ^ in2[24];
    assign G[101] = in[23] & in2[23];
    assign P[101] = in[23] ^ in2[23];
    assign G[102] = in[22] & in2[22];
    assign P[102] = in[22] ^ in2[22];
    assign G[103] = in[21] & in2[21];
    assign P[103] = in[21] ^ in2[21];
    assign G[104] = in[20] & in2[20];
    assign P[104] = in[20] ^ in2[20];
    assign G[105] = in[19] & in2[19];
    assign P[105] = in[19] ^ in2[19];
    assign G[106] = in[18] & in2[18];
    assign P[106] = in[18] ^ in2[18];
    assign G[107] = in[17] & in2[17];
    assign P[107] = in[17] ^ in2[17];
    assign G[108] = in[16] & in2[16];
    assign P[108] = in[16] ^ in2[16];
    assign G[109] = in[15] & in2[15];
    assign P[109] = in[15] ^ in2[15];
    assign G[110] = in[14] & in2[14];
    assign P[110] = in[14] ^ in2[14];
    assign G[111] = in[13] & in2[13];
    assign P[111] = in[13] ^ in2[13];
    assign G[112] = in[12] & in2[12];
    assign P[112] = in[12] ^ in2[12];
    assign G[113] = in[11] & in2[11];
    assign P[113] = in[11] ^ in2[11];
    assign G[114] = in[10] & in2[10];
    assign P[114] = in[10] ^ in2[10];
    assign G[115] = in[9] & in2[9];
    assign P[115] = in[9] ^ in2[9];
    assign G[116] = in[8] & in2[8];
    assign P[116] = in[8] ^ in2[8];
    assign G[117] = in[7] & in2[7];
    assign P[117] = in[7] ^ in2[7];
    assign G[118] = in[6] & in2[6];
    assign P[118] = in[6] ^ in2[6];
    assign G[119] = in[5] & in2[5];
    assign P[119] = in[5] ^ in2[5];
    assign G[120] = in[4] & in2[4];
    assign P[120] = in[4] ^ in2[4];
    assign G[121] = in[3] & in2[3];
    assign P[121] = in[3] ^ in2[3];
    assign G[122] = in[2] & in2[2];
    assign P[122] = in[2] ^ in2[2];
    assign G[123] = in[1] & in2[1];
    assign P[123] = in[1] ^ in2[1];
    assign G[124] = in[0] & in2[0];
    assign P[124] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign C[124] = G[123] | (P[123] & C[123]);
    assign cout = G[124] | (P[124] & C[124]);
    assign sum = P ^ C;
endmodule

module CLA124(output [123:0] sum, output cout, input [123:0] in1, input [123:0] in2;

    wire[123:0] G;
    wire[123:0] C;
    wire[123:0] P;

    assign G[0] = in[123] & in2[123];
    assign P[0] = in[123] ^ in2[123];
    assign G[1] = in[122] & in2[122];
    assign P[1] = in[122] ^ in2[122];
    assign G[2] = in[121] & in2[121];
    assign P[2] = in[121] ^ in2[121];
    assign G[3] = in[120] & in2[120];
    assign P[3] = in[120] ^ in2[120];
    assign G[4] = in[119] & in2[119];
    assign P[4] = in[119] ^ in2[119];
    assign G[5] = in[118] & in2[118];
    assign P[5] = in[118] ^ in2[118];
    assign G[6] = in[117] & in2[117];
    assign P[6] = in[117] ^ in2[117];
    assign G[7] = in[116] & in2[116];
    assign P[7] = in[116] ^ in2[116];
    assign G[8] = in[115] & in2[115];
    assign P[8] = in[115] ^ in2[115];
    assign G[9] = in[114] & in2[114];
    assign P[9] = in[114] ^ in2[114];
    assign G[10] = in[113] & in2[113];
    assign P[10] = in[113] ^ in2[113];
    assign G[11] = in[112] & in2[112];
    assign P[11] = in[112] ^ in2[112];
    assign G[12] = in[111] & in2[111];
    assign P[12] = in[111] ^ in2[111];
    assign G[13] = in[110] & in2[110];
    assign P[13] = in[110] ^ in2[110];
    assign G[14] = in[109] & in2[109];
    assign P[14] = in[109] ^ in2[109];
    assign G[15] = in[108] & in2[108];
    assign P[15] = in[108] ^ in2[108];
    assign G[16] = in[107] & in2[107];
    assign P[16] = in[107] ^ in2[107];
    assign G[17] = in[106] & in2[106];
    assign P[17] = in[106] ^ in2[106];
    assign G[18] = in[105] & in2[105];
    assign P[18] = in[105] ^ in2[105];
    assign G[19] = in[104] & in2[104];
    assign P[19] = in[104] ^ in2[104];
    assign G[20] = in[103] & in2[103];
    assign P[20] = in[103] ^ in2[103];
    assign G[21] = in[102] & in2[102];
    assign P[21] = in[102] ^ in2[102];
    assign G[22] = in[101] & in2[101];
    assign P[22] = in[101] ^ in2[101];
    assign G[23] = in[100] & in2[100];
    assign P[23] = in[100] ^ in2[100];
    assign G[24] = in[99] & in2[99];
    assign P[24] = in[99] ^ in2[99];
    assign G[25] = in[98] & in2[98];
    assign P[25] = in[98] ^ in2[98];
    assign G[26] = in[97] & in2[97];
    assign P[26] = in[97] ^ in2[97];
    assign G[27] = in[96] & in2[96];
    assign P[27] = in[96] ^ in2[96];
    assign G[28] = in[95] & in2[95];
    assign P[28] = in[95] ^ in2[95];
    assign G[29] = in[94] & in2[94];
    assign P[29] = in[94] ^ in2[94];
    assign G[30] = in[93] & in2[93];
    assign P[30] = in[93] ^ in2[93];
    assign G[31] = in[92] & in2[92];
    assign P[31] = in[92] ^ in2[92];
    assign G[32] = in[91] & in2[91];
    assign P[32] = in[91] ^ in2[91];
    assign G[33] = in[90] & in2[90];
    assign P[33] = in[90] ^ in2[90];
    assign G[34] = in[89] & in2[89];
    assign P[34] = in[89] ^ in2[89];
    assign G[35] = in[88] & in2[88];
    assign P[35] = in[88] ^ in2[88];
    assign G[36] = in[87] & in2[87];
    assign P[36] = in[87] ^ in2[87];
    assign G[37] = in[86] & in2[86];
    assign P[37] = in[86] ^ in2[86];
    assign G[38] = in[85] & in2[85];
    assign P[38] = in[85] ^ in2[85];
    assign G[39] = in[84] & in2[84];
    assign P[39] = in[84] ^ in2[84];
    assign G[40] = in[83] & in2[83];
    assign P[40] = in[83] ^ in2[83];
    assign G[41] = in[82] & in2[82];
    assign P[41] = in[82] ^ in2[82];
    assign G[42] = in[81] & in2[81];
    assign P[42] = in[81] ^ in2[81];
    assign G[43] = in[80] & in2[80];
    assign P[43] = in[80] ^ in2[80];
    assign G[44] = in[79] & in2[79];
    assign P[44] = in[79] ^ in2[79];
    assign G[45] = in[78] & in2[78];
    assign P[45] = in[78] ^ in2[78];
    assign G[46] = in[77] & in2[77];
    assign P[46] = in[77] ^ in2[77];
    assign G[47] = in[76] & in2[76];
    assign P[47] = in[76] ^ in2[76];
    assign G[48] = in[75] & in2[75];
    assign P[48] = in[75] ^ in2[75];
    assign G[49] = in[74] & in2[74];
    assign P[49] = in[74] ^ in2[74];
    assign G[50] = in[73] & in2[73];
    assign P[50] = in[73] ^ in2[73];
    assign G[51] = in[72] & in2[72];
    assign P[51] = in[72] ^ in2[72];
    assign G[52] = in[71] & in2[71];
    assign P[52] = in[71] ^ in2[71];
    assign G[53] = in[70] & in2[70];
    assign P[53] = in[70] ^ in2[70];
    assign G[54] = in[69] & in2[69];
    assign P[54] = in[69] ^ in2[69];
    assign G[55] = in[68] & in2[68];
    assign P[55] = in[68] ^ in2[68];
    assign G[56] = in[67] & in2[67];
    assign P[56] = in[67] ^ in2[67];
    assign G[57] = in[66] & in2[66];
    assign P[57] = in[66] ^ in2[66];
    assign G[58] = in[65] & in2[65];
    assign P[58] = in[65] ^ in2[65];
    assign G[59] = in[64] & in2[64];
    assign P[59] = in[64] ^ in2[64];
    assign G[60] = in[63] & in2[63];
    assign P[60] = in[63] ^ in2[63];
    assign G[61] = in[62] & in2[62];
    assign P[61] = in[62] ^ in2[62];
    assign G[62] = in[61] & in2[61];
    assign P[62] = in[61] ^ in2[61];
    assign G[63] = in[60] & in2[60];
    assign P[63] = in[60] ^ in2[60];
    assign G[64] = in[59] & in2[59];
    assign P[64] = in[59] ^ in2[59];
    assign G[65] = in[58] & in2[58];
    assign P[65] = in[58] ^ in2[58];
    assign G[66] = in[57] & in2[57];
    assign P[66] = in[57] ^ in2[57];
    assign G[67] = in[56] & in2[56];
    assign P[67] = in[56] ^ in2[56];
    assign G[68] = in[55] & in2[55];
    assign P[68] = in[55] ^ in2[55];
    assign G[69] = in[54] & in2[54];
    assign P[69] = in[54] ^ in2[54];
    assign G[70] = in[53] & in2[53];
    assign P[70] = in[53] ^ in2[53];
    assign G[71] = in[52] & in2[52];
    assign P[71] = in[52] ^ in2[52];
    assign G[72] = in[51] & in2[51];
    assign P[72] = in[51] ^ in2[51];
    assign G[73] = in[50] & in2[50];
    assign P[73] = in[50] ^ in2[50];
    assign G[74] = in[49] & in2[49];
    assign P[74] = in[49] ^ in2[49];
    assign G[75] = in[48] & in2[48];
    assign P[75] = in[48] ^ in2[48];
    assign G[76] = in[47] & in2[47];
    assign P[76] = in[47] ^ in2[47];
    assign G[77] = in[46] & in2[46];
    assign P[77] = in[46] ^ in2[46];
    assign G[78] = in[45] & in2[45];
    assign P[78] = in[45] ^ in2[45];
    assign G[79] = in[44] & in2[44];
    assign P[79] = in[44] ^ in2[44];
    assign G[80] = in[43] & in2[43];
    assign P[80] = in[43] ^ in2[43];
    assign G[81] = in[42] & in2[42];
    assign P[81] = in[42] ^ in2[42];
    assign G[82] = in[41] & in2[41];
    assign P[82] = in[41] ^ in2[41];
    assign G[83] = in[40] & in2[40];
    assign P[83] = in[40] ^ in2[40];
    assign G[84] = in[39] & in2[39];
    assign P[84] = in[39] ^ in2[39];
    assign G[85] = in[38] & in2[38];
    assign P[85] = in[38] ^ in2[38];
    assign G[86] = in[37] & in2[37];
    assign P[86] = in[37] ^ in2[37];
    assign G[87] = in[36] & in2[36];
    assign P[87] = in[36] ^ in2[36];
    assign G[88] = in[35] & in2[35];
    assign P[88] = in[35] ^ in2[35];
    assign G[89] = in[34] & in2[34];
    assign P[89] = in[34] ^ in2[34];
    assign G[90] = in[33] & in2[33];
    assign P[90] = in[33] ^ in2[33];
    assign G[91] = in[32] & in2[32];
    assign P[91] = in[32] ^ in2[32];
    assign G[92] = in[31] & in2[31];
    assign P[92] = in[31] ^ in2[31];
    assign G[93] = in[30] & in2[30];
    assign P[93] = in[30] ^ in2[30];
    assign G[94] = in[29] & in2[29];
    assign P[94] = in[29] ^ in2[29];
    assign G[95] = in[28] & in2[28];
    assign P[95] = in[28] ^ in2[28];
    assign G[96] = in[27] & in2[27];
    assign P[96] = in[27] ^ in2[27];
    assign G[97] = in[26] & in2[26];
    assign P[97] = in[26] ^ in2[26];
    assign G[98] = in[25] & in2[25];
    assign P[98] = in[25] ^ in2[25];
    assign G[99] = in[24] & in2[24];
    assign P[99] = in[24] ^ in2[24];
    assign G[100] = in[23] & in2[23];
    assign P[100] = in[23] ^ in2[23];
    assign G[101] = in[22] & in2[22];
    assign P[101] = in[22] ^ in2[22];
    assign G[102] = in[21] & in2[21];
    assign P[102] = in[21] ^ in2[21];
    assign G[103] = in[20] & in2[20];
    assign P[103] = in[20] ^ in2[20];
    assign G[104] = in[19] & in2[19];
    assign P[104] = in[19] ^ in2[19];
    assign G[105] = in[18] & in2[18];
    assign P[105] = in[18] ^ in2[18];
    assign G[106] = in[17] & in2[17];
    assign P[106] = in[17] ^ in2[17];
    assign G[107] = in[16] & in2[16];
    assign P[107] = in[16] ^ in2[16];
    assign G[108] = in[15] & in2[15];
    assign P[108] = in[15] ^ in2[15];
    assign G[109] = in[14] & in2[14];
    assign P[109] = in[14] ^ in2[14];
    assign G[110] = in[13] & in2[13];
    assign P[110] = in[13] ^ in2[13];
    assign G[111] = in[12] & in2[12];
    assign P[111] = in[12] ^ in2[12];
    assign G[112] = in[11] & in2[11];
    assign P[112] = in[11] ^ in2[11];
    assign G[113] = in[10] & in2[10];
    assign P[113] = in[10] ^ in2[10];
    assign G[114] = in[9] & in2[9];
    assign P[114] = in[9] ^ in2[9];
    assign G[115] = in[8] & in2[8];
    assign P[115] = in[8] ^ in2[8];
    assign G[116] = in[7] & in2[7];
    assign P[116] = in[7] ^ in2[7];
    assign G[117] = in[6] & in2[6];
    assign P[117] = in[6] ^ in2[6];
    assign G[118] = in[5] & in2[5];
    assign P[118] = in[5] ^ in2[5];
    assign G[119] = in[4] & in2[4];
    assign P[119] = in[4] ^ in2[4];
    assign G[120] = in[3] & in2[3];
    assign P[120] = in[3] ^ in2[3];
    assign G[121] = in[2] & in2[2];
    assign P[121] = in[2] ^ in2[2];
    assign G[122] = in[1] & in2[1];
    assign P[122] = in[1] ^ in2[1];
    assign G[123] = in[0] & in2[0];
    assign P[123] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign C[123] = G[122] | (P[122] & C[122]);
    assign cout = G[123] | (P[123] & C[123]);
    assign sum = P ^ C;
endmodule

module CLA123(output [122:0] sum, output cout, input [122:0] in1, input [122:0] in2;

    wire[122:0] G;
    wire[122:0] C;
    wire[122:0] P;

    assign G[0] = in[122] & in2[122];
    assign P[0] = in[122] ^ in2[122];
    assign G[1] = in[121] & in2[121];
    assign P[1] = in[121] ^ in2[121];
    assign G[2] = in[120] & in2[120];
    assign P[2] = in[120] ^ in2[120];
    assign G[3] = in[119] & in2[119];
    assign P[3] = in[119] ^ in2[119];
    assign G[4] = in[118] & in2[118];
    assign P[4] = in[118] ^ in2[118];
    assign G[5] = in[117] & in2[117];
    assign P[5] = in[117] ^ in2[117];
    assign G[6] = in[116] & in2[116];
    assign P[6] = in[116] ^ in2[116];
    assign G[7] = in[115] & in2[115];
    assign P[7] = in[115] ^ in2[115];
    assign G[8] = in[114] & in2[114];
    assign P[8] = in[114] ^ in2[114];
    assign G[9] = in[113] & in2[113];
    assign P[9] = in[113] ^ in2[113];
    assign G[10] = in[112] & in2[112];
    assign P[10] = in[112] ^ in2[112];
    assign G[11] = in[111] & in2[111];
    assign P[11] = in[111] ^ in2[111];
    assign G[12] = in[110] & in2[110];
    assign P[12] = in[110] ^ in2[110];
    assign G[13] = in[109] & in2[109];
    assign P[13] = in[109] ^ in2[109];
    assign G[14] = in[108] & in2[108];
    assign P[14] = in[108] ^ in2[108];
    assign G[15] = in[107] & in2[107];
    assign P[15] = in[107] ^ in2[107];
    assign G[16] = in[106] & in2[106];
    assign P[16] = in[106] ^ in2[106];
    assign G[17] = in[105] & in2[105];
    assign P[17] = in[105] ^ in2[105];
    assign G[18] = in[104] & in2[104];
    assign P[18] = in[104] ^ in2[104];
    assign G[19] = in[103] & in2[103];
    assign P[19] = in[103] ^ in2[103];
    assign G[20] = in[102] & in2[102];
    assign P[20] = in[102] ^ in2[102];
    assign G[21] = in[101] & in2[101];
    assign P[21] = in[101] ^ in2[101];
    assign G[22] = in[100] & in2[100];
    assign P[22] = in[100] ^ in2[100];
    assign G[23] = in[99] & in2[99];
    assign P[23] = in[99] ^ in2[99];
    assign G[24] = in[98] & in2[98];
    assign P[24] = in[98] ^ in2[98];
    assign G[25] = in[97] & in2[97];
    assign P[25] = in[97] ^ in2[97];
    assign G[26] = in[96] & in2[96];
    assign P[26] = in[96] ^ in2[96];
    assign G[27] = in[95] & in2[95];
    assign P[27] = in[95] ^ in2[95];
    assign G[28] = in[94] & in2[94];
    assign P[28] = in[94] ^ in2[94];
    assign G[29] = in[93] & in2[93];
    assign P[29] = in[93] ^ in2[93];
    assign G[30] = in[92] & in2[92];
    assign P[30] = in[92] ^ in2[92];
    assign G[31] = in[91] & in2[91];
    assign P[31] = in[91] ^ in2[91];
    assign G[32] = in[90] & in2[90];
    assign P[32] = in[90] ^ in2[90];
    assign G[33] = in[89] & in2[89];
    assign P[33] = in[89] ^ in2[89];
    assign G[34] = in[88] & in2[88];
    assign P[34] = in[88] ^ in2[88];
    assign G[35] = in[87] & in2[87];
    assign P[35] = in[87] ^ in2[87];
    assign G[36] = in[86] & in2[86];
    assign P[36] = in[86] ^ in2[86];
    assign G[37] = in[85] & in2[85];
    assign P[37] = in[85] ^ in2[85];
    assign G[38] = in[84] & in2[84];
    assign P[38] = in[84] ^ in2[84];
    assign G[39] = in[83] & in2[83];
    assign P[39] = in[83] ^ in2[83];
    assign G[40] = in[82] & in2[82];
    assign P[40] = in[82] ^ in2[82];
    assign G[41] = in[81] & in2[81];
    assign P[41] = in[81] ^ in2[81];
    assign G[42] = in[80] & in2[80];
    assign P[42] = in[80] ^ in2[80];
    assign G[43] = in[79] & in2[79];
    assign P[43] = in[79] ^ in2[79];
    assign G[44] = in[78] & in2[78];
    assign P[44] = in[78] ^ in2[78];
    assign G[45] = in[77] & in2[77];
    assign P[45] = in[77] ^ in2[77];
    assign G[46] = in[76] & in2[76];
    assign P[46] = in[76] ^ in2[76];
    assign G[47] = in[75] & in2[75];
    assign P[47] = in[75] ^ in2[75];
    assign G[48] = in[74] & in2[74];
    assign P[48] = in[74] ^ in2[74];
    assign G[49] = in[73] & in2[73];
    assign P[49] = in[73] ^ in2[73];
    assign G[50] = in[72] & in2[72];
    assign P[50] = in[72] ^ in2[72];
    assign G[51] = in[71] & in2[71];
    assign P[51] = in[71] ^ in2[71];
    assign G[52] = in[70] & in2[70];
    assign P[52] = in[70] ^ in2[70];
    assign G[53] = in[69] & in2[69];
    assign P[53] = in[69] ^ in2[69];
    assign G[54] = in[68] & in2[68];
    assign P[54] = in[68] ^ in2[68];
    assign G[55] = in[67] & in2[67];
    assign P[55] = in[67] ^ in2[67];
    assign G[56] = in[66] & in2[66];
    assign P[56] = in[66] ^ in2[66];
    assign G[57] = in[65] & in2[65];
    assign P[57] = in[65] ^ in2[65];
    assign G[58] = in[64] & in2[64];
    assign P[58] = in[64] ^ in2[64];
    assign G[59] = in[63] & in2[63];
    assign P[59] = in[63] ^ in2[63];
    assign G[60] = in[62] & in2[62];
    assign P[60] = in[62] ^ in2[62];
    assign G[61] = in[61] & in2[61];
    assign P[61] = in[61] ^ in2[61];
    assign G[62] = in[60] & in2[60];
    assign P[62] = in[60] ^ in2[60];
    assign G[63] = in[59] & in2[59];
    assign P[63] = in[59] ^ in2[59];
    assign G[64] = in[58] & in2[58];
    assign P[64] = in[58] ^ in2[58];
    assign G[65] = in[57] & in2[57];
    assign P[65] = in[57] ^ in2[57];
    assign G[66] = in[56] & in2[56];
    assign P[66] = in[56] ^ in2[56];
    assign G[67] = in[55] & in2[55];
    assign P[67] = in[55] ^ in2[55];
    assign G[68] = in[54] & in2[54];
    assign P[68] = in[54] ^ in2[54];
    assign G[69] = in[53] & in2[53];
    assign P[69] = in[53] ^ in2[53];
    assign G[70] = in[52] & in2[52];
    assign P[70] = in[52] ^ in2[52];
    assign G[71] = in[51] & in2[51];
    assign P[71] = in[51] ^ in2[51];
    assign G[72] = in[50] & in2[50];
    assign P[72] = in[50] ^ in2[50];
    assign G[73] = in[49] & in2[49];
    assign P[73] = in[49] ^ in2[49];
    assign G[74] = in[48] & in2[48];
    assign P[74] = in[48] ^ in2[48];
    assign G[75] = in[47] & in2[47];
    assign P[75] = in[47] ^ in2[47];
    assign G[76] = in[46] & in2[46];
    assign P[76] = in[46] ^ in2[46];
    assign G[77] = in[45] & in2[45];
    assign P[77] = in[45] ^ in2[45];
    assign G[78] = in[44] & in2[44];
    assign P[78] = in[44] ^ in2[44];
    assign G[79] = in[43] & in2[43];
    assign P[79] = in[43] ^ in2[43];
    assign G[80] = in[42] & in2[42];
    assign P[80] = in[42] ^ in2[42];
    assign G[81] = in[41] & in2[41];
    assign P[81] = in[41] ^ in2[41];
    assign G[82] = in[40] & in2[40];
    assign P[82] = in[40] ^ in2[40];
    assign G[83] = in[39] & in2[39];
    assign P[83] = in[39] ^ in2[39];
    assign G[84] = in[38] & in2[38];
    assign P[84] = in[38] ^ in2[38];
    assign G[85] = in[37] & in2[37];
    assign P[85] = in[37] ^ in2[37];
    assign G[86] = in[36] & in2[36];
    assign P[86] = in[36] ^ in2[36];
    assign G[87] = in[35] & in2[35];
    assign P[87] = in[35] ^ in2[35];
    assign G[88] = in[34] & in2[34];
    assign P[88] = in[34] ^ in2[34];
    assign G[89] = in[33] & in2[33];
    assign P[89] = in[33] ^ in2[33];
    assign G[90] = in[32] & in2[32];
    assign P[90] = in[32] ^ in2[32];
    assign G[91] = in[31] & in2[31];
    assign P[91] = in[31] ^ in2[31];
    assign G[92] = in[30] & in2[30];
    assign P[92] = in[30] ^ in2[30];
    assign G[93] = in[29] & in2[29];
    assign P[93] = in[29] ^ in2[29];
    assign G[94] = in[28] & in2[28];
    assign P[94] = in[28] ^ in2[28];
    assign G[95] = in[27] & in2[27];
    assign P[95] = in[27] ^ in2[27];
    assign G[96] = in[26] & in2[26];
    assign P[96] = in[26] ^ in2[26];
    assign G[97] = in[25] & in2[25];
    assign P[97] = in[25] ^ in2[25];
    assign G[98] = in[24] & in2[24];
    assign P[98] = in[24] ^ in2[24];
    assign G[99] = in[23] & in2[23];
    assign P[99] = in[23] ^ in2[23];
    assign G[100] = in[22] & in2[22];
    assign P[100] = in[22] ^ in2[22];
    assign G[101] = in[21] & in2[21];
    assign P[101] = in[21] ^ in2[21];
    assign G[102] = in[20] & in2[20];
    assign P[102] = in[20] ^ in2[20];
    assign G[103] = in[19] & in2[19];
    assign P[103] = in[19] ^ in2[19];
    assign G[104] = in[18] & in2[18];
    assign P[104] = in[18] ^ in2[18];
    assign G[105] = in[17] & in2[17];
    assign P[105] = in[17] ^ in2[17];
    assign G[106] = in[16] & in2[16];
    assign P[106] = in[16] ^ in2[16];
    assign G[107] = in[15] & in2[15];
    assign P[107] = in[15] ^ in2[15];
    assign G[108] = in[14] & in2[14];
    assign P[108] = in[14] ^ in2[14];
    assign G[109] = in[13] & in2[13];
    assign P[109] = in[13] ^ in2[13];
    assign G[110] = in[12] & in2[12];
    assign P[110] = in[12] ^ in2[12];
    assign G[111] = in[11] & in2[11];
    assign P[111] = in[11] ^ in2[11];
    assign G[112] = in[10] & in2[10];
    assign P[112] = in[10] ^ in2[10];
    assign G[113] = in[9] & in2[9];
    assign P[113] = in[9] ^ in2[9];
    assign G[114] = in[8] & in2[8];
    assign P[114] = in[8] ^ in2[8];
    assign G[115] = in[7] & in2[7];
    assign P[115] = in[7] ^ in2[7];
    assign G[116] = in[6] & in2[6];
    assign P[116] = in[6] ^ in2[6];
    assign G[117] = in[5] & in2[5];
    assign P[117] = in[5] ^ in2[5];
    assign G[118] = in[4] & in2[4];
    assign P[118] = in[4] ^ in2[4];
    assign G[119] = in[3] & in2[3];
    assign P[119] = in[3] ^ in2[3];
    assign G[120] = in[2] & in2[2];
    assign P[120] = in[2] ^ in2[2];
    assign G[121] = in[1] & in2[1];
    assign P[121] = in[1] ^ in2[1];
    assign G[122] = in[0] & in2[0];
    assign P[122] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign C[122] = G[121] | (P[121] & C[121]);
    assign cout = G[122] | (P[122] & C[122]);
    assign sum = P ^ C;
endmodule

module CLA122(output [121:0] sum, output cout, input [121:0] in1, input [121:0] in2;

    wire[121:0] G;
    wire[121:0] C;
    wire[121:0] P;

    assign G[0] = in[121] & in2[121];
    assign P[0] = in[121] ^ in2[121];
    assign G[1] = in[120] & in2[120];
    assign P[1] = in[120] ^ in2[120];
    assign G[2] = in[119] & in2[119];
    assign P[2] = in[119] ^ in2[119];
    assign G[3] = in[118] & in2[118];
    assign P[3] = in[118] ^ in2[118];
    assign G[4] = in[117] & in2[117];
    assign P[4] = in[117] ^ in2[117];
    assign G[5] = in[116] & in2[116];
    assign P[5] = in[116] ^ in2[116];
    assign G[6] = in[115] & in2[115];
    assign P[6] = in[115] ^ in2[115];
    assign G[7] = in[114] & in2[114];
    assign P[7] = in[114] ^ in2[114];
    assign G[8] = in[113] & in2[113];
    assign P[8] = in[113] ^ in2[113];
    assign G[9] = in[112] & in2[112];
    assign P[9] = in[112] ^ in2[112];
    assign G[10] = in[111] & in2[111];
    assign P[10] = in[111] ^ in2[111];
    assign G[11] = in[110] & in2[110];
    assign P[11] = in[110] ^ in2[110];
    assign G[12] = in[109] & in2[109];
    assign P[12] = in[109] ^ in2[109];
    assign G[13] = in[108] & in2[108];
    assign P[13] = in[108] ^ in2[108];
    assign G[14] = in[107] & in2[107];
    assign P[14] = in[107] ^ in2[107];
    assign G[15] = in[106] & in2[106];
    assign P[15] = in[106] ^ in2[106];
    assign G[16] = in[105] & in2[105];
    assign P[16] = in[105] ^ in2[105];
    assign G[17] = in[104] & in2[104];
    assign P[17] = in[104] ^ in2[104];
    assign G[18] = in[103] & in2[103];
    assign P[18] = in[103] ^ in2[103];
    assign G[19] = in[102] & in2[102];
    assign P[19] = in[102] ^ in2[102];
    assign G[20] = in[101] & in2[101];
    assign P[20] = in[101] ^ in2[101];
    assign G[21] = in[100] & in2[100];
    assign P[21] = in[100] ^ in2[100];
    assign G[22] = in[99] & in2[99];
    assign P[22] = in[99] ^ in2[99];
    assign G[23] = in[98] & in2[98];
    assign P[23] = in[98] ^ in2[98];
    assign G[24] = in[97] & in2[97];
    assign P[24] = in[97] ^ in2[97];
    assign G[25] = in[96] & in2[96];
    assign P[25] = in[96] ^ in2[96];
    assign G[26] = in[95] & in2[95];
    assign P[26] = in[95] ^ in2[95];
    assign G[27] = in[94] & in2[94];
    assign P[27] = in[94] ^ in2[94];
    assign G[28] = in[93] & in2[93];
    assign P[28] = in[93] ^ in2[93];
    assign G[29] = in[92] & in2[92];
    assign P[29] = in[92] ^ in2[92];
    assign G[30] = in[91] & in2[91];
    assign P[30] = in[91] ^ in2[91];
    assign G[31] = in[90] & in2[90];
    assign P[31] = in[90] ^ in2[90];
    assign G[32] = in[89] & in2[89];
    assign P[32] = in[89] ^ in2[89];
    assign G[33] = in[88] & in2[88];
    assign P[33] = in[88] ^ in2[88];
    assign G[34] = in[87] & in2[87];
    assign P[34] = in[87] ^ in2[87];
    assign G[35] = in[86] & in2[86];
    assign P[35] = in[86] ^ in2[86];
    assign G[36] = in[85] & in2[85];
    assign P[36] = in[85] ^ in2[85];
    assign G[37] = in[84] & in2[84];
    assign P[37] = in[84] ^ in2[84];
    assign G[38] = in[83] & in2[83];
    assign P[38] = in[83] ^ in2[83];
    assign G[39] = in[82] & in2[82];
    assign P[39] = in[82] ^ in2[82];
    assign G[40] = in[81] & in2[81];
    assign P[40] = in[81] ^ in2[81];
    assign G[41] = in[80] & in2[80];
    assign P[41] = in[80] ^ in2[80];
    assign G[42] = in[79] & in2[79];
    assign P[42] = in[79] ^ in2[79];
    assign G[43] = in[78] & in2[78];
    assign P[43] = in[78] ^ in2[78];
    assign G[44] = in[77] & in2[77];
    assign P[44] = in[77] ^ in2[77];
    assign G[45] = in[76] & in2[76];
    assign P[45] = in[76] ^ in2[76];
    assign G[46] = in[75] & in2[75];
    assign P[46] = in[75] ^ in2[75];
    assign G[47] = in[74] & in2[74];
    assign P[47] = in[74] ^ in2[74];
    assign G[48] = in[73] & in2[73];
    assign P[48] = in[73] ^ in2[73];
    assign G[49] = in[72] & in2[72];
    assign P[49] = in[72] ^ in2[72];
    assign G[50] = in[71] & in2[71];
    assign P[50] = in[71] ^ in2[71];
    assign G[51] = in[70] & in2[70];
    assign P[51] = in[70] ^ in2[70];
    assign G[52] = in[69] & in2[69];
    assign P[52] = in[69] ^ in2[69];
    assign G[53] = in[68] & in2[68];
    assign P[53] = in[68] ^ in2[68];
    assign G[54] = in[67] & in2[67];
    assign P[54] = in[67] ^ in2[67];
    assign G[55] = in[66] & in2[66];
    assign P[55] = in[66] ^ in2[66];
    assign G[56] = in[65] & in2[65];
    assign P[56] = in[65] ^ in2[65];
    assign G[57] = in[64] & in2[64];
    assign P[57] = in[64] ^ in2[64];
    assign G[58] = in[63] & in2[63];
    assign P[58] = in[63] ^ in2[63];
    assign G[59] = in[62] & in2[62];
    assign P[59] = in[62] ^ in2[62];
    assign G[60] = in[61] & in2[61];
    assign P[60] = in[61] ^ in2[61];
    assign G[61] = in[60] & in2[60];
    assign P[61] = in[60] ^ in2[60];
    assign G[62] = in[59] & in2[59];
    assign P[62] = in[59] ^ in2[59];
    assign G[63] = in[58] & in2[58];
    assign P[63] = in[58] ^ in2[58];
    assign G[64] = in[57] & in2[57];
    assign P[64] = in[57] ^ in2[57];
    assign G[65] = in[56] & in2[56];
    assign P[65] = in[56] ^ in2[56];
    assign G[66] = in[55] & in2[55];
    assign P[66] = in[55] ^ in2[55];
    assign G[67] = in[54] & in2[54];
    assign P[67] = in[54] ^ in2[54];
    assign G[68] = in[53] & in2[53];
    assign P[68] = in[53] ^ in2[53];
    assign G[69] = in[52] & in2[52];
    assign P[69] = in[52] ^ in2[52];
    assign G[70] = in[51] & in2[51];
    assign P[70] = in[51] ^ in2[51];
    assign G[71] = in[50] & in2[50];
    assign P[71] = in[50] ^ in2[50];
    assign G[72] = in[49] & in2[49];
    assign P[72] = in[49] ^ in2[49];
    assign G[73] = in[48] & in2[48];
    assign P[73] = in[48] ^ in2[48];
    assign G[74] = in[47] & in2[47];
    assign P[74] = in[47] ^ in2[47];
    assign G[75] = in[46] & in2[46];
    assign P[75] = in[46] ^ in2[46];
    assign G[76] = in[45] & in2[45];
    assign P[76] = in[45] ^ in2[45];
    assign G[77] = in[44] & in2[44];
    assign P[77] = in[44] ^ in2[44];
    assign G[78] = in[43] & in2[43];
    assign P[78] = in[43] ^ in2[43];
    assign G[79] = in[42] & in2[42];
    assign P[79] = in[42] ^ in2[42];
    assign G[80] = in[41] & in2[41];
    assign P[80] = in[41] ^ in2[41];
    assign G[81] = in[40] & in2[40];
    assign P[81] = in[40] ^ in2[40];
    assign G[82] = in[39] & in2[39];
    assign P[82] = in[39] ^ in2[39];
    assign G[83] = in[38] & in2[38];
    assign P[83] = in[38] ^ in2[38];
    assign G[84] = in[37] & in2[37];
    assign P[84] = in[37] ^ in2[37];
    assign G[85] = in[36] & in2[36];
    assign P[85] = in[36] ^ in2[36];
    assign G[86] = in[35] & in2[35];
    assign P[86] = in[35] ^ in2[35];
    assign G[87] = in[34] & in2[34];
    assign P[87] = in[34] ^ in2[34];
    assign G[88] = in[33] & in2[33];
    assign P[88] = in[33] ^ in2[33];
    assign G[89] = in[32] & in2[32];
    assign P[89] = in[32] ^ in2[32];
    assign G[90] = in[31] & in2[31];
    assign P[90] = in[31] ^ in2[31];
    assign G[91] = in[30] & in2[30];
    assign P[91] = in[30] ^ in2[30];
    assign G[92] = in[29] & in2[29];
    assign P[92] = in[29] ^ in2[29];
    assign G[93] = in[28] & in2[28];
    assign P[93] = in[28] ^ in2[28];
    assign G[94] = in[27] & in2[27];
    assign P[94] = in[27] ^ in2[27];
    assign G[95] = in[26] & in2[26];
    assign P[95] = in[26] ^ in2[26];
    assign G[96] = in[25] & in2[25];
    assign P[96] = in[25] ^ in2[25];
    assign G[97] = in[24] & in2[24];
    assign P[97] = in[24] ^ in2[24];
    assign G[98] = in[23] & in2[23];
    assign P[98] = in[23] ^ in2[23];
    assign G[99] = in[22] & in2[22];
    assign P[99] = in[22] ^ in2[22];
    assign G[100] = in[21] & in2[21];
    assign P[100] = in[21] ^ in2[21];
    assign G[101] = in[20] & in2[20];
    assign P[101] = in[20] ^ in2[20];
    assign G[102] = in[19] & in2[19];
    assign P[102] = in[19] ^ in2[19];
    assign G[103] = in[18] & in2[18];
    assign P[103] = in[18] ^ in2[18];
    assign G[104] = in[17] & in2[17];
    assign P[104] = in[17] ^ in2[17];
    assign G[105] = in[16] & in2[16];
    assign P[105] = in[16] ^ in2[16];
    assign G[106] = in[15] & in2[15];
    assign P[106] = in[15] ^ in2[15];
    assign G[107] = in[14] & in2[14];
    assign P[107] = in[14] ^ in2[14];
    assign G[108] = in[13] & in2[13];
    assign P[108] = in[13] ^ in2[13];
    assign G[109] = in[12] & in2[12];
    assign P[109] = in[12] ^ in2[12];
    assign G[110] = in[11] & in2[11];
    assign P[110] = in[11] ^ in2[11];
    assign G[111] = in[10] & in2[10];
    assign P[111] = in[10] ^ in2[10];
    assign G[112] = in[9] & in2[9];
    assign P[112] = in[9] ^ in2[9];
    assign G[113] = in[8] & in2[8];
    assign P[113] = in[8] ^ in2[8];
    assign G[114] = in[7] & in2[7];
    assign P[114] = in[7] ^ in2[7];
    assign G[115] = in[6] & in2[6];
    assign P[115] = in[6] ^ in2[6];
    assign G[116] = in[5] & in2[5];
    assign P[116] = in[5] ^ in2[5];
    assign G[117] = in[4] & in2[4];
    assign P[117] = in[4] ^ in2[4];
    assign G[118] = in[3] & in2[3];
    assign P[118] = in[3] ^ in2[3];
    assign G[119] = in[2] & in2[2];
    assign P[119] = in[2] ^ in2[2];
    assign G[120] = in[1] & in2[1];
    assign P[120] = in[1] ^ in2[1];
    assign G[121] = in[0] & in2[0];
    assign P[121] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign C[121] = G[120] | (P[120] & C[120]);
    assign cout = G[121] | (P[121] & C[121]);
    assign sum = P ^ C;
endmodule

module CLA121(output [120:0] sum, output cout, input [120:0] in1, input [120:0] in2;

    wire[120:0] G;
    wire[120:0] C;
    wire[120:0] P;

    assign G[0] = in[120] & in2[120];
    assign P[0] = in[120] ^ in2[120];
    assign G[1] = in[119] & in2[119];
    assign P[1] = in[119] ^ in2[119];
    assign G[2] = in[118] & in2[118];
    assign P[2] = in[118] ^ in2[118];
    assign G[3] = in[117] & in2[117];
    assign P[3] = in[117] ^ in2[117];
    assign G[4] = in[116] & in2[116];
    assign P[4] = in[116] ^ in2[116];
    assign G[5] = in[115] & in2[115];
    assign P[5] = in[115] ^ in2[115];
    assign G[6] = in[114] & in2[114];
    assign P[6] = in[114] ^ in2[114];
    assign G[7] = in[113] & in2[113];
    assign P[7] = in[113] ^ in2[113];
    assign G[8] = in[112] & in2[112];
    assign P[8] = in[112] ^ in2[112];
    assign G[9] = in[111] & in2[111];
    assign P[9] = in[111] ^ in2[111];
    assign G[10] = in[110] & in2[110];
    assign P[10] = in[110] ^ in2[110];
    assign G[11] = in[109] & in2[109];
    assign P[11] = in[109] ^ in2[109];
    assign G[12] = in[108] & in2[108];
    assign P[12] = in[108] ^ in2[108];
    assign G[13] = in[107] & in2[107];
    assign P[13] = in[107] ^ in2[107];
    assign G[14] = in[106] & in2[106];
    assign P[14] = in[106] ^ in2[106];
    assign G[15] = in[105] & in2[105];
    assign P[15] = in[105] ^ in2[105];
    assign G[16] = in[104] & in2[104];
    assign P[16] = in[104] ^ in2[104];
    assign G[17] = in[103] & in2[103];
    assign P[17] = in[103] ^ in2[103];
    assign G[18] = in[102] & in2[102];
    assign P[18] = in[102] ^ in2[102];
    assign G[19] = in[101] & in2[101];
    assign P[19] = in[101] ^ in2[101];
    assign G[20] = in[100] & in2[100];
    assign P[20] = in[100] ^ in2[100];
    assign G[21] = in[99] & in2[99];
    assign P[21] = in[99] ^ in2[99];
    assign G[22] = in[98] & in2[98];
    assign P[22] = in[98] ^ in2[98];
    assign G[23] = in[97] & in2[97];
    assign P[23] = in[97] ^ in2[97];
    assign G[24] = in[96] & in2[96];
    assign P[24] = in[96] ^ in2[96];
    assign G[25] = in[95] & in2[95];
    assign P[25] = in[95] ^ in2[95];
    assign G[26] = in[94] & in2[94];
    assign P[26] = in[94] ^ in2[94];
    assign G[27] = in[93] & in2[93];
    assign P[27] = in[93] ^ in2[93];
    assign G[28] = in[92] & in2[92];
    assign P[28] = in[92] ^ in2[92];
    assign G[29] = in[91] & in2[91];
    assign P[29] = in[91] ^ in2[91];
    assign G[30] = in[90] & in2[90];
    assign P[30] = in[90] ^ in2[90];
    assign G[31] = in[89] & in2[89];
    assign P[31] = in[89] ^ in2[89];
    assign G[32] = in[88] & in2[88];
    assign P[32] = in[88] ^ in2[88];
    assign G[33] = in[87] & in2[87];
    assign P[33] = in[87] ^ in2[87];
    assign G[34] = in[86] & in2[86];
    assign P[34] = in[86] ^ in2[86];
    assign G[35] = in[85] & in2[85];
    assign P[35] = in[85] ^ in2[85];
    assign G[36] = in[84] & in2[84];
    assign P[36] = in[84] ^ in2[84];
    assign G[37] = in[83] & in2[83];
    assign P[37] = in[83] ^ in2[83];
    assign G[38] = in[82] & in2[82];
    assign P[38] = in[82] ^ in2[82];
    assign G[39] = in[81] & in2[81];
    assign P[39] = in[81] ^ in2[81];
    assign G[40] = in[80] & in2[80];
    assign P[40] = in[80] ^ in2[80];
    assign G[41] = in[79] & in2[79];
    assign P[41] = in[79] ^ in2[79];
    assign G[42] = in[78] & in2[78];
    assign P[42] = in[78] ^ in2[78];
    assign G[43] = in[77] & in2[77];
    assign P[43] = in[77] ^ in2[77];
    assign G[44] = in[76] & in2[76];
    assign P[44] = in[76] ^ in2[76];
    assign G[45] = in[75] & in2[75];
    assign P[45] = in[75] ^ in2[75];
    assign G[46] = in[74] & in2[74];
    assign P[46] = in[74] ^ in2[74];
    assign G[47] = in[73] & in2[73];
    assign P[47] = in[73] ^ in2[73];
    assign G[48] = in[72] & in2[72];
    assign P[48] = in[72] ^ in2[72];
    assign G[49] = in[71] & in2[71];
    assign P[49] = in[71] ^ in2[71];
    assign G[50] = in[70] & in2[70];
    assign P[50] = in[70] ^ in2[70];
    assign G[51] = in[69] & in2[69];
    assign P[51] = in[69] ^ in2[69];
    assign G[52] = in[68] & in2[68];
    assign P[52] = in[68] ^ in2[68];
    assign G[53] = in[67] & in2[67];
    assign P[53] = in[67] ^ in2[67];
    assign G[54] = in[66] & in2[66];
    assign P[54] = in[66] ^ in2[66];
    assign G[55] = in[65] & in2[65];
    assign P[55] = in[65] ^ in2[65];
    assign G[56] = in[64] & in2[64];
    assign P[56] = in[64] ^ in2[64];
    assign G[57] = in[63] & in2[63];
    assign P[57] = in[63] ^ in2[63];
    assign G[58] = in[62] & in2[62];
    assign P[58] = in[62] ^ in2[62];
    assign G[59] = in[61] & in2[61];
    assign P[59] = in[61] ^ in2[61];
    assign G[60] = in[60] & in2[60];
    assign P[60] = in[60] ^ in2[60];
    assign G[61] = in[59] & in2[59];
    assign P[61] = in[59] ^ in2[59];
    assign G[62] = in[58] & in2[58];
    assign P[62] = in[58] ^ in2[58];
    assign G[63] = in[57] & in2[57];
    assign P[63] = in[57] ^ in2[57];
    assign G[64] = in[56] & in2[56];
    assign P[64] = in[56] ^ in2[56];
    assign G[65] = in[55] & in2[55];
    assign P[65] = in[55] ^ in2[55];
    assign G[66] = in[54] & in2[54];
    assign P[66] = in[54] ^ in2[54];
    assign G[67] = in[53] & in2[53];
    assign P[67] = in[53] ^ in2[53];
    assign G[68] = in[52] & in2[52];
    assign P[68] = in[52] ^ in2[52];
    assign G[69] = in[51] & in2[51];
    assign P[69] = in[51] ^ in2[51];
    assign G[70] = in[50] & in2[50];
    assign P[70] = in[50] ^ in2[50];
    assign G[71] = in[49] & in2[49];
    assign P[71] = in[49] ^ in2[49];
    assign G[72] = in[48] & in2[48];
    assign P[72] = in[48] ^ in2[48];
    assign G[73] = in[47] & in2[47];
    assign P[73] = in[47] ^ in2[47];
    assign G[74] = in[46] & in2[46];
    assign P[74] = in[46] ^ in2[46];
    assign G[75] = in[45] & in2[45];
    assign P[75] = in[45] ^ in2[45];
    assign G[76] = in[44] & in2[44];
    assign P[76] = in[44] ^ in2[44];
    assign G[77] = in[43] & in2[43];
    assign P[77] = in[43] ^ in2[43];
    assign G[78] = in[42] & in2[42];
    assign P[78] = in[42] ^ in2[42];
    assign G[79] = in[41] & in2[41];
    assign P[79] = in[41] ^ in2[41];
    assign G[80] = in[40] & in2[40];
    assign P[80] = in[40] ^ in2[40];
    assign G[81] = in[39] & in2[39];
    assign P[81] = in[39] ^ in2[39];
    assign G[82] = in[38] & in2[38];
    assign P[82] = in[38] ^ in2[38];
    assign G[83] = in[37] & in2[37];
    assign P[83] = in[37] ^ in2[37];
    assign G[84] = in[36] & in2[36];
    assign P[84] = in[36] ^ in2[36];
    assign G[85] = in[35] & in2[35];
    assign P[85] = in[35] ^ in2[35];
    assign G[86] = in[34] & in2[34];
    assign P[86] = in[34] ^ in2[34];
    assign G[87] = in[33] & in2[33];
    assign P[87] = in[33] ^ in2[33];
    assign G[88] = in[32] & in2[32];
    assign P[88] = in[32] ^ in2[32];
    assign G[89] = in[31] & in2[31];
    assign P[89] = in[31] ^ in2[31];
    assign G[90] = in[30] & in2[30];
    assign P[90] = in[30] ^ in2[30];
    assign G[91] = in[29] & in2[29];
    assign P[91] = in[29] ^ in2[29];
    assign G[92] = in[28] & in2[28];
    assign P[92] = in[28] ^ in2[28];
    assign G[93] = in[27] & in2[27];
    assign P[93] = in[27] ^ in2[27];
    assign G[94] = in[26] & in2[26];
    assign P[94] = in[26] ^ in2[26];
    assign G[95] = in[25] & in2[25];
    assign P[95] = in[25] ^ in2[25];
    assign G[96] = in[24] & in2[24];
    assign P[96] = in[24] ^ in2[24];
    assign G[97] = in[23] & in2[23];
    assign P[97] = in[23] ^ in2[23];
    assign G[98] = in[22] & in2[22];
    assign P[98] = in[22] ^ in2[22];
    assign G[99] = in[21] & in2[21];
    assign P[99] = in[21] ^ in2[21];
    assign G[100] = in[20] & in2[20];
    assign P[100] = in[20] ^ in2[20];
    assign G[101] = in[19] & in2[19];
    assign P[101] = in[19] ^ in2[19];
    assign G[102] = in[18] & in2[18];
    assign P[102] = in[18] ^ in2[18];
    assign G[103] = in[17] & in2[17];
    assign P[103] = in[17] ^ in2[17];
    assign G[104] = in[16] & in2[16];
    assign P[104] = in[16] ^ in2[16];
    assign G[105] = in[15] & in2[15];
    assign P[105] = in[15] ^ in2[15];
    assign G[106] = in[14] & in2[14];
    assign P[106] = in[14] ^ in2[14];
    assign G[107] = in[13] & in2[13];
    assign P[107] = in[13] ^ in2[13];
    assign G[108] = in[12] & in2[12];
    assign P[108] = in[12] ^ in2[12];
    assign G[109] = in[11] & in2[11];
    assign P[109] = in[11] ^ in2[11];
    assign G[110] = in[10] & in2[10];
    assign P[110] = in[10] ^ in2[10];
    assign G[111] = in[9] & in2[9];
    assign P[111] = in[9] ^ in2[9];
    assign G[112] = in[8] & in2[8];
    assign P[112] = in[8] ^ in2[8];
    assign G[113] = in[7] & in2[7];
    assign P[113] = in[7] ^ in2[7];
    assign G[114] = in[6] & in2[6];
    assign P[114] = in[6] ^ in2[6];
    assign G[115] = in[5] & in2[5];
    assign P[115] = in[5] ^ in2[5];
    assign G[116] = in[4] & in2[4];
    assign P[116] = in[4] ^ in2[4];
    assign G[117] = in[3] & in2[3];
    assign P[117] = in[3] ^ in2[3];
    assign G[118] = in[2] & in2[2];
    assign P[118] = in[2] ^ in2[2];
    assign G[119] = in[1] & in2[1];
    assign P[119] = in[1] ^ in2[1];
    assign G[120] = in[0] & in2[0];
    assign P[120] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign C[120] = G[119] | (P[119] & C[119]);
    assign cout = G[120] | (P[120] & C[120]);
    assign sum = P ^ C;
endmodule

module CLA120(output [119:0] sum, output cout, input [119:0] in1, input [119:0] in2;

    wire[119:0] G;
    wire[119:0] C;
    wire[119:0] P;

    assign G[0] = in[119] & in2[119];
    assign P[0] = in[119] ^ in2[119];
    assign G[1] = in[118] & in2[118];
    assign P[1] = in[118] ^ in2[118];
    assign G[2] = in[117] & in2[117];
    assign P[2] = in[117] ^ in2[117];
    assign G[3] = in[116] & in2[116];
    assign P[3] = in[116] ^ in2[116];
    assign G[4] = in[115] & in2[115];
    assign P[4] = in[115] ^ in2[115];
    assign G[5] = in[114] & in2[114];
    assign P[5] = in[114] ^ in2[114];
    assign G[6] = in[113] & in2[113];
    assign P[6] = in[113] ^ in2[113];
    assign G[7] = in[112] & in2[112];
    assign P[7] = in[112] ^ in2[112];
    assign G[8] = in[111] & in2[111];
    assign P[8] = in[111] ^ in2[111];
    assign G[9] = in[110] & in2[110];
    assign P[9] = in[110] ^ in2[110];
    assign G[10] = in[109] & in2[109];
    assign P[10] = in[109] ^ in2[109];
    assign G[11] = in[108] & in2[108];
    assign P[11] = in[108] ^ in2[108];
    assign G[12] = in[107] & in2[107];
    assign P[12] = in[107] ^ in2[107];
    assign G[13] = in[106] & in2[106];
    assign P[13] = in[106] ^ in2[106];
    assign G[14] = in[105] & in2[105];
    assign P[14] = in[105] ^ in2[105];
    assign G[15] = in[104] & in2[104];
    assign P[15] = in[104] ^ in2[104];
    assign G[16] = in[103] & in2[103];
    assign P[16] = in[103] ^ in2[103];
    assign G[17] = in[102] & in2[102];
    assign P[17] = in[102] ^ in2[102];
    assign G[18] = in[101] & in2[101];
    assign P[18] = in[101] ^ in2[101];
    assign G[19] = in[100] & in2[100];
    assign P[19] = in[100] ^ in2[100];
    assign G[20] = in[99] & in2[99];
    assign P[20] = in[99] ^ in2[99];
    assign G[21] = in[98] & in2[98];
    assign P[21] = in[98] ^ in2[98];
    assign G[22] = in[97] & in2[97];
    assign P[22] = in[97] ^ in2[97];
    assign G[23] = in[96] & in2[96];
    assign P[23] = in[96] ^ in2[96];
    assign G[24] = in[95] & in2[95];
    assign P[24] = in[95] ^ in2[95];
    assign G[25] = in[94] & in2[94];
    assign P[25] = in[94] ^ in2[94];
    assign G[26] = in[93] & in2[93];
    assign P[26] = in[93] ^ in2[93];
    assign G[27] = in[92] & in2[92];
    assign P[27] = in[92] ^ in2[92];
    assign G[28] = in[91] & in2[91];
    assign P[28] = in[91] ^ in2[91];
    assign G[29] = in[90] & in2[90];
    assign P[29] = in[90] ^ in2[90];
    assign G[30] = in[89] & in2[89];
    assign P[30] = in[89] ^ in2[89];
    assign G[31] = in[88] & in2[88];
    assign P[31] = in[88] ^ in2[88];
    assign G[32] = in[87] & in2[87];
    assign P[32] = in[87] ^ in2[87];
    assign G[33] = in[86] & in2[86];
    assign P[33] = in[86] ^ in2[86];
    assign G[34] = in[85] & in2[85];
    assign P[34] = in[85] ^ in2[85];
    assign G[35] = in[84] & in2[84];
    assign P[35] = in[84] ^ in2[84];
    assign G[36] = in[83] & in2[83];
    assign P[36] = in[83] ^ in2[83];
    assign G[37] = in[82] & in2[82];
    assign P[37] = in[82] ^ in2[82];
    assign G[38] = in[81] & in2[81];
    assign P[38] = in[81] ^ in2[81];
    assign G[39] = in[80] & in2[80];
    assign P[39] = in[80] ^ in2[80];
    assign G[40] = in[79] & in2[79];
    assign P[40] = in[79] ^ in2[79];
    assign G[41] = in[78] & in2[78];
    assign P[41] = in[78] ^ in2[78];
    assign G[42] = in[77] & in2[77];
    assign P[42] = in[77] ^ in2[77];
    assign G[43] = in[76] & in2[76];
    assign P[43] = in[76] ^ in2[76];
    assign G[44] = in[75] & in2[75];
    assign P[44] = in[75] ^ in2[75];
    assign G[45] = in[74] & in2[74];
    assign P[45] = in[74] ^ in2[74];
    assign G[46] = in[73] & in2[73];
    assign P[46] = in[73] ^ in2[73];
    assign G[47] = in[72] & in2[72];
    assign P[47] = in[72] ^ in2[72];
    assign G[48] = in[71] & in2[71];
    assign P[48] = in[71] ^ in2[71];
    assign G[49] = in[70] & in2[70];
    assign P[49] = in[70] ^ in2[70];
    assign G[50] = in[69] & in2[69];
    assign P[50] = in[69] ^ in2[69];
    assign G[51] = in[68] & in2[68];
    assign P[51] = in[68] ^ in2[68];
    assign G[52] = in[67] & in2[67];
    assign P[52] = in[67] ^ in2[67];
    assign G[53] = in[66] & in2[66];
    assign P[53] = in[66] ^ in2[66];
    assign G[54] = in[65] & in2[65];
    assign P[54] = in[65] ^ in2[65];
    assign G[55] = in[64] & in2[64];
    assign P[55] = in[64] ^ in2[64];
    assign G[56] = in[63] & in2[63];
    assign P[56] = in[63] ^ in2[63];
    assign G[57] = in[62] & in2[62];
    assign P[57] = in[62] ^ in2[62];
    assign G[58] = in[61] & in2[61];
    assign P[58] = in[61] ^ in2[61];
    assign G[59] = in[60] & in2[60];
    assign P[59] = in[60] ^ in2[60];
    assign G[60] = in[59] & in2[59];
    assign P[60] = in[59] ^ in2[59];
    assign G[61] = in[58] & in2[58];
    assign P[61] = in[58] ^ in2[58];
    assign G[62] = in[57] & in2[57];
    assign P[62] = in[57] ^ in2[57];
    assign G[63] = in[56] & in2[56];
    assign P[63] = in[56] ^ in2[56];
    assign G[64] = in[55] & in2[55];
    assign P[64] = in[55] ^ in2[55];
    assign G[65] = in[54] & in2[54];
    assign P[65] = in[54] ^ in2[54];
    assign G[66] = in[53] & in2[53];
    assign P[66] = in[53] ^ in2[53];
    assign G[67] = in[52] & in2[52];
    assign P[67] = in[52] ^ in2[52];
    assign G[68] = in[51] & in2[51];
    assign P[68] = in[51] ^ in2[51];
    assign G[69] = in[50] & in2[50];
    assign P[69] = in[50] ^ in2[50];
    assign G[70] = in[49] & in2[49];
    assign P[70] = in[49] ^ in2[49];
    assign G[71] = in[48] & in2[48];
    assign P[71] = in[48] ^ in2[48];
    assign G[72] = in[47] & in2[47];
    assign P[72] = in[47] ^ in2[47];
    assign G[73] = in[46] & in2[46];
    assign P[73] = in[46] ^ in2[46];
    assign G[74] = in[45] & in2[45];
    assign P[74] = in[45] ^ in2[45];
    assign G[75] = in[44] & in2[44];
    assign P[75] = in[44] ^ in2[44];
    assign G[76] = in[43] & in2[43];
    assign P[76] = in[43] ^ in2[43];
    assign G[77] = in[42] & in2[42];
    assign P[77] = in[42] ^ in2[42];
    assign G[78] = in[41] & in2[41];
    assign P[78] = in[41] ^ in2[41];
    assign G[79] = in[40] & in2[40];
    assign P[79] = in[40] ^ in2[40];
    assign G[80] = in[39] & in2[39];
    assign P[80] = in[39] ^ in2[39];
    assign G[81] = in[38] & in2[38];
    assign P[81] = in[38] ^ in2[38];
    assign G[82] = in[37] & in2[37];
    assign P[82] = in[37] ^ in2[37];
    assign G[83] = in[36] & in2[36];
    assign P[83] = in[36] ^ in2[36];
    assign G[84] = in[35] & in2[35];
    assign P[84] = in[35] ^ in2[35];
    assign G[85] = in[34] & in2[34];
    assign P[85] = in[34] ^ in2[34];
    assign G[86] = in[33] & in2[33];
    assign P[86] = in[33] ^ in2[33];
    assign G[87] = in[32] & in2[32];
    assign P[87] = in[32] ^ in2[32];
    assign G[88] = in[31] & in2[31];
    assign P[88] = in[31] ^ in2[31];
    assign G[89] = in[30] & in2[30];
    assign P[89] = in[30] ^ in2[30];
    assign G[90] = in[29] & in2[29];
    assign P[90] = in[29] ^ in2[29];
    assign G[91] = in[28] & in2[28];
    assign P[91] = in[28] ^ in2[28];
    assign G[92] = in[27] & in2[27];
    assign P[92] = in[27] ^ in2[27];
    assign G[93] = in[26] & in2[26];
    assign P[93] = in[26] ^ in2[26];
    assign G[94] = in[25] & in2[25];
    assign P[94] = in[25] ^ in2[25];
    assign G[95] = in[24] & in2[24];
    assign P[95] = in[24] ^ in2[24];
    assign G[96] = in[23] & in2[23];
    assign P[96] = in[23] ^ in2[23];
    assign G[97] = in[22] & in2[22];
    assign P[97] = in[22] ^ in2[22];
    assign G[98] = in[21] & in2[21];
    assign P[98] = in[21] ^ in2[21];
    assign G[99] = in[20] & in2[20];
    assign P[99] = in[20] ^ in2[20];
    assign G[100] = in[19] & in2[19];
    assign P[100] = in[19] ^ in2[19];
    assign G[101] = in[18] & in2[18];
    assign P[101] = in[18] ^ in2[18];
    assign G[102] = in[17] & in2[17];
    assign P[102] = in[17] ^ in2[17];
    assign G[103] = in[16] & in2[16];
    assign P[103] = in[16] ^ in2[16];
    assign G[104] = in[15] & in2[15];
    assign P[104] = in[15] ^ in2[15];
    assign G[105] = in[14] & in2[14];
    assign P[105] = in[14] ^ in2[14];
    assign G[106] = in[13] & in2[13];
    assign P[106] = in[13] ^ in2[13];
    assign G[107] = in[12] & in2[12];
    assign P[107] = in[12] ^ in2[12];
    assign G[108] = in[11] & in2[11];
    assign P[108] = in[11] ^ in2[11];
    assign G[109] = in[10] & in2[10];
    assign P[109] = in[10] ^ in2[10];
    assign G[110] = in[9] & in2[9];
    assign P[110] = in[9] ^ in2[9];
    assign G[111] = in[8] & in2[8];
    assign P[111] = in[8] ^ in2[8];
    assign G[112] = in[7] & in2[7];
    assign P[112] = in[7] ^ in2[7];
    assign G[113] = in[6] & in2[6];
    assign P[113] = in[6] ^ in2[6];
    assign G[114] = in[5] & in2[5];
    assign P[114] = in[5] ^ in2[5];
    assign G[115] = in[4] & in2[4];
    assign P[115] = in[4] ^ in2[4];
    assign G[116] = in[3] & in2[3];
    assign P[116] = in[3] ^ in2[3];
    assign G[117] = in[2] & in2[2];
    assign P[117] = in[2] ^ in2[2];
    assign G[118] = in[1] & in2[1];
    assign P[118] = in[1] ^ in2[1];
    assign G[119] = in[0] & in2[0];
    assign P[119] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign C[119] = G[118] | (P[118] & C[118]);
    assign cout = G[119] | (P[119] & C[119]);
    assign sum = P ^ C;
endmodule

module CLA119(output [118:0] sum, output cout, input [118:0] in1, input [118:0] in2;

    wire[118:0] G;
    wire[118:0] C;
    wire[118:0] P;

    assign G[0] = in[118] & in2[118];
    assign P[0] = in[118] ^ in2[118];
    assign G[1] = in[117] & in2[117];
    assign P[1] = in[117] ^ in2[117];
    assign G[2] = in[116] & in2[116];
    assign P[2] = in[116] ^ in2[116];
    assign G[3] = in[115] & in2[115];
    assign P[3] = in[115] ^ in2[115];
    assign G[4] = in[114] & in2[114];
    assign P[4] = in[114] ^ in2[114];
    assign G[5] = in[113] & in2[113];
    assign P[5] = in[113] ^ in2[113];
    assign G[6] = in[112] & in2[112];
    assign P[6] = in[112] ^ in2[112];
    assign G[7] = in[111] & in2[111];
    assign P[7] = in[111] ^ in2[111];
    assign G[8] = in[110] & in2[110];
    assign P[8] = in[110] ^ in2[110];
    assign G[9] = in[109] & in2[109];
    assign P[9] = in[109] ^ in2[109];
    assign G[10] = in[108] & in2[108];
    assign P[10] = in[108] ^ in2[108];
    assign G[11] = in[107] & in2[107];
    assign P[11] = in[107] ^ in2[107];
    assign G[12] = in[106] & in2[106];
    assign P[12] = in[106] ^ in2[106];
    assign G[13] = in[105] & in2[105];
    assign P[13] = in[105] ^ in2[105];
    assign G[14] = in[104] & in2[104];
    assign P[14] = in[104] ^ in2[104];
    assign G[15] = in[103] & in2[103];
    assign P[15] = in[103] ^ in2[103];
    assign G[16] = in[102] & in2[102];
    assign P[16] = in[102] ^ in2[102];
    assign G[17] = in[101] & in2[101];
    assign P[17] = in[101] ^ in2[101];
    assign G[18] = in[100] & in2[100];
    assign P[18] = in[100] ^ in2[100];
    assign G[19] = in[99] & in2[99];
    assign P[19] = in[99] ^ in2[99];
    assign G[20] = in[98] & in2[98];
    assign P[20] = in[98] ^ in2[98];
    assign G[21] = in[97] & in2[97];
    assign P[21] = in[97] ^ in2[97];
    assign G[22] = in[96] & in2[96];
    assign P[22] = in[96] ^ in2[96];
    assign G[23] = in[95] & in2[95];
    assign P[23] = in[95] ^ in2[95];
    assign G[24] = in[94] & in2[94];
    assign P[24] = in[94] ^ in2[94];
    assign G[25] = in[93] & in2[93];
    assign P[25] = in[93] ^ in2[93];
    assign G[26] = in[92] & in2[92];
    assign P[26] = in[92] ^ in2[92];
    assign G[27] = in[91] & in2[91];
    assign P[27] = in[91] ^ in2[91];
    assign G[28] = in[90] & in2[90];
    assign P[28] = in[90] ^ in2[90];
    assign G[29] = in[89] & in2[89];
    assign P[29] = in[89] ^ in2[89];
    assign G[30] = in[88] & in2[88];
    assign P[30] = in[88] ^ in2[88];
    assign G[31] = in[87] & in2[87];
    assign P[31] = in[87] ^ in2[87];
    assign G[32] = in[86] & in2[86];
    assign P[32] = in[86] ^ in2[86];
    assign G[33] = in[85] & in2[85];
    assign P[33] = in[85] ^ in2[85];
    assign G[34] = in[84] & in2[84];
    assign P[34] = in[84] ^ in2[84];
    assign G[35] = in[83] & in2[83];
    assign P[35] = in[83] ^ in2[83];
    assign G[36] = in[82] & in2[82];
    assign P[36] = in[82] ^ in2[82];
    assign G[37] = in[81] & in2[81];
    assign P[37] = in[81] ^ in2[81];
    assign G[38] = in[80] & in2[80];
    assign P[38] = in[80] ^ in2[80];
    assign G[39] = in[79] & in2[79];
    assign P[39] = in[79] ^ in2[79];
    assign G[40] = in[78] & in2[78];
    assign P[40] = in[78] ^ in2[78];
    assign G[41] = in[77] & in2[77];
    assign P[41] = in[77] ^ in2[77];
    assign G[42] = in[76] & in2[76];
    assign P[42] = in[76] ^ in2[76];
    assign G[43] = in[75] & in2[75];
    assign P[43] = in[75] ^ in2[75];
    assign G[44] = in[74] & in2[74];
    assign P[44] = in[74] ^ in2[74];
    assign G[45] = in[73] & in2[73];
    assign P[45] = in[73] ^ in2[73];
    assign G[46] = in[72] & in2[72];
    assign P[46] = in[72] ^ in2[72];
    assign G[47] = in[71] & in2[71];
    assign P[47] = in[71] ^ in2[71];
    assign G[48] = in[70] & in2[70];
    assign P[48] = in[70] ^ in2[70];
    assign G[49] = in[69] & in2[69];
    assign P[49] = in[69] ^ in2[69];
    assign G[50] = in[68] & in2[68];
    assign P[50] = in[68] ^ in2[68];
    assign G[51] = in[67] & in2[67];
    assign P[51] = in[67] ^ in2[67];
    assign G[52] = in[66] & in2[66];
    assign P[52] = in[66] ^ in2[66];
    assign G[53] = in[65] & in2[65];
    assign P[53] = in[65] ^ in2[65];
    assign G[54] = in[64] & in2[64];
    assign P[54] = in[64] ^ in2[64];
    assign G[55] = in[63] & in2[63];
    assign P[55] = in[63] ^ in2[63];
    assign G[56] = in[62] & in2[62];
    assign P[56] = in[62] ^ in2[62];
    assign G[57] = in[61] & in2[61];
    assign P[57] = in[61] ^ in2[61];
    assign G[58] = in[60] & in2[60];
    assign P[58] = in[60] ^ in2[60];
    assign G[59] = in[59] & in2[59];
    assign P[59] = in[59] ^ in2[59];
    assign G[60] = in[58] & in2[58];
    assign P[60] = in[58] ^ in2[58];
    assign G[61] = in[57] & in2[57];
    assign P[61] = in[57] ^ in2[57];
    assign G[62] = in[56] & in2[56];
    assign P[62] = in[56] ^ in2[56];
    assign G[63] = in[55] & in2[55];
    assign P[63] = in[55] ^ in2[55];
    assign G[64] = in[54] & in2[54];
    assign P[64] = in[54] ^ in2[54];
    assign G[65] = in[53] & in2[53];
    assign P[65] = in[53] ^ in2[53];
    assign G[66] = in[52] & in2[52];
    assign P[66] = in[52] ^ in2[52];
    assign G[67] = in[51] & in2[51];
    assign P[67] = in[51] ^ in2[51];
    assign G[68] = in[50] & in2[50];
    assign P[68] = in[50] ^ in2[50];
    assign G[69] = in[49] & in2[49];
    assign P[69] = in[49] ^ in2[49];
    assign G[70] = in[48] & in2[48];
    assign P[70] = in[48] ^ in2[48];
    assign G[71] = in[47] & in2[47];
    assign P[71] = in[47] ^ in2[47];
    assign G[72] = in[46] & in2[46];
    assign P[72] = in[46] ^ in2[46];
    assign G[73] = in[45] & in2[45];
    assign P[73] = in[45] ^ in2[45];
    assign G[74] = in[44] & in2[44];
    assign P[74] = in[44] ^ in2[44];
    assign G[75] = in[43] & in2[43];
    assign P[75] = in[43] ^ in2[43];
    assign G[76] = in[42] & in2[42];
    assign P[76] = in[42] ^ in2[42];
    assign G[77] = in[41] & in2[41];
    assign P[77] = in[41] ^ in2[41];
    assign G[78] = in[40] & in2[40];
    assign P[78] = in[40] ^ in2[40];
    assign G[79] = in[39] & in2[39];
    assign P[79] = in[39] ^ in2[39];
    assign G[80] = in[38] & in2[38];
    assign P[80] = in[38] ^ in2[38];
    assign G[81] = in[37] & in2[37];
    assign P[81] = in[37] ^ in2[37];
    assign G[82] = in[36] & in2[36];
    assign P[82] = in[36] ^ in2[36];
    assign G[83] = in[35] & in2[35];
    assign P[83] = in[35] ^ in2[35];
    assign G[84] = in[34] & in2[34];
    assign P[84] = in[34] ^ in2[34];
    assign G[85] = in[33] & in2[33];
    assign P[85] = in[33] ^ in2[33];
    assign G[86] = in[32] & in2[32];
    assign P[86] = in[32] ^ in2[32];
    assign G[87] = in[31] & in2[31];
    assign P[87] = in[31] ^ in2[31];
    assign G[88] = in[30] & in2[30];
    assign P[88] = in[30] ^ in2[30];
    assign G[89] = in[29] & in2[29];
    assign P[89] = in[29] ^ in2[29];
    assign G[90] = in[28] & in2[28];
    assign P[90] = in[28] ^ in2[28];
    assign G[91] = in[27] & in2[27];
    assign P[91] = in[27] ^ in2[27];
    assign G[92] = in[26] & in2[26];
    assign P[92] = in[26] ^ in2[26];
    assign G[93] = in[25] & in2[25];
    assign P[93] = in[25] ^ in2[25];
    assign G[94] = in[24] & in2[24];
    assign P[94] = in[24] ^ in2[24];
    assign G[95] = in[23] & in2[23];
    assign P[95] = in[23] ^ in2[23];
    assign G[96] = in[22] & in2[22];
    assign P[96] = in[22] ^ in2[22];
    assign G[97] = in[21] & in2[21];
    assign P[97] = in[21] ^ in2[21];
    assign G[98] = in[20] & in2[20];
    assign P[98] = in[20] ^ in2[20];
    assign G[99] = in[19] & in2[19];
    assign P[99] = in[19] ^ in2[19];
    assign G[100] = in[18] & in2[18];
    assign P[100] = in[18] ^ in2[18];
    assign G[101] = in[17] & in2[17];
    assign P[101] = in[17] ^ in2[17];
    assign G[102] = in[16] & in2[16];
    assign P[102] = in[16] ^ in2[16];
    assign G[103] = in[15] & in2[15];
    assign P[103] = in[15] ^ in2[15];
    assign G[104] = in[14] & in2[14];
    assign P[104] = in[14] ^ in2[14];
    assign G[105] = in[13] & in2[13];
    assign P[105] = in[13] ^ in2[13];
    assign G[106] = in[12] & in2[12];
    assign P[106] = in[12] ^ in2[12];
    assign G[107] = in[11] & in2[11];
    assign P[107] = in[11] ^ in2[11];
    assign G[108] = in[10] & in2[10];
    assign P[108] = in[10] ^ in2[10];
    assign G[109] = in[9] & in2[9];
    assign P[109] = in[9] ^ in2[9];
    assign G[110] = in[8] & in2[8];
    assign P[110] = in[8] ^ in2[8];
    assign G[111] = in[7] & in2[7];
    assign P[111] = in[7] ^ in2[7];
    assign G[112] = in[6] & in2[6];
    assign P[112] = in[6] ^ in2[6];
    assign G[113] = in[5] & in2[5];
    assign P[113] = in[5] ^ in2[5];
    assign G[114] = in[4] & in2[4];
    assign P[114] = in[4] ^ in2[4];
    assign G[115] = in[3] & in2[3];
    assign P[115] = in[3] ^ in2[3];
    assign G[116] = in[2] & in2[2];
    assign P[116] = in[2] ^ in2[2];
    assign G[117] = in[1] & in2[1];
    assign P[117] = in[1] ^ in2[1];
    assign G[118] = in[0] & in2[0];
    assign P[118] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign C[118] = G[117] | (P[117] & C[117]);
    assign cout = G[118] | (P[118] & C[118]);
    assign sum = P ^ C;
endmodule

module CLA118(output [117:0] sum, output cout, input [117:0] in1, input [117:0] in2;

    wire[117:0] G;
    wire[117:0] C;
    wire[117:0] P;

    assign G[0] = in[117] & in2[117];
    assign P[0] = in[117] ^ in2[117];
    assign G[1] = in[116] & in2[116];
    assign P[1] = in[116] ^ in2[116];
    assign G[2] = in[115] & in2[115];
    assign P[2] = in[115] ^ in2[115];
    assign G[3] = in[114] & in2[114];
    assign P[3] = in[114] ^ in2[114];
    assign G[4] = in[113] & in2[113];
    assign P[4] = in[113] ^ in2[113];
    assign G[5] = in[112] & in2[112];
    assign P[5] = in[112] ^ in2[112];
    assign G[6] = in[111] & in2[111];
    assign P[6] = in[111] ^ in2[111];
    assign G[7] = in[110] & in2[110];
    assign P[7] = in[110] ^ in2[110];
    assign G[8] = in[109] & in2[109];
    assign P[8] = in[109] ^ in2[109];
    assign G[9] = in[108] & in2[108];
    assign P[9] = in[108] ^ in2[108];
    assign G[10] = in[107] & in2[107];
    assign P[10] = in[107] ^ in2[107];
    assign G[11] = in[106] & in2[106];
    assign P[11] = in[106] ^ in2[106];
    assign G[12] = in[105] & in2[105];
    assign P[12] = in[105] ^ in2[105];
    assign G[13] = in[104] & in2[104];
    assign P[13] = in[104] ^ in2[104];
    assign G[14] = in[103] & in2[103];
    assign P[14] = in[103] ^ in2[103];
    assign G[15] = in[102] & in2[102];
    assign P[15] = in[102] ^ in2[102];
    assign G[16] = in[101] & in2[101];
    assign P[16] = in[101] ^ in2[101];
    assign G[17] = in[100] & in2[100];
    assign P[17] = in[100] ^ in2[100];
    assign G[18] = in[99] & in2[99];
    assign P[18] = in[99] ^ in2[99];
    assign G[19] = in[98] & in2[98];
    assign P[19] = in[98] ^ in2[98];
    assign G[20] = in[97] & in2[97];
    assign P[20] = in[97] ^ in2[97];
    assign G[21] = in[96] & in2[96];
    assign P[21] = in[96] ^ in2[96];
    assign G[22] = in[95] & in2[95];
    assign P[22] = in[95] ^ in2[95];
    assign G[23] = in[94] & in2[94];
    assign P[23] = in[94] ^ in2[94];
    assign G[24] = in[93] & in2[93];
    assign P[24] = in[93] ^ in2[93];
    assign G[25] = in[92] & in2[92];
    assign P[25] = in[92] ^ in2[92];
    assign G[26] = in[91] & in2[91];
    assign P[26] = in[91] ^ in2[91];
    assign G[27] = in[90] & in2[90];
    assign P[27] = in[90] ^ in2[90];
    assign G[28] = in[89] & in2[89];
    assign P[28] = in[89] ^ in2[89];
    assign G[29] = in[88] & in2[88];
    assign P[29] = in[88] ^ in2[88];
    assign G[30] = in[87] & in2[87];
    assign P[30] = in[87] ^ in2[87];
    assign G[31] = in[86] & in2[86];
    assign P[31] = in[86] ^ in2[86];
    assign G[32] = in[85] & in2[85];
    assign P[32] = in[85] ^ in2[85];
    assign G[33] = in[84] & in2[84];
    assign P[33] = in[84] ^ in2[84];
    assign G[34] = in[83] & in2[83];
    assign P[34] = in[83] ^ in2[83];
    assign G[35] = in[82] & in2[82];
    assign P[35] = in[82] ^ in2[82];
    assign G[36] = in[81] & in2[81];
    assign P[36] = in[81] ^ in2[81];
    assign G[37] = in[80] & in2[80];
    assign P[37] = in[80] ^ in2[80];
    assign G[38] = in[79] & in2[79];
    assign P[38] = in[79] ^ in2[79];
    assign G[39] = in[78] & in2[78];
    assign P[39] = in[78] ^ in2[78];
    assign G[40] = in[77] & in2[77];
    assign P[40] = in[77] ^ in2[77];
    assign G[41] = in[76] & in2[76];
    assign P[41] = in[76] ^ in2[76];
    assign G[42] = in[75] & in2[75];
    assign P[42] = in[75] ^ in2[75];
    assign G[43] = in[74] & in2[74];
    assign P[43] = in[74] ^ in2[74];
    assign G[44] = in[73] & in2[73];
    assign P[44] = in[73] ^ in2[73];
    assign G[45] = in[72] & in2[72];
    assign P[45] = in[72] ^ in2[72];
    assign G[46] = in[71] & in2[71];
    assign P[46] = in[71] ^ in2[71];
    assign G[47] = in[70] & in2[70];
    assign P[47] = in[70] ^ in2[70];
    assign G[48] = in[69] & in2[69];
    assign P[48] = in[69] ^ in2[69];
    assign G[49] = in[68] & in2[68];
    assign P[49] = in[68] ^ in2[68];
    assign G[50] = in[67] & in2[67];
    assign P[50] = in[67] ^ in2[67];
    assign G[51] = in[66] & in2[66];
    assign P[51] = in[66] ^ in2[66];
    assign G[52] = in[65] & in2[65];
    assign P[52] = in[65] ^ in2[65];
    assign G[53] = in[64] & in2[64];
    assign P[53] = in[64] ^ in2[64];
    assign G[54] = in[63] & in2[63];
    assign P[54] = in[63] ^ in2[63];
    assign G[55] = in[62] & in2[62];
    assign P[55] = in[62] ^ in2[62];
    assign G[56] = in[61] & in2[61];
    assign P[56] = in[61] ^ in2[61];
    assign G[57] = in[60] & in2[60];
    assign P[57] = in[60] ^ in2[60];
    assign G[58] = in[59] & in2[59];
    assign P[58] = in[59] ^ in2[59];
    assign G[59] = in[58] & in2[58];
    assign P[59] = in[58] ^ in2[58];
    assign G[60] = in[57] & in2[57];
    assign P[60] = in[57] ^ in2[57];
    assign G[61] = in[56] & in2[56];
    assign P[61] = in[56] ^ in2[56];
    assign G[62] = in[55] & in2[55];
    assign P[62] = in[55] ^ in2[55];
    assign G[63] = in[54] & in2[54];
    assign P[63] = in[54] ^ in2[54];
    assign G[64] = in[53] & in2[53];
    assign P[64] = in[53] ^ in2[53];
    assign G[65] = in[52] & in2[52];
    assign P[65] = in[52] ^ in2[52];
    assign G[66] = in[51] & in2[51];
    assign P[66] = in[51] ^ in2[51];
    assign G[67] = in[50] & in2[50];
    assign P[67] = in[50] ^ in2[50];
    assign G[68] = in[49] & in2[49];
    assign P[68] = in[49] ^ in2[49];
    assign G[69] = in[48] & in2[48];
    assign P[69] = in[48] ^ in2[48];
    assign G[70] = in[47] & in2[47];
    assign P[70] = in[47] ^ in2[47];
    assign G[71] = in[46] & in2[46];
    assign P[71] = in[46] ^ in2[46];
    assign G[72] = in[45] & in2[45];
    assign P[72] = in[45] ^ in2[45];
    assign G[73] = in[44] & in2[44];
    assign P[73] = in[44] ^ in2[44];
    assign G[74] = in[43] & in2[43];
    assign P[74] = in[43] ^ in2[43];
    assign G[75] = in[42] & in2[42];
    assign P[75] = in[42] ^ in2[42];
    assign G[76] = in[41] & in2[41];
    assign P[76] = in[41] ^ in2[41];
    assign G[77] = in[40] & in2[40];
    assign P[77] = in[40] ^ in2[40];
    assign G[78] = in[39] & in2[39];
    assign P[78] = in[39] ^ in2[39];
    assign G[79] = in[38] & in2[38];
    assign P[79] = in[38] ^ in2[38];
    assign G[80] = in[37] & in2[37];
    assign P[80] = in[37] ^ in2[37];
    assign G[81] = in[36] & in2[36];
    assign P[81] = in[36] ^ in2[36];
    assign G[82] = in[35] & in2[35];
    assign P[82] = in[35] ^ in2[35];
    assign G[83] = in[34] & in2[34];
    assign P[83] = in[34] ^ in2[34];
    assign G[84] = in[33] & in2[33];
    assign P[84] = in[33] ^ in2[33];
    assign G[85] = in[32] & in2[32];
    assign P[85] = in[32] ^ in2[32];
    assign G[86] = in[31] & in2[31];
    assign P[86] = in[31] ^ in2[31];
    assign G[87] = in[30] & in2[30];
    assign P[87] = in[30] ^ in2[30];
    assign G[88] = in[29] & in2[29];
    assign P[88] = in[29] ^ in2[29];
    assign G[89] = in[28] & in2[28];
    assign P[89] = in[28] ^ in2[28];
    assign G[90] = in[27] & in2[27];
    assign P[90] = in[27] ^ in2[27];
    assign G[91] = in[26] & in2[26];
    assign P[91] = in[26] ^ in2[26];
    assign G[92] = in[25] & in2[25];
    assign P[92] = in[25] ^ in2[25];
    assign G[93] = in[24] & in2[24];
    assign P[93] = in[24] ^ in2[24];
    assign G[94] = in[23] & in2[23];
    assign P[94] = in[23] ^ in2[23];
    assign G[95] = in[22] & in2[22];
    assign P[95] = in[22] ^ in2[22];
    assign G[96] = in[21] & in2[21];
    assign P[96] = in[21] ^ in2[21];
    assign G[97] = in[20] & in2[20];
    assign P[97] = in[20] ^ in2[20];
    assign G[98] = in[19] & in2[19];
    assign P[98] = in[19] ^ in2[19];
    assign G[99] = in[18] & in2[18];
    assign P[99] = in[18] ^ in2[18];
    assign G[100] = in[17] & in2[17];
    assign P[100] = in[17] ^ in2[17];
    assign G[101] = in[16] & in2[16];
    assign P[101] = in[16] ^ in2[16];
    assign G[102] = in[15] & in2[15];
    assign P[102] = in[15] ^ in2[15];
    assign G[103] = in[14] & in2[14];
    assign P[103] = in[14] ^ in2[14];
    assign G[104] = in[13] & in2[13];
    assign P[104] = in[13] ^ in2[13];
    assign G[105] = in[12] & in2[12];
    assign P[105] = in[12] ^ in2[12];
    assign G[106] = in[11] & in2[11];
    assign P[106] = in[11] ^ in2[11];
    assign G[107] = in[10] & in2[10];
    assign P[107] = in[10] ^ in2[10];
    assign G[108] = in[9] & in2[9];
    assign P[108] = in[9] ^ in2[9];
    assign G[109] = in[8] & in2[8];
    assign P[109] = in[8] ^ in2[8];
    assign G[110] = in[7] & in2[7];
    assign P[110] = in[7] ^ in2[7];
    assign G[111] = in[6] & in2[6];
    assign P[111] = in[6] ^ in2[6];
    assign G[112] = in[5] & in2[5];
    assign P[112] = in[5] ^ in2[5];
    assign G[113] = in[4] & in2[4];
    assign P[113] = in[4] ^ in2[4];
    assign G[114] = in[3] & in2[3];
    assign P[114] = in[3] ^ in2[3];
    assign G[115] = in[2] & in2[2];
    assign P[115] = in[2] ^ in2[2];
    assign G[116] = in[1] & in2[1];
    assign P[116] = in[1] ^ in2[1];
    assign G[117] = in[0] & in2[0];
    assign P[117] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign C[117] = G[116] | (P[116] & C[116]);
    assign cout = G[117] | (P[117] & C[117]);
    assign sum = P ^ C;
endmodule

module CLA117(output [116:0] sum, output cout, input [116:0] in1, input [116:0] in2;

    wire[116:0] G;
    wire[116:0] C;
    wire[116:0] P;

    assign G[0] = in[116] & in2[116];
    assign P[0] = in[116] ^ in2[116];
    assign G[1] = in[115] & in2[115];
    assign P[1] = in[115] ^ in2[115];
    assign G[2] = in[114] & in2[114];
    assign P[2] = in[114] ^ in2[114];
    assign G[3] = in[113] & in2[113];
    assign P[3] = in[113] ^ in2[113];
    assign G[4] = in[112] & in2[112];
    assign P[4] = in[112] ^ in2[112];
    assign G[5] = in[111] & in2[111];
    assign P[5] = in[111] ^ in2[111];
    assign G[6] = in[110] & in2[110];
    assign P[6] = in[110] ^ in2[110];
    assign G[7] = in[109] & in2[109];
    assign P[7] = in[109] ^ in2[109];
    assign G[8] = in[108] & in2[108];
    assign P[8] = in[108] ^ in2[108];
    assign G[9] = in[107] & in2[107];
    assign P[9] = in[107] ^ in2[107];
    assign G[10] = in[106] & in2[106];
    assign P[10] = in[106] ^ in2[106];
    assign G[11] = in[105] & in2[105];
    assign P[11] = in[105] ^ in2[105];
    assign G[12] = in[104] & in2[104];
    assign P[12] = in[104] ^ in2[104];
    assign G[13] = in[103] & in2[103];
    assign P[13] = in[103] ^ in2[103];
    assign G[14] = in[102] & in2[102];
    assign P[14] = in[102] ^ in2[102];
    assign G[15] = in[101] & in2[101];
    assign P[15] = in[101] ^ in2[101];
    assign G[16] = in[100] & in2[100];
    assign P[16] = in[100] ^ in2[100];
    assign G[17] = in[99] & in2[99];
    assign P[17] = in[99] ^ in2[99];
    assign G[18] = in[98] & in2[98];
    assign P[18] = in[98] ^ in2[98];
    assign G[19] = in[97] & in2[97];
    assign P[19] = in[97] ^ in2[97];
    assign G[20] = in[96] & in2[96];
    assign P[20] = in[96] ^ in2[96];
    assign G[21] = in[95] & in2[95];
    assign P[21] = in[95] ^ in2[95];
    assign G[22] = in[94] & in2[94];
    assign P[22] = in[94] ^ in2[94];
    assign G[23] = in[93] & in2[93];
    assign P[23] = in[93] ^ in2[93];
    assign G[24] = in[92] & in2[92];
    assign P[24] = in[92] ^ in2[92];
    assign G[25] = in[91] & in2[91];
    assign P[25] = in[91] ^ in2[91];
    assign G[26] = in[90] & in2[90];
    assign P[26] = in[90] ^ in2[90];
    assign G[27] = in[89] & in2[89];
    assign P[27] = in[89] ^ in2[89];
    assign G[28] = in[88] & in2[88];
    assign P[28] = in[88] ^ in2[88];
    assign G[29] = in[87] & in2[87];
    assign P[29] = in[87] ^ in2[87];
    assign G[30] = in[86] & in2[86];
    assign P[30] = in[86] ^ in2[86];
    assign G[31] = in[85] & in2[85];
    assign P[31] = in[85] ^ in2[85];
    assign G[32] = in[84] & in2[84];
    assign P[32] = in[84] ^ in2[84];
    assign G[33] = in[83] & in2[83];
    assign P[33] = in[83] ^ in2[83];
    assign G[34] = in[82] & in2[82];
    assign P[34] = in[82] ^ in2[82];
    assign G[35] = in[81] & in2[81];
    assign P[35] = in[81] ^ in2[81];
    assign G[36] = in[80] & in2[80];
    assign P[36] = in[80] ^ in2[80];
    assign G[37] = in[79] & in2[79];
    assign P[37] = in[79] ^ in2[79];
    assign G[38] = in[78] & in2[78];
    assign P[38] = in[78] ^ in2[78];
    assign G[39] = in[77] & in2[77];
    assign P[39] = in[77] ^ in2[77];
    assign G[40] = in[76] & in2[76];
    assign P[40] = in[76] ^ in2[76];
    assign G[41] = in[75] & in2[75];
    assign P[41] = in[75] ^ in2[75];
    assign G[42] = in[74] & in2[74];
    assign P[42] = in[74] ^ in2[74];
    assign G[43] = in[73] & in2[73];
    assign P[43] = in[73] ^ in2[73];
    assign G[44] = in[72] & in2[72];
    assign P[44] = in[72] ^ in2[72];
    assign G[45] = in[71] & in2[71];
    assign P[45] = in[71] ^ in2[71];
    assign G[46] = in[70] & in2[70];
    assign P[46] = in[70] ^ in2[70];
    assign G[47] = in[69] & in2[69];
    assign P[47] = in[69] ^ in2[69];
    assign G[48] = in[68] & in2[68];
    assign P[48] = in[68] ^ in2[68];
    assign G[49] = in[67] & in2[67];
    assign P[49] = in[67] ^ in2[67];
    assign G[50] = in[66] & in2[66];
    assign P[50] = in[66] ^ in2[66];
    assign G[51] = in[65] & in2[65];
    assign P[51] = in[65] ^ in2[65];
    assign G[52] = in[64] & in2[64];
    assign P[52] = in[64] ^ in2[64];
    assign G[53] = in[63] & in2[63];
    assign P[53] = in[63] ^ in2[63];
    assign G[54] = in[62] & in2[62];
    assign P[54] = in[62] ^ in2[62];
    assign G[55] = in[61] & in2[61];
    assign P[55] = in[61] ^ in2[61];
    assign G[56] = in[60] & in2[60];
    assign P[56] = in[60] ^ in2[60];
    assign G[57] = in[59] & in2[59];
    assign P[57] = in[59] ^ in2[59];
    assign G[58] = in[58] & in2[58];
    assign P[58] = in[58] ^ in2[58];
    assign G[59] = in[57] & in2[57];
    assign P[59] = in[57] ^ in2[57];
    assign G[60] = in[56] & in2[56];
    assign P[60] = in[56] ^ in2[56];
    assign G[61] = in[55] & in2[55];
    assign P[61] = in[55] ^ in2[55];
    assign G[62] = in[54] & in2[54];
    assign P[62] = in[54] ^ in2[54];
    assign G[63] = in[53] & in2[53];
    assign P[63] = in[53] ^ in2[53];
    assign G[64] = in[52] & in2[52];
    assign P[64] = in[52] ^ in2[52];
    assign G[65] = in[51] & in2[51];
    assign P[65] = in[51] ^ in2[51];
    assign G[66] = in[50] & in2[50];
    assign P[66] = in[50] ^ in2[50];
    assign G[67] = in[49] & in2[49];
    assign P[67] = in[49] ^ in2[49];
    assign G[68] = in[48] & in2[48];
    assign P[68] = in[48] ^ in2[48];
    assign G[69] = in[47] & in2[47];
    assign P[69] = in[47] ^ in2[47];
    assign G[70] = in[46] & in2[46];
    assign P[70] = in[46] ^ in2[46];
    assign G[71] = in[45] & in2[45];
    assign P[71] = in[45] ^ in2[45];
    assign G[72] = in[44] & in2[44];
    assign P[72] = in[44] ^ in2[44];
    assign G[73] = in[43] & in2[43];
    assign P[73] = in[43] ^ in2[43];
    assign G[74] = in[42] & in2[42];
    assign P[74] = in[42] ^ in2[42];
    assign G[75] = in[41] & in2[41];
    assign P[75] = in[41] ^ in2[41];
    assign G[76] = in[40] & in2[40];
    assign P[76] = in[40] ^ in2[40];
    assign G[77] = in[39] & in2[39];
    assign P[77] = in[39] ^ in2[39];
    assign G[78] = in[38] & in2[38];
    assign P[78] = in[38] ^ in2[38];
    assign G[79] = in[37] & in2[37];
    assign P[79] = in[37] ^ in2[37];
    assign G[80] = in[36] & in2[36];
    assign P[80] = in[36] ^ in2[36];
    assign G[81] = in[35] & in2[35];
    assign P[81] = in[35] ^ in2[35];
    assign G[82] = in[34] & in2[34];
    assign P[82] = in[34] ^ in2[34];
    assign G[83] = in[33] & in2[33];
    assign P[83] = in[33] ^ in2[33];
    assign G[84] = in[32] & in2[32];
    assign P[84] = in[32] ^ in2[32];
    assign G[85] = in[31] & in2[31];
    assign P[85] = in[31] ^ in2[31];
    assign G[86] = in[30] & in2[30];
    assign P[86] = in[30] ^ in2[30];
    assign G[87] = in[29] & in2[29];
    assign P[87] = in[29] ^ in2[29];
    assign G[88] = in[28] & in2[28];
    assign P[88] = in[28] ^ in2[28];
    assign G[89] = in[27] & in2[27];
    assign P[89] = in[27] ^ in2[27];
    assign G[90] = in[26] & in2[26];
    assign P[90] = in[26] ^ in2[26];
    assign G[91] = in[25] & in2[25];
    assign P[91] = in[25] ^ in2[25];
    assign G[92] = in[24] & in2[24];
    assign P[92] = in[24] ^ in2[24];
    assign G[93] = in[23] & in2[23];
    assign P[93] = in[23] ^ in2[23];
    assign G[94] = in[22] & in2[22];
    assign P[94] = in[22] ^ in2[22];
    assign G[95] = in[21] & in2[21];
    assign P[95] = in[21] ^ in2[21];
    assign G[96] = in[20] & in2[20];
    assign P[96] = in[20] ^ in2[20];
    assign G[97] = in[19] & in2[19];
    assign P[97] = in[19] ^ in2[19];
    assign G[98] = in[18] & in2[18];
    assign P[98] = in[18] ^ in2[18];
    assign G[99] = in[17] & in2[17];
    assign P[99] = in[17] ^ in2[17];
    assign G[100] = in[16] & in2[16];
    assign P[100] = in[16] ^ in2[16];
    assign G[101] = in[15] & in2[15];
    assign P[101] = in[15] ^ in2[15];
    assign G[102] = in[14] & in2[14];
    assign P[102] = in[14] ^ in2[14];
    assign G[103] = in[13] & in2[13];
    assign P[103] = in[13] ^ in2[13];
    assign G[104] = in[12] & in2[12];
    assign P[104] = in[12] ^ in2[12];
    assign G[105] = in[11] & in2[11];
    assign P[105] = in[11] ^ in2[11];
    assign G[106] = in[10] & in2[10];
    assign P[106] = in[10] ^ in2[10];
    assign G[107] = in[9] & in2[9];
    assign P[107] = in[9] ^ in2[9];
    assign G[108] = in[8] & in2[8];
    assign P[108] = in[8] ^ in2[8];
    assign G[109] = in[7] & in2[7];
    assign P[109] = in[7] ^ in2[7];
    assign G[110] = in[6] & in2[6];
    assign P[110] = in[6] ^ in2[6];
    assign G[111] = in[5] & in2[5];
    assign P[111] = in[5] ^ in2[5];
    assign G[112] = in[4] & in2[4];
    assign P[112] = in[4] ^ in2[4];
    assign G[113] = in[3] & in2[3];
    assign P[113] = in[3] ^ in2[3];
    assign G[114] = in[2] & in2[2];
    assign P[114] = in[2] ^ in2[2];
    assign G[115] = in[1] & in2[1];
    assign P[115] = in[1] ^ in2[1];
    assign G[116] = in[0] & in2[0];
    assign P[116] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign C[116] = G[115] | (P[115] & C[115]);
    assign cout = G[116] | (P[116] & C[116]);
    assign sum = P ^ C;
endmodule

module CLA116(output [115:0] sum, output cout, input [115:0] in1, input [115:0] in2;

    wire[115:0] G;
    wire[115:0] C;
    wire[115:0] P;

    assign G[0] = in[115] & in2[115];
    assign P[0] = in[115] ^ in2[115];
    assign G[1] = in[114] & in2[114];
    assign P[1] = in[114] ^ in2[114];
    assign G[2] = in[113] & in2[113];
    assign P[2] = in[113] ^ in2[113];
    assign G[3] = in[112] & in2[112];
    assign P[3] = in[112] ^ in2[112];
    assign G[4] = in[111] & in2[111];
    assign P[4] = in[111] ^ in2[111];
    assign G[5] = in[110] & in2[110];
    assign P[5] = in[110] ^ in2[110];
    assign G[6] = in[109] & in2[109];
    assign P[6] = in[109] ^ in2[109];
    assign G[7] = in[108] & in2[108];
    assign P[7] = in[108] ^ in2[108];
    assign G[8] = in[107] & in2[107];
    assign P[8] = in[107] ^ in2[107];
    assign G[9] = in[106] & in2[106];
    assign P[9] = in[106] ^ in2[106];
    assign G[10] = in[105] & in2[105];
    assign P[10] = in[105] ^ in2[105];
    assign G[11] = in[104] & in2[104];
    assign P[11] = in[104] ^ in2[104];
    assign G[12] = in[103] & in2[103];
    assign P[12] = in[103] ^ in2[103];
    assign G[13] = in[102] & in2[102];
    assign P[13] = in[102] ^ in2[102];
    assign G[14] = in[101] & in2[101];
    assign P[14] = in[101] ^ in2[101];
    assign G[15] = in[100] & in2[100];
    assign P[15] = in[100] ^ in2[100];
    assign G[16] = in[99] & in2[99];
    assign P[16] = in[99] ^ in2[99];
    assign G[17] = in[98] & in2[98];
    assign P[17] = in[98] ^ in2[98];
    assign G[18] = in[97] & in2[97];
    assign P[18] = in[97] ^ in2[97];
    assign G[19] = in[96] & in2[96];
    assign P[19] = in[96] ^ in2[96];
    assign G[20] = in[95] & in2[95];
    assign P[20] = in[95] ^ in2[95];
    assign G[21] = in[94] & in2[94];
    assign P[21] = in[94] ^ in2[94];
    assign G[22] = in[93] & in2[93];
    assign P[22] = in[93] ^ in2[93];
    assign G[23] = in[92] & in2[92];
    assign P[23] = in[92] ^ in2[92];
    assign G[24] = in[91] & in2[91];
    assign P[24] = in[91] ^ in2[91];
    assign G[25] = in[90] & in2[90];
    assign P[25] = in[90] ^ in2[90];
    assign G[26] = in[89] & in2[89];
    assign P[26] = in[89] ^ in2[89];
    assign G[27] = in[88] & in2[88];
    assign P[27] = in[88] ^ in2[88];
    assign G[28] = in[87] & in2[87];
    assign P[28] = in[87] ^ in2[87];
    assign G[29] = in[86] & in2[86];
    assign P[29] = in[86] ^ in2[86];
    assign G[30] = in[85] & in2[85];
    assign P[30] = in[85] ^ in2[85];
    assign G[31] = in[84] & in2[84];
    assign P[31] = in[84] ^ in2[84];
    assign G[32] = in[83] & in2[83];
    assign P[32] = in[83] ^ in2[83];
    assign G[33] = in[82] & in2[82];
    assign P[33] = in[82] ^ in2[82];
    assign G[34] = in[81] & in2[81];
    assign P[34] = in[81] ^ in2[81];
    assign G[35] = in[80] & in2[80];
    assign P[35] = in[80] ^ in2[80];
    assign G[36] = in[79] & in2[79];
    assign P[36] = in[79] ^ in2[79];
    assign G[37] = in[78] & in2[78];
    assign P[37] = in[78] ^ in2[78];
    assign G[38] = in[77] & in2[77];
    assign P[38] = in[77] ^ in2[77];
    assign G[39] = in[76] & in2[76];
    assign P[39] = in[76] ^ in2[76];
    assign G[40] = in[75] & in2[75];
    assign P[40] = in[75] ^ in2[75];
    assign G[41] = in[74] & in2[74];
    assign P[41] = in[74] ^ in2[74];
    assign G[42] = in[73] & in2[73];
    assign P[42] = in[73] ^ in2[73];
    assign G[43] = in[72] & in2[72];
    assign P[43] = in[72] ^ in2[72];
    assign G[44] = in[71] & in2[71];
    assign P[44] = in[71] ^ in2[71];
    assign G[45] = in[70] & in2[70];
    assign P[45] = in[70] ^ in2[70];
    assign G[46] = in[69] & in2[69];
    assign P[46] = in[69] ^ in2[69];
    assign G[47] = in[68] & in2[68];
    assign P[47] = in[68] ^ in2[68];
    assign G[48] = in[67] & in2[67];
    assign P[48] = in[67] ^ in2[67];
    assign G[49] = in[66] & in2[66];
    assign P[49] = in[66] ^ in2[66];
    assign G[50] = in[65] & in2[65];
    assign P[50] = in[65] ^ in2[65];
    assign G[51] = in[64] & in2[64];
    assign P[51] = in[64] ^ in2[64];
    assign G[52] = in[63] & in2[63];
    assign P[52] = in[63] ^ in2[63];
    assign G[53] = in[62] & in2[62];
    assign P[53] = in[62] ^ in2[62];
    assign G[54] = in[61] & in2[61];
    assign P[54] = in[61] ^ in2[61];
    assign G[55] = in[60] & in2[60];
    assign P[55] = in[60] ^ in2[60];
    assign G[56] = in[59] & in2[59];
    assign P[56] = in[59] ^ in2[59];
    assign G[57] = in[58] & in2[58];
    assign P[57] = in[58] ^ in2[58];
    assign G[58] = in[57] & in2[57];
    assign P[58] = in[57] ^ in2[57];
    assign G[59] = in[56] & in2[56];
    assign P[59] = in[56] ^ in2[56];
    assign G[60] = in[55] & in2[55];
    assign P[60] = in[55] ^ in2[55];
    assign G[61] = in[54] & in2[54];
    assign P[61] = in[54] ^ in2[54];
    assign G[62] = in[53] & in2[53];
    assign P[62] = in[53] ^ in2[53];
    assign G[63] = in[52] & in2[52];
    assign P[63] = in[52] ^ in2[52];
    assign G[64] = in[51] & in2[51];
    assign P[64] = in[51] ^ in2[51];
    assign G[65] = in[50] & in2[50];
    assign P[65] = in[50] ^ in2[50];
    assign G[66] = in[49] & in2[49];
    assign P[66] = in[49] ^ in2[49];
    assign G[67] = in[48] & in2[48];
    assign P[67] = in[48] ^ in2[48];
    assign G[68] = in[47] & in2[47];
    assign P[68] = in[47] ^ in2[47];
    assign G[69] = in[46] & in2[46];
    assign P[69] = in[46] ^ in2[46];
    assign G[70] = in[45] & in2[45];
    assign P[70] = in[45] ^ in2[45];
    assign G[71] = in[44] & in2[44];
    assign P[71] = in[44] ^ in2[44];
    assign G[72] = in[43] & in2[43];
    assign P[72] = in[43] ^ in2[43];
    assign G[73] = in[42] & in2[42];
    assign P[73] = in[42] ^ in2[42];
    assign G[74] = in[41] & in2[41];
    assign P[74] = in[41] ^ in2[41];
    assign G[75] = in[40] & in2[40];
    assign P[75] = in[40] ^ in2[40];
    assign G[76] = in[39] & in2[39];
    assign P[76] = in[39] ^ in2[39];
    assign G[77] = in[38] & in2[38];
    assign P[77] = in[38] ^ in2[38];
    assign G[78] = in[37] & in2[37];
    assign P[78] = in[37] ^ in2[37];
    assign G[79] = in[36] & in2[36];
    assign P[79] = in[36] ^ in2[36];
    assign G[80] = in[35] & in2[35];
    assign P[80] = in[35] ^ in2[35];
    assign G[81] = in[34] & in2[34];
    assign P[81] = in[34] ^ in2[34];
    assign G[82] = in[33] & in2[33];
    assign P[82] = in[33] ^ in2[33];
    assign G[83] = in[32] & in2[32];
    assign P[83] = in[32] ^ in2[32];
    assign G[84] = in[31] & in2[31];
    assign P[84] = in[31] ^ in2[31];
    assign G[85] = in[30] & in2[30];
    assign P[85] = in[30] ^ in2[30];
    assign G[86] = in[29] & in2[29];
    assign P[86] = in[29] ^ in2[29];
    assign G[87] = in[28] & in2[28];
    assign P[87] = in[28] ^ in2[28];
    assign G[88] = in[27] & in2[27];
    assign P[88] = in[27] ^ in2[27];
    assign G[89] = in[26] & in2[26];
    assign P[89] = in[26] ^ in2[26];
    assign G[90] = in[25] & in2[25];
    assign P[90] = in[25] ^ in2[25];
    assign G[91] = in[24] & in2[24];
    assign P[91] = in[24] ^ in2[24];
    assign G[92] = in[23] & in2[23];
    assign P[92] = in[23] ^ in2[23];
    assign G[93] = in[22] & in2[22];
    assign P[93] = in[22] ^ in2[22];
    assign G[94] = in[21] & in2[21];
    assign P[94] = in[21] ^ in2[21];
    assign G[95] = in[20] & in2[20];
    assign P[95] = in[20] ^ in2[20];
    assign G[96] = in[19] & in2[19];
    assign P[96] = in[19] ^ in2[19];
    assign G[97] = in[18] & in2[18];
    assign P[97] = in[18] ^ in2[18];
    assign G[98] = in[17] & in2[17];
    assign P[98] = in[17] ^ in2[17];
    assign G[99] = in[16] & in2[16];
    assign P[99] = in[16] ^ in2[16];
    assign G[100] = in[15] & in2[15];
    assign P[100] = in[15] ^ in2[15];
    assign G[101] = in[14] & in2[14];
    assign P[101] = in[14] ^ in2[14];
    assign G[102] = in[13] & in2[13];
    assign P[102] = in[13] ^ in2[13];
    assign G[103] = in[12] & in2[12];
    assign P[103] = in[12] ^ in2[12];
    assign G[104] = in[11] & in2[11];
    assign P[104] = in[11] ^ in2[11];
    assign G[105] = in[10] & in2[10];
    assign P[105] = in[10] ^ in2[10];
    assign G[106] = in[9] & in2[9];
    assign P[106] = in[9] ^ in2[9];
    assign G[107] = in[8] & in2[8];
    assign P[107] = in[8] ^ in2[8];
    assign G[108] = in[7] & in2[7];
    assign P[108] = in[7] ^ in2[7];
    assign G[109] = in[6] & in2[6];
    assign P[109] = in[6] ^ in2[6];
    assign G[110] = in[5] & in2[5];
    assign P[110] = in[5] ^ in2[5];
    assign G[111] = in[4] & in2[4];
    assign P[111] = in[4] ^ in2[4];
    assign G[112] = in[3] & in2[3];
    assign P[112] = in[3] ^ in2[3];
    assign G[113] = in[2] & in2[2];
    assign P[113] = in[2] ^ in2[2];
    assign G[114] = in[1] & in2[1];
    assign P[114] = in[1] ^ in2[1];
    assign G[115] = in[0] & in2[0];
    assign P[115] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign C[115] = G[114] | (P[114] & C[114]);
    assign cout = G[115] | (P[115] & C[115]);
    assign sum = P ^ C;
endmodule

module CLA115(output [114:0] sum, output cout, input [114:0] in1, input [114:0] in2;

    wire[114:0] G;
    wire[114:0] C;
    wire[114:0] P;

    assign G[0] = in[114] & in2[114];
    assign P[0] = in[114] ^ in2[114];
    assign G[1] = in[113] & in2[113];
    assign P[1] = in[113] ^ in2[113];
    assign G[2] = in[112] & in2[112];
    assign P[2] = in[112] ^ in2[112];
    assign G[3] = in[111] & in2[111];
    assign P[3] = in[111] ^ in2[111];
    assign G[4] = in[110] & in2[110];
    assign P[4] = in[110] ^ in2[110];
    assign G[5] = in[109] & in2[109];
    assign P[5] = in[109] ^ in2[109];
    assign G[6] = in[108] & in2[108];
    assign P[6] = in[108] ^ in2[108];
    assign G[7] = in[107] & in2[107];
    assign P[7] = in[107] ^ in2[107];
    assign G[8] = in[106] & in2[106];
    assign P[8] = in[106] ^ in2[106];
    assign G[9] = in[105] & in2[105];
    assign P[9] = in[105] ^ in2[105];
    assign G[10] = in[104] & in2[104];
    assign P[10] = in[104] ^ in2[104];
    assign G[11] = in[103] & in2[103];
    assign P[11] = in[103] ^ in2[103];
    assign G[12] = in[102] & in2[102];
    assign P[12] = in[102] ^ in2[102];
    assign G[13] = in[101] & in2[101];
    assign P[13] = in[101] ^ in2[101];
    assign G[14] = in[100] & in2[100];
    assign P[14] = in[100] ^ in2[100];
    assign G[15] = in[99] & in2[99];
    assign P[15] = in[99] ^ in2[99];
    assign G[16] = in[98] & in2[98];
    assign P[16] = in[98] ^ in2[98];
    assign G[17] = in[97] & in2[97];
    assign P[17] = in[97] ^ in2[97];
    assign G[18] = in[96] & in2[96];
    assign P[18] = in[96] ^ in2[96];
    assign G[19] = in[95] & in2[95];
    assign P[19] = in[95] ^ in2[95];
    assign G[20] = in[94] & in2[94];
    assign P[20] = in[94] ^ in2[94];
    assign G[21] = in[93] & in2[93];
    assign P[21] = in[93] ^ in2[93];
    assign G[22] = in[92] & in2[92];
    assign P[22] = in[92] ^ in2[92];
    assign G[23] = in[91] & in2[91];
    assign P[23] = in[91] ^ in2[91];
    assign G[24] = in[90] & in2[90];
    assign P[24] = in[90] ^ in2[90];
    assign G[25] = in[89] & in2[89];
    assign P[25] = in[89] ^ in2[89];
    assign G[26] = in[88] & in2[88];
    assign P[26] = in[88] ^ in2[88];
    assign G[27] = in[87] & in2[87];
    assign P[27] = in[87] ^ in2[87];
    assign G[28] = in[86] & in2[86];
    assign P[28] = in[86] ^ in2[86];
    assign G[29] = in[85] & in2[85];
    assign P[29] = in[85] ^ in2[85];
    assign G[30] = in[84] & in2[84];
    assign P[30] = in[84] ^ in2[84];
    assign G[31] = in[83] & in2[83];
    assign P[31] = in[83] ^ in2[83];
    assign G[32] = in[82] & in2[82];
    assign P[32] = in[82] ^ in2[82];
    assign G[33] = in[81] & in2[81];
    assign P[33] = in[81] ^ in2[81];
    assign G[34] = in[80] & in2[80];
    assign P[34] = in[80] ^ in2[80];
    assign G[35] = in[79] & in2[79];
    assign P[35] = in[79] ^ in2[79];
    assign G[36] = in[78] & in2[78];
    assign P[36] = in[78] ^ in2[78];
    assign G[37] = in[77] & in2[77];
    assign P[37] = in[77] ^ in2[77];
    assign G[38] = in[76] & in2[76];
    assign P[38] = in[76] ^ in2[76];
    assign G[39] = in[75] & in2[75];
    assign P[39] = in[75] ^ in2[75];
    assign G[40] = in[74] & in2[74];
    assign P[40] = in[74] ^ in2[74];
    assign G[41] = in[73] & in2[73];
    assign P[41] = in[73] ^ in2[73];
    assign G[42] = in[72] & in2[72];
    assign P[42] = in[72] ^ in2[72];
    assign G[43] = in[71] & in2[71];
    assign P[43] = in[71] ^ in2[71];
    assign G[44] = in[70] & in2[70];
    assign P[44] = in[70] ^ in2[70];
    assign G[45] = in[69] & in2[69];
    assign P[45] = in[69] ^ in2[69];
    assign G[46] = in[68] & in2[68];
    assign P[46] = in[68] ^ in2[68];
    assign G[47] = in[67] & in2[67];
    assign P[47] = in[67] ^ in2[67];
    assign G[48] = in[66] & in2[66];
    assign P[48] = in[66] ^ in2[66];
    assign G[49] = in[65] & in2[65];
    assign P[49] = in[65] ^ in2[65];
    assign G[50] = in[64] & in2[64];
    assign P[50] = in[64] ^ in2[64];
    assign G[51] = in[63] & in2[63];
    assign P[51] = in[63] ^ in2[63];
    assign G[52] = in[62] & in2[62];
    assign P[52] = in[62] ^ in2[62];
    assign G[53] = in[61] & in2[61];
    assign P[53] = in[61] ^ in2[61];
    assign G[54] = in[60] & in2[60];
    assign P[54] = in[60] ^ in2[60];
    assign G[55] = in[59] & in2[59];
    assign P[55] = in[59] ^ in2[59];
    assign G[56] = in[58] & in2[58];
    assign P[56] = in[58] ^ in2[58];
    assign G[57] = in[57] & in2[57];
    assign P[57] = in[57] ^ in2[57];
    assign G[58] = in[56] & in2[56];
    assign P[58] = in[56] ^ in2[56];
    assign G[59] = in[55] & in2[55];
    assign P[59] = in[55] ^ in2[55];
    assign G[60] = in[54] & in2[54];
    assign P[60] = in[54] ^ in2[54];
    assign G[61] = in[53] & in2[53];
    assign P[61] = in[53] ^ in2[53];
    assign G[62] = in[52] & in2[52];
    assign P[62] = in[52] ^ in2[52];
    assign G[63] = in[51] & in2[51];
    assign P[63] = in[51] ^ in2[51];
    assign G[64] = in[50] & in2[50];
    assign P[64] = in[50] ^ in2[50];
    assign G[65] = in[49] & in2[49];
    assign P[65] = in[49] ^ in2[49];
    assign G[66] = in[48] & in2[48];
    assign P[66] = in[48] ^ in2[48];
    assign G[67] = in[47] & in2[47];
    assign P[67] = in[47] ^ in2[47];
    assign G[68] = in[46] & in2[46];
    assign P[68] = in[46] ^ in2[46];
    assign G[69] = in[45] & in2[45];
    assign P[69] = in[45] ^ in2[45];
    assign G[70] = in[44] & in2[44];
    assign P[70] = in[44] ^ in2[44];
    assign G[71] = in[43] & in2[43];
    assign P[71] = in[43] ^ in2[43];
    assign G[72] = in[42] & in2[42];
    assign P[72] = in[42] ^ in2[42];
    assign G[73] = in[41] & in2[41];
    assign P[73] = in[41] ^ in2[41];
    assign G[74] = in[40] & in2[40];
    assign P[74] = in[40] ^ in2[40];
    assign G[75] = in[39] & in2[39];
    assign P[75] = in[39] ^ in2[39];
    assign G[76] = in[38] & in2[38];
    assign P[76] = in[38] ^ in2[38];
    assign G[77] = in[37] & in2[37];
    assign P[77] = in[37] ^ in2[37];
    assign G[78] = in[36] & in2[36];
    assign P[78] = in[36] ^ in2[36];
    assign G[79] = in[35] & in2[35];
    assign P[79] = in[35] ^ in2[35];
    assign G[80] = in[34] & in2[34];
    assign P[80] = in[34] ^ in2[34];
    assign G[81] = in[33] & in2[33];
    assign P[81] = in[33] ^ in2[33];
    assign G[82] = in[32] & in2[32];
    assign P[82] = in[32] ^ in2[32];
    assign G[83] = in[31] & in2[31];
    assign P[83] = in[31] ^ in2[31];
    assign G[84] = in[30] & in2[30];
    assign P[84] = in[30] ^ in2[30];
    assign G[85] = in[29] & in2[29];
    assign P[85] = in[29] ^ in2[29];
    assign G[86] = in[28] & in2[28];
    assign P[86] = in[28] ^ in2[28];
    assign G[87] = in[27] & in2[27];
    assign P[87] = in[27] ^ in2[27];
    assign G[88] = in[26] & in2[26];
    assign P[88] = in[26] ^ in2[26];
    assign G[89] = in[25] & in2[25];
    assign P[89] = in[25] ^ in2[25];
    assign G[90] = in[24] & in2[24];
    assign P[90] = in[24] ^ in2[24];
    assign G[91] = in[23] & in2[23];
    assign P[91] = in[23] ^ in2[23];
    assign G[92] = in[22] & in2[22];
    assign P[92] = in[22] ^ in2[22];
    assign G[93] = in[21] & in2[21];
    assign P[93] = in[21] ^ in2[21];
    assign G[94] = in[20] & in2[20];
    assign P[94] = in[20] ^ in2[20];
    assign G[95] = in[19] & in2[19];
    assign P[95] = in[19] ^ in2[19];
    assign G[96] = in[18] & in2[18];
    assign P[96] = in[18] ^ in2[18];
    assign G[97] = in[17] & in2[17];
    assign P[97] = in[17] ^ in2[17];
    assign G[98] = in[16] & in2[16];
    assign P[98] = in[16] ^ in2[16];
    assign G[99] = in[15] & in2[15];
    assign P[99] = in[15] ^ in2[15];
    assign G[100] = in[14] & in2[14];
    assign P[100] = in[14] ^ in2[14];
    assign G[101] = in[13] & in2[13];
    assign P[101] = in[13] ^ in2[13];
    assign G[102] = in[12] & in2[12];
    assign P[102] = in[12] ^ in2[12];
    assign G[103] = in[11] & in2[11];
    assign P[103] = in[11] ^ in2[11];
    assign G[104] = in[10] & in2[10];
    assign P[104] = in[10] ^ in2[10];
    assign G[105] = in[9] & in2[9];
    assign P[105] = in[9] ^ in2[9];
    assign G[106] = in[8] & in2[8];
    assign P[106] = in[8] ^ in2[8];
    assign G[107] = in[7] & in2[7];
    assign P[107] = in[7] ^ in2[7];
    assign G[108] = in[6] & in2[6];
    assign P[108] = in[6] ^ in2[6];
    assign G[109] = in[5] & in2[5];
    assign P[109] = in[5] ^ in2[5];
    assign G[110] = in[4] & in2[4];
    assign P[110] = in[4] ^ in2[4];
    assign G[111] = in[3] & in2[3];
    assign P[111] = in[3] ^ in2[3];
    assign G[112] = in[2] & in2[2];
    assign P[112] = in[2] ^ in2[2];
    assign G[113] = in[1] & in2[1];
    assign P[113] = in[1] ^ in2[1];
    assign G[114] = in[0] & in2[0];
    assign P[114] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign C[114] = G[113] | (P[113] & C[113]);
    assign cout = G[114] | (P[114] & C[114]);
    assign sum = P ^ C;
endmodule

module CLA114(output [113:0] sum, output cout, input [113:0] in1, input [113:0] in2;

    wire[113:0] G;
    wire[113:0] C;
    wire[113:0] P;

    assign G[0] = in[113] & in2[113];
    assign P[0] = in[113] ^ in2[113];
    assign G[1] = in[112] & in2[112];
    assign P[1] = in[112] ^ in2[112];
    assign G[2] = in[111] & in2[111];
    assign P[2] = in[111] ^ in2[111];
    assign G[3] = in[110] & in2[110];
    assign P[3] = in[110] ^ in2[110];
    assign G[4] = in[109] & in2[109];
    assign P[4] = in[109] ^ in2[109];
    assign G[5] = in[108] & in2[108];
    assign P[5] = in[108] ^ in2[108];
    assign G[6] = in[107] & in2[107];
    assign P[6] = in[107] ^ in2[107];
    assign G[7] = in[106] & in2[106];
    assign P[7] = in[106] ^ in2[106];
    assign G[8] = in[105] & in2[105];
    assign P[8] = in[105] ^ in2[105];
    assign G[9] = in[104] & in2[104];
    assign P[9] = in[104] ^ in2[104];
    assign G[10] = in[103] & in2[103];
    assign P[10] = in[103] ^ in2[103];
    assign G[11] = in[102] & in2[102];
    assign P[11] = in[102] ^ in2[102];
    assign G[12] = in[101] & in2[101];
    assign P[12] = in[101] ^ in2[101];
    assign G[13] = in[100] & in2[100];
    assign P[13] = in[100] ^ in2[100];
    assign G[14] = in[99] & in2[99];
    assign P[14] = in[99] ^ in2[99];
    assign G[15] = in[98] & in2[98];
    assign P[15] = in[98] ^ in2[98];
    assign G[16] = in[97] & in2[97];
    assign P[16] = in[97] ^ in2[97];
    assign G[17] = in[96] & in2[96];
    assign P[17] = in[96] ^ in2[96];
    assign G[18] = in[95] & in2[95];
    assign P[18] = in[95] ^ in2[95];
    assign G[19] = in[94] & in2[94];
    assign P[19] = in[94] ^ in2[94];
    assign G[20] = in[93] & in2[93];
    assign P[20] = in[93] ^ in2[93];
    assign G[21] = in[92] & in2[92];
    assign P[21] = in[92] ^ in2[92];
    assign G[22] = in[91] & in2[91];
    assign P[22] = in[91] ^ in2[91];
    assign G[23] = in[90] & in2[90];
    assign P[23] = in[90] ^ in2[90];
    assign G[24] = in[89] & in2[89];
    assign P[24] = in[89] ^ in2[89];
    assign G[25] = in[88] & in2[88];
    assign P[25] = in[88] ^ in2[88];
    assign G[26] = in[87] & in2[87];
    assign P[26] = in[87] ^ in2[87];
    assign G[27] = in[86] & in2[86];
    assign P[27] = in[86] ^ in2[86];
    assign G[28] = in[85] & in2[85];
    assign P[28] = in[85] ^ in2[85];
    assign G[29] = in[84] & in2[84];
    assign P[29] = in[84] ^ in2[84];
    assign G[30] = in[83] & in2[83];
    assign P[30] = in[83] ^ in2[83];
    assign G[31] = in[82] & in2[82];
    assign P[31] = in[82] ^ in2[82];
    assign G[32] = in[81] & in2[81];
    assign P[32] = in[81] ^ in2[81];
    assign G[33] = in[80] & in2[80];
    assign P[33] = in[80] ^ in2[80];
    assign G[34] = in[79] & in2[79];
    assign P[34] = in[79] ^ in2[79];
    assign G[35] = in[78] & in2[78];
    assign P[35] = in[78] ^ in2[78];
    assign G[36] = in[77] & in2[77];
    assign P[36] = in[77] ^ in2[77];
    assign G[37] = in[76] & in2[76];
    assign P[37] = in[76] ^ in2[76];
    assign G[38] = in[75] & in2[75];
    assign P[38] = in[75] ^ in2[75];
    assign G[39] = in[74] & in2[74];
    assign P[39] = in[74] ^ in2[74];
    assign G[40] = in[73] & in2[73];
    assign P[40] = in[73] ^ in2[73];
    assign G[41] = in[72] & in2[72];
    assign P[41] = in[72] ^ in2[72];
    assign G[42] = in[71] & in2[71];
    assign P[42] = in[71] ^ in2[71];
    assign G[43] = in[70] & in2[70];
    assign P[43] = in[70] ^ in2[70];
    assign G[44] = in[69] & in2[69];
    assign P[44] = in[69] ^ in2[69];
    assign G[45] = in[68] & in2[68];
    assign P[45] = in[68] ^ in2[68];
    assign G[46] = in[67] & in2[67];
    assign P[46] = in[67] ^ in2[67];
    assign G[47] = in[66] & in2[66];
    assign P[47] = in[66] ^ in2[66];
    assign G[48] = in[65] & in2[65];
    assign P[48] = in[65] ^ in2[65];
    assign G[49] = in[64] & in2[64];
    assign P[49] = in[64] ^ in2[64];
    assign G[50] = in[63] & in2[63];
    assign P[50] = in[63] ^ in2[63];
    assign G[51] = in[62] & in2[62];
    assign P[51] = in[62] ^ in2[62];
    assign G[52] = in[61] & in2[61];
    assign P[52] = in[61] ^ in2[61];
    assign G[53] = in[60] & in2[60];
    assign P[53] = in[60] ^ in2[60];
    assign G[54] = in[59] & in2[59];
    assign P[54] = in[59] ^ in2[59];
    assign G[55] = in[58] & in2[58];
    assign P[55] = in[58] ^ in2[58];
    assign G[56] = in[57] & in2[57];
    assign P[56] = in[57] ^ in2[57];
    assign G[57] = in[56] & in2[56];
    assign P[57] = in[56] ^ in2[56];
    assign G[58] = in[55] & in2[55];
    assign P[58] = in[55] ^ in2[55];
    assign G[59] = in[54] & in2[54];
    assign P[59] = in[54] ^ in2[54];
    assign G[60] = in[53] & in2[53];
    assign P[60] = in[53] ^ in2[53];
    assign G[61] = in[52] & in2[52];
    assign P[61] = in[52] ^ in2[52];
    assign G[62] = in[51] & in2[51];
    assign P[62] = in[51] ^ in2[51];
    assign G[63] = in[50] & in2[50];
    assign P[63] = in[50] ^ in2[50];
    assign G[64] = in[49] & in2[49];
    assign P[64] = in[49] ^ in2[49];
    assign G[65] = in[48] & in2[48];
    assign P[65] = in[48] ^ in2[48];
    assign G[66] = in[47] & in2[47];
    assign P[66] = in[47] ^ in2[47];
    assign G[67] = in[46] & in2[46];
    assign P[67] = in[46] ^ in2[46];
    assign G[68] = in[45] & in2[45];
    assign P[68] = in[45] ^ in2[45];
    assign G[69] = in[44] & in2[44];
    assign P[69] = in[44] ^ in2[44];
    assign G[70] = in[43] & in2[43];
    assign P[70] = in[43] ^ in2[43];
    assign G[71] = in[42] & in2[42];
    assign P[71] = in[42] ^ in2[42];
    assign G[72] = in[41] & in2[41];
    assign P[72] = in[41] ^ in2[41];
    assign G[73] = in[40] & in2[40];
    assign P[73] = in[40] ^ in2[40];
    assign G[74] = in[39] & in2[39];
    assign P[74] = in[39] ^ in2[39];
    assign G[75] = in[38] & in2[38];
    assign P[75] = in[38] ^ in2[38];
    assign G[76] = in[37] & in2[37];
    assign P[76] = in[37] ^ in2[37];
    assign G[77] = in[36] & in2[36];
    assign P[77] = in[36] ^ in2[36];
    assign G[78] = in[35] & in2[35];
    assign P[78] = in[35] ^ in2[35];
    assign G[79] = in[34] & in2[34];
    assign P[79] = in[34] ^ in2[34];
    assign G[80] = in[33] & in2[33];
    assign P[80] = in[33] ^ in2[33];
    assign G[81] = in[32] & in2[32];
    assign P[81] = in[32] ^ in2[32];
    assign G[82] = in[31] & in2[31];
    assign P[82] = in[31] ^ in2[31];
    assign G[83] = in[30] & in2[30];
    assign P[83] = in[30] ^ in2[30];
    assign G[84] = in[29] & in2[29];
    assign P[84] = in[29] ^ in2[29];
    assign G[85] = in[28] & in2[28];
    assign P[85] = in[28] ^ in2[28];
    assign G[86] = in[27] & in2[27];
    assign P[86] = in[27] ^ in2[27];
    assign G[87] = in[26] & in2[26];
    assign P[87] = in[26] ^ in2[26];
    assign G[88] = in[25] & in2[25];
    assign P[88] = in[25] ^ in2[25];
    assign G[89] = in[24] & in2[24];
    assign P[89] = in[24] ^ in2[24];
    assign G[90] = in[23] & in2[23];
    assign P[90] = in[23] ^ in2[23];
    assign G[91] = in[22] & in2[22];
    assign P[91] = in[22] ^ in2[22];
    assign G[92] = in[21] & in2[21];
    assign P[92] = in[21] ^ in2[21];
    assign G[93] = in[20] & in2[20];
    assign P[93] = in[20] ^ in2[20];
    assign G[94] = in[19] & in2[19];
    assign P[94] = in[19] ^ in2[19];
    assign G[95] = in[18] & in2[18];
    assign P[95] = in[18] ^ in2[18];
    assign G[96] = in[17] & in2[17];
    assign P[96] = in[17] ^ in2[17];
    assign G[97] = in[16] & in2[16];
    assign P[97] = in[16] ^ in2[16];
    assign G[98] = in[15] & in2[15];
    assign P[98] = in[15] ^ in2[15];
    assign G[99] = in[14] & in2[14];
    assign P[99] = in[14] ^ in2[14];
    assign G[100] = in[13] & in2[13];
    assign P[100] = in[13] ^ in2[13];
    assign G[101] = in[12] & in2[12];
    assign P[101] = in[12] ^ in2[12];
    assign G[102] = in[11] & in2[11];
    assign P[102] = in[11] ^ in2[11];
    assign G[103] = in[10] & in2[10];
    assign P[103] = in[10] ^ in2[10];
    assign G[104] = in[9] & in2[9];
    assign P[104] = in[9] ^ in2[9];
    assign G[105] = in[8] & in2[8];
    assign P[105] = in[8] ^ in2[8];
    assign G[106] = in[7] & in2[7];
    assign P[106] = in[7] ^ in2[7];
    assign G[107] = in[6] & in2[6];
    assign P[107] = in[6] ^ in2[6];
    assign G[108] = in[5] & in2[5];
    assign P[108] = in[5] ^ in2[5];
    assign G[109] = in[4] & in2[4];
    assign P[109] = in[4] ^ in2[4];
    assign G[110] = in[3] & in2[3];
    assign P[110] = in[3] ^ in2[3];
    assign G[111] = in[2] & in2[2];
    assign P[111] = in[2] ^ in2[2];
    assign G[112] = in[1] & in2[1];
    assign P[112] = in[1] ^ in2[1];
    assign G[113] = in[0] & in2[0];
    assign P[113] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign C[113] = G[112] | (P[112] & C[112]);
    assign cout = G[113] | (P[113] & C[113]);
    assign sum = P ^ C;
endmodule

module CLA113(output [112:0] sum, output cout, input [112:0] in1, input [112:0] in2;

    wire[112:0] G;
    wire[112:0] C;
    wire[112:0] P;

    assign G[0] = in[112] & in2[112];
    assign P[0] = in[112] ^ in2[112];
    assign G[1] = in[111] & in2[111];
    assign P[1] = in[111] ^ in2[111];
    assign G[2] = in[110] & in2[110];
    assign P[2] = in[110] ^ in2[110];
    assign G[3] = in[109] & in2[109];
    assign P[3] = in[109] ^ in2[109];
    assign G[4] = in[108] & in2[108];
    assign P[4] = in[108] ^ in2[108];
    assign G[5] = in[107] & in2[107];
    assign P[5] = in[107] ^ in2[107];
    assign G[6] = in[106] & in2[106];
    assign P[6] = in[106] ^ in2[106];
    assign G[7] = in[105] & in2[105];
    assign P[7] = in[105] ^ in2[105];
    assign G[8] = in[104] & in2[104];
    assign P[8] = in[104] ^ in2[104];
    assign G[9] = in[103] & in2[103];
    assign P[9] = in[103] ^ in2[103];
    assign G[10] = in[102] & in2[102];
    assign P[10] = in[102] ^ in2[102];
    assign G[11] = in[101] & in2[101];
    assign P[11] = in[101] ^ in2[101];
    assign G[12] = in[100] & in2[100];
    assign P[12] = in[100] ^ in2[100];
    assign G[13] = in[99] & in2[99];
    assign P[13] = in[99] ^ in2[99];
    assign G[14] = in[98] & in2[98];
    assign P[14] = in[98] ^ in2[98];
    assign G[15] = in[97] & in2[97];
    assign P[15] = in[97] ^ in2[97];
    assign G[16] = in[96] & in2[96];
    assign P[16] = in[96] ^ in2[96];
    assign G[17] = in[95] & in2[95];
    assign P[17] = in[95] ^ in2[95];
    assign G[18] = in[94] & in2[94];
    assign P[18] = in[94] ^ in2[94];
    assign G[19] = in[93] & in2[93];
    assign P[19] = in[93] ^ in2[93];
    assign G[20] = in[92] & in2[92];
    assign P[20] = in[92] ^ in2[92];
    assign G[21] = in[91] & in2[91];
    assign P[21] = in[91] ^ in2[91];
    assign G[22] = in[90] & in2[90];
    assign P[22] = in[90] ^ in2[90];
    assign G[23] = in[89] & in2[89];
    assign P[23] = in[89] ^ in2[89];
    assign G[24] = in[88] & in2[88];
    assign P[24] = in[88] ^ in2[88];
    assign G[25] = in[87] & in2[87];
    assign P[25] = in[87] ^ in2[87];
    assign G[26] = in[86] & in2[86];
    assign P[26] = in[86] ^ in2[86];
    assign G[27] = in[85] & in2[85];
    assign P[27] = in[85] ^ in2[85];
    assign G[28] = in[84] & in2[84];
    assign P[28] = in[84] ^ in2[84];
    assign G[29] = in[83] & in2[83];
    assign P[29] = in[83] ^ in2[83];
    assign G[30] = in[82] & in2[82];
    assign P[30] = in[82] ^ in2[82];
    assign G[31] = in[81] & in2[81];
    assign P[31] = in[81] ^ in2[81];
    assign G[32] = in[80] & in2[80];
    assign P[32] = in[80] ^ in2[80];
    assign G[33] = in[79] & in2[79];
    assign P[33] = in[79] ^ in2[79];
    assign G[34] = in[78] & in2[78];
    assign P[34] = in[78] ^ in2[78];
    assign G[35] = in[77] & in2[77];
    assign P[35] = in[77] ^ in2[77];
    assign G[36] = in[76] & in2[76];
    assign P[36] = in[76] ^ in2[76];
    assign G[37] = in[75] & in2[75];
    assign P[37] = in[75] ^ in2[75];
    assign G[38] = in[74] & in2[74];
    assign P[38] = in[74] ^ in2[74];
    assign G[39] = in[73] & in2[73];
    assign P[39] = in[73] ^ in2[73];
    assign G[40] = in[72] & in2[72];
    assign P[40] = in[72] ^ in2[72];
    assign G[41] = in[71] & in2[71];
    assign P[41] = in[71] ^ in2[71];
    assign G[42] = in[70] & in2[70];
    assign P[42] = in[70] ^ in2[70];
    assign G[43] = in[69] & in2[69];
    assign P[43] = in[69] ^ in2[69];
    assign G[44] = in[68] & in2[68];
    assign P[44] = in[68] ^ in2[68];
    assign G[45] = in[67] & in2[67];
    assign P[45] = in[67] ^ in2[67];
    assign G[46] = in[66] & in2[66];
    assign P[46] = in[66] ^ in2[66];
    assign G[47] = in[65] & in2[65];
    assign P[47] = in[65] ^ in2[65];
    assign G[48] = in[64] & in2[64];
    assign P[48] = in[64] ^ in2[64];
    assign G[49] = in[63] & in2[63];
    assign P[49] = in[63] ^ in2[63];
    assign G[50] = in[62] & in2[62];
    assign P[50] = in[62] ^ in2[62];
    assign G[51] = in[61] & in2[61];
    assign P[51] = in[61] ^ in2[61];
    assign G[52] = in[60] & in2[60];
    assign P[52] = in[60] ^ in2[60];
    assign G[53] = in[59] & in2[59];
    assign P[53] = in[59] ^ in2[59];
    assign G[54] = in[58] & in2[58];
    assign P[54] = in[58] ^ in2[58];
    assign G[55] = in[57] & in2[57];
    assign P[55] = in[57] ^ in2[57];
    assign G[56] = in[56] & in2[56];
    assign P[56] = in[56] ^ in2[56];
    assign G[57] = in[55] & in2[55];
    assign P[57] = in[55] ^ in2[55];
    assign G[58] = in[54] & in2[54];
    assign P[58] = in[54] ^ in2[54];
    assign G[59] = in[53] & in2[53];
    assign P[59] = in[53] ^ in2[53];
    assign G[60] = in[52] & in2[52];
    assign P[60] = in[52] ^ in2[52];
    assign G[61] = in[51] & in2[51];
    assign P[61] = in[51] ^ in2[51];
    assign G[62] = in[50] & in2[50];
    assign P[62] = in[50] ^ in2[50];
    assign G[63] = in[49] & in2[49];
    assign P[63] = in[49] ^ in2[49];
    assign G[64] = in[48] & in2[48];
    assign P[64] = in[48] ^ in2[48];
    assign G[65] = in[47] & in2[47];
    assign P[65] = in[47] ^ in2[47];
    assign G[66] = in[46] & in2[46];
    assign P[66] = in[46] ^ in2[46];
    assign G[67] = in[45] & in2[45];
    assign P[67] = in[45] ^ in2[45];
    assign G[68] = in[44] & in2[44];
    assign P[68] = in[44] ^ in2[44];
    assign G[69] = in[43] & in2[43];
    assign P[69] = in[43] ^ in2[43];
    assign G[70] = in[42] & in2[42];
    assign P[70] = in[42] ^ in2[42];
    assign G[71] = in[41] & in2[41];
    assign P[71] = in[41] ^ in2[41];
    assign G[72] = in[40] & in2[40];
    assign P[72] = in[40] ^ in2[40];
    assign G[73] = in[39] & in2[39];
    assign P[73] = in[39] ^ in2[39];
    assign G[74] = in[38] & in2[38];
    assign P[74] = in[38] ^ in2[38];
    assign G[75] = in[37] & in2[37];
    assign P[75] = in[37] ^ in2[37];
    assign G[76] = in[36] & in2[36];
    assign P[76] = in[36] ^ in2[36];
    assign G[77] = in[35] & in2[35];
    assign P[77] = in[35] ^ in2[35];
    assign G[78] = in[34] & in2[34];
    assign P[78] = in[34] ^ in2[34];
    assign G[79] = in[33] & in2[33];
    assign P[79] = in[33] ^ in2[33];
    assign G[80] = in[32] & in2[32];
    assign P[80] = in[32] ^ in2[32];
    assign G[81] = in[31] & in2[31];
    assign P[81] = in[31] ^ in2[31];
    assign G[82] = in[30] & in2[30];
    assign P[82] = in[30] ^ in2[30];
    assign G[83] = in[29] & in2[29];
    assign P[83] = in[29] ^ in2[29];
    assign G[84] = in[28] & in2[28];
    assign P[84] = in[28] ^ in2[28];
    assign G[85] = in[27] & in2[27];
    assign P[85] = in[27] ^ in2[27];
    assign G[86] = in[26] & in2[26];
    assign P[86] = in[26] ^ in2[26];
    assign G[87] = in[25] & in2[25];
    assign P[87] = in[25] ^ in2[25];
    assign G[88] = in[24] & in2[24];
    assign P[88] = in[24] ^ in2[24];
    assign G[89] = in[23] & in2[23];
    assign P[89] = in[23] ^ in2[23];
    assign G[90] = in[22] & in2[22];
    assign P[90] = in[22] ^ in2[22];
    assign G[91] = in[21] & in2[21];
    assign P[91] = in[21] ^ in2[21];
    assign G[92] = in[20] & in2[20];
    assign P[92] = in[20] ^ in2[20];
    assign G[93] = in[19] & in2[19];
    assign P[93] = in[19] ^ in2[19];
    assign G[94] = in[18] & in2[18];
    assign P[94] = in[18] ^ in2[18];
    assign G[95] = in[17] & in2[17];
    assign P[95] = in[17] ^ in2[17];
    assign G[96] = in[16] & in2[16];
    assign P[96] = in[16] ^ in2[16];
    assign G[97] = in[15] & in2[15];
    assign P[97] = in[15] ^ in2[15];
    assign G[98] = in[14] & in2[14];
    assign P[98] = in[14] ^ in2[14];
    assign G[99] = in[13] & in2[13];
    assign P[99] = in[13] ^ in2[13];
    assign G[100] = in[12] & in2[12];
    assign P[100] = in[12] ^ in2[12];
    assign G[101] = in[11] & in2[11];
    assign P[101] = in[11] ^ in2[11];
    assign G[102] = in[10] & in2[10];
    assign P[102] = in[10] ^ in2[10];
    assign G[103] = in[9] & in2[9];
    assign P[103] = in[9] ^ in2[9];
    assign G[104] = in[8] & in2[8];
    assign P[104] = in[8] ^ in2[8];
    assign G[105] = in[7] & in2[7];
    assign P[105] = in[7] ^ in2[7];
    assign G[106] = in[6] & in2[6];
    assign P[106] = in[6] ^ in2[6];
    assign G[107] = in[5] & in2[5];
    assign P[107] = in[5] ^ in2[5];
    assign G[108] = in[4] & in2[4];
    assign P[108] = in[4] ^ in2[4];
    assign G[109] = in[3] & in2[3];
    assign P[109] = in[3] ^ in2[3];
    assign G[110] = in[2] & in2[2];
    assign P[110] = in[2] ^ in2[2];
    assign G[111] = in[1] & in2[1];
    assign P[111] = in[1] ^ in2[1];
    assign G[112] = in[0] & in2[0];
    assign P[112] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign C[112] = G[111] | (P[111] & C[111]);
    assign cout = G[112] | (P[112] & C[112]);
    assign sum = P ^ C;
endmodule

module CLA112(output [111:0] sum, output cout, input [111:0] in1, input [111:0] in2;

    wire[111:0] G;
    wire[111:0] C;
    wire[111:0] P;

    assign G[0] = in[111] & in2[111];
    assign P[0] = in[111] ^ in2[111];
    assign G[1] = in[110] & in2[110];
    assign P[1] = in[110] ^ in2[110];
    assign G[2] = in[109] & in2[109];
    assign P[2] = in[109] ^ in2[109];
    assign G[3] = in[108] & in2[108];
    assign P[3] = in[108] ^ in2[108];
    assign G[4] = in[107] & in2[107];
    assign P[4] = in[107] ^ in2[107];
    assign G[5] = in[106] & in2[106];
    assign P[5] = in[106] ^ in2[106];
    assign G[6] = in[105] & in2[105];
    assign P[6] = in[105] ^ in2[105];
    assign G[7] = in[104] & in2[104];
    assign P[7] = in[104] ^ in2[104];
    assign G[8] = in[103] & in2[103];
    assign P[8] = in[103] ^ in2[103];
    assign G[9] = in[102] & in2[102];
    assign P[9] = in[102] ^ in2[102];
    assign G[10] = in[101] & in2[101];
    assign P[10] = in[101] ^ in2[101];
    assign G[11] = in[100] & in2[100];
    assign P[11] = in[100] ^ in2[100];
    assign G[12] = in[99] & in2[99];
    assign P[12] = in[99] ^ in2[99];
    assign G[13] = in[98] & in2[98];
    assign P[13] = in[98] ^ in2[98];
    assign G[14] = in[97] & in2[97];
    assign P[14] = in[97] ^ in2[97];
    assign G[15] = in[96] & in2[96];
    assign P[15] = in[96] ^ in2[96];
    assign G[16] = in[95] & in2[95];
    assign P[16] = in[95] ^ in2[95];
    assign G[17] = in[94] & in2[94];
    assign P[17] = in[94] ^ in2[94];
    assign G[18] = in[93] & in2[93];
    assign P[18] = in[93] ^ in2[93];
    assign G[19] = in[92] & in2[92];
    assign P[19] = in[92] ^ in2[92];
    assign G[20] = in[91] & in2[91];
    assign P[20] = in[91] ^ in2[91];
    assign G[21] = in[90] & in2[90];
    assign P[21] = in[90] ^ in2[90];
    assign G[22] = in[89] & in2[89];
    assign P[22] = in[89] ^ in2[89];
    assign G[23] = in[88] & in2[88];
    assign P[23] = in[88] ^ in2[88];
    assign G[24] = in[87] & in2[87];
    assign P[24] = in[87] ^ in2[87];
    assign G[25] = in[86] & in2[86];
    assign P[25] = in[86] ^ in2[86];
    assign G[26] = in[85] & in2[85];
    assign P[26] = in[85] ^ in2[85];
    assign G[27] = in[84] & in2[84];
    assign P[27] = in[84] ^ in2[84];
    assign G[28] = in[83] & in2[83];
    assign P[28] = in[83] ^ in2[83];
    assign G[29] = in[82] & in2[82];
    assign P[29] = in[82] ^ in2[82];
    assign G[30] = in[81] & in2[81];
    assign P[30] = in[81] ^ in2[81];
    assign G[31] = in[80] & in2[80];
    assign P[31] = in[80] ^ in2[80];
    assign G[32] = in[79] & in2[79];
    assign P[32] = in[79] ^ in2[79];
    assign G[33] = in[78] & in2[78];
    assign P[33] = in[78] ^ in2[78];
    assign G[34] = in[77] & in2[77];
    assign P[34] = in[77] ^ in2[77];
    assign G[35] = in[76] & in2[76];
    assign P[35] = in[76] ^ in2[76];
    assign G[36] = in[75] & in2[75];
    assign P[36] = in[75] ^ in2[75];
    assign G[37] = in[74] & in2[74];
    assign P[37] = in[74] ^ in2[74];
    assign G[38] = in[73] & in2[73];
    assign P[38] = in[73] ^ in2[73];
    assign G[39] = in[72] & in2[72];
    assign P[39] = in[72] ^ in2[72];
    assign G[40] = in[71] & in2[71];
    assign P[40] = in[71] ^ in2[71];
    assign G[41] = in[70] & in2[70];
    assign P[41] = in[70] ^ in2[70];
    assign G[42] = in[69] & in2[69];
    assign P[42] = in[69] ^ in2[69];
    assign G[43] = in[68] & in2[68];
    assign P[43] = in[68] ^ in2[68];
    assign G[44] = in[67] & in2[67];
    assign P[44] = in[67] ^ in2[67];
    assign G[45] = in[66] & in2[66];
    assign P[45] = in[66] ^ in2[66];
    assign G[46] = in[65] & in2[65];
    assign P[46] = in[65] ^ in2[65];
    assign G[47] = in[64] & in2[64];
    assign P[47] = in[64] ^ in2[64];
    assign G[48] = in[63] & in2[63];
    assign P[48] = in[63] ^ in2[63];
    assign G[49] = in[62] & in2[62];
    assign P[49] = in[62] ^ in2[62];
    assign G[50] = in[61] & in2[61];
    assign P[50] = in[61] ^ in2[61];
    assign G[51] = in[60] & in2[60];
    assign P[51] = in[60] ^ in2[60];
    assign G[52] = in[59] & in2[59];
    assign P[52] = in[59] ^ in2[59];
    assign G[53] = in[58] & in2[58];
    assign P[53] = in[58] ^ in2[58];
    assign G[54] = in[57] & in2[57];
    assign P[54] = in[57] ^ in2[57];
    assign G[55] = in[56] & in2[56];
    assign P[55] = in[56] ^ in2[56];
    assign G[56] = in[55] & in2[55];
    assign P[56] = in[55] ^ in2[55];
    assign G[57] = in[54] & in2[54];
    assign P[57] = in[54] ^ in2[54];
    assign G[58] = in[53] & in2[53];
    assign P[58] = in[53] ^ in2[53];
    assign G[59] = in[52] & in2[52];
    assign P[59] = in[52] ^ in2[52];
    assign G[60] = in[51] & in2[51];
    assign P[60] = in[51] ^ in2[51];
    assign G[61] = in[50] & in2[50];
    assign P[61] = in[50] ^ in2[50];
    assign G[62] = in[49] & in2[49];
    assign P[62] = in[49] ^ in2[49];
    assign G[63] = in[48] & in2[48];
    assign P[63] = in[48] ^ in2[48];
    assign G[64] = in[47] & in2[47];
    assign P[64] = in[47] ^ in2[47];
    assign G[65] = in[46] & in2[46];
    assign P[65] = in[46] ^ in2[46];
    assign G[66] = in[45] & in2[45];
    assign P[66] = in[45] ^ in2[45];
    assign G[67] = in[44] & in2[44];
    assign P[67] = in[44] ^ in2[44];
    assign G[68] = in[43] & in2[43];
    assign P[68] = in[43] ^ in2[43];
    assign G[69] = in[42] & in2[42];
    assign P[69] = in[42] ^ in2[42];
    assign G[70] = in[41] & in2[41];
    assign P[70] = in[41] ^ in2[41];
    assign G[71] = in[40] & in2[40];
    assign P[71] = in[40] ^ in2[40];
    assign G[72] = in[39] & in2[39];
    assign P[72] = in[39] ^ in2[39];
    assign G[73] = in[38] & in2[38];
    assign P[73] = in[38] ^ in2[38];
    assign G[74] = in[37] & in2[37];
    assign P[74] = in[37] ^ in2[37];
    assign G[75] = in[36] & in2[36];
    assign P[75] = in[36] ^ in2[36];
    assign G[76] = in[35] & in2[35];
    assign P[76] = in[35] ^ in2[35];
    assign G[77] = in[34] & in2[34];
    assign P[77] = in[34] ^ in2[34];
    assign G[78] = in[33] & in2[33];
    assign P[78] = in[33] ^ in2[33];
    assign G[79] = in[32] & in2[32];
    assign P[79] = in[32] ^ in2[32];
    assign G[80] = in[31] & in2[31];
    assign P[80] = in[31] ^ in2[31];
    assign G[81] = in[30] & in2[30];
    assign P[81] = in[30] ^ in2[30];
    assign G[82] = in[29] & in2[29];
    assign P[82] = in[29] ^ in2[29];
    assign G[83] = in[28] & in2[28];
    assign P[83] = in[28] ^ in2[28];
    assign G[84] = in[27] & in2[27];
    assign P[84] = in[27] ^ in2[27];
    assign G[85] = in[26] & in2[26];
    assign P[85] = in[26] ^ in2[26];
    assign G[86] = in[25] & in2[25];
    assign P[86] = in[25] ^ in2[25];
    assign G[87] = in[24] & in2[24];
    assign P[87] = in[24] ^ in2[24];
    assign G[88] = in[23] & in2[23];
    assign P[88] = in[23] ^ in2[23];
    assign G[89] = in[22] & in2[22];
    assign P[89] = in[22] ^ in2[22];
    assign G[90] = in[21] & in2[21];
    assign P[90] = in[21] ^ in2[21];
    assign G[91] = in[20] & in2[20];
    assign P[91] = in[20] ^ in2[20];
    assign G[92] = in[19] & in2[19];
    assign P[92] = in[19] ^ in2[19];
    assign G[93] = in[18] & in2[18];
    assign P[93] = in[18] ^ in2[18];
    assign G[94] = in[17] & in2[17];
    assign P[94] = in[17] ^ in2[17];
    assign G[95] = in[16] & in2[16];
    assign P[95] = in[16] ^ in2[16];
    assign G[96] = in[15] & in2[15];
    assign P[96] = in[15] ^ in2[15];
    assign G[97] = in[14] & in2[14];
    assign P[97] = in[14] ^ in2[14];
    assign G[98] = in[13] & in2[13];
    assign P[98] = in[13] ^ in2[13];
    assign G[99] = in[12] & in2[12];
    assign P[99] = in[12] ^ in2[12];
    assign G[100] = in[11] & in2[11];
    assign P[100] = in[11] ^ in2[11];
    assign G[101] = in[10] & in2[10];
    assign P[101] = in[10] ^ in2[10];
    assign G[102] = in[9] & in2[9];
    assign P[102] = in[9] ^ in2[9];
    assign G[103] = in[8] & in2[8];
    assign P[103] = in[8] ^ in2[8];
    assign G[104] = in[7] & in2[7];
    assign P[104] = in[7] ^ in2[7];
    assign G[105] = in[6] & in2[6];
    assign P[105] = in[6] ^ in2[6];
    assign G[106] = in[5] & in2[5];
    assign P[106] = in[5] ^ in2[5];
    assign G[107] = in[4] & in2[4];
    assign P[107] = in[4] ^ in2[4];
    assign G[108] = in[3] & in2[3];
    assign P[108] = in[3] ^ in2[3];
    assign G[109] = in[2] & in2[2];
    assign P[109] = in[2] ^ in2[2];
    assign G[110] = in[1] & in2[1];
    assign P[110] = in[1] ^ in2[1];
    assign G[111] = in[0] & in2[0];
    assign P[111] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign C[111] = G[110] | (P[110] & C[110]);
    assign cout = G[111] | (P[111] & C[111]);
    assign sum = P ^ C;
endmodule

module CLA111(output [110:0] sum, output cout, input [110:0] in1, input [110:0] in2;

    wire[110:0] G;
    wire[110:0] C;
    wire[110:0] P;

    assign G[0] = in[110] & in2[110];
    assign P[0] = in[110] ^ in2[110];
    assign G[1] = in[109] & in2[109];
    assign P[1] = in[109] ^ in2[109];
    assign G[2] = in[108] & in2[108];
    assign P[2] = in[108] ^ in2[108];
    assign G[3] = in[107] & in2[107];
    assign P[3] = in[107] ^ in2[107];
    assign G[4] = in[106] & in2[106];
    assign P[4] = in[106] ^ in2[106];
    assign G[5] = in[105] & in2[105];
    assign P[5] = in[105] ^ in2[105];
    assign G[6] = in[104] & in2[104];
    assign P[6] = in[104] ^ in2[104];
    assign G[7] = in[103] & in2[103];
    assign P[7] = in[103] ^ in2[103];
    assign G[8] = in[102] & in2[102];
    assign P[8] = in[102] ^ in2[102];
    assign G[9] = in[101] & in2[101];
    assign P[9] = in[101] ^ in2[101];
    assign G[10] = in[100] & in2[100];
    assign P[10] = in[100] ^ in2[100];
    assign G[11] = in[99] & in2[99];
    assign P[11] = in[99] ^ in2[99];
    assign G[12] = in[98] & in2[98];
    assign P[12] = in[98] ^ in2[98];
    assign G[13] = in[97] & in2[97];
    assign P[13] = in[97] ^ in2[97];
    assign G[14] = in[96] & in2[96];
    assign P[14] = in[96] ^ in2[96];
    assign G[15] = in[95] & in2[95];
    assign P[15] = in[95] ^ in2[95];
    assign G[16] = in[94] & in2[94];
    assign P[16] = in[94] ^ in2[94];
    assign G[17] = in[93] & in2[93];
    assign P[17] = in[93] ^ in2[93];
    assign G[18] = in[92] & in2[92];
    assign P[18] = in[92] ^ in2[92];
    assign G[19] = in[91] & in2[91];
    assign P[19] = in[91] ^ in2[91];
    assign G[20] = in[90] & in2[90];
    assign P[20] = in[90] ^ in2[90];
    assign G[21] = in[89] & in2[89];
    assign P[21] = in[89] ^ in2[89];
    assign G[22] = in[88] & in2[88];
    assign P[22] = in[88] ^ in2[88];
    assign G[23] = in[87] & in2[87];
    assign P[23] = in[87] ^ in2[87];
    assign G[24] = in[86] & in2[86];
    assign P[24] = in[86] ^ in2[86];
    assign G[25] = in[85] & in2[85];
    assign P[25] = in[85] ^ in2[85];
    assign G[26] = in[84] & in2[84];
    assign P[26] = in[84] ^ in2[84];
    assign G[27] = in[83] & in2[83];
    assign P[27] = in[83] ^ in2[83];
    assign G[28] = in[82] & in2[82];
    assign P[28] = in[82] ^ in2[82];
    assign G[29] = in[81] & in2[81];
    assign P[29] = in[81] ^ in2[81];
    assign G[30] = in[80] & in2[80];
    assign P[30] = in[80] ^ in2[80];
    assign G[31] = in[79] & in2[79];
    assign P[31] = in[79] ^ in2[79];
    assign G[32] = in[78] & in2[78];
    assign P[32] = in[78] ^ in2[78];
    assign G[33] = in[77] & in2[77];
    assign P[33] = in[77] ^ in2[77];
    assign G[34] = in[76] & in2[76];
    assign P[34] = in[76] ^ in2[76];
    assign G[35] = in[75] & in2[75];
    assign P[35] = in[75] ^ in2[75];
    assign G[36] = in[74] & in2[74];
    assign P[36] = in[74] ^ in2[74];
    assign G[37] = in[73] & in2[73];
    assign P[37] = in[73] ^ in2[73];
    assign G[38] = in[72] & in2[72];
    assign P[38] = in[72] ^ in2[72];
    assign G[39] = in[71] & in2[71];
    assign P[39] = in[71] ^ in2[71];
    assign G[40] = in[70] & in2[70];
    assign P[40] = in[70] ^ in2[70];
    assign G[41] = in[69] & in2[69];
    assign P[41] = in[69] ^ in2[69];
    assign G[42] = in[68] & in2[68];
    assign P[42] = in[68] ^ in2[68];
    assign G[43] = in[67] & in2[67];
    assign P[43] = in[67] ^ in2[67];
    assign G[44] = in[66] & in2[66];
    assign P[44] = in[66] ^ in2[66];
    assign G[45] = in[65] & in2[65];
    assign P[45] = in[65] ^ in2[65];
    assign G[46] = in[64] & in2[64];
    assign P[46] = in[64] ^ in2[64];
    assign G[47] = in[63] & in2[63];
    assign P[47] = in[63] ^ in2[63];
    assign G[48] = in[62] & in2[62];
    assign P[48] = in[62] ^ in2[62];
    assign G[49] = in[61] & in2[61];
    assign P[49] = in[61] ^ in2[61];
    assign G[50] = in[60] & in2[60];
    assign P[50] = in[60] ^ in2[60];
    assign G[51] = in[59] & in2[59];
    assign P[51] = in[59] ^ in2[59];
    assign G[52] = in[58] & in2[58];
    assign P[52] = in[58] ^ in2[58];
    assign G[53] = in[57] & in2[57];
    assign P[53] = in[57] ^ in2[57];
    assign G[54] = in[56] & in2[56];
    assign P[54] = in[56] ^ in2[56];
    assign G[55] = in[55] & in2[55];
    assign P[55] = in[55] ^ in2[55];
    assign G[56] = in[54] & in2[54];
    assign P[56] = in[54] ^ in2[54];
    assign G[57] = in[53] & in2[53];
    assign P[57] = in[53] ^ in2[53];
    assign G[58] = in[52] & in2[52];
    assign P[58] = in[52] ^ in2[52];
    assign G[59] = in[51] & in2[51];
    assign P[59] = in[51] ^ in2[51];
    assign G[60] = in[50] & in2[50];
    assign P[60] = in[50] ^ in2[50];
    assign G[61] = in[49] & in2[49];
    assign P[61] = in[49] ^ in2[49];
    assign G[62] = in[48] & in2[48];
    assign P[62] = in[48] ^ in2[48];
    assign G[63] = in[47] & in2[47];
    assign P[63] = in[47] ^ in2[47];
    assign G[64] = in[46] & in2[46];
    assign P[64] = in[46] ^ in2[46];
    assign G[65] = in[45] & in2[45];
    assign P[65] = in[45] ^ in2[45];
    assign G[66] = in[44] & in2[44];
    assign P[66] = in[44] ^ in2[44];
    assign G[67] = in[43] & in2[43];
    assign P[67] = in[43] ^ in2[43];
    assign G[68] = in[42] & in2[42];
    assign P[68] = in[42] ^ in2[42];
    assign G[69] = in[41] & in2[41];
    assign P[69] = in[41] ^ in2[41];
    assign G[70] = in[40] & in2[40];
    assign P[70] = in[40] ^ in2[40];
    assign G[71] = in[39] & in2[39];
    assign P[71] = in[39] ^ in2[39];
    assign G[72] = in[38] & in2[38];
    assign P[72] = in[38] ^ in2[38];
    assign G[73] = in[37] & in2[37];
    assign P[73] = in[37] ^ in2[37];
    assign G[74] = in[36] & in2[36];
    assign P[74] = in[36] ^ in2[36];
    assign G[75] = in[35] & in2[35];
    assign P[75] = in[35] ^ in2[35];
    assign G[76] = in[34] & in2[34];
    assign P[76] = in[34] ^ in2[34];
    assign G[77] = in[33] & in2[33];
    assign P[77] = in[33] ^ in2[33];
    assign G[78] = in[32] & in2[32];
    assign P[78] = in[32] ^ in2[32];
    assign G[79] = in[31] & in2[31];
    assign P[79] = in[31] ^ in2[31];
    assign G[80] = in[30] & in2[30];
    assign P[80] = in[30] ^ in2[30];
    assign G[81] = in[29] & in2[29];
    assign P[81] = in[29] ^ in2[29];
    assign G[82] = in[28] & in2[28];
    assign P[82] = in[28] ^ in2[28];
    assign G[83] = in[27] & in2[27];
    assign P[83] = in[27] ^ in2[27];
    assign G[84] = in[26] & in2[26];
    assign P[84] = in[26] ^ in2[26];
    assign G[85] = in[25] & in2[25];
    assign P[85] = in[25] ^ in2[25];
    assign G[86] = in[24] & in2[24];
    assign P[86] = in[24] ^ in2[24];
    assign G[87] = in[23] & in2[23];
    assign P[87] = in[23] ^ in2[23];
    assign G[88] = in[22] & in2[22];
    assign P[88] = in[22] ^ in2[22];
    assign G[89] = in[21] & in2[21];
    assign P[89] = in[21] ^ in2[21];
    assign G[90] = in[20] & in2[20];
    assign P[90] = in[20] ^ in2[20];
    assign G[91] = in[19] & in2[19];
    assign P[91] = in[19] ^ in2[19];
    assign G[92] = in[18] & in2[18];
    assign P[92] = in[18] ^ in2[18];
    assign G[93] = in[17] & in2[17];
    assign P[93] = in[17] ^ in2[17];
    assign G[94] = in[16] & in2[16];
    assign P[94] = in[16] ^ in2[16];
    assign G[95] = in[15] & in2[15];
    assign P[95] = in[15] ^ in2[15];
    assign G[96] = in[14] & in2[14];
    assign P[96] = in[14] ^ in2[14];
    assign G[97] = in[13] & in2[13];
    assign P[97] = in[13] ^ in2[13];
    assign G[98] = in[12] & in2[12];
    assign P[98] = in[12] ^ in2[12];
    assign G[99] = in[11] & in2[11];
    assign P[99] = in[11] ^ in2[11];
    assign G[100] = in[10] & in2[10];
    assign P[100] = in[10] ^ in2[10];
    assign G[101] = in[9] & in2[9];
    assign P[101] = in[9] ^ in2[9];
    assign G[102] = in[8] & in2[8];
    assign P[102] = in[8] ^ in2[8];
    assign G[103] = in[7] & in2[7];
    assign P[103] = in[7] ^ in2[7];
    assign G[104] = in[6] & in2[6];
    assign P[104] = in[6] ^ in2[6];
    assign G[105] = in[5] & in2[5];
    assign P[105] = in[5] ^ in2[5];
    assign G[106] = in[4] & in2[4];
    assign P[106] = in[4] ^ in2[4];
    assign G[107] = in[3] & in2[3];
    assign P[107] = in[3] ^ in2[3];
    assign G[108] = in[2] & in2[2];
    assign P[108] = in[2] ^ in2[2];
    assign G[109] = in[1] & in2[1];
    assign P[109] = in[1] ^ in2[1];
    assign G[110] = in[0] & in2[0];
    assign P[110] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign C[110] = G[109] | (P[109] & C[109]);
    assign cout = G[110] | (P[110] & C[110]);
    assign sum = P ^ C;
endmodule

module CLA110(output [109:0] sum, output cout, input [109:0] in1, input [109:0] in2;

    wire[109:0] G;
    wire[109:0] C;
    wire[109:0] P;

    assign G[0] = in[109] & in2[109];
    assign P[0] = in[109] ^ in2[109];
    assign G[1] = in[108] & in2[108];
    assign P[1] = in[108] ^ in2[108];
    assign G[2] = in[107] & in2[107];
    assign P[2] = in[107] ^ in2[107];
    assign G[3] = in[106] & in2[106];
    assign P[3] = in[106] ^ in2[106];
    assign G[4] = in[105] & in2[105];
    assign P[4] = in[105] ^ in2[105];
    assign G[5] = in[104] & in2[104];
    assign P[5] = in[104] ^ in2[104];
    assign G[6] = in[103] & in2[103];
    assign P[6] = in[103] ^ in2[103];
    assign G[7] = in[102] & in2[102];
    assign P[7] = in[102] ^ in2[102];
    assign G[8] = in[101] & in2[101];
    assign P[8] = in[101] ^ in2[101];
    assign G[9] = in[100] & in2[100];
    assign P[9] = in[100] ^ in2[100];
    assign G[10] = in[99] & in2[99];
    assign P[10] = in[99] ^ in2[99];
    assign G[11] = in[98] & in2[98];
    assign P[11] = in[98] ^ in2[98];
    assign G[12] = in[97] & in2[97];
    assign P[12] = in[97] ^ in2[97];
    assign G[13] = in[96] & in2[96];
    assign P[13] = in[96] ^ in2[96];
    assign G[14] = in[95] & in2[95];
    assign P[14] = in[95] ^ in2[95];
    assign G[15] = in[94] & in2[94];
    assign P[15] = in[94] ^ in2[94];
    assign G[16] = in[93] & in2[93];
    assign P[16] = in[93] ^ in2[93];
    assign G[17] = in[92] & in2[92];
    assign P[17] = in[92] ^ in2[92];
    assign G[18] = in[91] & in2[91];
    assign P[18] = in[91] ^ in2[91];
    assign G[19] = in[90] & in2[90];
    assign P[19] = in[90] ^ in2[90];
    assign G[20] = in[89] & in2[89];
    assign P[20] = in[89] ^ in2[89];
    assign G[21] = in[88] & in2[88];
    assign P[21] = in[88] ^ in2[88];
    assign G[22] = in[87] & in2[87];
    assign P[22] = in[87] ^ in2[87];
    assign G[23] = in[86] & in2[86];
    assign P[23] = in[86] ^ in2[86];
    assign G[24] = in[85] & in2[85];
    assign P[24] = in[85] ^ in2[85];
    assign G[25] = in[84] & in2[84];
    assign P[25] = in[84] ^ in2[84];
    assign G[26] = in[83] & in2[83];
    assign P[26] = in[83] ^ in2[83];
    assign G[27] = in[82] & in2[82];
    assign P[27] = in[82] ^ in2[82];
    assign G[28] = in[81] & in2[81];
    assign P[28] = in[81] ^ in2[81];
    assign G[29] = in[80] & in2[80];
    assign P[29] = in[80] ^ in2[80];
    assign G[30] = in[79] & in2[79];
    assign P[30] = in[79] ^ in2[79];
    assign G[31] = in[78] & in2[78];
    assign P[31] = in[78] ^ in2[78];
    assign G[32] = in[77] & in2[77];
    assign P[32] = in[77] ^ in2[77];
    assign G[33] = in[76] & in2[76];
    assign P[33] = in[76] ^ in2[76];
    assign G[34] = in[75] & in2[75];
    assign P[34] = in[75] ^ in2[75];
    assign G[35] = in[74] & in2[74];
    assign P[35] = in[74] ^ in2[74];
    assign G[36] = in[73] & in2[73];
    assign P[36] = in[73] ^ in2[73];
    assign G[37] = in[72] & in2[72];
    assign P[37] = in[72] ^ in2[72];
    assign G[38] = in[71] & in2[71];
    assign P[38] = in[71] ^ in2[71];
    assign G[39] = in[70] & in2[70];
    assign P[39] = in[70] ^ in2[70];
    assign G[40] = in[69] & in2[69];
    assign P[40] = in[69] ^ in2[69];
    assign G[41] = in[68] & in2[68];
    assign P[41] = in[68] ^ in2[68];
    assign G[42] = in[67] & in2[67];
    assign P[42] = in[67] ^ in2[67];
    assign G[43] = in[66] & in2[66];
    assign P[43] = in[66] ^ in2[66];
    assign G[44] = in[65] & in2[65];
    assign P[44] = in[65] ^ in2[65];
    assign G[45] = in[64] & in2[64];
    assign P[45] = in[64] ^ in2[64];
    assign G[46] = in[63] & in2[63];
    assign P[46] = in[63] ^ in2[63];
    assign G[47] = in[62] & in2[62];
    assign P[47] = in[62] ^ in2[62];
    assign G[48] = in[61] & in2[61];
    assign P[48] = in[61] ^ in2[61];
    assign G[49] = in[60] & in2[60];
    assign P[49] = in[60] ^ in2[60];
    assign G[50] = in[59] & in2[59];
    assign P[50] = in[59] ^ in2[59];
    assign G[51] = in[58] & in2[58];
    assign P[51] = in[58] ^ in2[58];
    assign G[52] = in[57] & in2[57];
    assign P[52] = in[57] ^ in2[57];
    assign G[53] = in[56] & in2[56];
    assign P[53] = in[56] ^ in2[56];
    assign G[54] = in[55] & in2[55];
    assign P[54] = in[55] ^ in2[55];
    assign G[55] = in[54] & in2[54];
    assign P[55] = in[54] ^ in2[54];
    assign G[56] = in[53] & in2[53];
    assign P[56] = in[53] ^ in2[53];
    assign G[57] = in[52] & in2[52];
    assign P[57] = in[52] ^ in2[52];
    assign G[58] = in[51] & in2[51];
    assign P[58] = in[51] ^ in2[51];
    assign G[59] = in[50] & in2[50];
    assign P[59] = in[50] ^ in2[50];
    assign G[60] = in[49] & in2[49];
    assign P[60] = in[49] ^ in2[49];
    assign G[61] = in[48] & in2[48];
    assign P[61] = in[48] ^ in2[48];
    assign G[62] = in[47] & in2[47];
    assign P[62] = in[47] ^ in2[47];
    assign G[63] = in[46] & in2[46];
    assign P[63] = in[46] ^ in2[46];
    assign G[64] = in[45] & in2[45];
    assign P[64] = in[45] ^ in2[45];
    assign G[65] = in[44] & in2[44];
    assign P[65] = in[44] ^ in2[44];
    assign G[66] = in[43] & in2[43];
    assign P[66] = in[43] ^ in2[43];
    assign G[67] = in[42] & in2[42];
    assign P[67] = in[42] ^ in2[42];
    assign G[68] = in[41] & in2[41];
    assign P[68] = in[41] ^ in2[41];
    assign G[69] = in[40] & in2[40];
    assign P[69] = in[40] ^ in2[40];
    assign G[70] = in[39] & in2[39];
    assign P[70] = in[39] ^ in2[39];
    assign G[71] = in[38] & in2[38];
    assign P[71] = in[38] ^ in2[38];
    assign G[72] = in[37] & in2[37];
    assign P[72] = in[37] ^ in2[37];
    assign G[73] = in[36] & in2[36];
    assign P[73] = in[36] ^ in2[36];
    assign G[74] = in[35] & in2[35];
    assign P[74] = in[35] ^ in2[35];
    assign G[75] = in[34] & in2[34];
    assign P[75] = in[34] ^ in2[34];
    assign G[76] = in[33] & in2[33];
    assign P[76] = in[33] ^ in2[33];
    assign G[77] = in[32] & in2[32];
    assign P[77] = in[32] ^ in2[32];
    assign G[78] = in[31] & in2[31];
    assign P[78] = in[31] ^ in2[31];
    assign G[79] = in[30] & in2[30];
    assign P[79] = in[30] ^ in2[30];
    assign G[80] = in[29] & in2[29];
    assign P[80] = in[29] ^ in2[29];
    assign G[81] = in[28] & in2[28];
    assign P[81] = in[28] ^ in2[28];
    assign G[82] = in[27] & in2[27];
    assign P[82] = in[27] ^ in2[27];
    assign G[83] = in[26] & in2[26];
    assign P[83] = in[26] ^ in2[26];
    assign G[84] = in[25] & in2[25];
    assign P[84] = in[25] ^ in2[25];
    assign G[85] = in[24] & in2[24];
    assign P[85] = in[24] ^ in2[24];
    assign G[86] = in[23] & in2[23];
    assign P[86] = in[23] ^ in2[23];
    assign G[87] = in[22] & in2[22];
    assign P[87] = in[22] ^ in2[22];
    assign G[88] = in[21] & in2[21];
    assign P[88] = in[21] ^ in2[21];
    assign G[89] = in[20] & in2[20];
    assign P[89] = in[20] ^ in2[20];
    assign G[90] = in[19] & in2[19];
    assign P[90] = in[19] ^ in2[19];
    assign G[91] = in[18] & in2[18];
    assign P[91] = in[18] ^ in2[18];
    assign G[92] = in[17] & in2[17];
    assign P[92] = in[17] ^ in2[17];
    assign G[93] = in[16] & in2[16];
    assign P[93] = in[16] ^ in2[16];
    assign G[94] = in[15] & in2[15];
    assign P[94] = in[15] ^ in2[15];
    assign G[95] = in[14] & in2[14];
    assign P[95] = in[14] ^ in2[14];
    assign G[96] = in[13] & in2[13];
    assign P[96] = in[13] ^ in2[13];
    assign G[97] = in[12] & in2[12];
    assign P[97] = in[12] ^ in2[12];
    assign G[98] = in[11] & in2[11];
    assign P[98] = in[11] ^ in2[11];
    assign G[99] = in[10] & in2[10];
    assign P[99] = in[10] ^ in2[10];
    assign G[100] = in[9] & in2[9];
    assign P[100] = in[9] ^ in2[9];
    assign G[101] = in[8] & in2[8];
    assign P[101] = in[8] ^ in2[8];
    assign G[102] = in[7] & in2[7];
    assign P[102] = in[7] ^ in2[7];
    assign G[103] = in[6] & in2[6];
    assign P[103] = in[6] ^ in2[6];
    assign G[104] = in[5] & in2[5];
    assign P[104] = in[5] ^ in2[5];
    assign G[105] = in[4] & in2[4];
    assign P[105] = in[4] ^ in2[4];
    assign G[106] = in[3] & in2[3];
    assign P[106] = in[3] ^ in2[3];
    assign G[107] = in[2] & in2[2];
    assign P[107] = in[2] ^ in2[2];
    assign G[108] = in[1] & in2[1];
    assign P[108] = in[1] ^ in2[1];
    assign G[109] = in[0] & in2[0];
    assign P[109] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign C[109] = G[108] | (P[108] & C[108]);
    assign cout = G[109] | (P[109] & C[109]);
    assign sum = P ^ C;
endmodule

module CLA109(output [108:0] sum, output cout, input [108:0] in1, input [108:0] in2;

    wire[108:0] G;
    wire[108:0] C;
    wire[108:0] P;

    assign G[0] = in[108] & in2[108];
    assign P[0] = in[108] ^ in2[108];
    assign G[1] = in[107] & in2[107];
    assign P[1] = in[107] ^ in2[107];
    assign G[2] = in[106] & in2[106];
    assign P[2] = in[106] ^ in2[106];
    assign G[3] = in[105] & in2[105];
    assign P[3] = in[105] ^ in2[105];
    assign G[4] = in[104] & in2[104];
    assign P[4] = in[104] ^ in2[104];
    assign G[5] = in[103] & in2[103];
    assign P[5] = in[103] ^ in2[103];
    assign G[6] = in[102] & in2[102];
    assign P[6] = in[102] ^ in2[102];
    assign G[7] = in[101] & in2[101];
    assign P[7] = in[101] ^ in2[101];
    assign G[8] = in[100] & in2[100];
    assign P[8] = in[100] ^ in2[100];
    assign G[9] = in[99] & in2[99];
    assign P[9] = in[99] ^ in2[99];
    assign G[10] = in[98] & in2[98];
    assign P[10] = in[98] ^ in2[98];
    assign G[11] = in[97] & in2[97];
    assign P[11] = in[97] ^ in2[97];
    assign G[12] = in[96] & in2[96];
    assign P[12] = in[96] ^ in2[96];
    assign G[13] = in[95] & in2[95];
    assign P[13] = in[95] ^ in2[95];
    assign G[14] = in[94] & in2[94];
    assign P[14] = in[94] ^ in2[94];
    assign G[15] = in[93] & in2[93];
    assign P[15] = in[93] ^ in2[93];
    assign G[16] = in[92] & in2[92];
    assign P[16] = in[92] ^ in2[92];
    assign G[17] = in[91] & in2[91];
    assign P[17] = in[91] ^ in2[91];
    assign G[18] = in[90] & in2[90];
    assign P[18] = in[90] ^ in2[90];
    assign G[19] = in[89] & in2[89];
    assign P[19] = in[89] ^ in2[89];
    assign G[20] = in[88] & in2[88];
    assign P[20] = in[88] ^ in2[88];
    assign G[21] = in[87] & in2[87];
    assign P[21] = in[87] ^ in2[87];
    assign G[22] = in[86] & in2[86];
    assign P[22] = in[86] ^ in2[86];
    assign G[23] = in[85] & in2[85];
    assign P[23] = in[85] ^ in2[85];
    assign G[24] = in[84] & in2[84];
    assign P[24] = in[84] ^ in2[84];
    assign G[25] = in[83] & in2[83];
    assign P[25] = in[83] ^ in2[83];
    assign G[26] = in[82] & in2[82];
    assign P[26] = in[82] ^ in2[82];
    assign G[27] = in[81] & in2[81];
    assign P[27] = in[81] ^ in2[81];
    assign G[28] = in[80] & in2[80];
    assign P[28] = in[80] ^ in2[80];
    assign G[29] = in[79] & in2[79];
    assign P[29] = in[79] ^ in2[79];
    assign G[30] = in[78] & in2[78];
    assign P[30] = in[78] ^ in2[78];
    assign G[31] = in[77] & in2[77];
    assign P[31] = in[77] ^ in2[77];
    assign G[32] = in[76] & in2[76];
    assign P[32] = in[76] ^ in2[76];
    assign G[33] = in[75] & in2[75];
    assign P[33] = in[75] ^ in2[75];
    assign G[34] = in[74] & in2[74];
    assign P[34] = in[74] ^ in2[74];
    assign G[35] = in[73] & in2[73];
    assign P[35] = in[73] ^ in2[73];
    assign G[36] = in[72] & in2[72];
    assign P[36] = in[72] ^ in2[72];
    assign G[37] = in[71] & in2[71];
    assign P[37] = in[71] ^ in2[71];
    assign G[38] = in[70] & in2[70];
    assign P[38] = in[70] ^ in2[70];
    assign G[39] = in[69] & in2[69];
    assign P[39] = in[69] ^ in2[69];
    assign G[40] = in[68] & in2[68];
    assign P[40] = in[68] ^ in2[68];
    assign G[41] = in[67] & in2[67];
    assign P[41] = in[67] ^ in2[67];
    assign G[42] = in[66] & in2[66];
    assign P[42] = in[66] ^ in2[66];
    assign G[43] = in[65] & in2[65];
    assign P[43] = in[65] ^ in2[65];
    assign G[44] = in[64] & in2[64];
    assign P[44] = in[64] ^ in2[64];
    assign G[45] = in[63] & in2[63];
    assign P[45] = in[63] ^ in2[63];
    assign G[46] = in[62] & in2[62];
    assign P[46] = in[62] ^ in2[62];
    assign G[47] = in[61] & in2[61];
    assign P[47] = in[61] ^ in2[61];
    assign G[48] = in[60] & in2[60];
    assign P[48] = in[60] ^ in2[60];
    assign G[49] = in[59] & in2[59];
    assign P[49] = in[59] ^ in2[59];
    assign G[50] = in[58] & in2[58];
    assign P[50] = in[58] ^ in2[58];
    assign G[51] = in[57] & in2[57];
    assign P[51] = in[57] ^ in2[57];
    assign G[52] = in[56] & in2[56];
    assign P[52] = in[56] ^ in2[56];
    assign G[53] = in[55] & in2[55];
    assign P[53] = in[55] ^ in2[55];
    assign G[54] = in[54] & in2[54];
    assign P[54] = in[54] ^ in2[54];
    assign G[55] = in[53] & in2[53];
    assign P[55] = in[53] ^ in2[53];
    assign G[56] = in[52] & in2[52];
    assign P[56] = in[52] ^ in2[52];
    assign G[57] = in[51] & in2[51];
    assign P[57] = in[51] ^ in2[51];
    assign G[58] = in[50] & in2[50];
    assign P[58] = in[50] ^ in2[50];
    assign G[59] = in[49] & in2[49];
    assign P[59] = in[49] ^ in2[49];
    assign G[60] = in[48] & in2[48];
    assign P[60] = in[48] ^ in2[48];
    assign G[61] = in[47] & in2[47];
    assign P[61] = in[47] ^ in2[47];
    assign G[62] = in[46] & in2[46];
    assign P[62] = in[46] ^ in2[46];
    assign G[63] = in[45] & in2[45];
    assign P[63] = in[45] ^ in2[45];
    assign G[64] = in[44] & in2[44];
    assign P[64] = in[44] ^ in2[44];
    assign G[65] = in[43] & in2[43];
    assign P[65] = in[43] ^ in2[43];
    assign G[66] = in[42] & in2[42];
    assign P[66] = in[42] ^ in2[42];
    assign G[67] = in[41] & in2[41];
    assign P[67] = in[41] ^ in2[41];
    assign G[68] = in[40] & in2[40];
    assign P[68] = in[40] ^ in2[40];
    assign G[69] = in[39] & in2[39];
    assign P[69] = in[39] ^ in2[39];
    assign G[70] = in[38] & in2[38];
    assign P[70] = in[38] ^ in2[38];
    assign G[71] = in[37] & in2[37];
    assign P[71] = in[37] ^ in2[37];
    assign G[72] = in[36] & in2[36];
    assign P[72] = in[36] ^ in2[36];
    assign G[73] = in[35] & in2[35];
    assign P[73] = in[35] ^ in2[35];
    assign G[74] = in[34] & in2[34];
    assign P[74] = in[34] ^ in2[34];
    assign G[75] = in[33] & in2[33];
    assign P[75] = in[33] ^ in2[33];
    assign G[76] = in[32] & in2[32];
    assign P[76] = in[32] ^ in2[32];
    assign G[77] = in[31] & in2[31];
    assign P[77] = in[31] ^ in2[31];
    assign G[78] = in[30] & in2[30];
    assign P[78] = in[30] ^ in2[30];
    assign G[79] = in[29] & in2[29];
    assign P[79] = in[29] ^ in2[29];
    assign G[80] = in[28] & in2[28];
    assign P[80] = in[28] ^ in2[28];
    assign G[81] = in[27] & in2[27];
    assign P[81] = in[27] ^ in2[27];
    assign G[82] = in[26] & in2[26];
    assign P[82] = in[26] ^ in2[26];
    assign G[83] = in[25] & in2[25];
    assign P[83] = in[25] ^ in2[25];
    assign G[84] = in[24] & in2[24];
    assign P[84] = in[24] ^ in2[24];
    assign G[85] = in[23] & in2[23];
    assign P[85] = in[23] ^ in2[23];
    assign G[86] = in[22] & in2[22];
    assign P[86] = in[22] ^ in2[22];
    assign G[87] = in[21] & in2[21];
    assign P[87] = in[21] ^ in2[21];
    assign G[88] = in[20] & in2[20];
    assign P[88] = in[20] ^ in2[20];
    assign G[89] = in[19] & in2[19];
    assign P[89] = in[19] ^ in2[19];
    assign G[90] = in[18] & in2[18];
    assign P[90] = in[18] ^ in2[18];
    assign G[91] = in[17] & in2[17];
    assign P[91] = in[17] ^ in2[17];
    assign G[92] = in[16] & in2[16];
    assign P[92] = in[16] ^ in2[16];
    assign G[93] = in[15] & in2[15];
    assign P[93] = in[15] ^ in2[15];
    assign G[94] = in[14] & in2[14];
    assign P[94] = in[14] ^ in2[14];
    assign G[95] = in[13] & in2[13];
    assign P[95] = in[13] ^ in2[13];
    assign G[96] = in[12] & in2[12];
    assign P[96] = in[12] ^ in2[12];
    assign G[97] = in[11] & in2[11];
    assign P[97] = in[11] ^ in2[11];
    assign G[98] = in[10] & in2[10];
    assign P[98] = in[10] ^ in2[10];
    assign G[99] = in[9] & in2[9];
    assign P[99] = in[9] ^ in2[9];
    assign G[100] = in[8] & in2[8];
    assign P[100] = in[8] ^ in2[8];
    assign G[101] = in[7] & in2[7];
    assign P[101] = in[7] ^ in2[7];
    assign G[102] = in[6] & in2[6];
    assign P[102] = in[6] ^ in2[6];
    assign G[103] = in[5] & in2[5];
    assign P[103] = in[5] ^ in2[5];
    assign G[104] = in[4] & in2[4];
    assign P[104] = in[4] ^ in2[4];
    assign G[105] = in[3] & in2[3];
    assign P[105] = in[3] ^ in2[3];
    assign G[106] = in[2] & in2[2];
    assign P[106] = in[2] ^ in2[2];
    assign G[107] = in[1] & in2[1];
    assign P[107] = in[1] ^ in2[1];
    assign G[108] = in[0] & in2[0];
    assign P[108] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign C[108] = G[107] | (P[107] & C[107]);
    assign cout = G[108] | (P[108] & C[108]);
    assign sum = P ^ C;
endmodule

module CLA108(output [107:0] sum, output cout, input [107:0] in1, input [107:0] in2;

    wire[107:0] G;
    wire[107:0] C;
    wire[107:0] P;

    assign G[0] = in[107] & in2[107];
    assign P[0] = in[107] ^ in2[107];
    assign G[1] = in[106] & in2[106];
    assign P[1] = in[106] ^ in2[106];
    assign G[2] = in[105] & in2[105];
    assign P[2] = in[105] ^ in2[105];
    assign G[3] = in[104] & in2[104];
    assign P[3] = in[104] ^ in2[104];
    assign G[4] = in[103] & in2[103];
    assign P[4] = in[103] ^ in2[103];
    assign G[5] = in[102] & in2[102];
    assign P[5] = in[102] ^ in2[102];
    assign G[6] = in[101] & in2[101];
    assign P[6] = in[101] ^ in2[101];
    assign G[7] = in[100] & in2[100];
    assign P[7] = in[100] ^ in2[100];
    assign G[8] = in[99] & in2[99];
    assign P[8] = in[99] ^ in2[99];
    assign G[9] = in[98] & in2[98];
    assign P[9] = in[98] ^ in2[98];
    assign G[10] = in[97] & in2[97];
    assign P[10] = in[97] ^ in2[97];
    assign G[11] = in[96] & in2[96];
    assign P[11] = in[96] ^ in2[96];
    assign G[12] = in[95] & in2[95];
    assign P[12] = in[95] ^ in2[95];
    assign G[13] = in[94] & in2[94];
    assign P[13] = in[94] ^ in2[94];
    assign G[14] = in[93] & in2[93];
    assign P[14] = in[93] ^ in2[93];
    assign G[15] = in[92] & in2[92];
    assign P[15] = in[92] ^ in2[92];
    assign G[16] = in[91] & in2[91];
    assign P[16] = in[91] ^ in2[91];
    assign G[17] = in[90] & in2[90];
    assign P[17] = in[90] ^ in2[90];
    assign G[18] = in[89] & in2[89];
    assign P[18] = in[89] ^ in2[89];
    assign G[19] = in[88] & in2[88];
    assign P[19] = in[88] ^ in2[88];
    assign G[20] = in[87] & in2[87];
    assign P[20] = in[87] ^ in2[87];
    assign G[21] = in[86] & in2[86];
    assign P[21] = in[86] ^ in2[86];
    assign G[22] = in[85] & in2[85];
    assign P[22] = in[85] ^ in2[85];
    assign G[23] = in[84] & in2[84];
    assign P[23] = in[84] ^ in2[84];
    assign G[24] = in[83] & in2[83];
    assign P[24] = in[83] ^ in2[83];
    assign G[25] = in[82] & in2[82];
    assign P[25] = in[82] ^ in2[82];
    assign G[26] = in[81] & in2[81];
    assign P[26] = in[81] ^ in2[81];
    assign G[27] = in[80] & in2[80];
    assign P[27] = in[80] ^ in2[80];
    assign G[28] = in[79] & in2[79];
    assign P[28] = in[79] ^ in2[79];
    assign G[29] = in[78] & in2[78];
    assign P[29] = in[78] ^ in2[78];
    assign G[30] = in[77] & in2[77];
    assign P[30] = in[77] ^ in2[77];
    assign G[31] = in[76] & in2[76];
    assign P[31] = in[76] ^ in2[76];
    assign G[32] = in[75] & in2[75];
    assign P[32] = in[75] ^ in2[75];
    assign G[33] = in[74] & in2[74];
    assign P[33] = in[74] ^ in2[74];
    assign G[34] = in[73] & in2[73];
    assign P[34] = in[73] ^ in2[73];
    assign G[35] = in[72] & in2[72];
    assign P[35] = in[72] ^ in2[72];
    assign G[36] = in[71] & in2[71];
    assign P[36] = in[71] ^ in2[71];
    assign G[37] = in[70] & in2[70];
    assign P[37] = in[70] ^ in2[70];
    assign G[38] = in[69] & in2[69];
    assign P[38] = in[69] ^ in2[69];
    assign G[39] = in[68] & in2[68];
    assign P[39] = in[68] ^ in2[68];
    assign G[40] = in[67] & in2[67];
    assign P[40] = in[67] ^ in2[67];
    assign G[41] = in[66] & in2[66];
    assign P[41] = in[66] ^ in2[66];
    assign G[42] = in[65] & in2[65];
    assign P[42] = in[65] ^ in2[65];
    assign G[43] = in[64] & in2[64];
    assign P[43] = in[64] ^ in2[64];
    assign G[44] = in[63] & in2[63];
    assign P[44] = in[63] ^ in2[63];
    assign G[45] = in[62] & in2[62];
    assign P[45] = in[62] ^ in2[62];
    assign G[46] = in[61] & in2[61];
    assign P[46] = in[61] ^ in2[61];
    assign G[47] = in[60] & in2[60];
    assign P[47] = in[60] ^ in2[60];
    assign G[48] = in[59] & in2[59];
    assign P[48] = in[59] ^ in2[59];
    assign G[49] = in[58] & in2[58];
    assign P[49] = in[58] ^ in2[58];
    assign G[50] = in[57] & in2[57];
    assign P[50] = in[57] ^ in2[57];
    assign G[51] = in[56] & in2[56];
    assign P[51] = in[56] ^ in2[56];
    assign G[52] = in[55] & in2[55];
    assign P[52] = in[55] ^ in2[55];
    assign G[53] = in[54] & in2[54];
    assign P[53] = in[54] ^ in2[54];
    assign G[54] = in[53] & in2[53];
    assign P[54] = in[53] ^ in2[53];
    assign G[55] = in[52] & in2[52];
    assign P[55] = in[52] ^ in2[52];
    assign G[56] = in[51] & in2[51];
    assign P[56] = in[51] ^ in2[51];
    assign G[57] = in[50] & in2[50];
    assign P[57] = in[50] ^ in2[50];
    assign G[58] = in[49] & in2[49];
    assign P[58] = in[49] ^ in2[49];
    assign G[59] = in[48] & in2[48];
    assign P[59] = in[48] ^ in2[48];
    assign G[60] = in[47] & in2[47];
    assign P[60] = in[47] ^ in2[47];
    assign G[61] = in[46] & in2[46];
    assign P[61] = in[46] ^ in2[46];
    assign G[62] = in[45] & in2[45];
    assign P[62] = in[45] ^ in2[45];
    assign G[63] = in[44] & in2[44];
    assign P[63] = in[44] ^ in2[44];
    assign G[64] = in[43] & in2[43];
    assign P[64] = in[43] ^ in2[43];
    assign G[65] = in[42] & in2[42];
    assign P[65] = in[42] ^ in2[42];
    assign G[66] = in[41] & in2[41];
    assign P[66] = in[41] ^ in2[41];
    assign G[67] = in[40] & in2[40];
    assign P[67] = in[40] ^ in2[40];
    assign G[68] = in[39] & in2[39];
    assign P[68] = in[39] ^ in2[39];
    assign G[69] = in[38] & in2[38];
    assign P[69] = in[38] ^ in2[38];
    assign G[70] = in[37] & in2[37];
    assign P[70] = in[37] ^ in2[37];
    assign G[71] = in[36] & in2[36];
    assign P[71] = in[36] ^ in2[36];
    assign G[72] = in[35] & in2[35];
    assign P[72] = in[35] ^ in2[35];
    assign G[73] = in[34] & in2[34];
    assign P[73] = in[34] ^ in2[34];
    assign G[74] = in[33] & in2[33];
    assign P[74] = in[33] ^ in2[33];
    assign G[75] = in[32] & in2[32];
    assign P[75] = in[32] ^ in2[32];
    assign G[76] = in[31] & in2[31];
    assign P[76] = in[31] ^ in2[31];
    assign G[77] = in[30] & in2[30];
    assign P[77] = in[30] ^ in2[30];
    assign G[78] = in[29] & in2[29];
    assign P[78] = in[29] ^ in2[29];
    assign G[79] = in[28] & in2[28];
    assign P[79] = in[28] ^ in2[28];
    assign G[80] = in[27] & in2[27];
    assign P[80] = in[27] ^ in2[27];
    assign G[81] = in[26] & in2[26];
    assign P[81] = in[26] ^ in2[26];
    assign G[82] = in[25] & in2[25];
    assign P[82] = in[25] ^ in2[25];
    assign G[83] = in[24] & in2[24];
    assign P[83] = in[24] ^ in2[24];
    assign G[84] = in[23] & in2[23];
    assign P[84] = in[23] ^ in2[23];
    assign G[85] = in[22] & in2[22];
    assign P[85] = in[22] ^ in2[22];
    assign G[86] = in[21] & in2[21];
    assign P[86] = in[21] ^ in2[21];
    assign G[87] = in[20] & in2[20];
    assign P[87] = in[20] ^ in2[20];
    assign G[88] = in[19] & in2[19];
    assign P[88] = in[19] ^ in2[19];
    assign G[89] = in[18] & in2[18];
    assign P[89] = in[18] ^ in2[18];
    assign G[90] = in[17] & in2[17];
    assign P[90] = in[17] ^ in2[17];
    assign G[91] = in[16] & in2[16];
    assign P[91] = in[16] ^ in2[16];
    assign G[92] = in[15] & in2[15];
    assign P[92] = in[15] ^ in2[15];
    assign G[93] = in[14] & in2[14];
    assign P[93] = in[14] ^ in2[14];
    assign G[94] = in[13] & in2[13];
    assign P[94] = in[13] ^ in2[13];
    assign G[95] = in[12] & in2[12];
    assign P[95] = in[12] ^ in2[12];
    assign G[96] = in[11] & in2[11];
    assign P[96] = in[11] ^ in2[11];
    assign G[97] = in[10] & in2[10];
    assign P[97] = in[10] ^ in2[10];
    assign G[98] = in[9] & in2[9];
    assign P[98] = in[9] ^ in2[9];
    assign G[99] = in[8] & in2[8];
    assign P[99] = in[8] ^ in2[8];
    assign G[100] = in[7] & in2[7];
    assign P[100] = in[7] ^ in2[7];
    assign G[101] = in[6] & in2[6];
    assign P[101] = in[6] ^ in2[6];
    assign G[102] = in[5] & in2[5];
    assign P[102] = in[5] ^ in2[5];
    assign G[103] = in[4] & in2[4];
    assign P[103] = in[4] ^ in2[4];
    assign G[104] = in[3] & in2[3];
    assign P[104] = in[3] ^ in2[3];
    assign G[105] = in[2] & in2[2];
    assign P[105] = in[2] ^ in2[2];
    assign G[106] = in[1] & in2[1];
    assign P[106] = in[1] ^ in2[1];
    assign G[107] = in[0] & in2[0];
    assign P[107] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign C[107] = G[106] | (P[106] & C[106]);
    assign cout = G[107] | (P[107] & C[107]);
    assign sum = P ^ C;
endmodule

module CLA107(output [106:0] sum, output cout, input [106:0] in1, input [106:0] in2;

    wire[106:0] G;
    wire[106:0] C;
    wire[106:0] P;

    assign G[0] = in[106] & in2[106];
    assign P[0] = in[106] ^ in2[106];
    assign G[1] = in[105] & in2[105];
    assign P[1] = in[105] ^ in2[105];
    assign G[2] = in[104] & in2[104];
    assign P[2] = in[104] ^ in2[104];
    assign G[3] = in[103] & in2[103];
    assign P[3] = in[103] ^ in2[103];
    assign G[4] = in[102] & in2[102];
    assign P[4] = in[102] ^ in2[102];
    assign G[5] = in[101] & in2[101];
    assign P[5] = in[101] ^ in2[101];
    assign G[6] = in[100] & in2[100];
    assign P[6] = in[100] ^ in2[100];
    assign G[7] = in[99] & in2[99];
    assign P[7] = in[99] ^ in2[99];
    assign G[8] = in[98] & in2[98];
    assign P[8] = in[98] ^ in2[98];
    assign G[9] = in[97] & in2[97];
    assign P[9] = in[97] ^ in2[97];
    assign G[10] = in[96] & in2[96];
    assign P[10] = in[96] ^ in2[96];
    assign G[11] = in[95] & in2[95];
    assign P[11] = in[95] ^ in2[95];
    assign G[12] = in[94] & in2[94];
    assign P[12] = in[94] ^ in2[94];
    assign G[13] = in[93] & in2[93];
    assign P[13] = in[93] ^ in2[93];
    assign G[14] = in[92] & in2[92];
    assign P[14] = in[92] ^ in2[92];
    assign G[15] = in[91] & in2[91];
    assign P[15] = in[91] ^ in2[91];
    assign G[16] = in[90] & in2[90];
    assign P[16] = in[90] ^ in2[90];
    assign G[17] = in[89] & in2[89];
    assign P[17] = in[89] ^ in2[89];
    assign G[18] = in[88] & in2[88];
    assign P[18] = in[88] ^ in2[88];
    assign G[19] = in[87] & in2[87];
    assign P[19] = in[87] ^ in2[87];
    assign G[20] = in[86] & in2[86];
    assign P[20] = in[86] ^ in2[86];
    assign G[21] = in[85] & in2[85];
    assign P[21] = in[85] ^ in2[85];
    assign G[22] = in[84] & in2[84];
    assign P[22] = in[84] ^ in2[84];
    assign G[23] = in[83] & in2[83];
    assign P[23] = in[83] ^ in2[83];
    assign G[24] = in[82] & in2[82];
    assign P[24] = in[82] ^ in2[82];
    assign G[25] = in[81] & in2[81];
    assign P[25] = in[81] ^ in2[81];
    assign G[26] = in[80] & in2[80];
    assign P[26] = in[80] ^ in2[80];
    assign G[27] = in[79] & in2[79];
    assign P[27] = in[79] ^ in2[79];
    assign G[28] = in[78] & in2[78];
    assign P[28] = in[78] ^ in2[78];
    assign G[29] = in[77] & in2[77];
    assign P[29] = in[77] ^ in2[77];
    assign G[30] = in[76] & in2[76];
    assign P[30] = in[76] ^ in2[76];
    assign G[31] = in[75] & in2[75];
    assign P[31] = in[75] ^ in2[75];
    assign G[32] = in[74] & in2[74];
    assign P[32] = in[74] ^ in2[74];
    assign G[33] = in[73] & in2[73];
    assign P[33] = in[73] ^ in2[73];
    assign G[34] = in[72] & in2[72];
    assign P[34] = in[72] ^ in2[72];
    assign G[35] = in[71] & in2[71];
    assign P[35] = in[71] ^ in2[71];
    assign G[36] = in[70] & in2[70];
    assign P[36] = in[70] ^ in2[70];
    assign G[37] = in[69] & in2[69];
    assign P[37] = in[69] ^ in2[69];
    assign G[38] = in[68] & in2[68];
    assign P[38] = in[68] ^ in2[68];
    assign G[39] = in[67] & in2[67];
    assign P[39] = in[67] ^ in2[67];
    assign G[40] = in[66] & in2[66];
    assign P[40] = in[66] ^ in2[66];
    assign G[41] = in[65] & in2[65];
    assign P[41] = in[65] ^ in2[65];
    assign G[42] = in[64] & in2[64];
    assign P[42] = in[64] ^ in2[64];
    assign G[43] = in[63] & in2[63];
    assign P[43] = in[63] ^ in2[63];
    assign G[44] = in[62] & in2[62];
    assign P[44] = in[62] ^ in2[62];
    assign G[45] = in[61] & in2[61];
    assign P[45] = in[61] ^ in2[61];
    assign G[46] = in[60] & in2[60];
    assign P[46] = in[60] ^ in2[60];
    assign G[47] = in[59] & in2[59];
    assign P[47] = in[59] ^ in2[59];
    assign G[48] = in[58] & in2[58];
    assign P[48] = in[58] ^ in2[58];
    assign G[49] = in[57] & in2[57];
    assign P[49] = in[57] ^ in2[57];
    assign G[50] = in[56] & in2[56];
    assign P[50] = in[56] ^ in2[56];
    assign G[51] = in[55] & in2[55];
    assign P[51] = in[55] ^ in2[55];
    assign G[52] = in[54] & in2[54];
    assign P[52] = in[54] ^ in2[54];
    assign G[53] = in[53] & in2[53];
    assign P[53] = in[53] ^ in2[53];
    assign G[54] = in[52] & in2[52];
    assign P[54] = in[52] ^ in2[52];
    assign G[55] = in[51] & in2[51];
    assign P[55] = in[51] ^ in2[51];
    assign G[56] = in[50] & in2[50];
    assign P[56] = in[50] ^ in2[50];
    assign G[57] = in[49] & in2[49];
    assign P[57] = in[49] ^ in2[49];
    assign G[58] = in[48] & in2[48];
    assign P[58] = in[48] ^ in2[48];
    assign G[59] = in[47] & in2[47];
    assign P[59] = in[47] ^ in2[47];
    assign G[60] = in[46] & in2[46];
    assign P[60] = in[46] ^ in2[46];
    assign G[61] = in[45] & in2[45];
    assign P[61] = in[45] ^ in2[45];
    assign G[62] = in[44] & in2[44];
    assign P[62] = in[44] ^ in2[44];
    assign G[63] = in[43] & in2[43];
    assign P[63] = in[43] ^ in2[43];
    assign G[64] = in[42] & in2[42];
    assign P[64] = in[42] ^ in2[42];
    assign G[65] = in[41] & in2[41];
    assign P[65] = in[41] ^ in2[41];
    assign G[66] = in[40] & in2[40];
    assign P[66] = in[40] ^ in2[40];
    assign G[67] = in[39] & in2[39];
    assign P[67] = in[39] ^ in2[39];
    assign G[68] = in[38] & in2[38];
    assign P[68] = in[38] ^ in2[38];
    assign G[69] = in[37] & in2[37];
    assign P[69] = in[37] ^ in2[37];
    assign G[70] = in[36] & in2[36];
    assign P[70] = in[36] ^ in2[36];
    assign G[71] = in[35] & in2[35];
    assign P[71] = in[35] ^ in2[35];
    assign G[72] = in[34] & in2[34];
    assign P[72] = in[34] ^ in2[34];
    assign G[73] = in[33] & in2[33];
    assign P[73] = in[33] ^ in2[33];
    assign G[74] = in[32] & in2[32];
    assign P[74] = in[32] ^ in2[32];
    assign G[75] = in[31] & in2[31];
    assign P[75] = in[31] ^ in2[31];
    assign G[76] = in[30] & in2[30];
    assign P[76] = in[30] ^ in2[30];
    assign G[77] = in[29] & in2[29];
    assign P[77] = in[29] ^ in2[29];
    assign G[78] = in[28] & in2[28];
    assign P[78] = in[28] ^ in2[28];
    assign G[79] = in[27] & in2[27];
    assign P[79] = in[27] ^ in2[27];
    assign G[80] = in[26] & in2[26];
    assign P[80] = in[26] ^ in2[26];
    assign G[81] = in[25] & in2[25];
    assign P[81] = in[25] ^ in2[25];
    assign G[82] = in[24] & in2[24];
    assign P[82] = in[24] ^ in2[24];
    assign G[83] = in[23] & in2[23];
    assign P[83] = in[23] ^ in2[23];
    assign G[84] = in[22] & in2[22];
    assign P[84] = in[22] ^ in2[22];
    assign G[85] = in[21] & in2[21];
    assign P[85] = in[21] ^ in2[21];
    assign G[86] = in[20] & in2[20];
    assign P[86] = in[20] ^ in2[20];
    assign G[87] = in[19] & in2[19];
    assign P[87] = in[19] ^ in2[19];
    assign G[88] = in[18] & in2[18];
    assign P[88] = in[18] ^ in2[18];
    assign G[89] = in[17] & in2[17];
    assign P[89] = in[17] ^ in2[17];
    assign G[90] = in[16] & in2[16];
    assign P[90] = in[16] ^ in2[16];
    assign G[91] = in[15] & in2[15];
    assign P[91] = in[15] ^ in2[15];
    assign G[92] = in[14] & in2[14];
    assign P[92] = in[14] ^ in2[14];
    assign G[93] = in[13] & in2[13];
    assign P[93] = in[13] ^ in2[13];
    assign G[94] = in[12] & in2[12];
    assign P[94] = in[12] ^ in2[12];
    assign G[95] = in[11] & in2[11];
    assign P[95] = in[11] ^ in2[11];
    assign G[96] = in[10] & in2[10];
    assign P[96] = in[10] ^ in2[10];
    assign G[97] = in[9] & in2[9];
    assign P[97] = in[9] ^ in2[9];
    assign G[98] = in[8] & in2[8];
    assign P[98] = in[8] ^ in2[8];
    assign G[99] = in[7] & in2[7];
    assign P[99] = in[7] ^ in2[7];
    assign G[100] = in[6] & in2[6];
    assign P[100] = in[6] ^ in2[6];
    assign G[101] = in[5] & in2[5];
    assign P[101] = in[5] ^ in2[5];
    assign G[102] = in[4] & in2[4];
    assign P[102] = in[4] ^ in2[4];
    assign G[103] = in[3] & in2[3];
    assign P[103] = in[3] ^ in2[3];
    assign G[104] = in[2] & in2[2];
    assign P[104] = in[2] ^ in2[2];
    assign G[105] = in[1] & in2[1];
    assign P[105] = in[1] ^ in2[1];
    assign G[106] = in[0] & in2[0];
    assign P[106] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign C[106] = G[105] | (P[105] & C[105]);
    assign cout = G[106] | (P[106] & C[106]);
    assign sum = P ^ C;
endmodule

module CLA106(output [105:0] sum, output cout, input [105:0] in1, input [105:0] in2;

    wire[105:0] G;
    wire[105:0] C;
    wire[105:0] P;

    assign G[0] = in[105] & in2[105];
    assign P[0] = in[105] ^ in2[105];
    assign G[1] = in[104] & in2[104];
    assign P[1] = in[104] ^ in2[104];
    assign G[2] = in[103] & in2[103];
    assign P[2] = in[103] ^ in2[103];
    assign G[3] = in[102] & in2[102];
    assign P[3] = in[102] ^ in2[102];
    assign G[4] = in[101] & in2[101];
    assign P[4] = in[101] ^ in2[101];
    assign G[5] = in[100] & in2[100];
    assign P[5] = in[100] ^ in2[100];
    assign G[6] = in[99] & in2[99];
    assign P[6] = in[99] ^ in2[99];
    assign G[7] = in[98] & in2[98];
    assign P[7] = in[98] ^ in2[98];
    assign G[8] = in[97] & in2[97];
    assign P[8] = in[97] ^ in2[97];
    assign G[9] = in[96] & in2[96];
    assign P[9] = in[96] ^ in2[96];
    assign G[10] = in[95] & in2[95];
    assign P[10] = in[95] ^ in2[95];
    assign G[11] = in[94] & in2[94];
    assign P[11] = in[94] ^ in2[94];
    assign G[12] = in[93] & in2[93];
    assign P[12] = in[93] ^ in2[93];
    assign G[13] = in[92] & in2[92];
    assign P[13] = in[92] ^ in2[92];
    assign G[14] = in[91] & in2[91];
    assign P[14] = in[91] ^ in2[91];
    assign G[15] = in[90] & in2[90];
    assign P[15] = in[90] ^ in2[90];
    assign G[16] = in[89] & in2[89];
    assign P[16] = in[89] ^ in2[89];
    assign G[17] = in[88] & in2[88];
    assign P[17] = in[88] ^ in2[88];
    assign G[18] = in[87] & in2[87];
    assign P[18] = in[87] ^ in2[87];
    assign G[19] = in[86] & in2[86];
    assign P[19] = in[86] ^ in2[86];
    assign G[20] = in[85] & in2[85];
    assign P[20] = in[85] ^ in2[85];
    assign G[21] = in[84] & in2[84];
    assign P[21] = in[84] ^ in2[84];
    assign G[22] = in[83] & in2[83];
    assign P[22] = in[83] ^ in2[83];
    assign G[23] = in[82] & in2[82];
    assign P[23] = in[82] ^ in2[82];
    assign G[24] = in[81] & in2[81];
    assign P[24] = in[81] ^ in2[81];
    assign G[25] = in[80] & in2[80];
    assign P[25] = in[80] ^ in2[80];
    assign G[26] = in[79] & in2[79];
    assign P[26] = in[79] ^ in2[79];
    assign G[27] = in[78] & in2[78];
    assign P[27] = in[78] ^ in2[78];
    assign G[28] = in[77] & in2[77];
    assign P[28] = in[77] ^ in2[77];
    assign G[29] = in[76] & in2[76];
    assign P[29] = in[76] ^ in2[76];
    assign G[30] = in[75] & in2[75];
    assign P[30] = in[75] ^ in2[75];
    assign G[31] = in[74] & in2[74];
    assign P[31] = in[74] ^ in2[74];
    assign G[32] = in[73] & in2[73];
    assign P[32] = in[73] ^ in2[73];
    assign G[33] = in[72] & in2[72];
    assign P[33] = in[72] ^ in2[72];
    assign G[34] = in[71] & in2[71];
    assign P[34] = in[71] ^ in2[71];
    assign G[35] = in[70] & in2[70];
    assign P[35] = in[70] ^ in2[70];
    assign G[36] = in[69] & in2[69];
    assign P[36] = in[69] ^ in2[69];
    assign G[37] = in[68] & in2[68];
    assign P[37] = in[68] ^ in2[68];
    assign G[38] = in[67] & in2[67];
    assign P[38] = in[67] ^ in2[67];
    assign G[39] = in[66] & in2[66];
    assign P[39] = in[66] ^ in2[66];
    assign G[40] = in[65] & in2[65];
    assign P[40] = in[65] ^ in2[65];
    assign G[41] = in[64] & in2[64];
    assign P[41] = in[64] ^ in2[64];
    assign G[42] = in[63] & in2[63];
    assign P[42] = in[63] ^ in2[63];
    assign G[43] = in[62] & in2[62];
    assign P[43] = in[62] ^ in2[62];
    assign G[44] = in[61] & in2[61];
    assign P[44] = in[61] ^ in2[61];
    assign G[45] = in[60] & in2[60];
    assign P[45] = in[60] ^ in2[60];
    assign G[46] = in[59] & in2[59];
    assign P[46] = in[59] ^ in2[59];
    assign G[47] = in[58] & in2[58];
    assign P[47] = in[58] ^ in2[58];
    assign G[48] = in[57] & in2[57];
    assign P[48] = in[57] ^ in2[57];
    assign G[49] = in[56] & in2[56];
    assign P[49] = in[56] ^ in2[56];
    assign G[50] = in[55] & in2[55];
    assign P[50] = in[55] ^ in2[55];
    assign G[51] = in[54] & in2[54];
    assign P[51] = in[54] ^ in2[54];
    assign G[52] = in[53] & in2[53];
    assign P[52] = in[53] ^ in2[53];
    assign G[53] = in[52] & in2[52];
    assign P[53] = in[52] ^ in2[52];
    assign G[54] = in[51] & in2[51];
    assign P[54] = in[51] ^ in2[51];
    assign G[55] = in[50] & in2[50];
    assign P[55] = in[50] ^ in2[50];
    assign G[56] = in[49] & in2[49];
    assign P[56] = in[49] ^ in2[49];
    assign G[57] = in[48] & in2[48];
    assign P[57] = in[48] ^ in2[48];
    assign G[58] = in[47] & in2[47];
    assign P[58] = in[47] ^ in2[47];
    assign G[59] = in[46] & in2[46];
    assign P[59] = in[46] ^ in2[46];
    assign G[60] = in[45] & in2[45];
    assign P[60] = in[45] ^ in2[45];
    assign G[61] = in[44] & in2[44];
    assign P[61] = in[44] ^ in2[44];
    assign G[62] = in[43] & in2[43];
    assign P[62] = in[43] ^ in2[43];
    assign G[63] = in[42] & in2[42];
    assign P[63] = in[42] ^ in2[42];
    assign G[64] = in[41] & in2[41];
    assign P[64] = in[41] ^ in2[41];
    assign G[65] = in[40] & in2[40];
    assign P[65] = in[40] ^ in2[40];
    assign G[66] = in[39] & in2[39];
    assign P[66] = in[39] ^ in2[39];
    assign G[67] = in[38] & in2[38];
    assign P[67] = in[38] ^ in2[38];
    assign G[68] = in[37] & in2[37];
    assign P[68] = in[37] ^ in2[37];
    assign G[69] = in[36] & in2[36];
    assign P[69] = in[36] ^ in2[36];
    assign G[70] = in[35] & in2[35];
    assign P[70] = in[35] ^ in2[35];
    assign G[71] = in[34] & in2[34];
    assign P[71] = in[34] ^ in2[34];
    assign G[72] = in[33] & in2[33];
    assign P[72] = in[33] ^ in2[33];
    assign G[73] = in[32] & in2[32];
    assign P[73] = in[32] ^ in2[32];
    assign G[74] = in[31] & in2[31];
    assign P[74] = in[31] ^ in2[31];
    assign G[75] = in[30] & in2[30];
    assign P[75] = in[30] ^ in2[30];
    assign G[76] = in[29] & in2[29];
    assign P[76] = in[29] ^ in2[29];
    assign G[77] = in[28] & in2[28];
    assign P[77] = in[28] ^ in2[28];
    assign G[78] = in[27] & in2[27];
    assign P[78] = in[27] ^ in2[27];
    assign G[79] = in[26] & in2[26];
    assign P[79] = in[26] ^ in2[26];
    assign G[80] = in[25] & in2[25];
    assign P[80] = in[25] ^ in2[25];
    assign G[81] = in[24] & in2[24];
    assign P[81] = in[24] ^ in2[24];
    assign G[82] = in[23] & in2[23];
    assign P[82] = in[23] ^ in2[23];
    assign G[83] = in[22] & in2[22];
    assign P[83] = in[22] ^ in2[22];
    assign G[84] = in[21] & in2[21];
    assign P[84] = in[21] ^ in2[21];
    assign G[85] = in[20] & in2[20];
    assign P[85] = in[20] ^ in2[20];
    assign G[86] = in[19] & in2[19];
    assign P[86] = in[19] ^ in2[19];
    assign G[87] = in[18] & in2[18];
    assign P[87] = in[18] ^ in2[18];
    assign G[88] = in[17] & in2[17];
    assign P[88] = in[17] ^ in2[17];
    assign G[89] = in[16] & in2[16];
    assign P[89] = in[16] ^ in2[16];
    assign G[90] = in[15] & in2[15];
    assign P[90] = in[15] ^ in2[15];
    assign G[91] = in[14] & in2[14];
    assign P[91] = in[14] ^ in2[14];
    assign G[92] = in[13] & in2[13];
    assign P[92] = in[13] ^ in2[13];
    assign G[93] = in[12] & in2[12];
    assign P[93] = in[12] ^ in2[12];
    assign G[94] = in[11] & in2[11];
    assign P[94] = in[11] ^ in2[11];
    assign G[95] = in[10] & in2[10];
    assign P[95] = in[10] ^ in2[10];
    assign G[96] = in[9] & in2[9];
    assign P[96] = in[9] ^ in2[9];
    assign G[97] = in[8] & in2[8];
    assign P[97] = in[8] ^ in2[8];
    assign G[98] = in[7] & in2[7];
    assign P[98] = in[7] ^ in2[7];
    assign G[99] = in[6] & in2[6];
    assign P[99] = in[6] ^ in2[6];
    assign G[100] = in[5] & in2[5];
    assign P[100] = in[5] ^ in2[5];
    assign G[101] = in[4] & in2[4];
    assign P[101] = in[4] ^ in2[4];
    assign G[102] = in[3] & in2[3];
    assign P[102] = in[3] ^ in2[3];
    assign G[103] = in[2] & in2[2];
    assign P[103] = in[2] ^ in2[2];
    assign G[104] = in[1] & in2[1];
    assign P[104] = in[1] ^ in2[1];
    assign G[105] = in[0] & in2[0];
    assign P[105] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign C[105] = G[104] | (P[104] & C[104]);
    assign cout = G[105] | (P[105] & C[105]);
    assign sum = P ^ C;
endmodule

module CLA105(output [104:0] sum, output cout, input [104:0] in1, input [104:0] in2;

    wire[104:0] G;
    wire[104:0] C;
    wire[104:0] P;

    assign G[0] = in[104] & in2[104];
    assign P[0] = in[104] ^ in2[104];
    assign G[1] = in[103] & in2[103];
    assign P[1] = in[103] ^ in2[103];
    assign G[2] = in[102] & in2[102];
    assign P[2] = in[102] ^ in2[102];
    assign G[3] = in[101] & in2[101];
    assign P[3] = in[101] ^ in2[101];
    assign G[4] = in[100] & in2[100];
    assign P[4] = in[100] ^ in2[100];
    assign G[5] = in[99] & in2[99];
    assign P[5] = in[99] ^ in2[99];
    assign G[6] = in[98] & in2[98];
    assign P[6] = in[98] ^ in2[98];
    assign G[7] = in[97] & in2[97];
    assign P[7] = in[97] ^ in2[97];
    assign G[8] = in[96] & in2[96];
    assign P[8] = in[96] ^ in2[96];
    assign G[9] = in[95] & in2[95];
    assign P[9] = in[95] ^ in2[95];
    assign G[10] = in[94] & in2[94];
    assign P[10] = in[94] ^ in2[94];
    assign G[11] = in[93] & in2[93];
    assign P[11] = in[93] ^ in2[93];
    assign G[12] = in[92] & in2[92];
    assign P[12] = in[92] ^ in2[92];
    assign G[13] = in[91] & in2[91];
    assign P[13] = in[91] ^ in2[91];
    assign G[14] = in[90] & in2[90];
    assign P[14] = in[90] ^ in2[90];
    assign G[15] = in[89] & in2[89];
    assign P[15] = in[89] ^ in2[89];
    assign G[16] = in[88] & in2[88];
    assign P[16] = in[88] ^ in2[88];
    assign G[17] = in[87] & in2[87];
    assign P[17] = in[87] ^ in2[87];
    assign G[18] = in[86] & in2[86];
    assign P[18] = in[86] ^ in2[86];
    assign G[19] = in[85] & in2[85];
    assign P[19] = in[85] ^ in2[85];
    assign G[20] = in[84] & in2[84];
    assign P[20] = in[84] ^ in2[84];
    assign G[21] = in[83] & in2[83];
    assign P[21] = in[83] ^ in2[83];
    assign G[22] = in[82] & in2[82];
    assign P[22] = in[82] ^ in2[82];
    assign G[23] = in[81] & in2[81];
    assign P[23] = in[81] ^ in2[81];
    assign G[24] = in[80] & in2[80];
    assign P[24] = in[80] ^ in2[80];
    assign G[25] = in[79] & in2[79];
    assign P[25] = in[79] ^ in2[79];
    assign G[26] = in[78] & in2[78];
    assign P[26] = in[78] ^ in2[78];
    assign G[27] = in[77] & in2[77];
    assign P[27] = in[77] ^ in2[77];
    assign G[28] = in[76] & in2[76];
    assign P[28] = in[76] ^ in2[76];
    assign G[29] = in[75] & in2[75];
    assign P[29] = in[75] ^ in2[75];
    assign G[30] = in[74] & in2[74];
    assign P[30] = in[74] ^ in2[74];
    assign G[31] = in[73] & in2[73];
    assign P[31] = in[73] ^ in2[73];
    assign G[32] = in[72] & in2[72];
    assign P[32] = in[72] ^ in2[72];
    assign G[33] = in[71] & in2[71];
    assign P[33] = in[71] ^ in2[71];
    assign G[34] = in[70] & in2[70];
    assign P[34] = in[70] ^ in2[70];
    assign G[35] = in[69] & in2[69];
    assign P[35] = in[69] ^ in2[69];
    assign G[36] = in[68] & in2[68];
    assign P[36] = in[68] ^ in2[68];
    assign G[37] = in[67] & in2[67];
    assign P[37] = in[67] ^ in2[67];
    assign G[38] = in[66] & in2[66];
    assign P[38] = in[66] ^ in2[66];
    assign G[39] = in[65] & in2[65];
    assign P[39] = in[65] ^ in2[65];
    assign G[40] = in[64] & in2[64];
    assign P[40] = in[64] ^ in2[64];
    assign G[41] = in[63] & in2[63];
    assign P[41] = in[63] ^ in2[63];
    assign G[42] = in[62] & in2[62];
    assign P[42] = in[62] ^ in2[62];
    assign G[43] = in[61] & in2[61];
    assign P[43] = in[61] ^ in2[61];
    assign G[44] = in[60] & in2[60];
    assign P[44] = in[60] ^ in2[60];
    assign G[45] = in[59] & in2[59];
    assign P[45] = in[59] ^ in2[59];
    assign G[46] = in[58] & in2[58];
    assign P[46] = in[58] ^ in2[58];
    assign G[47] = in[57] & in2[57];
    assign P[47] = in[57] ^ in2[57];
    assign G[48] = in[56] & in2[56];
    assign P[48] = in[56] ^ in2[56];
    assign G[49] = in[55] & in2[55];
    assign P[49] = in[55] ^ in2[55];
    assign G[50] = in[54] & in2[54];
    assign P[50] = in[54] ^ in2[54];
    assign G[51] = in[53] & in2[53];
    assign P[51] = in[53] ^ in2[53];
    assign G[52] = in[52] & in2[52];
    assign P[52] = in[52] ^ in2[52];
    assign G[53] = in[51] & in2[51];
    assign P[53] = in[51] ^ in2[51];
    assign G[54] = in[50] & in2[50];
    assign P[54] = in[50] ^ in2[50];
    assign G[55] = in[49] & in2[49];
    assign P[55] = in[49] ^ in2[49];
    assign G[56] = in[48] & in2[48];
    assign P[56] = in[48] ^ in2[48];
    assign G[57] = in[47] & in2[47];
    assign P[57] = in[47] ^ in2[47];
    assign G[58] = in[46] & in2[46];
    assign P[58] = in[46] ^ in2[46];
    assign G[59] = in[45] & in2[45];
    assign P[59] = in[45] ^ in2[45];
    assign G[60] = in[44] & in2[44];
    assign P[60] = in[44] ^ in2[44];
    assign G[61] = in[43] & in2[43];
    assign P[61] = in[43] ^ in2[43];
    assign G[62] = in[42] & in2[42];
    assign P[62] = in[42] ^ in2[42];
    assign G[63] = in[41] & in2[41];
    assign P[63] = in[41] ^ in2[41];
    assign G[64] = in[40] & in2[40];
    assign P[64] = in[40] ^ in2[40];
    assign G[65] = in[39] & in2[39];
    assign P[65] = in[39] ^ in2[39];
    assign G[66] = in[38] & in2[38];
    assign P[66] = in[38] ^ in2[38];
    assign G[67] = in[37] & in2[37];
    assign P[67] = in[37] ^ in2[37];
    assign G[68] = in[36] & in2[36];
    assign P[68] = in[36] ^ in2[36];
    assign G[69] = in[35] & in2[35];
    assign P[69] = in[35] ^ in2[35];
    assign G[70] = in[34] & in2[34];
    assign P[70] = in[34] ^ in2[34];
    assign G[71] = in[33] & in2[33];
    assign P[71] = in[33] ^ in2[33];
    assign G[72] = in[32] & in2[32];
    assign P[72] = in[32] ^ in2[32];
    assign G[73] = in[31] & in2[31];
    assign P[73] = in[31] ^ in2[31];
    assign G[74] = in[30] & in2[30];
    assign P[74] = in[30] ^ in2[30];
    assign G[75] = in[29] & in2[29];
    assign P[75] = in[29] ^ in2[29];
    assign G[76] = in[28] & in2[28];
    assign P[76] = in[28] ^ in2[28];
    assign G[77] = in[27] & in2[27];
    assign P[77] = in[27] ^ in2[27];
    assign G[78] = in[26] & in2[26];
    assign P[78] = in[26] ^ in2[26];
    assign G[79] = in[25] & in2[25];
    assign P[79] = in[25] ^ in2[25];
    assign G[80] = in[24] & in2[24];
    assign P[80] = in[24] ^ in2[24];
    assign G[81] = in[23] & in2[23];
    assign P[81] = in[23] ^ in2[23];
    assign G[82] = in[22] & in2[22];
    assign P[82] = in[22] ^ in2[22];
    assign G[83] = in[21] & in2[21];
    assign P[83] = in[21] ^ in2[21];
    assign G[84] = in[20] & in2[20];
    assign P[84] = in[20] ^ in2[20];
    assign G[85] = in[19] & in2[19];
    assign P[85] = in[19] ^ in2[19];
    assign G[86] = in[18] & in2[18];
    assign P[86] = in[18] ^ in2[18];
    assign G[87] = in[17] & in2[17];
    assign P[87] = in[17] ^ in2[17];
    assign G[88] = in[16] & in2[16];
    assign P[88] = in[16] ^ in2[16];
    assign G[89] = in[15] & in2[15];
    assign P[89] = in[15] ^ in2[15];
    assign G[90] = in[14] & in2[14];
    assign P[90] = in[14] ^ in2[14];
    assign G[91] = in[13] & in2[13];
    assign P[91] = in[13] ^ in2[13];
    assign G[92] = in[12] & in2[12];
    assign P[92] = in[12] ^ in2[12];
    assign G[93] = in[11] & in2[11];
    assign P[93] = in[11] ^ in2[11];
    assign G[94] = in[10] & in2[10];
    assign P[94] = in[10] ^ in2[10];
    assign G[95] = in[9] & in2[9];
    assign P[95] = in[9] ^ in2[9];
    assign G[96] = in[8] & in2[8];
    assign P[96] = in[8] ^ in2[8];
    assign G[97] = in[7] & in2[7];
    assign P[97] = in[7] ^ in2[7];
    assign G[98] = in[6] & in2[6];
    assign P[98] = in[6] ^ in2[6];
    assign G[99] = in[5] & in2[5];
    assign P[99] = in[5] ^ in2[5];
    assign G[100] = in[4] & in2[4];
    assign P[100] = in[4] ^ in2[4];
    assign G[101] = in[3] & in2[3];
    assign P[101] = in[3] ^ in2[3];
    assign G[102] = in[2] & in2[2];
    assign P[102] = in[2] ^ in2[2];
    assign G[103] = in[1] & in2[1];
    assign P[103] = in[1] ^ in2[1];
    assign G[104] = in[0] & in2[0];
    assign P[104] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign C[104] = G[103] | (P[103] & C[103]);
    assign cout = G[104] | (P[104] & C[104]);
    assign sum = P ^ C;
endmodule

module CLA104(output [103:0] sum, output cout, input [103:0] in1, input [103:0] in2;

    wire[103:0] G;
    wire[103:0] C;
    wire[103:0] P;

    assign G[0] = in[103] & in2[103];
    assign P[0] = in[103] ^ in2[103];
    assign G[1] = in[102] & in2[102];
    assign P[1] = in[102] ^ in2[102];
    assign G[2] = in[101] & in2[101];
    assign P[2] = in[101] ^ in2[101];
    assign G[3] = in[100] & in2[100];
    assign P[3] = in[100] ^ in2[100];
    assign G[4] = in[99] & in2[99];
    assign P[4] = in[99] ^ in2[99];
    assign G[5] = in[98] & in2[98];
    assign P[5] = in[98] ^ in2[98];
    assign G[6] = in[97] & in2[97];
    assign P[6] = in[97] ^ in2[97];
    assign G[7] = in[96] & in2[96];
    assign P[7] = in[96] ^ in2[96];
    assign G[8] = in[95] & in2[95];
    assign P[8] = in[95] ^ in2[95];
    assign G[9] = in[94] & in2[94];
    assign P[9] = in[94] ^ in2[94];
    assign G[10] = in[93] & in2[93];
    assign P[10] = in[93] ^ in2[93];
    assign G[11] = in[92] & in2[92];
    assign P[11] = in[92] ^ in2[92];
    assign G[12] = in[91] & in2[91];
    assign P[12] = in[91] ^ in2[91];
    assign G[13] = in[90] & in2[90];
    assign P[13] = in[90] ^ in2[90];
    assign G[14] = in[89] & in2[89];
    assign P[14] = in[89] ^ in2[89];
    assign G[15] = in[88] & in2[88];
    assign P[15] = in[88] ^ in2[88];
    assign G[16] = in[87] & in2[87];
    assign P[16] = in[87] ^ in2[87];
    assign G[17] = in[86] & in2[86];
    assign P[17] = in[86] ^ in2[86];
    assign G[18] = in[85] & in2[85];
    assign P[18] = in[85] ^ in2[85];
    assign G[19] = in[84] & in2[84];
    assign P[19] = in[84] ^ in2[84];
    assign G[20] = in[83] & in2[83];
    assign P[20] = in[83] ^ in2[83];
    assign G[21] = in[82] & in2[82];
    assign P[21] = in[82] ^ in2[82];
    assign G[22] = in[81] & in2[81];
    assign P[22] = in[81] ^ in2[81];
    assign G[23] = in[80] & in2[80];
    assign P[23] = in[80] ^ in2[80];
    assign G[24] = in[79] & in2[79];
    assign P[24] = in[79] ^ in2[79];
    assign G[25] = in[78] & in2[78];
    assign P[25] = in[78] ^ in2[78];
    assign G[26] = in[77] & in2[77];
    assign P[26] = in[77] ^ in2[77];
    assign G[27] = in[76] & in2[76];
    assign P[27] = in[76] ^ in2[76];
    assign G[28] = in[75] & in2[75];
    assign P[28] = in[75] ^ in2[75];
    assign G[29] = in[74] & in2[74];
    assign P[29] = in[74] ^ in2[74];
    assign G[30] = in[73] & in2[73];
    assign P[30] = in[73] ^ in2[73];
    assign G[31] = in[72] & in2[72];
    assign P[31] = in[72] ^ in2[72];
    assign G[32] = in[71] & in2[71];
    assign P[32] = in[71] ^ in2[71];
    assign G[33] = in[70] & in2[70];
    assign P[33] = in[70] ^ in2[70];
    assign G[34] = in[69] & in2[69];
    assign P[34] = in[69] ^ in2[69];
    assign G[35] = in[68] & in2[68];
    assign P[35] = in[68] ^ in2[68];
    assign G[36] = in[67] & in2[67];
    assign P[36] = in[67] ^ in2[67];
    assign G[37] = in[66] & in2[66];
    assign P[37] = in[66] ^ in2[66];
    assign G[38] = in[65] & in2[65];
    assign P[38] = in[65] ^ in2[65];
    assign G[39] = in[64] & in2[64];
    assign P[39] = in[64] ^ in2[64];
    assign G[40] = in[63] & in2[63];
    assign P[40] = in[63] ^ in2[63];
    assign G[41] = in[62] & in2[62];
    assign P[41] = in[62] ^ in2[62];
    assign G[42] = in[61] & in2[61];
    assign P[42] = in[61] ^ in2[61];
    assign G[43] = in[60] & in2[60];
    assign P[43] = in[60] ^ in2[60];
    assign G[44] = in[59] & in2[59];
    assign P[44] = in[59] ^ in2[59];
    assign G[45] = in[58] & in2[58];
    assign P[45] = in[58] ^ in2[58];
    assign G[46] = in[57] & in2[57];
    assign P[46] = in[57] ^ in2[57];
    assign G[47] = in[56] & in2[56];
    assign P[47] = in[56] ^ in2[56];
    assign G[48] = in[55] & in2[55];
    assign P[48] = in[55] ^ in2[55];
    assign G[49] = in[54] & in2[54];
    assign P[49] = in[54] ^ in2[54];
    assign G[50] = in[53] & in2[53];
    assign P[50] = in[53] ^ in2[53];
    assign G[51] = in[52] & in2[52];
    assign P[51] = in[52] ^ in2[52];
    assign G[52] = in[51] & in2[51];
    assign P[52] = in[51] ^ in2[51];
    assign G[53] = in[50] & in2[50];
    assign P[53] = in[50] ^ in2[50];
    assign G[54] = in[49] & in2[49];
    assign P[54] = in[49] ^ in2[49];
    assign G[55] = in[48] & in2[48];
    assign P[55] = in[48] ^ in2[48];
    assign G[56] = in[47] & in2[47];
    assign P[56] = in[47] ^ in2[47];
    assign G[57] = in[46] & in2[46];
    assign P[57] = in[46] ^ in2[46];
    assign G[58] = in[45] & in2[45];
    assign P[58] = in[45] ^ in2[45];
    assign G[59] = in[44] & in2[44];
    assign P[59] = in[44] ^ in2[44];
    assign G[60] = in[43] & in2[43];
    assign P[60] = in[43] ^ in2[43];
    assign G[61] = in[42] & in2[42];
    assign P[61] = in[42] ^ in2[42];
    assign G[62] = in[41] & in2[41];
    assign P[62] = in[41] ^ in2[41];
    assign G[63] = in[40] & in2[40];
    assign P[63] = in[40] ^ in2[40];
    assign G[64] = in[39] & in2[39];
    assign P[64] = in[39] ^ in2[39];
    assign G[65] = in[38] & in2[38];
    assign P[65] = in[38] ^ in2[38];
    assign G[66] = in[37] & in2[37];
    assign P[66] = in[37] ^ in2[37];
    assign G[67] = in[36] & in2[36];
    assign P[67] = in[36] ^ in2[36];
    assign G[68] = in[35] & in2[35];
    assign P[68] = in[35] ^ in2[35];
    assign G[69] = in[34] & in2[34];
    assign P[69] = in[34] ^ in2[34];
    assign G[70] = in[33] & in2[33];
    assign P[70] = in[33] ^ in2[33];
    assign G[71] = in[32] & in2[32];
    assign P[71] = in[32] ^ in2[32];
    assign G[72] = in[31] & in2[31];
    assign P[72] = in[31] ^ in2[31];
    assign G[73] = in[30] & in2[30];
    assign P[73] = in[30] ^ in2[30];
    assign G[74] = in[29] & in2[29];
    assign P[74] = in[29] ^ in2[29];
    assign G[75] = in[28] & in2[28];
    assign P[75] = in[28] ^ in2[28];
    assign G[76] = in[27] & in2[27];
    assign P[76] = in[27] ^ in2[27];
    assign G[77] = in[26] & in2[26];
    assign P[77] = in[26] ^ in2[26];
    assign G[78] = in[25] & in2[25];
    assign P[78] = in[25] ^ in2[25];
    assign G[79] = in[24] & in2[24];
    assign P[79] = in[24] ^ in2[24];
    assign G[80] = in[23] & in2[23];
    assign P[80] = in[23] ^ in2[23];
    assign G[81] = in[22] & in2[22];
    assign P[81] = in[22] ^ in2[22];
    assign G[82] = in[21] & in2[21];
    assign P[82] = in[21] ^ in2[21];
    assign G[83] = in[20] & in2[20];
    assign P[83] = in[20] ^ in2[20];
    assign G[84] = in[19] & in2[19];
    assign P[84] = in[19] ^ in2[19];
    assign G[85] = in[18] & in2[18];
    assign P[85] = in[18] ^ in2[18];
    assign G[86] = in[17] & in2[17];
    assign P[86] = in[17] ^ in2[17];
    assign G[87] = in[16] & in2[16];
    assign P[87] = in[16] ^ in2[16];
    assign G[88] = in[15] & in2[15];
    assign P[88] = in[15] ^ in2[15];
    assign G[89] = in[14] & in2[14];
    assign P[89] = in[14] ^ in2[14];
    assign G[90] = in[13] & in2[13];
    assign P[90] = in[13] ^ in2[13];
    assign G[91] = in[12] & in2[12];
    assign P[91] = in[12] ^ in2[12];
    assign G[92] = in[11] & in2[11];
    assign P[92] = in[11] ^ in2[11];
    assign G[93] = in[10] & in2[10];
    assign P[93] = in[10] ^ in2[10];
    assign G[94] = in[9] & in2[9];
    assign P[94] = in[9] ^ in2[9];
    assign G[95] = in[8] & in2[8];
    assign P[95] = in[8] ^ in2[8];
    assign G[96] = in[7] & in2[7];
    assign P[96] = in[7] ^ in2[7];
    assign G[97] = in[6] & in2[6];
    assign P[97] = in[6] ^ in2[6];
    assign G[98] = in[5] & in2[5];
    assign P[98] = in[5] ^ in2[5];
    assign G[99] = in[4] & in2[4];
    assign P[99] = in[4] ^ in2[4];
    assign G[100] = in[3] & in2[3];
    assign P[100] = in[3] ^ in2[3];
    assign G[101] = in[2] & in2[2];
    assign P[101] = in[2] ^ in2[2];
    assign G[102] = in[1] & in2[1];
    assign P[102] = in[1] ^ in2[1];
    assign G[103] = in[0] & in2[0];
    assign P[103] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign C[103] = G[102] | (P[102] & C[102]);
    assign cout = G[103] | (P[103] & C[103]);
    assign sum = P ^ C;
endmodule

module CLA103(output [102:0] sum, output cout, input [102:0] in1, input [102:0] in2;

    wire[102:0] G;
    wire[102:0] C;
    wire[102:0] P;

    assign G[0] = in[102] & in2[102];
    assign P[0] = in[102] ^ in2[102];
    assign G[1] = in[101] & in2[101];
    assign P[1] = in[101] ^ in2[101];
    assign G[2] = in[100] & in2[100];
    assign P[2] = in[100] ^ in2[100];
    assign G[3] = in[99] & in2[99];
    assign P[3] = in[99] ^ in2[99];
    assign G[4] = in[98] & in2[98];
    assign P[4] = in[98] ^ in2[98];
    assign G[5] = in[97] & in2[97];
    assign P[5] = in[97] ^ in2[97];
    assign G[6] = in[96] & in2[96];
    assign P[6] = in[96] ^ in2[96];
    assign G[7] = in[95] & in2[95];
    assign P[7] = in[95] ^ in2[95];
    assign G[8] = in[94] & in2[94];
    assign P[8] = in[94] ^ in2[94];
    assign G[9] = in[93] & in2[93];
    assign P[9] = in[93] ^ in2[93];
    assign G[10] = in[92] & in2[92];
    assign P[10] = in[92] ^ in2[92];
    assign G[11] = in[91] & in2[91];
    assign P[11] = in[91] ^ in2[91];
    assign G[12] = in[90] & in2[90];
    assign P[12] = in[90] ^ in2[90];
    assign G[13] = in[89] & in2[89];
    assign P[13] = in[89] ^ in2[89];
    assign G[14] = in[88] & in2[88];
    assign P[14] = in[88] ^ in2[88];
    assign G[15] = in[87] & in2[87];
    assign P[15] = in[87] ^ in2[87];
    assign G[16] = in[86] & in2[86];
    assign P[16] = in[86] ^ in2[86];
    assign G[17] = in[85] & in2[85];
    assign P[17] = in[85] ^ in2[85];
    assign G[18] = in[84] & in2[84];
    assign P[18] = in[84] ^ in2[84];
    assign G[19] = in[83] & in2[83];
    assign P[19] = in[83] ^ in2[83];
    assign G[20] = in[82] & in2[82];
    assign P[20] = in[82] ^ in2[82];
    assign G[21] = in[81] & in2[81];
    assign P[21] = in[81] ^ in2[81];
    assign G[22] = in[80] & in2[80];
    assign P[22] = in[80] ^ in2[80];
    assign G[23] = in[79] & in2[79];
    assign P[23] = in[79] ^ in2[79];
    assign G[24] = in[78] & in2[78];
    assign P[24] = in[78] ^ in2[78];
    assign G[25] = in[77] & in2[77];
    assign P[25] = in[77] ^ in2[77];
    assign G[26] = in[76] & in2[76];
    assign P[26] = in[76] ^ in2[76];
    assign G[27] = in[75] & in2[75];
    assign P[27] = in[75] ^ in2[75];
    assign G[28] = in[74] & in2[74];
    assign P[28] = in[74] ^ in2[74];
    assign G[29] = in[73] & in2[73];
    assign P[29] = in[73] ^ in2[73];
    assign G[30] = in[72] & in2[72];
    assign P[30] = in[72] ^ in2[72];
    assign G[31] = in[71] & in2[71];
    assign P[31] = in[71] ^ in2[71];
    assign G[32] = in[70] & in2[70];
    assign P[32] = in[70] ^ in2[70];
    assign G[33] = in[69] & in2[69];
    assign P[33] = in[69] ^ in2[69];
    assign G[34] = in[68] & in2[68];
    assign P[34] = in[68] ^ in2[68];
    assign G[35] = in[67] & in2[67];
    assign P[35] = in[67] ^ in2[67];
    assign G[36] = in[66] & in2[66];
    assign P[36] = in[66] ^ in2[66];
    assign G[37] = in[65] & in2[65];
    assign P[37] = in[65] ^ in2[65];
    assign G[38] = in[64] & in2[64];
    assign P[38] = in[64] ^ in2[64];
    assign G[39] = in[63] & in2[63];
    assign P[39] = in[63] ^ in2[63];
    assign G[40] = in[62] & in2[62];
    assign P[40] = in[62] ^ in2[62];
    assign G[41] = in[61] & in2[61];
    assign P[41] = in[61] ^ in2[61];
    assign G[42] = in[60] & in2[60];
    assign P[42] = in[60] ^ in2[60];
    assign G[43] = in[59] & in2[59];
    assign P[43] = in[59] ^ in2[59];
    assign G[44] = in[58] & in2[58];
    assign P[44] = in[58] ^ in2[58];
    assign G[45] = in[57] & in2[57];
    assign P[45] = in[57] ^ in2[57];
    assign G[46] = in[56] & in2[56];
    assign P[46] = in[56] ^ in2[56];
    assign G[47] = in[55] & in2[55];
    assign P[47] = in[55] ^ in2[55];
    assign G[48] = in[54] & in2[54];
    assign P[48] = in[54] ^ in2[54];
    assign G[49] = in[53] & in2[53];
    assign P[49] = in[53] ^ in2[53];
    assign G[50] = in[52] & in2[52];
    assign P[50] = in[52] ^ in2[52];
    assign G[51] = in[51] & in2[51];
    assign P[51] = in[51] ^ in2[51];
    assign G[52] = in[50] & in2[50];
    assign P[52] = in[50] ^ in2[50];
    assign G[53] = in[49] & in2[49];
    assign P[53] = in[49] ^ in2[49];
    assign G[54] = in[48] & in2[48];
    assign P[54] = in[48] ^ in2[48];
    assign G[55] = in[47] & in2[47];
    assign P[55] = in[47] ^ in2[47];
    assign G[56] = in[46] & in2[46];
    assign P[56] = in[46] ^ in2[46];
    assign G[57] = in[45] & in2[45];
    assign P[57] = in[45] ^ in2[45];
    assign G[58] = in[44] & in2[44];
    assign P[58] = in[44] ^ in2[44];
    assign G[59] = in[43] & in2[43];
    assign P[59] = in[43] ^ in2[43];
    assign G[60] = in[42] & in2[42];
    assign P[60] = in[42] ^ in2[42];
    assign G[61] = in[41] & in2[41];
    assign P[61] = in[41] ^ in2[41];
    assign G[62] = in[40] & in2[40];
    assign P[62] = in[40] ^ in2[40];
    assign G[63] = in[39] & in2[39];
    assign P[63] = in[39] ^ in2[39];
    assign G[64] = in[38] & in2[38];
    assign P[64] = in[38] ^ in2[38];
    assign G[65] = in[37] & in2[37];
    assign P[65] = in[37] ^ in2[37];
    assign G[66] = in[36] & in2[36];
    assign P[66] = in[36] ^ in2[36];
    assign G[67] = in[35] & in2[35];
    assign P[67] = in[35] ^ in2[35];
    assign G[68] = in[34] & in2[34];
    assign P[68] = in[34] ^ in2[34];
    assign G[69] = in[33] & in2[33];
    assign P[69] = in[33] ^ in2[33];
    assign G[70] = in[32] & in2[32];
    assign P[70] = in[32] ^ in2[32];
    assign G[71] = in[31] & in2[31];
    assign P[71] = in[31] ^ in2[31];
    assign G[72] = in[30] & in2[30];
    assign P[72] = in[30] ^ in2[30];
    assign G[73] = in[29] & in2[29];
    assign P[73] = in[29] ^ in2[29];
    assign G[74] = in[28] & in2[28];
    assign P[74] = in[28] ^ in2[28];
    assign G[75] = in[27] & in2[27];
    assign P[75] = in[27] ^ in2[27];
    assign G[76] = in[26] & in2[26];
    assign P[76] = in[26] ^ in2[26];
    assign G[77] = in[25] & in2[25];
    assign P[77] = in[25] ^ in2[25];
    assign G[78] = in[24] & in2[24];
    assign P[78] = in[24] ^ in2[24];
    assign G[79] = in[23] & in2[23];
    assign P[79] = in[23] ^ in2[23];
    assign G[80] = in[22] & in2[22];
    assign P[80] = in[22] ^ in2[22];
    assign G[81] = in[21] & in2[21];
    assign P[81] = in[21] ^ in2[21];
    assign G[82] = in[20] & in2[20];
    assign P[82] = in[20] ^ in2[20];
    assign G[83] = in[19] & in2[19];
    assign P[83] = in[19] ^ in2[19];
    assign G[84] = in[18] & in2[18];
    assign P[84] = in[18] ^ in2[18];
    assign G[85] = in[17] & in2[17];
    assign P[85] = in[17] ^ in2[17];
    assign G[86] = in[16] & in2[16];
    assign P[86] = in[16] ^ in2[16];
    assign G[87] = in[15] & in2[15];
    assign P[87] = in[15] ^ in2[15];
    assign G[88] = in[14] & in2[14];
    assign P[88] = in[14] ^ in2[14];
    assign G[89] = in[13] & in2[13];
    assign P[89] = in[13] ^ in2[13];
    assign G[90] = in[12] & in2[12];
    assign P[90] = in[12] ^ in2[12];
    assign G[91] = in[11] & in2[11];
    assign P[91] = in[11] ^ in2[11];
    assign G[92] = in[10] & in2[10];
    assign P[92] = in[10] ^ in2[10];
    assign G[93] = in[9] & in2[9];
    assign P[93] = in[9] ^ in2[9];
    assign G[94] = in[8] & in2[8];
    assign P[94] = in[8] ^ in2[8];
    assign G[95] = in[7] & in2[7];
    assign P[95] = in[7] ^ in2[7];
    assign G[96] = in[6] & in2[6];
    assign P[96] = in[6] ^ in2[6];
    assign G[97] = in[5] & in2[5];
    assign P[97] = in[5] ^ in2[5];
    assign G[98] = in[4] & in2[4];
    assign P[98] = in[4] ^ in2[4];
    assign G[99] = in[3] & in2[3];
    assign P[99] = in[3] ^ in2[3];
    assign G[100] = in[2] & in2[2];
    assign P[100] = in[2] ^ in2[2];
    assign G[101] = in[1] & in2[1];
    assign P[101] = in[1] ^ in2[1];
    assign G[102] = in[0] & in2[0];
    assign P[102] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign C[102] = G[101] | (P[101] & C[101]);
    assign cout = G[102] | (P[102] & C[102]);
    assign sum = P ^ C;
endmodule

module CLA102(output [101:0] sum, output cout, input [101:0] in1, input [101:0] in2;

    wire[101:0] G;
    wire[101:0] C;
    wire[101:0] P;

    assign G[0] = in[101] & in2[101];
    assign P[0] = in[101] ^ in2[101];
    assign G[1] = in[100] & in2[100];
    assign P[1] = in[100] ^ in2[100];
    assign G[2] = in[99] & in2[99];
    assign P[2] = in[99] ^ in2[99];
    assign G[3] = in[98] & in2[98];
    assign P[3] = in[98] ^ in2[98];
    assign G[4] = in[97] & in2[97];
    assign P[4] = in[97] ^ in2[97];
    assign G[5] = in[96] & in2[96];
    assign P[5] = in[96] ^ in2[96];
    assign G[6] = in[95] & in2[95];
    assign P[6] = in[95] ^ in2[95];
    assign G[7] = in[94] & in2[94];
    assign P[7] = in[94] ^ in2[94];
    assign G[8] = in[93] & in2[93];
    assign P[8] = in[93] ^ in2[93];
    assign G[9] = in[92] & in2[92];
    assign P[9] = in[92] ^ in2[92];
    assign G[10] = in[91] & in2[91];
    assign P[10] = in[91] ^ in2[91];
    assign G[11] = in[90] & in2[90];
    assign P[11] = in[90] ^ in2[90];
    assign G[12] = in[89] & in2[89];
    assign P[12] = in[89] ^ in2[89];
    assign G[13] = in[88] & in2[88];
    assign P[13] = in[88] ^ in2[88];
    assign G[14] = in[87] & in2[87];
    assign P[14] = in[87] ^ in2[87];
    assign G[15] = in[86] & in2[86];
    assign P[15] = in[86] ^ in2[86];
    assign G[16] = in[85] & in2[85];
    assign P[16] = in[85] ^ in2[85];
    assign G[17] = in[84] & in2[84];
    assign P[17] = in[84] ^ in2[84];
    assign G[18] = in[83] & in2[83];
    assign P[18] = in[83] ^ in2[83];
    assign G[19] = in[82] & in2[82];
    assign P[19] = in[82] ^ in2[82];
    assign G[20] = in[81] & in2[81];
    assign P[20] = in[81] ^ in2[81];
    assign G[21] = in[80] & in2[80];
    assign P[21] = in[80] ^ in2[80];
    assign G[22] = in[79] & in2[79];
    assign P[22] = in[79] ^ in2[79];
    assign G[23] = in[78] & in2[78];
    assign P[23] = in[78] ^ in2[78];
    assign G[24] = in[77] & in2[77];
    assign P[24] = in[77] ^ in2[77];
    assign G[25] = in[76] & in2[76];
    assign P[25] = in[76] ^ in2[76];
    assign G[26] = in[75] & in2[75];
    assign P[26] = in[75] ^ in2[75];
    assign G[27] = in[74] & in2[74];
    assign P[27] = in[74] ^ in2[74];
    assign G[28] = in[73] & in2[73];
    assign P[28] = in[73] ^ in2[73];
    assign G[29] = in[72] & in2[72];
    assign P[29] = in[72] ^ in2[72];
    assign G[30] = in[71] & in2[71];
    assign P[30] = in[71] ^ in2[71];
    assign G[31] = in[70] & in2[70];
    assign P[31] = in[70] ^ in2[70];
    assign G[32] = in[69] & in2[69];
    assign P[32] = in[69] ^ in2[69];
    assign G[33] = in[68] & in2[68];
    assign P[33] = in[68] ^ in2[68];
    assign G[34] = in[67] & in2[67];
    assign P[34] = in[67] ^ in2[67];
    assign G[35] = in[66] & in2[66];
    assign P[35] = in[66] ^ in2[66];
    assign G[36] = in[65] & in2[65];
    assign P[36] = in[65] ^ in2[65];
    assign G[37] = in[64] & in2[64];
    assign P[37] = in[64] ^ in2[64];
    assign G[38] = in[63] & in2[63];
    assign P[38] = in[63] ^ in2[63];
    assign G[39] = in[62] & in2[62];
    assign P[39] = in[62] ^ in2[62];
    assign G[40] = in[61] & in2[61];
    assign P[40] = in[61] ^ in2[61];
    assign G[41] = in[60] & in2[60];
    assign P[41] = in[60] ^ in2[60];
    assign G[42] = in[59] & in2[59];
    assign P[42] = in[59] ^ in2[59];
    assign G[43] = in[58] & in2[58];
    assign P[43] = in[58] ^ in2[58];
    assign G[44] = in[57] & in2[57];
    assign P[44] = in[57] ^ in2[57];
    assign G[45] = in[56] & in2[56];
    assign P[45] = in[56] ^ in2[56];
    assign G[46] = in[55] & in2[55];
    assign P[46] = in[55] ^ in2[55];
    assign G[47] = in[54] & in2[54];
    assign P[47] = in[54] ^ in2[54];
    assign G[48] = in[53] & in2[53];
    assign P[48] = in[53] ^ in2[53];
    assign G[49] = in[52] & in2[52];
    assign P[49] = in[52] ^ in2[52];
    assign G[50] = in[51] & in2[51];
    assign P[50] = in[51] ^ in2[51];
    assign G[51] = in[50] & in2[50];
    assign P[51] = in[50] ^ in2[50];
    assign G[52] = in[49] & in2[49];
    assign P[52] = in[49] ^ in2[49];
    assign G[53] = in[48] & in2[48];
    assign P[53] = in[48] ^ in2[48];
    assign G[54] = in[47] & in2[47];
    assign P[54] = in[47] ^ in2[47];
    assign G[55] = in[46] & in2[46];
    assign P[55] = in[46] ^ in2[46];
    assign G[56] = in[45] & in2[45];
    assign P[56] = in[45] ^ in2[45];
    assign G[57] = in[44] & in2[44];
    assign P[57] = in[44] ^ in2[44];
    assign G[58] = in[43] & in2[43];
    assign P[58] = in[43] ^ in2[43];
    assign G[59] = in[42] & in2[42];
    assign P[59] = in[42] ^ in2[42];
    assign G[60] = in[41] & in2[41];
    assign P[60] = in[41] ^ in2[41];
    assign G[61] = in[40] & in2[40];
    assign P[61] = in[40] ^ in2[40];
    assign G[62] = in[39] & in2[39];
    assign P[62] = in[39] ^ in2[39];
    assign G[63] = in[38] & in2[38];
    assign P[63] = in[38] ^ in2[38];
    assign G[64] = in[37] & in2[37];
    assign P[64] = in[37] ^ in2[37];
    assign G[65] = in[36] & in2[36];
    assign P[65] = in[36] ^ in2[36];
    assign G[66] = in[35] & in2[35];
    assign P[66] = in[35] ^ in2[35];
    assign G[67] = in[34] & in2[34];
    assign P[67] = in[34] ^ in2[34];
    assign G[68] = in[33] & in2[33];
    assign P[68] = in[33] ^ in2[33];
    assign G[69] = in[32] & in2[32];
    assign P[69] = in[32] ^ in2[32];
    assign G[70] = in[31] & in2[31];
    assign P[70] = in[31] ^ in2[31];
    assign G[71] = in[30] & in2[30];
    assign P[71] = in[30] ^ in2[30];
    assign G[72] = in[29] & in2[29];
    assign P[72] = in[29] ^ in2[29];
    assign G[73] = in[28] & in2[28];
    assign P[73] = in[28] ^ in2[28];
    assign G[74] = in[27] & in2[27];
    assign P[74] = in[27] ^ in2[27];
    assign G[75] = in[26] & in2[26];
    assign P[75] = in[26] ^ in2[26];
    assign G[76] = in[25] & in2[25];
    assign P[76] = in[25] ^ in2[25];
    assign G[77] = in[24] & in2[24];
    assign P[77] = in[24] ^ in2[24];
    assign G[78] = in[23] & in2[23];
    assign P[78] = in[23] ^ in2[23];
    assign G[79] = in[22] & in2[22];
    assign P[79] = in[22] ^ in2[22];
    assign G[80] = in[21] & in2[21];
    assign P[80] = in[21] ^ in2[21];
    assign G[81] = in[20] & in2[20];
    assign P[81] = in[20] ^ in2[20];
    assign G[82] = in[19] & in2[19];
    assign P[82] = in[19] ^ in2[19];
    assign G[83] = in[18] & in2[18];
    assign P[83] = in[18] ^ in2[18];
    assign G[84] = in[17] & in2[17];
    assign P[84] = in[17] ^ in2[17];
    assign G[85] = in[16] & in2[16];
    assign P[85] = in[16] ^ in2[16];
    assign G[86] = in[15] & in2[15];
    assign P[86] = in[15] ^ in2[15];
    assign G[87] = in[14] & in2[14];
    assign P[87] = in[14] ^ in2[14];
    assign G[88] = in[13] & in2[13];
    assign P[88] = in[13] ^ in2[13];
    assign G[89] = in[12] & in2[12];
    assign P[89] = in[12] ^ in2[12];
    assign G[90] = in[11] & in2[11];
    assign P[90] = in[11] ^ in2[11];
    assign G[91] = in[10] & in2[10];
    assign P[91] = in[10] ^ in2[10];
    assign G[92] = in[9] & in2[9];
    assign P[92] = in[9] ^ in2[9];
    assign G[93] = in[8] & in2[8];
    assign P[93] = in[8] ^ in2[8];
    assign G[94] = in[7] & in2[7];
    assign P[94] = in[7] ^ in2[7];
    assign G[95] = in[6] & in2[6];
    assign P[95] = in[6] ^ in2[6];
    assign G[96] = in[5] & in2[5];
    assign P[96] = in[5] ^ in2[5];
    assign G[97] = in[4] & in2[4];
    assign P[97] = in[4] ^ in2[4];
    assign G[98] = in[3] & in2[3];
    assign P[98] = in[3] ^ in2[3];
    assign G[99] = in[2] & in2[2];
    assign P[99] = in[2] ^ in2[2];
    assign G[100] = in[1] & in2[1];
    assign P[100] = in[1] ^ in2[1];
    assign G[101] = in[0] & in2[0];
    assign P[101] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign C[101] = G[100] | (P[100] & C[100]);
    assign cout = G[101] | (P[101] & C[101]);
    assign sum = P ^ C;
endmodule

module CLA101(output [100:0] sum, output cout, input [100:0] in1, input [100:0] in2;

    wire[100:0] G;
    wire[100:0] C;
    wire[100:0] P;

    assign G[0] = in[100] & in2[100];
    assign P[0] = in[100] ^ in2[100];
    assign G[1] = in[99] & in2[99];
    assign P[1] = in[99] ^ in2[99];
    assign G[2] = in[98] & in2[98];
    assign P[2] = in[98] ^ in2[98];
    assign G[3] = in[97] & in2[97];
    assign P[3] = in[97] ^ in2[97];
    assign G[4] = in[96] & in2[96];
    assign P[4] = in[96] ^ in2[96];
    assign G[5] = in[95] & in2[95];
    assign P[5] = in[95] ^ in2[95];
    assign G[6] = in[94] & in2[94];
    assign P[6] = in[94] ^ in2[94];
    assign G[7] = in[93] & in2[93];
    assign P[7] = in[93] ^ in2[93];
    assign G[8] = in[92] & in2[92];
    assign P[8] = in[92] ^ in2[92];
    assign G[9] = in[91] & in2[91];
    assign P[9] = in[91] ^ in2[91];
    assign G[10] = in[90] & in2[90];
    assign P[10] = in[90] ^ in2[90];
    assign G[11] = in[89] & in2[89];
    assign P[11] = in[89] ^ in2[89];
    assign G[12] = in[88] & in2[88];
    assign P[12] = in[88] ^ in2[88];
    assign G[13] = in[87] & in2[87];
    assign P[13] = in[87] ^ in2[87];
    assign G[14] = in[86] & in2[86];
    assign P[14] = in[86] ^ in2[86];
    assign G[15] = in[85] & in2[85];
    assign P[15] = in[85] ^ in2[85];
    assign G[16] = in[84] & in2[84];
    assign P[16] = in[84] ^ in2[84];
    assign G[17] = in[83] & in2[83];
    assign P[17] = in[83] ^ in2[83];
    assign G[18] = in[82] & in2[82];
    assign P[18] = in[82] ^ in2[82];
    assign G[19] = in[81] & in2[81];
    assign P[19] = in[81] ^ in2[81];
    assign G[20] = in[80] & in2[80];
    assign P[20] = in[80] ^ in2[80];
    assign G[21] = in[79] & in2[79];
    assign P[21] = in[79] ^ in2[79];
    assign G[22] = in[78] & in2[78];
    assign P[22] = in[78] ^ in2[78];
    assign G[23] = in[77] & in2[77];
    assign P[23] = in[77] ^ in2[77];
    assign G[24] = in[76] & in2[76];
    assign P[24] = in[76] ^ in2[76];
    assign G[25] = in[75] & in2[75];
    assign P[25] = in[75] ^ in2[75];
    assign G[26] = in[74] & in2[74];
    assign P[26] = in[74] ^ in2[74];
    assign G[27] = in[73] & in2[73];
    assign P[27] = in[73] ^ in2[73];
    assign G[28] = in[72] & in2[72];
    assign P[28] = in[72] ^ in2[72];
    assign G[29] = in[71] & in2[71];
    assign P[29] = in[71] ^ in2[71];
    assign G[30] = in[70] & in2[70];
    assign P[30] = in[70] ^ in2[70];
    assign G[31] = in[69] & in2[69];
    assign P[31] = in[69] ^ in2[69];
    assign G[32] = in[68] & in2[68];
    assign P[32] = in[68] ^ in2[68];
    assign G[33] = in[67] & in2[67];
    assign P[33] = in[67] ^ in2[67];
    assign G[34] = in[66] & in2[66];
    assign P[34] = in[66] ^ in2[66];
    assign G[35] = in[65] & in2[65];
    assign P[35] = in[65] ^ in2[65];
    assign G[36] = in[64] & in2[64];
    assign P[36] = in[64] ^ in2[64];
    assign G[37] = in[63] & in2[63];
    assign P[37] = in[63] ^ in2[63];
    assign G[38] = in[62] & in2[62];
    assign P[38] = in[62] ^ in2[62];
    assign G[39] = in[61] & in2[61];
    assign P[39] = in[61] ^ in2[61];
    assign G[40] = in[60] & in2[60];
    assign P[40] = in[60] ^ in2[60];
    assign G[41] = in[59] & in2[59];
    assign P[41] = in[59] ^ in2[59];
    assign G[42] = in[58] & in2[58];
    assign P[42] = in[58] ^ in2[58];
    assign G[43] = in[57] & in2[57];
    assign P[43] = in[57] ^ in2[57];
    assign G[44] = in[56] & in2[56];
    assign P[44] = in[56] ^ in2[56];
    assign G[45] = in[55] & in2[55];
    assign P[45] = in[55] ^ in2[55];
    assign G[46] = in[54] & in2[54];
    assign P[46] = in[54] ^ in2[54];
    assign G[47] = in[53] & in2[53];
    assign P[47] = in[53] ^ in2[53];
    assign G[48] = in[52] & in2[52];
    assign P[48] = in[52] ^ in2[52];
    assign G[49] = in[51] & in2[51];
    assign P[49] = in[51] ^ in2[51];
    assign G[50] = in[50] & in2[50];
    assign P[50] = in[50] ^ in2[50];
    assign G[51] = in[49] & in2[49];
    assign P[51] = in[49] ^ in2[49];
    assign G[52] = in[48] & in2[48];
    assign P[52] = in[48] ^ in2[48];
    assign G[53] = in[47] & in2[47];
    assign P[53] = in[47] ^ in2[47];
    assign G[54] = in[46] & in2[46];
    assign P[54] = in[46] ^ in2[46];
    assign G[55] = in[45] & in2[45];
    assign P[55] = in[45] ^ in2[45];
    assign G[56] = in[44] & in2[44];
    assign P[56] = in[44] ^ in2[44];
    assign G[57] = in[43] & in2[43];
    assign P[57] = in[43] ^ in2[43];
    assign G[58] = in[42] & in2[42];
    assign P[58] = in[42] ^ in2[42];
    assign G[59] = in[41] & in2[41];
    assign P[59] = in[41] ^ in2[41];
    assign G[60] = in[40] & in2[40];
    assign P[60] = in[40] ^ in2[40];
    assign G[61] = in[39] & in2[39];
    assign P[61] = in[39] ^ in2[39];
    assign G[62] = in[38] & in2[38];
    assign P[62] = in[38] ^ in2[38];
    assign G[63] = in[37] & in2[37];
    assign P[63] = in[37] ^ in2[37];
    assign G[64] = in[36] & in2[36];
    assign P[64] = in[36] ^ in2[36];
    assign G[65] = in[35] & in2[35];
    assign P[65] = in[35] ^ in2[35];
    assign G[66] = in[34] & in2[34];
    assign P[66] = in[34] ^ in2[34];
    assign G[67] = in[33] & in2[33];
    assign P[67] = in[33] ^ in2[33];
    assign G[68] = in[32] & in2[32];
    assign P[68] = in[32] ^ in2[32];
    assign G[69] = in[31] & in2[31];
    assign P[69] = in[31] ^ in2[31];
    assign G[70] = in[30] & in2[30];
    assign P[70] = in[30] ^ in2[30];
    assign G[71] = in[29] & in2[29];
    assign P[71] = in[29] ^ in2[29];
    assign G[72] = in[28] & in2[28];
    assign P[72] = in[28] ^ in2[28];
    assign G[73] = in[27] & in2[27];
    assign P[73] = in[27] ^ in2[27];
    assign G[74] = in[26] & in2[26];
    assign P[74] = in[26] ^ in2[26];
    assign G[75] = in[25] & in2[25];
    assign P[75] = in[25] ^ in2[25];
    assign G[76] = in[24] & in2[24];
    assign P[76] = in[24] ^ in2[24];
    assign G[77] = in[23] & in2[23];
    assign P[77] = in[23] ^ in2[23];
    assign G[78] = in[22] & in2[22];
    assign P[78] = in[22] ^ in2[22];
    assign G[79] = in[21] & in2[21];
    assign P[79] = in[21] ^ in2[21];
    assign G[80] = in[20] & in2[20];
    assign P[80] = in[20] ^ in2[20];
    assign G[81] = in[19] & in2[19];
    assign P[81] = in[19] ^ in2[19];
    assign G[82] = in[18] & in2[18];
    assign P[82] = in[18] ^ in2[18];
    assign G[83] = in[17] & in2[17];
    assign P[83] = in[17] ^ in2[17];
    assign G[84] = in[16] & in2[16];
    assign P[84] = in[16] ^ in2[16];
    assign G[85] = in[15] & in2[15];
    assign P[85] = in[15] ^ in2[15];
    assign G[86] = in[14] & in2[14];
    assign P[86] = in[14] ^ in2[14];
    assign G[87] = in[13] & in2[13];
    assign P[87] = in[13] ^ in2[13];
    assign G[88] = in[12] & in2[12];
    assign P[88] = in[12] ^ in2[12];
    assign G[89] = in[11] & in2[11];
    assign P[89] = in[11] ^ in2[11];
    assign G[90] = in[10] & in2[10];
    assign P[90] = in[10] ^ in2[10];
    assign G[91] = in[9] & in2[9];
    assign P[91] = in[9] ^ in2[9];
    assign G[92] = in[8] & in2[8];
    assign P[92] = in[8] ^ in2[8];
    assign G[93] = in[7] & in2[7];
    assign P[93] = in[7] ^ in2[7];
    assign G[94] = in[6] & in2[6];
    assign P[94] = in[6] ^ in2[6];
    assign G[95] = in[5] & in2[5];
    assign P[95] = in[5] ^ in2[5];
    assign G[96] = in[4] & in2[4];
    assign P[96] = in[4] ^ in2[4];
    assign G[97] = in[3] & in2[3];
    assign P[97] = in[3] ^ in2[3];
    assign G[98] = in[2] & in2[2];
    assign P[98] = in[2] ^ in2[2];
    assign G[99] = in[1] & in2[1];
    assign P[99] = in[1] ^ in2[1];
    assign G[100] = in[0] & in2[0];
    assign P[100] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign C[100] = G[99] | (P[99] & C[99]);
    assign cout = G[100] | (P[100] & C[100]);
    assign sum = P ^ C;
endmodule

module CLA100(output [99:0] sum, output cout, input [99:0] in1, input [99:0] in2;

    wire[99:0] G;
    wire[99:0] C;
    wire[99:0] P;

    assign G[0] = in[99] & in2[99];
    assign P[0] = in[99] ^ in2[99];
    assign G[1] = in[98] & in2[98];
    assign P[1] = in[98] ^ in2[98];
    assign G[2] = in[97] & in2[97];
    assign P[2] = in[97] ^ in2[97];
    assign G[3] = in[96] & in2[96];
    assign P[3] = in[96] ^ in2[96];
    assign G[4] = in[95] & in2[95];
    assign P[4] = in[95] ^ in2[95];
    assign G[5] = in[94] & in2[94];
    assign P[5] = in[94] ^ in2[94];
    assign G[6] = in[93] & in2[93];
    assign P[6] = in[93] ^ in2[93];
    assign G[7] = in[92] & in2[92];
    assign P[7] = in[92] ^ in2[92];
    assign G[8] = in[91] & in2[91];
    assign P[8] = in[91] ^ in2[91];
    assign G[9] = in[90] & in2[90];
    assign P[9] = in[90] ^ in2[90];
    assign G[10] = in[89] & in2[89];
    assign P[10] = in[89] ^ in2[89];
    assign G[11] = in[88] & in2[88];
    assign P[11] = in[88] ^ in2[88];
    assign G[12] = in[87] & in2[87];
    assign P[12] = in[87] ^ in2[87];
    assign G[13] = in[86] & in2[86];
    assign P[13] = in[86] ^ in2[86];
    assign G[14] = in[85] & in2[85];
    assign P[14] = in[85] ^ in2[85];
    assign G[15] = in[84] & in2[84];
    assign P[15] = in[84] ^ in2[84];
    assign G[16] = in[83] & in2[83];
    assign P[16] = in[83] ^ in2[83];
    assign G[17] = in[82] & in2[82];
    assign P[17] = in[82] ^ in2[82];
    assign G[18] = in[81] & in2[81];
    assign P[18] = in[81] ^ in2[81];
    assign G[19] = in[80] & in2[80];
    assign P[19] = in[80] ^ in2[80];
    assign G[20] = in[79] & in2[79];
    assign P[20] = in[79] ^ in2[79];
    assign G[21] = in[78] & in2[78];
    assign P[21] = in[78] ^ in2[78];
    assign G[22] = in[77] & in2[77];
    assign P[22] = in[77] ^ in2[77];
    assign G[23] = in[76] & in2[76];
    assign P[23] = in[76] ^ in2[76];
    assign G[24] = in[75] & in2[75];
    assign P[24] = in[75] ^ in2[75];
    assign G[25] = in[74] & in2[74];
    assign P[25] = in[74] ^ in2[74];
    assign G[26] = in[73] & in2[73];
    assign P[26] = in[73] ^ in2[73];
    assign G[27] = in[72] & in2[72];
    assign P[27] = in[72] ^ in2[72];
    assign G[28] = in[71] & in2[71];
    assign P[28] = in[71] ^ in2[71];
    assign G[29] = in[70] & in2[70];
    assign P[29] = in[70] ^ in2[70];
    assign G[30] = in[69] & in2[69];
    assign P[30] = in[69] ^ in2[69];
    assign G[31] = in[68] & in2[68];
    assign P[31] = in[68] ^ in2[68];
    assign G[32] = in[67] & in2[67];
    assign P[32] = in[67] ^ in2[67];
    assign G[33] = in[66] & in2[66];
    assign P[33] = in[66] ^ in2[66];
    assign G[34] = in[65] & in2[65];
    assign P[34] = in[65] ^ in2[65];
    assign G[35] = in[64] & in2[64];
    assign P[35] = in[64] ^ in2[64];
    assign G[36] = in[63] & in2[63];
    assign P[36] = in[63] ^ in2[63];
    assign G[37] = in[62] & in2[62];
    assign P[37] = in[62] ^ in2[62];
    assign G[38] = in[61] & in2[61];
    assign P[38] = in[61] ^ in2[61];
    assign G[39] = in[60] & in2[60];
    assign P[39] = in[60] ^ in2[60];
    assign G[40] = in[59] & in2[59];
    assign P[40] = in[59] ^ in2[59];
    assign G[41] = in[58] & in2[58];
    assign P[41] = in[58] ^ in2[58];
    assign G[42] = in[57] & in2[57];
    assign P[42] = in[57] ^ in2[57];
    assign G[43] = in[56] & in2[56];
    assign P[43] = in[56] ^ in2[56];
    assign G[44] = in[55] & in2[55];
    assign P[44] = in[55] ^ in2[55];
    assign G[45] = in[54] & in2[54];
    assign P[45] = in[54] ^ in2[54];
    assign G[46] = in[53] & in2[53];
    assign P[46] = in[53] ^ in2[53];
    assign G[47] = in[52] & in2[52];
    assign P[47] = in[52] ^ in2[52];
    assign G[48] = in[51] & in2[51];
    assign P[48] = in[51] ^ in2[51];
    assign G[49] = in[50] & in2[50];
    assign P[49] = in[50] ^ in2[50];
    assign G[50] = in[49] & in2[49];
    assign P[50] = in[49] ^ in2[49];
    assign G[51] = in[48] & in2[48];
    assign P[51] = in[48] ^ in2[48];
    assign G[52] = in[47] & in2[47];
    assign P[52] = in[47] ^ in2[47];
    assign G[53] = in[46] & in2[46];
    assign P[53] = in[46] ^ in2[46];
    assign G[54] = in[45] & in2[45];
    assign P[54] = in[45] ^ in2[45];
    assign G[55] = in[44] & in2[44];
    assign P[55] = in[44] ^ in2[44];
    assign G[56] = in[43] & in2[43];
    assign P[56] = in[43] ^ in2[43];
    assign G[57] = in[42] & in2[42];
    assign P[57] = in[42] ^ in2[42];
    assign G[58] = in[41] & in2[41];
    assign P[58] = in[41] ^ in2[41];
    assign G[59] = in[40] & in2[40];
    assign P[59] = in[40] ^ in2[40];
    assign G[60] = in[39] & in2[39];
    assign P[60] = in[39] ^ in2[39];
    assign G[61] = in[38] & in2[38];
    assign P[61] = in[38] ^ in2[38];
    assign G[62] = in[37] & in2[37];
    assign P[62] = in[37] ^ in2[37];
    assign G[63] = in[36] & in2[36];
    assign P[63] = in[36] ^ in2[36];
    assign G[64] = in[35] & in2[35];
    assign P[64] = in[35] ^ in2[35];
    assign G[65] = in[34] & in2[34];
    assign P[65] = in[34] ^ in2[34];
    assign G[66] = in[33] & in2[33];
    assign P[66] = in[33] ^ in2[33];
    assign G[67] = in[32] & in2[32];
    assign P[67] = in[32] ^ in2[32];
    assign G[68] = in[31] & in2[31];
    assign P[68] = in[31] ^ in2[31];
    assign G[69] = in[30] & in2[30];
    assign P[69] = in[30] ^ in2[30];
    assign G[70] = in[29] & in2[29];
    assign P[70] = in[29] ^ in2[29];
    assign G[71] = in[28] & in2[28];
    assign P[71] = in[28] ^ in2[28];
    assign G[72] = in[27] & in2[27];
    assign P[72] = in[27] ^ in2[27];
    assign G[73] = in[26] & in2[26];
    assign P[73] = in[26] ^ in2[26];
    assign G[74] = in[25] & in2[25];
    assign P[74] = in[25] ^ in2[25];
    assign G[75] = in[24] & in2[24];
    assign P[75] = in[24] ^ in2[24];
    assign G[76] = in[23] & in2[23];
    assign P[76] = in[23] ^ in2[23];
    assign G[77] = in[22] & in2[22];
    assign P[77] = in[22] ^ in2[22];
    assign G[78] = in[21] & in2[21];
    assign P[78] = in[21] ^ in2[21];
    assign G[79] = in[20] & in2[20];
    assign P[79] = in[20] ^ in2[20];
    assign G[80] = in[19] & in2[19];
    assign P[80] = in[19] ^ in2[19];
    assign G[81] = in[18] & in2[18];
    assign P[81] = in[18] ^ in2[18];
    assign G[82] = in[17] & in2[17];
    assign P[82] = in[17] ^ in2[17];
    assign G[83] = in[16] & in2[16];
    assign P[83] = in[16] ^ in2[16];
    assign G[84] = in[15] & in2[15];
    assign P[84] = in[15] ^ in2[15];
    assign G[85] = in[14] & in2[14];
    assign P[85] = in[14] ^ in2[14];
    assign G[86] = in[13] & in2[13];
    assign P[86] = in[13] ^ in2[13];
    assign G[87] = in[12] & in2[12];
    assign P[87] = in[12] ^ in2[12];
    assign G[88] = in[11] & in2[11];
    assign P[88] = in[11] ^ in2[11];
    assign G[89] = in[10] & in2[10];
    assign P[89] = in[10] ^ in2[10];
    assign G[90] = in[9] & in2[9];
    assign P[90] = in[9] ^ in2[9];
    assign G[91] = in[8] & in2[8];
    assign P[91] = in[8] ^ in2[8];
    assign G[92] = in[7] & in2[7];
    assign P[92] = in[7] ^ in2[7];
    assign G[93] = in[6] & in2[6];
    assign P[93] = in[6] ^ in2[6];
    assign G[94] = in[5] & in2[5];
    assign P[94] = in[5] ^ in2[5];
    assign G[95] = in[4] & in2[4];
    assign P[95] = in[4] ^ in2[4];
    assign G[96] = in[3] & in2[3];
    assign P[96] = in[3] ^ in2[3];
    assign G[97] = in[2] & in2[2];
    assign P[97] = in[2] ^ in2[2];
    assign G[98] = in[1] & in2[1];
    assign P[98] = in[1] ^ in2[1];
    assign G[99] = in[0] & in2[0];
    assign P[99] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign C[99] = G[98] | (P[98] & C[98]);
    assign cout = G[99] | (P[99] & C[99]);
    assign sum = P ^ C;
endmodule

module CLA99(output [98:0] sum, output cout, input [98:0] in1, input [98:0] in2;

    wire[98:0] G;
    wire[98:0] C;
    wire[98:0] P;

    assign G[0] = in[98] & in2[98];
    assign P[0] = in[98] ^ in2[98];
    assign G[1] = in[97] & in2[97];
    assign P[1] = in[97] ^ in2[97];
    assign G[2] = in[96] & in2[96];
    assign P[2] = in[96] ^ in2[96];
    assign G[3] = in[95] & in2[95];
    assign P[3] = in[95] ^ in2[95];
    assign G[4] = in[94] & in2[94];
    assign P[4] = in[94] ^ in2[94];
    assign G[5] = in[93] & in2[93];
    assign P[5] = in[93] ^ in2[93];
    assign G[6] = in[92] & in2[92];
    assign P[6] = in[92] ^ in2[92];
    assign G[7] = in[91] & in2[91];
    assign P[7] = in[91] ^ in2[91];
    assign G[8] = in[90] & in2[90];
    assign P[8] = in[90] ^ in2[90];
    assign G[9] = in[89] & in2[89];
    assign P[9] = in[89] ^ in2[89];
    assign G[10] = in[88] & in2[88];
    assign P[10] = in[88] ^ in2[88];
    assign G[11] = in[87] & in2[87];
    assign P[11] = in[87] ^ in2[87];
    assign G[12] = in[86] & in2[86];
    assign P[12] = in[86] ^ in2[86];
    assign G[13] = in[85] & in2[85];
    assign P[13] = in[85] ^ in2[85];
    assign G[14] = in[84] & in2[84];
    assign P[14] = in[84] ^ in2[84];
    assign G[15] = in[83] & in2[83];
    assign P[15] = in[83] ^ in2[83];
    assign G[16] = in[82] & in2[82];
    assign P[16] = in[82] ^ in2[82];
    assign G[17] = in[81] & in2[81];
    assign P[17] = in[81] ^ in2[81];
    assign G[18] = in[80] & in2[80];
    assign P[18] = in[80] ^ in2[80];
    assign G[19] = in[79] & in2[79];
    assign P[19] = in[79] ^ in2[79];
    assign G[20] = in[78] & in2[78];
    assign P[20] = in[78] ^ in2[78];
    assign G[21] = in[77] & in2[77];
    assign P[21] = in[77] ^ in2[77];
    assign G[22] = in[76] & in2[76];
    assign P[22] = in[76] ^ in2[76];
    assign G[23] = in[75] & in2[75];
    assign P[23] = in[75] ^ in2[75];
    assign G[24] = in[74] & in2[74];
    assign P[24] = in[74] ^ in2[74];
    assign G[25] = in[73] & in2[73];
    assign P[25] = in[73] ^ in2[73];
    assign G[26] = in[72] & in2[72];
    assign P[26] = in[72] ^ in2[72];
    assign G[27] = in[71] & in2[71];
    assign P[27] = in[71] ^ in2[71];
    assign G[28] = in[70] & in2[70];
    assign P[28] = in[70] ^ in2[70];
    assign G[29] = in[69] & in2[69];
    assign P[29] = in[69] ^ in2[69];
    assign G[30] = in[68] & in2[68];
    assign P[30] = in[68] ^ in2[68];
    assign G[31] = in[67] & in2[67];
    assign P[31] = in[67] ^ in2[67];
    assign G[32] = in[66] & in2[66];
    assign P[32] = in[66] ^ in2[66];
    assign G[33] = in[65] & in2[65];
    assign P[33] = in[65] ^ in2[65];
    assign G[34] = in[64] & in2[64];
    assign P[34] = in[64] ^ in2[64];
    assign G[35] = in[63] & in2[63];
    assign P[35] = in[63] ^ in2[63];
    assign G[36] = in[62] & in2[62];
    assign P[36] = in[62] ^ in2[62];
    assign G[37] = in[61] & in2[61];
    assign P[37] = in[61] ^ in2[61];
    assign G[38] = in[60] & in2[60];
    assign P[38] = in[60] ^ in2[60];
    assign G[39] = in[59] & in2[59];
    assign P[39] = in[59] ^ in2[59];
    assign G[40] = in[58] & in2[58];
    assign P[40] = in[58] ^ in2[58];
    assign G[41] = in[57] & in2[57];
    assign P[41] = in[57] ^ in2[57];
    assign G[42] = in[56] & in2[56];
    assign P[42] = in[56] ^ in2[56];
    assign G[43] = in[55] & in2[55];
    assign P[43] = in[55] ^ in2[55];
    assign G[44] = in[54] & in2[54];
    assign P[44] = in[54] ^ in2[54];
    assign G[45] = in[53] & in2[53];
    assign P[45] = in[53] ^ in2[53];
    assign G[46] = in[52] & in2[52];
    assign P[46] = in[52] ^ in2[52];
    assign G[47] = in[51] & in2[51];
    assign P[47] = in[51] ^ in2[51];
    assign G[48] = in[50] & in2[50];
    assign P[48] = in[50] ^ in2[50];
    assign G[49] = in[49] & in2[49];
    assign P[49] = in[49] ^ in2[49];
    assign G[50] = in[48] & in2[48];
    assign P[50] = in[48] ^ in2[48];
    assign G[51] = in[47] & in2[47];
    assign P[51] = in[47] ^ in2[47];
    assign G[52] = in[46] & in2[46];
    assign P[52] = in[46] ^ in2[46];
    assign G[53] = in[45] & in2[45];
    assign P[53] = in[45] ^ in2[45];
    assign G[54] = in[44] & in2[44];
    assign P[54] = in[44] ^ in2[44];
    assign G[55] = in[43] & in2[43];
    assign P[55] = in[43] ^ in2[43];
    assign G[56] = in[42] & in2[42];
    assign P[56] = in[42] ^ in2[42];
    assign G[57] = in[41] & in2[41];
    assign P[57] = in[41] ^ in2[41];
    assign G[58] = in[40] & in2[40];
    assign P[58] = in[40] ^ in2[40];
    assign G[59] = in[39] & in2[39];
    assign P[59] = in[39] ^ in2[39];
    assign G[60] = in[38] & in2[38];
    assign P[60] = in[38] ^ in2[38];
    assign G[61] = in[37] & in2[37];
    assign P[61] = in[37] ^ in2[37];
    assign G[62] = in[36] & in2[36];
    assign P[62] = in[36] ^ in2[36];
    assign G[63] = in[35] & in2[35];
    assign P[63] = in[35] ^ in2[35];
    assign G[64] = in[34] & in2[34];
    assign P[64] = in[34] ^ in2[34];
    assign G[65] = in[33] & in2[33];
    assign P[65] = in[33] ^ in2[33];
    assign G[66] = in[32] & in2[32];
    assign P[66] = in[32] ^ in2[32];
    assign G[67] = in[31] & in2[31];
    assign P[67] = in[31] ^ in2[31];
    assign G[68] = in[30] & in2[30];
    assign P[68] = in[30] ^ in2[30];
    assign G[69] = in[29] & in2[29];
    assign P[69] = in[29] ^ in2[29];
    assign G[70] = in[28] & in2[28];
    assign P[70] = in[28] ^ in2[28];
    assign G[71] = in[27] & in2[27];
    assign P[71] = in[27] ^ in2[27];
    assign G[72] = in[26] & in2[26];
    assign P[72] = in[26] ^ in2[26];
    assign G[73] = in[25] & in2[25];
    assign P[73] = in[25] ^ in2[25];
    assign G[74] = in[24] & in2[24];
    assign P[74] = in[24] ^ in2[24];
    assign G[75] = in[23] & in2[23];
    assign P[75] = in[23] ^ in2[23];
    assign G[76] = in[22] & in2[22];
    assign P[76] = in[22] ^ in2[22];
    assign G[77] = in[21] & in2[21];
    assign P[77] = in[21] ^ in2[21];
    assign G[78] = in[20] & in2[20];
    assign P[78] = in[20] ^ in2[20];
    assign G[79] = in[19] & in2[19];
    assign P[79] = in[19] ^ in2[19];
    assign G[80] = in[18] & in2[18];
    assign P[80] = in[18] ^ in2[18];
    assign G[81] = in[17] & in2[17];
    assign P[81] = in[17] ^ in2[17];
    assign G[82] = in[16] & in2[16];
    assign P[82] = in[16] ^ in2[16];
    assign G[83] = in[15] & in2[15];
    assign P[83] = in[15] ^ in2[15];
    assign G[84] = in[14] & in2[14];
    assign P[84] = in[14] ^ in2[14];
    assign G[85] = in[13] & in2[13];
    assign P[85] = in[13] ^ in2[13];
    assign G[86] = in[12] & in2[12];
    assign P[86] = in[12] ^ in2[12];
    assign G[87] = in[11] & in2[11];
    assign P[87] = in[11] ^ in2[11];
    assign G[88] = in[10] & in2[10];
    assign P[88] = in[10] ^ in2[10];
    assign G[89] = in[9] & in2[9];
    assign P[89] = in[9] ^ in2[9];
    assign G[90] = in[8] & in2[8];
    assign P[90] = in[8] ^ in2[8];
    assign G[91] = in[7] & in2[7];
    assign P[91] = in[7] ^ in2[7];
    assign G[92] = in[6] & in2[6];
    assign P[92] = in[6] ^ in2[6];
    assign G[93] = in[5] & in2[5];
    assign P[93] = in[5] ^ in2[5];
    assign G[94] = in[4] & in2[4];
    assign P[94] = in[4] ^ in2[4];
    assign G[95] = in[3] & in2[3];
    assign P[95] = in[3] ^ in2[3];
    assign G[96] = in[2] & in2[2];
    assign P[96] = in[2] ^ in2[2];
    assign G[97] = in[1] & in2[1];
    assign P[97] = in[1] ^ in2[1];
    assign G[98] = in[0] & in2[0];
    assign P[98] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign C[98] = G[97] | (P[97] & C[97]);
    assign cout = G[98] | (P[98] & C[98]);
    assign sum = P ^ C;
endmodule

module CLA98(output [97:0] sum, output cout, input [97:0] in1, input [97:0] in2;

    wire[97:0] G;
    wire[97:0] C;
    wire[97:0] P;

    assign G[0] = in[97] & in2[97];
    assign P[0] = in[97] ^ in2[97];
    assign G[1] = in[96] & in2[96];
    assign P[1] = in[96] ^ in2[96];
    assign G[2] = in[95] & in2[95];
    assign P[2] = in[95] ^ in2[95];
    assign G[3] = in[94] & in2[94];
    assign P[3] = in[94] ^ in2[94];
    assign G[4] = in[93] & in2[93];
    assign P[4] = in[93] ^ in2[93];
    assign G[5] = in[92] & in2[92];
    assign P[5] = in[92] ^ in2[92];
    assign G[6] = in[91] & in2[91];
    assign P[6] = in[91] ^ in2[91];
    assign G[7] = in[90] & in2[90];
    assign P[7] = in[90] ^ in2[90];
    assign G[8] = in[89] & in2[89];
    assign P[8] = in[89] ^ in2[89];
    assign G[9] = in[88] & in2[88];
    assign P[9] = in[88] ^ in2[88];
    assign G[10] = in[87] & in2[87];
    assign P[10] = in[87] ^ in2[87];
    assign G[11] = in[86] & in2[86];
    assign P[11] = in[86] ^ in2[86];
    assign G[12] = in[85] & in2[85];
    assign P[12] = in[85] ^ in2[85];
    assign G[13] = in[84] & in2[84];
    assign P[13] = in[84] ^ in2[84];
    assign G[14] = in[83] & in2[83];
    assign P[14] = in[83] ^ in2[83];
    assign G[15] = in[82] & in2[82];
    assign P[15] = in[82] ^ in2[82];
    assign G[16] = in[81] & in2[81];
    assign P[16] = in[81] ^ in2[81];
    assign G[17] = in[80] & in2[80];
    assign P[17] = in[80] ^ in2[80];
    assign G[18] = in[79] & in2[79];
    assign P[18] = in[79] ^ in2[79];
    assign G[19] = in[78] & in2[78];
    assign P[19] = in[78] ^ in2[78];
    assign G[20] = in[77] & in2[77];
    assign P[20] = in[77] ^ in2[77];
    assign G[21] = in[76] & in2[76];
    assign P[21] = in[76] ^ in2[76];
    assign G[22] = in[75] & in2[75];
    assign P[22] = in[75] ^ in2[75];
    assign G[23] = in[74] & in2[74];
    assign P[23] = in[74] ^ in2[74];
    assign G[24] = in[73] & in2[73];
    assign P[24] = in[73] ^ in2[73];
    assign G[25] = in[72] & in2[72];
    assign P[25] = in[72] ^ in2[72];
    assign G[26] = in[71] & in2[71];
    assign P[26] = in[71] ^ in2[71];
    assign G[27] = in[70] & in2[70];
    assign P[27] = in[70] ^ in2[70];
    assign G[28] = in[69] & in2[69];
    assign P[28] = in[69] ^ in2[69];
    assign G[29] = in[68] & in2[68];
    assign P[29] = in[68] ^ in2[68];
    assign G[30] = in[67] & in2[67];
    assign P[30] = in[67] ^ in2[67];
    assign G[31] = in[66] & in2[66];
    assign P[31] = in[66] ^ in2[66];
    assign G[32] = in[65] & in2[65];
    assign P[32] = in[65] ^ in2[65];
    assign G[33] = in[64] & in2[64];
    assign P[33] = in[64] ^ in2[64];
    assign G[34] = in[63] & in2[63];
    assign P[34] = in[63] ^ in2[63];
    assign G[35] = in[62] & in2[62];
    assign P[35] = in[62] ^ in2[62];
    assign G[36] = in[61] & in2[61];
    assign P[36] = in[61] ^ in2[61];
    assign G[37] = in[60] & in2[60];
    assign P[37] = in[60] ^ in2[60];
    assign G[38] = in[59] & in2[59];
    assign P[38] = in[59] ^ in2[59];
    assign G[39] = in[58] & in2[58];
    assign P[39] = in[58] ^ in2[58];
    assign G[40] = in[57] & in2[57];
    assign P[40] = in[57] ^ in2[57];
    assign G[41] = in[56] & in2[56];
    assign P[41] = in[56] ^ in2[56];
    assign G[42] = in[55] & in2[55];
    assign P[42] = in[55] ^ in2[55];
    assign G[43] = in[54] & in2[54];
    assign P[43] = in[54] ^ in2[54];
    assign G[44] = in[53] & in2[53];
    assign P[44] = in[53] ^ in2[53];
    assign G[45] = in[52] & in2[52];
    assign P[45] = in[52] ^ in2[52];
    assign G[46] = in[51] & in2[51];
    assign P[46] = in[51] ^ in2[51];
    assign G[47] = in[50] & in2[50];
    assign P[47] = in[50] ^ in2[50];
    assign G[48] = in[49] & in2[49];
    assign P[48] = in[49] ^ in2[49];
    assign G[49] = in[48] & in2[48];
    assign P[49] = in[48] ^ in2[48];
    assign G[50] = in[47] & in2[47];
    assign P[50] = in[47] ^ in2[47];
    assign G[51] = in[46] & in2[46];
    assign P[51] = in[46] ^ in2[46];
    assign G[52] = in[45] & in2[45];
    assign P[52] = in[45] ^ in2[45];
    assign G[53] = in[44] & in2[44];
    assign P[53] = in[44] ^ in2[44];
    assign G[54] = in[43] & in2[43];
    assign P[54] = in[43] ^ in2[43];
    assign G[55] = in[42] & in2[42];
    assign P[55] = in[42] ^ in2[42];
    assign G[56] = in[41] & in2[41];
    assign P[56] = in[41] ^ in2[41];
    assign G[57] = in[40] & in2[40];
    assign P[57] = in[40] ^ in2[40];
    assign G[58] = in[39] & in2[39];
    assign P[58] = in[39] ^ in2[39];
    assign G[59] = in[38] & in2[38];
    assign P[59] = in[38] ^ in2[38];
    assign G[60] = in[37] & in2[37];
    assign P[60] = in[37] ^ in2[37];
    assign G[61] = in[36] & in2[36];
    assign P[61] = in[36] ^ in2[36];
    assign G[62] = in[35] & in2[35];
    assign P[62] = in[35] ^ in2[35];
    assign G[63] = in[34] & in2[34];
    assign P[63] = in[34] ^ in2[34];
    assign G[64] = in[33] & in2[33];
    assign P[64] = in[33] ^ in2[33];
    assign G[65] = in[32] & in2[32];
    assign P[65] = in[32] ^ in2[32];
    assign G[66] = in[31] & in2[31];
    assign P[66] = in[31] ^ in2[31];
    assign G[67] = in[30] & in2[30];
    assign P[67] = in[30] ^ in2[30];
    assign G[68] = in[29] & in2[29];
    assign P[68] = in[29] ^ in2[29];
    assign G[69] = in[28] & in2[28];
    assign P[69] = in[28] ^ in2[28];
    assign G[70] = in[27] & in2[27];
    assign P[70] = in[27] ^ in2[27];
    assign G[71] = in[26] & in2[26];
    assign P[71] = in[26] ^ in2[26];
    assign G[72] = in[25] & in2[25];
    assign P[72] = in[25] ^ in2[25];
    assign G[73] = in[24] & in2[24];
    assign P[73] = in[24] ^ in2[24];
    assign G[74] = in[23] & in2[23];
    assign P[74] = in[23] ^ in2[23];
    assign G[75] = in[22] & in2[22];
    assign P[75] = in[22] ^ in2[22];
    assign G[76] = in[21] & in2[21];
    assign P[76] = in[21] ^ in2[21];
    assign G[77] = in[20] & in2[20];
    assign P[77] = in[20] ^ in2[20];
    assign G[78] = in[19] & in2[19];
    assign P[78] = in[19] ^ in2[19];
    assign G[79] = in[18] & in2[18];
    assign P[79] = in[18] ^ in2[18];
    assign G[80] = in[17] & in2[17];
    assign P[80] = in[17] ^ in2[17];
    assign G[81] = in[16] & in2[16];
    assign P[81] = in[16] ^ in2[16];
    assign G[82] = in[15] & in2[15];
    assign P[82] = in[15] ^ in2[15];
    assign G[83] = in[14] & in2[14];
    assign P[83] = in[14] ^ in2[14];
    assign G[84] = in[13] & in2[13];
    assign P[84] = in[13] ^ in2[13];
    assign G[85] = in[12] & in2[12];
    assign P[85] = in[12] ^ in2[12];
    assign G[86] = in[11] & in2[11];
    assign P[86] = in[11] ^ in2[11];
    assign G[87] = in[10] & in2[10];
    assign P[87] = in[10] ^ in2[10];
    assign G[88] = in[9] & in2[9];
    assign P[88] = in[9] ^ in2[9];
    assign G[89] = in[8] & in2[8];
    assign P[89] = in[8] ^ in2[8];
    assign G[90] = in[7] & in2[7];
    assign P[90] = in[7] ^ in2[7];
    assign G[91] = in[6] & in2[6];
    assign P[91] = in[6] ^ in2[6];
    assign G[92] = in[5] & in2[5];
    assign P[92] = in[5] ^ in2[5];
    assign G[93] = in[4] & in2[4];
    assign P[93] = in[4] ^ in2[4];
    assign G[94] = in[3] & in2[3];
    assign P[94] = in[3] ^ in2[3];
    assign G[95] = in[2] & in2[2];
    assign P[95] = in[2] ^ in2[2];
    assign G[96] = in[1] & in2[1];
    assign P[96] = in[1] ^ in2[1];
    assign G[97] = in[0] & in2[0];
    assign P[97] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign C[97] = G[96] | (P[96] & C[96]);
    assign cout = G[97] | (P[97] & C[97]);
    assign sum = P ^ C;
endmodule

module CLA97(output [96:0] sum, output cout, input [96:0] in1, input [96:0] in2;

    wire[96:0] G;
    wire[96:0] C;
    wire[96:0] P;

    assign G[0] = in[96] & in2[96];
    assign P[0] = in[96] ^ in2[96];
    assign G[1] = in[95] & in2[95];
    assign P[1] = in[95] ^ in2[95];
    assign G[2] = in[94] & in2[94];
    assign P[2] = in[94] ^ in2[94];
    assign G[3] = in[93] & in2[93];
    assign P[3] = in[93] ^ in2[93];
    assign G[4] = in[92] & in2[92];
    assign P[4] = in[92] ^ in2[92];
    assign G[5] = in[91] & in2[91];
    assign P[5] = in[91] ^ in2[91];
    assign G[6] = in[90] & in2[90];
    assign P[6] = in[90] ^ in2[90];
    assign G[7] = in[89] & in2[89];
    assign P[7] = in[89] ^ in2[89];
    assign G[8] = in[88] & in2[88];
    assign P[8] = in[88] ^ in2[88];
    assign G[9] = in[87] & in2[87];
    assign P[9] = in[87] ^ in2[87];
    assign G[10] = in[86] & in2[86];
    assign P[10] = in[86] ^ in2[86];
    assign G[11] = in[85] & in2[85];
    assign P[11] = in[85] ^ in2[85];
    assign G[12] = in[84] & in2[84];
    assign P[12] = in[84] ^ in2[84];
    assign G[13] = in[83] & in2[83];
    assign P[13] = in[83] ^ in2[83];
    assign G[14] = in[82] & in2[82];
    assign P[14] = in[82] ^ in2[82];
    assign G[15] = in[81] & in2[81];
    assign P[15] = in[81] ^ in2[81];
    assign G[16] = in[80] & in2[80];
    assign P[16] = in[80] ^ in2[80];
    assign G[17] = in[79] & in2[79];
    assign P[17] = in[79] ^ in2[79];
    assign G[18] = in[78] & in2[78];
    assign P[18] = in[78] ^ in2[78];
    assign G[19] = in[77] & in2[77];
    assign P[19] = in[77] ^ in2[77];
    assign G[20] = in[76] & in2[76];
    assign P[20] = in[76] ^ in2[76];
    assign G[21] = in[75] & in2[75];
    assign P[21] = in[75] ^ in2[75];
    assign G[22] = in[74] & in2[74];
    assign P[22] = in[74] ^ in2[74];
    assign G[23] = in[73] & in2[73];
    assign P[23] = in[73] ^ in2[73];
    assign G[24] = in[72] & in2[72];
    assign P[24] = in[72] ^ in2[72];
    assign G[25] = in[71] & in2[71];
    assign P[25] = in[71] ^ in2[71];
    assign G[26] = in[70] & in2[70];
    assign P[26] = in[70] ^ in2[70];
    assign G[27] = in[69] & in2[69];
    assign P[27] = in[69] ^ in2[69];
    assign G[28] = in[68] & in2[68];
    assign P[28] = in[68] ^ in2[68];
    assign G[29] = in[67] & in2[67];
    assign P[29] = in[67] ^ in2[67];
    assign G[30] = in[66] & in2[66];
    assign P[30] = in[66] ^ in2[66];
    assign G[31] = in[65] & in2[65];
    assign P[31] = in[65] ^ in2[65];
    assign G[32] = in[64] & in2[64];
    assign P[32] = in[64] ^ in2[64];
    assign G[33] = in[63] & in2[63];
    assign P[33] = in[63] ^ in2[63];
    assign G[34] = in[62] & in2[62];
    assign P[34] = in[62] ^ in2[62];
    assign G[35] = in[61] & in2[61];
    assign P[35] = in[61] ^ in2[61];
    assign G[36] = in[60] & in2[60];
    assign P[36] = in[60] ^ in2[60];
    assign G[37] = in[59] & in2[59];
    assign P[37] = in[59] ^ in2[59];
    assign G[38] = in[58] & in2[58];
    assign P[38] = in[58] ^ in2[58];
    assign G[39] = in[57] & in2[57];
    assign P[39] = in[57] ^ in2[57];
    assign G[40] = in[56] & in2[56];
    assign P[40] = in[56] ^ in2[56];
    assign G[41] = in[55] & in2[55];
    assign P[41] = in[55] ^ in2[55];
    assign G[42] = in[54] & in2[54];
    assign P[42] = in[54] ^ in2[54];
    assign G[43] = in[53] & in2[53];
    assign P[43] = in[53] ^ in2[53];
    assign G[44] = in[52] & in2[52];
    assign P[44] = in[52] ^ in2[52];
    assign G[45] = in[51] & in2[51];
    assign P[45] = in[51] ^ in2[51];
    assign G[46] = in[50] & in2[50];
    assign P[46] = in[50] ^ in2[50];
    assign G[47] = in[49] & in2[49];
    assign P[47] = in[49] ^ in2[49];
    assign G[48] = in[48] & in2[48];
    assign P[48] = in[48] ^ in2[48];
    assign G[49] = in[47] & in2[47];
    assign P[49] = in[47] ^ in2[47];
    assign G[50] = in[46] & in2[46];
    assign P[50] = in[46] ^ in2[46];
    assign G[51] = in[45] & in2[45];
    assign P[51] = in[45] ^ in2[45];
    assign G[52] = in[44] & in2[44];
    assign P[52] = in[44] ^ in2[44];
    assign G[53] = in[43] & in2[43];
    assign P[53] = in[43] ^ in2[43];
    assign G[54] = in[42] & in2[42];
    assign P[54] = in[42] ^ in2[42];
    assign G[55] = in[41] & in2[41];
    assign P[55] = in[41] ^ in2[41];
    assign G[56] = in[40] & in2[40];
    assign P[56] = in[40] ^ in2[40];
    assign G[57] = in[39] & in2[39];
    assign P[57] = in[39] ^ in2[39];
    assign G[58] = in[38] & in2[38];
    assign P[58] = in[38] ^ in2[38];
    assign G[59] = in[37] & in2[37];
    assign P[59] = in[37] ^ in2[37];
    assign G[60] = in[36] & in2[36];
    assign P[60] = in[36] ^ in2[36];
    assign G[61] = in[35] & in2[35];
    assign P[61] = in[35] ^ in2[35];
    assign G[62] = in[34] & in2[34];
    assign P[62] = in[34] ^ in2[34];
    assign G[63] = in[33] & in2[33];
    assign P[63] = in[33] ^ in2[33];
    assign G[64] = in[32] & in2[32];
    assign P[64] = in[32] ^ in2[32];
    assign G[65] = in[31] & in2[31];
    assign P[65] = in[31] ^ in2[31];
    assign G[66] = in[30] & in2[30];
    assign P[66] = in[30] ^ in2[30];
    assign G[67] = in[29] & in2[29];
    assign P[67] = in[29] ^ in2[29];
    assign G[68] = in[28] & in2[28];
    assign P[68] = in[28] ^ in2[28];
    assign G[69] = in[27] & in2[27];
    assign P[69] = in[27] ^ in2[27];
    assign G[70] = in[26] & in2[26];
    assign P[70] = in[26] ^ in2[26];
    assign G[71] = in[25] & in2[25];
    assign P[71] = in[25] ^ in2[25];
    assign G[72] = in[24] & in2[24];
    assign P[72] = in[24] ^ in2[24];
    assign G[73] = in[23] & in2[23];
    assign P[73] = in[23] ^ in2[23];
    assign G[74] = in[22] & in2[22];
    assign P[74] = in[22] ^ in2[22];
    assign G[75] = in[21] & in2[21];
    assign P[75] = in[21] ^ in2[21];
    assign G[76] = in[20] & in2[20];
    assign P[76] = in[20] ^ in2[20];
    assign G[77] = in[19] & in2[19];
    assign P[77] = in[19] ^ in2[19];
    assign G[78] = in[18] & in2[18];
    assign P[78] = in[18] ^ in2[18];
    assign G[79] = in[17] & in2[17];
    assign P[79] = in[17] ^ in2[17];
    assign G[80] = in[16] & in2[16];
    assign P[80] = in[16] ^ in2[16];
    assign G[81] = in[15] & in2[15];
    assign P[81] = in[15] ^ in2[15];
    assign G[82] = in[14] & in2[14];
    assign P[82] = in[14] ^ in2[14];
    assign G[83] = in[13] & in2[13];
    assign P[83] = in[13] ^ in2[13];
    assign G[84] = in[12] & in2[12];
    assign P[84] = in[12] ^ in2[12];
    assign G[85] = in[11] & in2[11];
    assign P[85] = in[11] ^ in2[11];
    assign G[86] = in[10] & in2[10];
    assign P[86] = in[10] ^ in2[10];
    assign G[87] = in[9] & in2[9];
    assign P[87] = in[9] ^ in2[9];
    assign G[88] = in[8] & in2[8];
    assign P[88] = in[8] ^ in2[8];
    assign G[89] = in[7] & in2[7];
    assign P[89] = in[7] ^ in2[7];
    assign G[90] = in[6] & in2[6];
    assign P[90] = in[6] ^ in2[6];
    assign G[91] = in[5] & in2[5];
    assign P[91] = in[5] ^ in2[5];
    assign G[92] = in[4] & in2[4];
    assign P[92] = in[4] ^ in2[4];
    assign G[93] = in[3] & in2[3];
    assign P[93] = in[3] ^ in2[3];
    assign G[94] = in[2] & in2[2];
    assign P[94] = in[2] ^ in2[2];
    assign G[95] = in[1] & in2[1];
    assign P[95] = in[1] ^ in2[1];
    assign G[96] = in[0] & in2[0];
    assign P[96] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign C[96] = G[95] | (P[95] & C[95]);
    assign cout = G[96] | (P[96] & C[96]);
    assign sum = P ^ C;
endmodule

module CLA96(output [95:0] sum, output cout, input [95:0] in1, input [95:0] in2;

    wire[95:0] G;
    wire[95:0] C;
    wire[95:0] P;

    assign G[0] = in[95] & in2[95];
    assign P[0] = in[95] ^ in2[95];
    assign G[1] = in[94] & in2[94];
    assign P[1] = in[94] ^ in2[94];
    assign G[2] = in[93] & in2[93];
    assign P[2] = in[93] ^ in2[93];
    assign G[3] = in[92] & in2[92];
    assign P[3] = in[92] ^ in2[92];
    assign G[4] = in[91] & in2[91];
    assign P[4] = in[91] ^ in2[91];
    assign G[5] = in[90] & in2[90];
    assign P[5] = in[90] ^ in2[90];
    assign G[6] = in[89] & in2[89];
    assign P[6] = in[89] ^ in2[89];
    assign G[7] = in[88] & in2[88];
    assign P[7] = in[88] ^ in2[88];
    assign G[8] = in[87] & in2[87];
    assign P[8] = in[87] ^ in2[87];
    assign G[9] = in[86] & in2[86];
    assign P[9] = in[86] ^ in2[86];
    assign G[10] = in[85] & in2[85];
    assign P[10] = in[85] ^ in2[85];
    assign G[11] = in[84] & in2[84];
    assign P[11] = in[84] ^ in2[84];
    assign G[12] = in[83] & in2[83];
    assign P[12] = in[83] ^ in2[83];
    assign G[13] = in[82] & in2[82];
    assign P[13] = in[82] ^ in2[82];
    assign G[14] = in[81] & in2[81];
    assign P[14] = in[81] ^ in2[81];
    assign G[15] = in[80] & in2[80];
    assign P[15] = in[80] ^ in2[80];
    assign G[16] = in[79] & in2[79];
    assign P[16] = in[79] ^ in2[79];
    assign G[17] = in[78] & in2[78];
    assign P[17] = in[78] ^ in2[78];
    assign G[18] = in[77] & in2[77];
    assign P[18] = in[77] ^ in2[77];
    assign G[19] = in[76] & in2[76];
    assign P[19] = in[76] ^ in2[76];
    assign G[20] = in[75] & in2[75];
    assign P[20] = in[75] ^ in2[75];
    assign G[21] = in[74] & in2[74];
    assign P[21] = in[74] ^ in2[74];
    assign G[22] = in[73] & in2[73];
    assign P[22] = in[73] ^ in2[73];
    assign G[23] = in[72] & in2[72];
    assign P[23] = in[72] ^ in2[72];
    assign G[24] = in[71] & in2[71];
    assign P[24] = in[71] ^ in2[71];
    assign G[25] = in[70] & in2[70];
    assign P[25] = in[70] ^ in2[70];
    assign G[26] = in[69] & in2[69];
    assign P[26] = in[69] ^ in2[69];
    assign G[27] = in[68] & in2[68];
    assign P[27] = in[68] ^ in2[68];
    assign G[28] = in[67] & in2[67];
    assign P[28] = in[67] ^ in2[67];
    assign G[29] = in[66] & in2[66];
    assign P[29] = in[66] ^ in2[66];
    assign G[30] = in[65] & in2[65];
    assign P[30] = in[65] ^ in2[65];
    assign G[31] = in[64] & in2[64];
    assign P[31] = in[64] ^ in2[64];
    assign G[32] = in[63] & in2[63];
    assign P[32] = in[63] ^ in2[63];
    assign G[33] = in[62] & in2[62];
    assign P[33] = in[62] ^ in2[62];
    assign G[34] = in[61] & in2[61];
    assign P[34] = in[61] ^ in2[61];
    assign G[35] = in[60] & in2[60];
    assign P[35] = in[60] ^ in2[60];
    assign G[36] = in[59] & in2[59];
    assign P[36] = in[59] ^ in2[59];
    assign G[37] = in[58] & in2[58];
    assign P[37] = in[58] ^ in2[58];
    assign G[38] = in[57] & in2[57];
    assign P[38] = in[57] ^ in2[57];
    assign G[39] = in[56] & in2[56];
    assign P[39] = in[56] ^ in2[56];
    assign G[40] = in[55] & in2[55];
    assign P[40] = in[55] ^ in2[55];
    assign G[41] = in[54] & in2[54];
    assign P[41] = in[54] ^ in2[54];
    assign G[42] = in[53] & in2[53];
    assign P[42] = in[53] ^ in2[53];
    assign G[43] = in[52] & in2[52];
    assign P[43] = in[52] ^ in2[52];
    assign G[44] = in[51] & in2[51];
    assign P[44] = in[51] ^ in2[51];
    assign G[45] = in[50] & in2[50];
    assign P[45] = in[50] ^ in2[50];
    assign G[46] = in[49] & in2[49];
    assign P[46] = in[49] ^ in2[49];
    assign G[47] = in[48] & in2[48];
    assign P[47] = in[48] ^ in2[48];
    assign G[48] = in[47] & in2[47];
    assign P[48] = in[47] ^ in2[47];
    assign G[49] = in[46] & in2[46];
    assign P[49] = in[46] ^ in2[46];
    assign G[50] = in[45] & in2[45];
    assign P[50] = in[45] ^ in2[45];
    assign G[51] = in[44] & in2[44];
    assign P[51] = in[44] ^ in2[44];
    assign G[52] = in[43] & in2[43];
    assign P[52] = in[43] ^ in2[43];
    assign G[53] = in[42] & in2[42];
    assign P[53] = in[42] ^ in2[42];
    assign G[54] = in[41] & in2[41];
    assign P[54] = in[41] ^ in2[41];
    assign G[55] = in[40] & in2[40];
    assign P[55] = in[40] ^ in2[40];
    assign G[56] = in[39] & in2[39];
    assign P[56] = in[39] ^ in2[39];
    assign G[57] = in[38] & in2[38];
    assign P[57] = in[38] ^ in2[38];
    assign G[58] = in[37] & in2[37];
    assign P[58] = in[37] ^ in2[37];
    assign G[59] = in[36] & in2[36];
    assign P[59] = in[36] ^ in2[36];
    assign G[60] = in[35] & in2[35];
    assign P[60] = in[35] ^ in2[35];
    assign G[61] = in[34] & in2[34];
    assign P[61] = in[34] ^ in2[34];
    assign G[62] = in[33] & in2[33];
    assign P[62] = in[33] ^ in2[33];
    assign G[63] = in[32] & in2[32];
    assign P[63] = in[32] ^ in2[32];
    assign G[64] = in[31] & in2[31];
    assign P[64] = in[31] ^ in2[31];
    assign G[65] = in[30] & in2[30];
    assign P[65] = in[30] ^ in2[30];
    assign G[66] = in[29] & in2[29];
    assign P[66] = in[29] ^ in2[29];
    assign G[67] = in[28] & in2[28];
    assign P[67] = in[28] ^ in2[28];
    assign G[68] = in[27] & in2[27];
    assign P[68] = in[27] ^ in2[27];
    assign G[69] = in[26] & in2[26];
    assign P[69] = in[26] ^ in2[26];
    assign G[70] = in[25] & in2[25];
    assign P[70] = in[25] ^ in2[25];
    assign G[71] = in[24] & in2[24];
    assign P[71] = in[24] ^ in2[24];
    assign G[72] = in[23] & in2[23];
    assign P[72] = in[23] ^ in2[23];
    assign G[73] = in[22] & in2[22];
    assign P[73] = in[22] ^ in2[22];
    assign G[74] = in[21] & in2[21];
    assign P[74] = in[21] ^ in2[21];
    assign G[75] = in[20] & in2[20];
    assign P[75] = in[20] ^ in2[20];
    assign G[76] = in[19] & in2[19];
    assign P[76] = in[19] ^ in2[19];
    assign G[77] = in[18] & in2[18];
    assign P[77] = in[18] ^ in2[18];
    assign G[78] = in[17] & in2[17];
    assign P[78] = in[17] ^ in2[17];
    assign G[79] = in[16] & in2[16];
    assign P[79] = in[16] ^ in2[16];
    assign G[80] = in[15] & in2[15];
    assign P[80] = in[15] ^ in2[15];
    assign G[81] = in[14] & in2[14];
    assign P[81] = in[14] ^ in2[14];
    assign G[82] = in[13] & in2[13];
    assign P[82] = in[13] ^ in2[13];
    assign G[83] = in[12] & in2[12];
    assign P[83] = in[12] ^ in2[12];
    assign G[84] = in[11] & in2[11];
    assign P[84] = in[11] ^ in2[11];
    assign G[85] = in[10] & in2[10];
    assign P[85] = in[10] ^ in2[10];
    assign G[86] = in[9] & in2[9];
    assign P[86] = in[9] ^ in2[9];
    assign G[87] = in[8] & in2[8];
    assign P[87] = in[8] ^ in2[8];
    assign G[88] = in[7] & in2[7];
    assign P[88] = in[7] ^ in2[7];
    assign G[89] = in[6] & in2[6];
    assign P[89] = in[6] ^ in2[6];
    assign G[90] = in[5] & in2[5];
    assign P[90] = in[5] ^ in2[5];
    assign G[91] = in[4] & in2[4];
    assign P[91] = in[4] ^ in2[4];
    assign G[92] = in[3] & in2[3];
    assign P[92] = in[3] ^ in2[3];
    assign G[93] = in[2] & in2[2];
    assign P[93] = in[2] ^ in2[2];
    assign G[94] = in[1] & in2[1];
    assign P[94] = in[1] ^ in2[1];
    assign G[95] = in[0] & in2[0];
    assign P[95] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign C[95] = G[94] | (P[94] & C[94]);
    assign cout = G[95] | (P[95] & C[95]);
    assign sum = P ^ C;
endmodule

module CLA95(output [94:0] sum, output cout, input [94:0] in1, input [94:0] in2;

    wire[94:0] G;
    wire[94:0] C;
    wire[94:0] P;

    assign G[0] = in[94] & in2[94];
    assign P[0] = in[94] ^ in2[94];
    assign G[1] = in[93] & in2[93];
    assign P[1] = in[93] ^ in2[93];
    assign G[2] = in[92] & in2[92];
    assign P[2] = in[92] ^ in2[92];
    assign G[3] = in[91] & in2[91];
    assign P[3] = in[91] ^ in2[91];
    assign G[4] = in[90] & in2[90];
    assign P[4] = in[90] ^ in2[90];
    assign G[5] = in[89] & in2[89];
    assign P[5] = in[89] ^ in2[89];
    assign G[6] = in[88] & in2[88];
    assign P[6] = in[88] ^ in2[88];
    assign G[7] = in[87] & in2[87];
    assign P[7] = in[87] ^ in2[87];
    assign G[8] = in[86] & in2[86];
    assign P[8] = in[86] ^ in2[86];
    assign G[9] = in[85] & in2[85];
    assign P[9] = in[85] ^ in2[85];
    assign G[10] = in[84] & in2[84];
    assign P[10] = in[84] ^ in2[84];
    assign G[11] = in[83] & in2[83];
    assign P[11] = in[83] ^ in2[83];
    assign G[12] = in[82] & in2[82];
    assign P[12] = in[82] ^ in2[82];
    assign G[13] = in[81] & in2[81];
    assign P[13] = in[81] ^ in2[81];
    assign G[14] = in[80] & in2[80];
    assign P[14] = in[80] ^ in2[80];
    assign G[15] = in[79] & in2[79];
    assign P[15] = in[79] ^ in2[79];
    assign G[16] = in[78] & in2[78];
    assign P[16] = in[78] ^ in2[78];
    assign G[17] = in[77] & in2[77];
    assign P[17] = in[77] ^ in2[77];
    assign G[18] = in[76] & in2[76];
    assign P[18] = in[76] ^ in2[76];
    assign G[19] = in[75] & in2[75];
    assign P[19] = in[75] ^ in2[75];
    assign G[20] = in[74] & in2[74];
    assign P[20] = in[74] ^ in2[74];
    assign G[21] = in[73] & in2[73];
    assign P[21] = in[73] ^ in2[73];
    assign G[22] = in[72] & in2[72];
    assign P[22] = in[72] ^ in2[72];
    assign G[23] = in[71] & in2[71];
    assign P[23] = in[71] ^ in2[71];
    assign G[24] = in[70] & in2[70];
    assign P[24] = in[70] ^ in2[70];
    assign G[25] = in[69] & in2[69];
    assign P[25] = in[69] ^ in2[69];
    assign G[26] = in[68] & in2[68];
    assign P[26] = in[68] ^ in2[68];
    assign G[27] = in[67] & in2[67];
    assign P[27] = in[67] ^ in2[67];
    assign G[28] = in[66] & in2[66];
    assign P[28] = in[66] ^ in2[66];
    assign G[29] = in[65] & in2[65];
    assign P[29] = in[65] ^ in2[65];
    assign G[30] = in[64] & in2[64];
    assign P[30] = in[64] ^ in2[64];
    assign G[31] = in[63] & in2[63];
    assign P[31] = in[63] ^ in2[63];
    assign G[32] = in[62] & in2[62];
    assign P[32] = in[62] ^ in2[62];
    assign G[33] = in[61] & in2[61];
    assign P[33] = in[61] ^ in2[61];
    assign G[34] = in[60] & in2[60];
    assign P[34] = in[60] ^ in2[60];
    assign G[35] = in[59] & in2[59];
    assign P[35] = in[59] ^ in2[59];
    assign G[36] = in[58] & in2[58];
    assign P[36] = in[58] ^ in2[58];
    assign G[37] = in[57] & in2[57];
    assign P[37] = in[57] ^ in2[57];
    assign G[38] = in[56] & in2[56];
    assign P[38] = in[56] ^ in2[56];
    assign G[39] = in[55] & in2[55];
    assign P[39] = in[55] ^ in2[55];
    assign G[40] = in[54] & in2[54];
    assign P[40] = in[54] ^ in2[54];
    assign G[41] = in[53] & in2[53];
    assign P[41] = in[53] ^ in2[53];
    assign G[42] = in[52] & in2[52];
    assign P[42] = in[52] ^ in2[52];
    assign G[43] = in[51] & in2[51];
    assign P[43] = in[51] ^ in2[51];
    assign G[44] = in[50] & in2[50];
    assign P[44] = in[50] ^ in2[50];
    assign G[45] = in[49] & in2[49];
    assign P[45] = in[49] ^ in2[49];
    assign G[46] = in[48] & in2[48];
    assign P[46] = in[48] ^ in2[48];
    assign G[47] = in[47] & in2[47];
    assign P[47] = in[47] ^ in2[47];
    assign G[48] = in[46] & in2[46];
    assign P[48] = in[46] ^ in2[46];
    assign G[49] = in[45] & in2[45];
    assign P[49] = in[45] ^ in2[45];
    assign G[50] = in[44] & in2[44];
    assign P[50] = in[44] ^ in2[44];
    assign G[51] = in[43] & in2[43];
    assign P[51] = in[43] ^ in2[43];
    assign G[52] = in[42] & in2[42];
    assign P[52] = in[42] ^ in2[42];
    assign G[53] = in[41] & in2[41];
    assign P[53] = in[41] ^ in2[41];
    assign G[54] = in[40] & in2[40];
    assign P[54] = in[40] ^ in2[40];
    assign G[55] = in[39] & in2[39];
    assign P[55] = in[39] ^ in2[39];
    assign G[56] = in[38] & in2[38];
    assign P[56] = in[38] ^ in2[38];
    assign G[57] = in[37] & in2[37];
    assign P[57] = in[37] ^ in2[37];
    assign G[58] = in[36] & in2[36];
    assign P[58] = in[36] ^ in2[36];
    assign G[59] = in[35] & in2[35];
    assign P[59] = in[35] ^ in2[35];
    assign G[60] = in[34] & in2[34];
    assign P[60] = in[34] ^ in2[34];
    assign G[61] = in[33] & in2[33];
    assign P[61] = in[33] ^ in2[33];
    assign G[62] = in[32] & in2[32];
    assign P[62] = in[32] ^ in2[32];
    assign G[63] = in[31] & in2[31];
    assign P[63] = in[31] ^ in2[31];
    assign G[64] = in[30] & in2[30];
    assign P[64] = in[30] ^ in2[30];
    assign G[65] = in[29] & in2[29];
    assign P[65] = in[29] ^ in2[29];
    assign G[66] = in[28] & in2[28];
    assign P[66] = in[28] ^ in2[28];
    assign G[67] = in[27] & in2[27];
    assign P[67] = in[27] ^ in2[27];
    assign G[68] = in[26] & in2[26];
    assign P[68] = in[26] ^ in2[26];
    assign G[69] = in[25] & in2[25];
    assign P[69] = in[25] ^ in2[25];
    assign G[70] = in[24] & in2[24];
    assign P[70] = in[24] ^ in2[24];
    assign G[71] = in[23] & in2[23];
    assign P[71] = in[23] ^ in2[23];
    assign G[72] = in[22] & in2[22];
    assign P[72] = in[22] ^ in2[22];
    assign G[73] = in[21] & in2[21];
    assign P[73] = in[21] ^ in2[21];
    assign G[74] = in[20] & in2[20];
    assign P[74] = in[20] ^ in2[20];
    assign G[75] = in[19] & in2[19];
    assign P[75] = in[19] ^ in2[19];
    assign G[76] = in[18] & in2[18];
    assign P[76] = in[18] ^ in2[18];
    assign G[77] = in[17] & in2[17];
    assign P[77] = in[17] ^ in2[17];
    assign G[78] = in[16] & in2[16];
    assign P[78] = in[16] ^ in2[16];
    assign G[79] = in[15] & in2[15];
    assign P[79] = in[15] ^ in2[15];
    assign G[80] = in[14] & in2[14];
    assign P[80] = in[14] ^ in2[14];
    assign G[81] = in[13] & in2[13];
    assign P[81] = in[13] ^ in2[13];
    assign G[82] = in[12] & in2[12];
    assign P[82] = in[12] ^ in2[12];
    assign G[83] = in[11] & in2[11];
    assign P[83] = in[11] ^ in2[11];
    assign G[84] = in[10] & in2[10];
    assign P[84] = in[10] ^ in2[10];
    assign G[85] = in[9] & in2[9];
    assign P[85] = in[9] ^ in2[9];
    assign G[86] = in[8] & in2[8];
    assign P[86] = in[8] ^ in2[8];
    assign G[87] = in[7] & in2[7];
    assign P[87] = in[7] ^ in2[7];
    assign G[88] = in[6] & in2[6];
    assign P[88] = in[6] ^ in2[6];
    assign G[89] = in[5] & in2[5];
    assign P[89] = in[5] ^ in2[5];
    assign G[90] = in[4] & in2[4];
    assign P[90] = in[4] ^ in2[4];
    assign G[91] = in[3] & in2[3];
    assign P[91] = in[3] ^ in2[3];
    assign G[92] = in[2] & in2[2];
    assign P[92] = in[2] ^ in2[2];
    assign G[93] = in[1] & in2[1];
    assign P[93] = in[1] ^ in2[1];
    assign G[94] = in[0] & in2[0];
    assign P[94] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign C[94] = G[93] | (P[93] & C[93]);
    assign cout = G[94] | (P[94] & C[94]);
    assign sum = P ^ C;
endmodule

module CLA94(output [93:0] sum, output cout, input [93:0] in1, input [93:0] in2;

    wire[93:0] G;
    wire[93:0] C;
    wire[93:0] P;

    assign G[0] = in[93] & in2[93];
    assign P[0] = in[93] ^ in2[93];
    assign G[1] = in[92] & in2[92];
    assign P[1] = in[92] ^ in2[92];
    assign G[2] = in[91] & in2[91];
    assign P[2] = in[91] ^ in2[91];
    assign G[3] = in[90] & in2[90];
    assign P[3] = in[90] ^ in2[90];
    assign G[4] = in[89] & in2[89];
    assign P[4] = in[89] ^ in2[89];
    assign G[5] = in[88] & in2[88];
    assign P[5] = in[88] ^ in2[88];
    assign G[6] = in[87] & in2[87];
    assign P[6] = in[87] ^ in2[87];
    assign G[7] = in[86] & in2[86];
    assign P[7] = in[86] ^ in2[86];
    assign G[8] = in[85] & in2[85];
    assign P[8] = in[85] ^ in2[85];
    assign G[9] = in[84] & in2[84];
    assign P[9] = in[84] ^ in2[84];
    assign G[10] = in[83] & in2[83];
    assign P[10] = in[83] ^ in2[83];
    assign G[11] = in[82] & in2[82];
    assign P[11] = in[82] ^ in2[82];
    assign G[12] = in[81] & in2[81];
    assign P[12] = in[81] ^ in2[81];
    assign G[13] = in[80] & in2[80];
    assign P[13] = in[80] ^ in2[80];
    assign G[14] = in[79] & in2[79];
    assign P[14] = in[79] ^ in2[79];
    assign G[15] = in[78] & in2[78];
    assign P[15] = in[78] ^ in2[78];
    assign G[16] = in[77] & in2[77];
    assign P[16] = in[77] ^ in2[77];
    assign G[17] = in[76] & in2[76];
    assign P[17] = in[76] ^ in2[76];
    assign G[18] = in[75] & in2[75];
    assign P[18] = in[75] ^ in2[75];
    assign G[19] = in[74] & in2[74];
    assign P[19] = in[74] ^ in2[74];
    assign G[20] = in[73] & in2[73];
    assign P[20] = in[73] ^ in2[73];
    assign G[21] = in[72] & in2[72];
    assign P[21] = in[72] ^ in2[72];
    assign G[22] = in[71] & in2[71];
    assign P[22] = in[71] ^ in2[71];
    assign G[23] = in[70] & in2[70];
    assign P[23] = in[70] ^ in2[70];
    assign G[24] = in[69] & in2[69];
    assign P[24] = in[69] ^ in2[69];
    assign G[25] = in[68] & in2[68];
    assign P[25] = in[68] ^ in2[68];
    assign G[26] = in[67] & in2[67];
    assign P[26] = in[67] ^ in2[67];
    assign G[27] = in[66] & in2[66];
    assign P[27] = in[66] ^ in2[66];
    assign G[28] = in[65] & in2[65];
    assign P[28] = in[65] ^ in2[65];
    assign G[29] = in[64] & in2[64];
    assign P[29] = in[64] ^ in2[64];
    assign G[30] = in[63] & in2[63];
    assign P[30] = in[63] ^ in2[63];
    assign G[31] = in[62] & in2[62];
    assign P[31] = in[62] ^ in2[62];
    assign G[32] = in[61] & in2[61];
    assign P[32] = in[61] ^ in2[61];
    assign G[33] = in[60] & in2[60];
    assign P[33] = in[60] ^ in2[60];
    assign G[34] = in[59] & in2[59];
    assign P[34] = in[59] ^ in2[59];
    assign G[35] = in[58] & in2[58];
    assign P[35] = in[58] ^ in2[58];
    assign G[36] = in[57] & in2[57];
    assign P[36] = in[57] ^ in2[57];
    assign G[37] = in[56] & in2[56];
    assign P[37] = in[56] ^ in2[56];
    assign G[38] = in[55] & in2[55];
    assign P[38] = in[55] ^ in2[55];
    assign G[39] = in[54] & in2[54];
    assign P[39] = in[54] ^ in2[54];
    assign G[40] = in[53] & in2[53];
    assign P[40] = in[53] ^ in2[53];
    assign G[41] = in[52] & in2[52];
    assign P[41] = in[52] ^ in2[52];
    assign G[42] = in[51] & in2[51];
    assign P[42] = in[51] ^ in2[51];
    assign G[43] = in[50] & in2[50];
    assign P[43] = in[50] ^ in2[50];
    assign G[44] = in[49] & in2[49];
    assign P[44] = in[49] ^ in2[49];
    assign G[45] = in[48] & in2[48];
    assign P[45] = in[48] ^ in2[48];
    assign G[46] = in[47] & in2[47];
    assign P[46] = in[47] ^ in2[47];
    assign G[47] = in[46] & in2[46];
    assign P[47] = in[46] ^ in2[46];
    assign G[48] = in[45] & in2[45];
    assign P[48] = in[45] ^ in2[45];
    assign G[49] = in[44] & in2[44];
    assign P[49] = in[44] ^ in2[44];
    assign G[50] = in[43] & in2[43];
    assign P[50] = in[43] ^ in2[43];
    assign G[51] = in[42] & in2[42];
    assign P[51] = in[42] ^ in2[42];
    assign G[52] = in[41] & in2[41];
    assign P[52] = in[41] ^ in2[41];
    assign G[53] = in[40] & in2[40];
    assign P[53] = in[40] ^ in2[40];
    assign G[54] = in[39] & in2[39];
    assign P[54] = in[39] ^ in2[39];
    assign G[55] = in[38] & in2[38];
    assign P[55] = in[38] ^ in2[38];
    assign G[56] = in[37] & in2[37];
    assign P[56] = in[37] ^ in2[37];
    assign G[57] = in[36] & in2[36];
    assign P[57] = in[36] ^ in2[36];
    assign G[58] = in[35] & in2[35];
    assign P[58] = in[35] ^ in2[35];
    assign G[59] = in[34] & in2[34];
    assign P[59] = in[34] ^ in2[34];
    assign G[60] = in[33] & in2[33];
    assign P[60] = in[33] ^ in2[33];
    assign G[61] = in[32] & in2[32];
    assign P[61] = in[32] ^ in2[32];
    assign G[62] = in[31] & in2[31];
    assign P[62] = in[31] ^ in2[31];
    assign G[63] = in[30] & in2[30];
    assign P[63] = in[30] ^ in2[30];
    assign G[64] = in[29] & in2[29];
    assign P[64] = in[29] ^ in2[29];
    assign G[65] = in[28] & in2[28];
    assign P[65] = in[28] ^ in2[28];
    assign G[66] = in[27] & in2[27];
    assign P[66] = in[27] ^ in2[27];
    assign G[67] = in[26] & in2[26];
    assign P[67] = in[26] ^ in2[26];
    assign G[68] = in[25] & in2[25];
    assign P[68] = in[25] ^ in2[25];
    assign G[69] = in[24] & in2[24];
    assign P[69] = in[24] ^ in2[24];
    assign G[70] = in[23] & in2[23];
    assign P[70] = in[23] ^ in2[23];
    assign G[71] = in[22] & in2[22];
    assign P[71] = in[22] ^ in2[22];
    assign G[72] = in[21] & in2[21];
    assign P[72] = in[21] ^ in2[21];
    assign G[73] = in[20] & in2[20];
    assign P[73] = in[20] ^ in2[20];
    assign G[74] = in[19] & in2[19];
    assign P[74] = in[19] ^ in2[19];
    assign G[75] = in[18] & in2[18];
    assign P[75] = in[18] ^ in2[18];
    assign G[76] = in[17] & in2[17];
    assign P[76] = in[17] ^ in2[17];
    assign G[77] = in[16] & in2[16];
    assign P[77] = in[16] ^ in2[16];
    assign G[78] = in[15] & in2[15];
    assign P[78] = in[15] ^ in2[15];
    assign G[79] = in[14] & in2[14];
    assign P[79] = in[14] ^ in2[14];
    assign G[80] = in[13] & in2[13];
    assign P[80] = in[13] ^ in2[13];
    assign G[81] = in[12] & in2[12];
    assign P[81] = in[12] ^ in2[12];
    assign G[82] = in[11] & in2[11];
    assign P[82] = in[11] ^ in2[11];
    assign G[83] = in[10] & in2[10];
    assign P[83] = in[10] ^ in2[10];
    assign G[84] = in[9] & in2[9];
    assign P[84] = in[9] ^ in2[9];
    assign G[85] = in[8] & in2[8];
    assign P[85] = in[8] ^ in2[8];
    assign G[86] = in[7] & in2[7];
    assign P[86] = in[7] ^ in2[7];
    assign G[87] = in[6] & in2[6];
    assign P[87] = in[6] ^ in2[6];
    assign G[88] = in[5] & in2[5];
    assign P[88] = in[5] ^ in2[5];
    assign G[89] = in[4] & in2[4];
    assign P[89] = in[4] ^ in2[4];
    assign G[90] = in[3] & in2[3];
    assign P[90] = in[3] ^ in2[3];
    assign G[91] = in[2] & in2[2];
    assign P[91] = in[2] ^ in2[2];
    assign G[92] = in[1] & in2[1];
    assign P[92] = in[1] ^ in2[1];
    assign G[93] = in[0] & in2[0];
    assign P[93] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign C[93] = G[92] | (P[92] & C[92]);
    assign cout = G[93] | (P[93] & C[93]);
    assign sum = P ^ C;
endmodule

module CLA93(output [92:0] sum, output cout, input [92:0] in1, input [92:0] in2;

    wire[92:0] G;
    wire[92:0] C;
    wire[92:0] P;

    assign G[0] = in[92] & in2[92];
    assign P[0] = in[92] ^ in2[92];
    assign G[1] = in[91] & in2[91];
    assign P[1] = in[91] ^ in2[91];
    assign G[2] = in[90] & in2[90];
    assign P[2] = in[90] ^ in2[90];
    assign G[3] = in[89] & in2[89];
    assign P[3] = in[89] ^ in2[89];
    assign G[4] = in[88] & in2[88];
    assign P[4] = in[88] ^ in2[88];
    assign G[5] = in[87] & in2[87];
    assign P[5] = in[87] ^ in2[87];
    assign G[6] = in[86] & in2[86];
    assign P[6] = in[86] ^ in2[86];
    assign G[7] = in[85] & in2[85];
    assign P[7] = in[85] ^ in2[85];
    assign G[8] = in[84] & in2[84];
    assign P[8] = in[84] ^ in2[84];
    assign G[9] = in[83] & in2[83];
    assign P[9] = in[83] ^ in2[83];
    assign G[10] = in[82] & in2[82];
    assign P[10] = in[82] ^ in2[82];
    assign G[11] = in[81] & in2[81];
    assign P[11] = in[81] ^ in2[81];
    assign G[12] = in[80] & in2[80];
    assign P[12] = in[80] ^ in2[80];
    assign G[13] = in[79] & in2[79];
    assign P[13] = in[79] ^ in2[79];
    assign G[14] = in[78] & in2[78];
    assign P[14] = in[78] ^ in2[78];
    assign G[15] = in[77] & in2[77];
    assign P[15] = in[77] ^ in2[77];
    assign G[16] = in[76] & in2[76];
    assign P[16] = in[76] ^ in2[76];
    assign G[17] = in[75] & in2[75];
    assign P[17] = in[75] ^ in2[75];
    assign G[18] = in[74] & in2[74];
    assign P[18] = in[74] ^ in2[74];
    assign G[19] = in[73] & in2[73];
    assign P[19] = in[73] ^ in2[73];
    assign G[20] = in[72] & in2[72];
    assign P[20] = in[72] ^ in2[72];
    assign G[21] = in[71] & in2[71];
    assign P[21] = in[71] ^ in2[71];
    assign G[22] = in[70] & in2[70];
    assign P[22] = in[70] ^ in2[70];
    assign G[23] = in[69] & in2[69];
    assign P[23] = in[69] ^ in2[69];
    assign G[24] = in[68] & in2[68];
    assign P[24] = in[68] ^ in2[68];
    assign G[25] = in[67] & in2[67];
    assign P[25] = in[67] ^ in2[67];
    assign G[26] = in[66] & in2[66];
    assign P[26] = in[66] ^ in2[66];
    assign G[27] = in[65] & in2[65];
    assign P[27] = in[65] ^ in2[65];
    assign G[28] = in[64] & in2[64];
    assign P[28] = in[64] ^ in2[64];
    assign G[29] = in[63] & in2[63];
    assign P[29] = in[63] ^ in2[63];
    assign G[30] = in[62] & in2[62];
    assign P[30] = in[62] ^ in2[62];
    assign G[31] = in[61] & in2[61];
    assign P[31] = in[61] ^ in2[61];
    assign G[32] = in[60] & in2[60];
    assign P[32] = in[60] ^ in2[60];
    assign G[33] = in[59] & in2[59];
    assign P[33] = in[59] ^ in2[59];
    assign G[34] = in[58] & in2[58];
    assign P[34] = in[58] ^ in2[58];
    assign G[35] = in[57] & in2[57];
    assign P[35] = in[57] ^ in2[57];
    assign G[36] = in[56] & in2[56];
    assign P[36] = in[56] ^ in2[56];
    assign G[37] = in[55] & in2[55];
    assign P[37] = in[55] ^ in2[55];
    assign G[38] = in[54] & in2[54];
    assign P[38] = in[54] ^ in2[54];
    assign G[39] = in[53] & in2[53];
    assign P[39] = in[53] ^ in2[53];
    assign G[40] = in[52] & in2[52];
    assign P[40] = in[52] ^ in2[52];
    assign G[41] = in[51] & in2[51];
    assign P[41] = in[51] ^ in2[51];
    assign G[42] = in[50] & in2[50];
    assign P[42] = in[50] ^ in2[50];
    assign G[43] = in[49] & in2[49];
    assign P[43] = in[49] ^ in2[49];
    assign G[44] = in[48] & in2[48];
    assign P[44] = in[48] ^ in2[48];
    assign G[45] = in[47] & in2[47];
    assign P[45] = in[47] ^ in2[47];
    assign G[46] = in[46] & in2[46];
    assign P[46] = in[46] ^ in2[46];
    assign G[47] = in[45] & in2[45];
    assign P[47] = in[45] ^ in2[45];
    assign G[48] = in[44] & in2[44];
    assign P[48] = in[44] ^ in2[44];
    assign G[49] = in[43] & in2[43];
    assign P[49] = in[43] ^ in2[43];
    assign G[50] = in[42] & in2[42];
    assign P[50] = in[42] ^ in2[42];
    assign G[51] = in[41] & in2[41];
    assign P[51] = in[41] ^ in2[41];
    assign G[52] = in[40] & in2[40];
    assign P[52] = in[40] ^ in2[40];
    assign G[53] = in[39] & in2[39];
    assign P[53] = in[39] ^ in2[39];
    assign G[54] = in[38] & in2[38];
    assign P[54] = in[38] ^ in2[38];
    assign G[55] = in[37] & in2[37];
    assign P[55] = in[37] ^ in2[37];
    assign G[56] = in[36] & in2[36];
    assign P[56] = in[36] ^ in2[36];
    assign G[57] = in[35] & in2[35];
    assign P[57] = in[35] ^ in2[35];
    assign G[58] = in[34] & in2[34];
    assign P[58] = in[34] ^ in2[34];
    assign G[59] = in[33] & in2[33];
    assign P[59] = in[33] ^ in2[33];
    assign G[60] = in[32] & in2[32];
    assign P[60] = in[32] ^ in2[32];
    assign G[61] = in[31] & in2[31];
    assign P[61] = in[31] ^ in2[31];
    assign G[62] = in[30] & in2[30];
    assign P[62] = in[30] ^ in2[30];
    assign G[63] = in[29] & in2[29];
    assign P[63] = in[29] ^ in2[29];
    assign G[64] = in[28] & in2[28];
    assign P[64] = in[28] ^ in2[28];
    assign G[65] = in[27] & in2[27];
    assign P[65] = in[27] ^ in2[27];
    assign G[66] = in[26] & in2[26];
    assign P[66] = in[26] ^ in2[26];
    assign G[67] = in[25] & in2[25];
    assign P[67] = in[25] ^ in2[25];
    assign G[68] = in[24] & in2[24];
    assign P[68] = in[24] ^ in2[24];
    assign G[69] = in[23] & in2[23];
    assign P[69] = in[23] ^ in2[23];
    assign G[70] = in[22] & in2[22];
    assign P[70] = in[22] ^ in2[22];
    assign G[71] = in[21] & in2[21];
    assign P[71] = in[21] ^ in2[21];
    assign G[72] = in[20] & in2[20];
    assign P[72] = in[20] ^ in2[20];
    assign G[73] = in[19] & in2[19];
    assign P[73] = in[19] ^ in2[19];
    assign G[74] = in[18] & in2[18];
    assign P[74] = in[18] ^ in2[18];
    assign G[75] = in[17] & in2[17];
    assign P[75] = in[17] ^ in2[17];
    assign G[76] = in[16] & in2[16];
    assign P[76] = in[16] ^ in2[16];
    assign G[77] = in[15] & in2[15];
    assign P[77] = in[15] ^ in2[15];
    assign G[78] = in[14] & in2[14];
    assign P[78] = in[14] ^ in2[14];
    assign G[79] = in[13] & in2[13];
    assign P[79] = in[13] ^ in2[13];
    assign G[80] = in[12] & in2[12];
    assign P[80] = in[12] ^ in2[12];
    assign G[81] = in[11] & in2[11];
    assign P[81] = in[11] ^ in2[11];
    assign G[82] = in[10] & in2[10];
    assign P[82] = in[10] ^ in2[10];
    assign G[83] = in[9] & in2[9];
    assign P[83] = in[9] ^ in2[9];
    assign G[84] = in[8] & in2[8];
    assign P[84] = in[8] ^ in2[8];
    assign G[85] = in[7] & in2[7];
    assign P[85] = in[7] ^ in2[7];
    assign G[86] = in[6] & in2[6];
    assign P[86] = in[6] ^ in2[6];
    assign G[87] = in[5] & in2[5];
    assign P[87] = in[5] ^ in2[5];
    assign G[88] = in[4] & in2[4];
    assign P[88] = in[4] ^ in2[4];
    assign G[89] = in[3] & in2[3];
    assign P[89] = in[3] ^ in2[3];
    assign G[90] = in[2] & in2[2];
    assign P[90] = in[2] ^ in2[2];
    assign G[91] = in[1] & in2[1];
    assign P[91] = in[1] ^ in2[1];
    assign G[92] = in[0] & in2[0];
    assign P[92] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign C[92] = G[91] | (P[91] & C[91]);
    assign cout = G[92] | (P[92] & C[92]);
    assign sum = P ^ C;
endmodule

module CLA92(output [91:0] sum, output cout, input [91:0] in1, input [91:0] in2;

    wire[91:0] G;
    wire[91:0] C;
    wire[91:0] P;

    assign G[0] = in[91] & in2[91];
    assign P[0] = in[91] ^ in2[91];
    assign G[1] = in[90] & in2[90];
    assign P[1] = in[90] ^ in2[90];
    assign G[2] = in[89] & in2[89];
    assign P[2] = in[89] ^ in2[89];
    assign G[3] = in[88] & in2[88];
    assign P[3] = in[88] ^ in2[88];
    assign G[4] = in[87] & in2[87];
    assign P[4] = in[87] ^ in2[87];
    assign G[5] = in[86] & in2[86];
    assign P[5] = in[86] ^ in2[86];
    assign G[6] = in[85] & in2[85];
    assign P[6] = in[85] ^ in2[85];
    assign G[7] = in[84] & in2[84];
    assign P[7] = in[84] ^ in2[84];
    assign G[8] = in[83] & in2[83];
    assign P[8] = in[83] ^ in2[83];
    assign G[9] = in[82] & in2[82];
    assign P[9] = in[82] ^ in2[82];
    assign G[10] = in[81] & in2[81];
    assign P[10] = in[81] ^ in2[81];
    assign G[11] = in[80] & in2[80];
    assign P[11] = in[80] ^ in2[80];
    assign G[12] = in[79] & in2[79];
    assign P[12] = in[79] ^ in2[79];
    assign G[13] = in[78] & in2[78];
    assign P[13] = in[78] ^ in2[78];
    assign G[14] = in[77] & in2[77];
    assign P[14] = in[77] ^ in2[77];
    assign G[15] = in[76] & in2[76];
    assign P[15] = in[76] ^ in2[76];
    assign G[16] = in[75] & in2[75];
    assign P[16] = in[75] ^ in2[75];
    assign G[17] = in[74] & in2[74];
    assign P[17] = in[74] ^ in2[74];
    assign G[18] = in[73] & in2[73];
    assign P[18] = in[73] ^ in2[73];
    assign G[19] = in[72] & in2[72];
    assign P[19] = in[72] ^ in2[72];
    assign G[20] = in[71] & in2[71];
    assign P[20] = in[71] ^ in2[71];
    assign G[21] = in[70] & in2[70];
    assign P[21] = in[70] ^ in2[70];
    assign G[22] = in[69] & in2[69];
    assign P[22] = in[69] ^ in2[69];
    assign G[23] = in[68] & in2[68];
    assign P[23] = in[68] ^ in2[68];
    assign G[24] = in[67] & in2[67];
    assign P[24] = in[67] ^ in2[67];
    assign G[25] = in[66] & in2[66];
    assign P[25] = in[66] ^ in2[66];
    assign G[26] = in[65] & in2[65];
    assign P[26] = in[65] ^ in2[65];
    assign G[27] = in[64] & in2[64];
    assign P[27] = in[64] ^ in2[64];
    assign G[28] = in[63] & in2[63];
    assign P[28] = in[63] ^ in2[63];
    assign G[29] = in[62] & in2[62];
    assign P[29] = in[62] ^ in2[62];
    assign G[30] = in[61] & in2[61];
    assign P[30] = in[61] ^ in2[61];
    assign G[31] = in[60] & in2[60];
    assign P[31] = in[60] ^ in2[60];
    assign G[32] = in[59] & in2[59];
    assign P[32] = in[59] ^ in2[59];
    assign G[33] = in[58] & in2[58];
    assign P[33] = in[58] ^ in2[58];
    assign G[34] = in[57] & in2[57];
    assign P[34] = in[57] ^ in2[57];
    assign G[35] = in[56] & in2[56];
    assign P[35] = in[56] ^ in2[56];
    assign G[36] = in[55] & in2[55];
    assign P[36] = in[55] ^ in2[55];
    assign G[37] = in[54] & in2[54];
    assign P[37] = in[54] ^ in2[54];
    assign G[38] = in[53] & in2[53];
    assign P[38] = in[53] ^ in2[53];
    assign G[39] = in[52] & in2[52];
    assign P[39] = in[52] ^ in2[52];
    assign G[40] = in[51] & in2[51];
    assign P[40] = in[51] ^ in2[51];
    assign G[41] = in[50] & in2[50];
    assign P[41] = in[50] ^ in2[50];
    assign G[42] = in[49] & in2[49];
    assign P[42] = in[49] ^ in2[49];
    assign G[43] = in[48] & in2[48];
    assign P[43] = in[48] ^ in2[48];
    assign G[44] = in[47] & in2[47];
    assign P[44] = in[47] ^ in2[47];
    assign G[45] = in[46] & in2[46];
    assign P[45] = in[46] ^ in2[46];
    assign G[46] = in[45] & in2[45];
    assign P[46] = in[45] ^ in2[45];
    assign G[47] = in[44] & in2[44];
    assign P[47] = in[44] ^ in2[44];
    assign G[48] = in[43] & in2[43];
    assign P[48] = in[43] ^ in2[43];
    assign G[49] = in[42] & in2[42];
    assign P[49] = in[42] ^ in2[42];
    assign G[50] = in[41] & in2[41];
    assign P[50] = in[41] ^ in2[41];
    assign G[51] = in[40] & in2[40];
    assign P[51] = in[40] ^ in2[40];
    assign G[52] = in[39] & in2[39];
    assign P[52] = in[39] ^ in2[39];
    assign G[53] = in[38] & in2[38];
    assign P[53] = in[38] ^ in2[38];
    assign G[54] = in[37] & in2[37];
    assign P[54] = in[37] ^ in2[37];
    assign G[55] = in[36] & in2[36];
    assign P[55] = in[36] ^ in2[36];
    assign G[56] = in[35] & in2[35];
    assign P[56] = in[35] ^ in2[35];
    assign G[57] = in[34] & in2[34];
    assign P[57] = in[34] ^ in2[34];
    assign G[58] = in[33] & in2[33];
    assign P[58] = in[33] ^ in2[33];
    assign G[59] = in[32] & in2[32];
    assign P[59] = in[32] ^ in2[32];
    assign G[60] = in[31] & in2[31];
    assign P[60] = in[31] ^ in2[31];
    assign G[61] = in[30] & in2[30];
    assign P[61] = in[30] ^ in2[30];
    assign G[62] = in[29] & in2[29];
    assign P[62] = in[29] ^ in2[29];
    assign G[63] = in[28] & in2[28];
    assign P[63] = in[28] ^ in2[28];
    assign G[64] = in[27] & in2[27];
    assign P[64] = in[27] ^ in2[27];
    assign G[65] = in[26] & in2[26];
    assign P[65] = in[26] ^ in2[26];
    assign G[66] = in[25] & in2[25];
    assign P[66] = in[25] ^ in2[25];
    assign G[67] = in[24] & in2[24];
    assign P[67] = in[24] ^ in2[24];
    assign G[68] = in[23] & in2[23];
    assign P[68] = in[23] ^ in2[23];
    assign G[69] = in[22] & in2[22];
    assign P[69] = in[22] ^ in2[22];
    assign G[70] = in[21] & in2[21];
    assign P[70] = in[21] ^ in2[21];
    assign G[71] = in[20] & in2[20];
    assign P[71] = in[20] ^ in2[20];
    assign G[72] = in[19] & in2[19];
    assign P[72] = in[19] ^ in2[19];
    assign G[73] = in[18] & in2[18];
    assign P[73] = in[18] ^ in2[18];
    assign G[74] = in[17] & in2[17];
    assign P[74] = in[17] ^ in2[17];
    assign G[75] = in[16] & in2[16];
    assign P[75] = in[16] ^ in2[16];
    assign G[76] = in[15] & in2[15];
    assign P[76] = in[15] ^ in2[15];
    assign G[77] = in[14] & in2[14];
    assign P[77] = in[14] ^ in2[14];
    assign G[78] = in[13] & in2[13];
    assign P[78] = in[13] ^ in2[13];
    assign G[79] = in[12] & in2[12];
    assign P[79] = in[12] ^ in2[12];
    assign G[80] = in[11] & in2[11];
    assign P[80] = in[11] ^ in2[11];
    assign G[81] = in[10] & in2[10];
    assign P[81] = in[10] ^ in2[10];
    assign G[82] = in[9] & in2[9];
    assign P[82] = in[9] ^ in2[9];
    assign G[83] = in[8] & in2[8];
    assign P[83] = in[8] ^ in2[8];
    assign G[84] = in[7] & in2[7];
    assign P[84] = in[7] ^ in2[7];
    assign G[85] = in[6] & in2[6];
    assign P[85] = in[6] ^ in2[6];
    assign G[86] = in[5] & in2[5];
    assign P[86] = in[5] ^ in2[5];
    assign G[87] = in[4] & in2[4];
    assign P[87] = in[4] ^ in2[4];
    assign G[88] = in[3] & in2[3];
    assign P[88] = in[3] ^ in2[3];
    assign G[89] = in[2] & in2[2];
    assign P[89] = in[2] ^ in2[2];
    assign G[90] = in[1] & in2[1];
    assign P[90] = in[1] ^ in2[1];
    assign G[91] = in[0] & in2[0];
    assign P[91] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign C[91] = G[90] | (P[90] & C[90]);
    assign cout = G[91] | (P[91] & C[91]);
    assign sum = P ^ C;
endmodule

module CLA91(output [90:0] sum, output cout, input [90:0] in1, input [90:0] in2;

    wire[90:0] G;
    wire[90:0] C;
    wire[90:0] P;

    assign G[0] = in[90] & in2[90];
    assign P[0] = in[90] ^ in2[90];
    assign G[1] = in[89] & in2[89];
    assign P[1] = in[89] ^ in2[89];
    assign G[2] = in[88] & in2[88];
    assign P[2] = in[88] ^ in2[88];
    assign G[3] = in[87] & in2[87];
    assign P[3] = in[87] ^ in2[87];
    assign G[4] = in[86] & in2[86];
    assign P[4] = in[86] ^ in2[86];
    assign G[5] = in[85] & in2[85];
    assign P[5] = in[85] ^ in2[85];
    assign G[6] = in[84] & in2[84];
    assign P[6] = in[84] ^ in2[84];
    assign G[7] = in[83] & in2[83];
    assign P[7] = in[83] ^ in2[83];
    assign G[8] = in[82] & in2[82];
    assign P[8] = in[82] ^ in2[82];
    assign G[9] = in[81] & in2[81];
    assign P[9] = in[81] ^ in2[81];
    assign G[10] = in[80] & in2[80];
    assign P[10] = in[80] ^ in2[80];
    assign G[11] = in[79] & in2[79];
    assign P[11] = in[79] ^ in2[79];
    assign G[12] = in[78] & in2[78];
    assign P[12] = in[78] ^ in2[78];
    assign G[13] = in[77] & in2[77];
    assign P[13] = in[77] ^ in2[77];
    assign G[14] = in[76] & in2[76];
    assign P[14] = in[76] ^ in2[76];
    assign G[15] = in[75] & in2[75];
    assign P[15] = in[75] ^ in2[75];
    assign G[16] = in[74] & in2[74];
    assign P[16] = in[74] ^ in2[74];
    assign G[17] = in[73] & in2[73];
    assign P[17] = in[73] ^ in2[73];
    assign G[18] = in[72] & in2[72];
    assign P[18] = in[72] ^ in2[72];
    assign G[19] = in[71] & in2[71];
    assign P[19] = in[71] ^ in2[71];
    assign G[20] = in[70] & in2[70];
    assign P[20] = in[70] ^ in2[70];
    assign G[21] = in[69] & in2[69];
    assign P[21] = in[69] ^ in2[69];
    assign G[22] = in[68] & in2[68];
    assign P[22] = in[68] ^ in2[68];
    assign G[23] = in[67] & in2[67];
    assign P[23] = in[67] ^ in2[67];
    assign G[24] = in[66] & in2[66];
    assign P[24] = in[66] ^ in2[66];
    assign G[25] = in[65] & in2[65];
    assign P[25] = in[65] ^ in2[65];
    assign G[26] = in[64] & in2[64];
    assign P[26] = in[64] ^ in2[64];
    assign G[27] = in[63] & in2[63];
    assign P[27] = in[63] ^ in2[63];
    assign G[28] = in[62] & in2[62];
    assign P[28] = in[62] ^ in2[62];
    assign G[29] = in[61] & in2[61];
    assign P[29] = in[61] ^ in2[61];
    assign G[30] = in[60] & in2[60];
    assign P[30] = in[60] ^ in2[60];
    assign G[31] = in[59] & in2[59];
    assign P[31] = in[59] ^ in2[59];
    assign G[32] = in[58] & in2[58];
    assign P[32] = in[58] ^ in2[58];
    assign G[33] = in[57] & in2[57];
    assign P[33] = in[57] ^ in2[57];
    assign G[34] = in[56] & in2[56];
    assign P[34] = in[56] ^ in2[56];
    assign G[35] = in[55] & in2[55];
    assign P[35] = in[55] ^ in2[55];
    assign G[36] = in[54] & in2[54];
    assign P[36] = in[54] ^ in2[54];
    assign G[37] = in[53] & in2[53];
    assign P[37] = in[53] ^ in2[53];
    assign G[38] = in[52] & in2[52];
    assign P[38] = in[52] ^ in2[52];
    assign G[39] = in[51] & in2[51];
    assign P[39] = in[51] ^ in2[51];
    assign G[40] = in[50] & in2[50];
    assign P[40] = in[50] ^ in2[50];
    assign G[41] = in[49] & in2[49];
    assign P[41] = in[49] ^ in2[49];
    assign G[42] = in[48] & in2[48];
    assign P[42] = in[48] ^ in2[48];
    assign G[43] = in[47] & in2[47];
    assign P[43] = in[47] ^ in2[47];
    assign G[44] = in[46] & in2[46];
    assign P[44] = in[46] ^ in2[46];
    assign G[45] = in[45] & in2[45];
    assign P[45] = in[45] ^ in2[45];
    assign G[46] = in[44] & in2[44];
    assign P[46] = in[44] ^ in2[44];
    assign G[47] = in[43] & in2[43];
    assign P[47] = in[43] ^ in2[43];
    assign G[48] = in[42] & in2[42];
    assign P[48] = in[42] ^ in2[42];
    assign G[49] = in[41] & in2[41];
    assign P[49] = in[41] ^ in2[41];
    assign G[50] = in[40] & in2[40];
    assign P[50] = in[40] ^ in2[40];
    assign G[51] = in[39] & in2[39];
    assign P[51] = in[39] ^ in2[39];
    assign G[52] = in[38] & in2[38];
    assign P[52] = in[38] ^ in2[38];
    assign G[53] = in[37] & in2[37];
    assign P[53] = in[37] ^ in2[37];
    assign G[54] = in[36] & in2[36];
    assign P[54] = in[36] ^ in2[36];
    assign G[55] = in[35] & in2[35];
    assign P[55] = in[35] ^ in2[35];
    assign G[56] = in[34] & in2[34];
    assign P[56] = in[34] ^ in2[34];
    assign G[57] = in[33] & in2[33];
    assign P[57] = in[33] ^ in2[33];
    assign G[58] = in[32] & in2[32];
    assign P[58] = in[32] ^ in2[32];
    assign G[59] = in[31] & in2[31];
    assign P[59] = in[31] ^ in2[31];
    assign G[60] = in[30] & in2[30];
    assign P[60] = in[30] ^ in2[30];
    assign G[61] = in[29] & in2[29];
    assign P[61] = in[29] ^ in2[29];
    assign G[62] = in[28] & in2[28];
    assign P[62] = in[28] ^ in2[28];
    assign G[63] = in[27] & in2[27];
    assign P[63] = in[27] ^ in2[27];
    assign G[64] = in[26] & in2[26];
    assign P[64] = in[26] ^ in2[26];
    assign G[65] = in[25] & in2[25];
    assign P[65] = in[25] ^ in2[25];
    assign G[66] = in[24] & in2[24];
    assign P[66] = in[24] ^ in2[24];
    assign G[67] = in[23] & in2[23];
    assign P[67] = in[23] ^ in2[23];
    assign G[68] = in[22] & in2[22];
    assign P[68] = in[22] ^ in2[22];
    assign G[69] = in[21] & in2[21];
    assign P[69] = in[21] ^ in2[21];
    assign G[70] = in[20] & in2[20];
    assign P[70] = in[20] ^ in2[20];
    assign G[71] = in[19] & in2[19];
    assign P[71] = in[19] ^ in2[19];
    assign G[72] = in[18] & in2[18];
    assign P[72] = in[18] ^ in2[18];
    assign G[73] = in[17] & in2[17];
    assign P[73] = in[17] ^ in2[17];
    assign G[74] = in[16] & in2[16];
    assign P[74] = in[16] ^ in2[16];
    assign G[75] = in[15] & in2[15];
    assign P[75] = in[15] ^ in2[15];
    assign G[76] = in[14] & in2[14];
    assign P[76] = in[14] ^ in2[14];
    assign G[77] = in[13] & in2[13];
    assign P[77] = in[13] ^ in2[13];
    assign G[78] = in[12] & in2[12];
    assign P[78] = in[12] ^ in2[12];
    assign G[79] = in[11] & in2[11];
    assign P[79] = in[11] ^ in2[11];
    assign G[80] = in[10] & in2[10];
    assign P[80] = in[10] ^ in2[10];
    assign G[81] = in[9] & in2[9];
    assign P[81] = in[9] ^ in2[9];
    assign G[82] = in[8] & in2[8];
    assign P[82] = in[8] ^ in2[8];
    assign G[83] = in[7] & in2[7];
    assign P[83] = in[7] ^ in2[7];
    assign G[84] = in[6] & in2[6];
    assign P[84] = in[6] ^ in2[6];
    assign G[85] = in[5] & in2[5];
    assign P[85] = in[5] ^ in2[5];
    assign G[86] = in[4] & in2[4];
    assign P[86] = in[4] ^ in2[4];
    assign G[87] = in[3] & in2[3];
    assign P[87] = in[3] ^ in2[3];
    assign G[88] = in[2] & in2[2];
    assign P[88] = in[2] ^ in2[2];
    assign G[89] = in[1] & in2[1];
    assign P[89] = in[1] ^ in2[1];
    assign G[90] = in[0] & in2[0];
    assign P[90] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign C[90] = G[89] | (P[89] & C[89]);
    assign cout = G[90] | (P[90] & C[90]);
    assign sum = P ^ C;
endmodule

module CLA90(output [89:0] sum, output cout, input [89:0] in1, input [89:0] in2;

    wire[89:0] G;
    wire[89:0] C;
    wire[89:0] P;

    assign G[0] = in[89] & in2[89];
    assign P[0] = in[89] ^ in2[89];
    assign G[1] = in[88] & in2[88];
    assign P[1] = in[88] ^ in2[88];
    assign G[2] = in[87] & in2[87];
    assign P[2] = in[87] ^ in2[87];
    assign G[3] = in[86] & in2[86];
    assign P[3] = in[86] ^ in2[86];
    assign G[4] = in[85] & in2[85];
    assign P[4] = in[85] ^ in2[85];
    assign G[5] = in[84] & in2[84];
    assign P[5] = in[84] ^ in2[84];
    assign G[6] = in[83] & in2[83];
    assign P[6] = in[83] ^ in2[83];
    assign G[7] = in[82] & in2[82];
    assign P[7] = in[82] ^ in2[82];
    assign G[8] = in[81] & in2[81];
    assign P[8] = in[81] ^ in2[81];
    assign G[9] = in[80] & in2[80];
    assign P[9] = in[80] ^ in2[80];
    assign G[10] = in[79] & in2[79];
    assign P[10] = in[79] ^ in2[79];
    assign G[11] = in[78] & in2[78];
    assign P[11] = in[78] ^ in2[78];
    assign G[12] = in[77] & in2[77];
    assign P[12] = in[77] ^ in2[77];
    assign G[13] = in[76] & in2[76];
    assign P[13] = in[76] ^ in2[76];
    assign G[14] = in[75] & in2[75];
    assign P[14] = in[75] ^ in2[75];
    assign G[15] = in[74] & in2[74];
    assign P[15] = in[74] ^ in2[74];
    assign G[16] = in[73] & in2[73];
    assign P[16] = in[73] ^ in2[73];
    assign G[17] = in[72] & in2[72];
    assign P[17] = in[72] ^ in2[72];
    assign G[18] = in[71] & in2[71];
    assign P[18] = in[71] ^ in2[71];
    assign G[19] = in[70] & in2[70];
    assign P[19] = in[70] ^ in2[70];
    assign G[20] = in[69] & in2[69];
    assign P[20] = in[69] ^ in2[69];
    assign G[21] = in[68] & in2[68];
    assign P[21] = in[68] ^ in2[68];
    assign G[22] = in[67] & in2[67];
    assign P[22] = in[67] ^ in2[67];
    assign G[23] = in[66] & in2[66];
    assign P[23] = in[66] ^ in2[66];
    assign G[24] = in[65] & in2[65];
    assign P[24] = in[65] ^ in2[65];
    assign G[25] = in[64] & in2[64];
    assign P[25] = in[64] ^ in2[64];
    assign G[26] = in[63] & in2[63];
    assign P[26] = in[63] ^ in2[63];
    assign G[27] = in[62] & in2[62];
    assign P[27] = in[62] ^ in2[62];
    assign G[28] = in[61] & in2[61];
    assign P[28] = in[61] ^ in2[61];
    assign G[29] = in[60] & in2[60];
    assign P[29] = in[60] ^ in2[60];
    assign G[30] = in[59] & in2[59];
    assign P[30] = in[59] ^ in2[59];
    assign G[31] = in[58] & in2[58];
    assign P[31] = in[58] ^ in2[58];
    assign G[32] = in[57] & in2[57];
    assign P[32] = in[57] ^ in2[57];
    assign G[33] = in[56] & in2[56];
    assign P[33] = in[56] ^ in2[56];
    assign G[34] = in[55] & in2[55];
    assign P[34] = in[55] ^ in2[55];
    assign G[35] = in[54] & in2[54];
    assign P[35] = in[54] ^ in2[54];
    assign G[36] = in[53] & in2[53];
    assign P[36] = in[53] ^ in2[53];
    assign G[37] = in[52] & in2[52];
    assign P[37] = in[52] ^ in2[52];
    assign G[38] = in[51] & in2[51];
    assign P[38] = in[51] ^ in2[51];
    assign G[39] = in[50] & in2[50];
    assign P[39] = in[50] ^ in2[50];
    assign G[40] = in[49] & in2[49];
    assign P[40] = in[49] ^ in2[49];
    assign G[41] = in[48] & in2[48];
    assign P[41] = in[48] ^ in2[48];
    assign G[42] = in[47] & in2[47];
    assign P[42] = in[47] ^ in2[47];
    assign G[43] = in[46] & in2[46];
    assign P[43] = in[46] ^ in2[46];
    assign G[44] = in[45] & in2[45];
    assign P[44] = in[45] ^ in2[45];
    assign G[45] = in[44] & in2[44];
    assign P[45] = in[44] ^ in2[44];
    assign G[46] = in[43] & in2[43];
    assign P[46] = in[43] ^ in2[43];
    assign G[47] = in[42] & in2[42];
    assign P[47] = in[42] ^ in2[42];
    assign G[48] = in[41] & in2[41];
    assign P[48] = in[41] ^ in2[41];
    assign G[49] = in[40] & in2[40];
    assign P[49] = in[40] ^ in2[40];
    assign G[50] = in[39] & in2[39];
    assign P[50] = in[39] ^ in2[39];
    assign G[51] = in[38] & in2[38];
    assign P[51] = in[38] ^ in2[38];
    assign G[52] = in[37] & in2[37];
    assign P[52] = in[37] ^ in2[37];
    assign G[53] = in[36] & in2[36];
    assign P[53] = in[36] ^ in2[36];
    assign G[54] = in[35] & in2[35];
    assign P[54] = in[35] ^ in2[35];
    assign G[55] = in[34] & in2[34];
    assign P[55] = in[34] ^ in2[34];
    assign G[56] = in[33] & in2[33];
    assign P[56] = in[33] ^ in2[33];
    assign G[57] = in[32] & in2[32];
    assign P[57] = in[32] ^ in2[32];
    assign G[58] = in[31] & in2[31];
    assign P[58] = in[31] ^ in2[31];
    assign G[59] = in[30] & in2[30];
    assign P[59] = in[30] ^ in2[30];
    assign G[60] = in[29] & in2[29];
    assign P[60] = in[29] ^ in2[29];
    assign G[61] = in[28] & in2[28];
    assign P[61] = in[28] ^ in2[28];
    assign G[62] = in[27] & in2[27];
    assign P[62] = in[27] ^ in2[27];
    assign G[63] = in[26] & in2[26];
    assign P[63] = in[26] ^ in2[26];
    assign G[64] = in[25] & in2[25];
    assign P[64] = in[25] ^ in2[25];
    assign G[65] = in[24] & in2[24];
    assign P[65] = in[24] ^ in2[24];
    assign G[66] = in[23] & in2[23];
    assign P[66] = in[23] ^ in2[23];
    assign G[67] = in[22] & in2[22];
    assign P[67] = in[22] ^ in2[22];
    assign G[68] = in[21] & in2[21];
    assign P[68] = in[21] ^ in2[21];
    assign G[69] = in[20] & in2[20];
    assign P[69] = in[20] ^ in2[20];
    assign G[70] = in[19] & in2[19];
    assign P[70] = in[19] ^ in2[19];
    assign G[71] = in[18] & in2[18];
    assign P[71] = in[18] ^ in2[18];
    assign G[72] = in[17] & in2[17];
    assign P[72] = in[17] ^ in2[17];
    assign G[73] = in[16] & in2[16];
    assign P[73] = in[16] ^ in2[16];
    assign G[74] = in[15] & in2[15];
    assign P[74] = in[15] ^ in2[15];
    assign G[75] = in[14] & in2[14];
    assign P[75] = in[14] ^ in2[14];
    assign G[76] = in[13] & in2[13];
    assign P[76] = in[13] ^ in2[13];
    assign G[77] = in[12] & in2[12];
    assign P[77] = in[12] ^ in2[12];
    assign G[78] = in[11] & in2[11];
    assign P[78] = in[11] ^ in2[11];
    assign G[79] = in[10] & in2[10];
    assign P[79] = in[10] ^ in2[10];
    assign G[80] = in[9] & in2[9];
    assign P[80] = in[9] ^ in2[9];
    assign G[81] = in[8] & in2[8];
    assign P[81] = in[8] ^ in2[8];
    assign G[82] = in[7] & in2[7];
    assign P[82] = in[7] ^ in2[7];
    assign G[83] = in[6] & in2[6];
    assign P[83] = in[6] ^ in2[6];
    assign G[84] = in[5] & in2[5];
    assign P[84] = in[5] ^ in2[5];
    assign G[85] = in[4] & in2[4];
    assign P[85] = in[4] ^ in2[4];
    assign G[86] = in[3] & in2[3];
    assign P[86] = in[3] ^ in2[3];
    assign G[87] = in[2] & in2[2];
    assign P[87] = in[2] ^ in2[2];
    assign G[88] = in[1] & in2[1];
    assign P[88] = in[1] ^ in2[1];
    assign G[89] = in[0] & in2[0];
    assign P[89] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign C[89] = G[88] | (P[88] & C[88]);
    assign cout = G[89] | (P[89] & C[89]);
    assign sum = P ^ C;
endmodule

module CLA89(output [88:0] sum, output cout, input [88:0] in1, input [88:0] in2;

    wire[88:0] G;
    wire[88:0] C;
    wire[88:0] P;

    assign G[0] = in[88] & in2[88];
    assign P[0] = in[88] ^ in2[88];
    assign G[1] = in[87] & in2[87];
    assign P[1] = in[87] ^ in2[87];
    assign G[2] = in[86] & in2[86];
    assign P[2] = in[86] ^ in2[86];
    assign G[3] = in[85] & in2[85];
    assign P[3] = in[85] ^ in2[85];
    assign G[4] = in[84] & in2[84];
    assign P[4] = in[84] ^ in2[84];
    assign G[5] = in[83] & in2[83];
    assign P[5] = in[83] ^ in2[83];
    assign G[6] = in[82] & in2[82];
    assign P[6] = in[82] ^ in2[82];
    assign G[7] = in[81] & in2[81];
    assign P[7] = in[81] ^ in2[81];
    assign G[8] = in[80] & in2[80];
    assign P[8] = in[80] ^ in2[80];
    assign G[9] = in[79] & in2[79];
    assign P[9] = in[79] ^ in2[79];
    assign G[10] = in[78] & in2[78];
    assign P[10] = in[78] ^ in2[78];
    assign G[11] = in[77] & in2[77];
    assign P[11] = in[77] ^ in2[77];
    assign G[12] = in[76] & in2[76];
    assign P[12] = in[76] ^ in2[76];
    assign G[13] = in[75] & in2[75];
    assign P[13] = in[75] ^ in2[75];
    assign G[14] = in[74] & in2[74];
    assign P[14] = in[74] ^ in2[74];
    assign G[15] = in[73] & in2[73];
    assign P[15] = in[73] ^ in2[73];
    assign G[16] = in[72] & in2[72];
    assign P[16] = in[72] ^ in2[72];
    assign G[17] = in[71] & in2[71];
    assign P[17] = in[71] ^ in2[71];
    assign G[18] = in[70] & in2[70];
    assign P[18] = in[70] ^ in2[70];
    assign G[19] = in[69] & in2[69];
    assign P[19] = in[69] ^ in2[69];
    assign G[20] = in[68] & in2[68];
    assign P[20] = in[68] ^ in2[68];
    assign G[21] = in[67] & in2[67];
    assign P[21] = in[67] ^ in2[67];
    assign G[22] = in[66] & in2[66];
    assign P[22] = in[66] ^ in2[66];
    assign G[23] = in[65] & in2[65];
    assign P[23] = in[65] ^ in2[65];
    assign G[24] = in[64] & in2[64];
    assign P[24] = in[64] ^ in2[64];
    assign G[25] = in[63] & in2[63];
    assign P[25] = in[63] ^ in2[63];
    assign G[26] = in[62] & in2[62];
    assign P[26] = in[62] ^ in2[62];
    assign G[27] = in[61] & in2[61];
    assign P[27] = in[61] ^ in2[61];
    assign G[28] = in[60] & in2[60];
    assign P[28] = in[60] ^ in2[60];
    assign G[29] = in[59] & in2[59];
    assign P[29] = in[59] ^ in2[59];
    assign G[30] = in[58] & in2[58];
    assign P[30] = in[58] ^ in2[58];
    assign G[31] = in[57] & in2[57];
    assign P[31] = in[57] ^ in2[57];
    assign G[32] = in[56] & in2[56];
    assign P[32] = in[56] ^ in2[56];
    assign G[33] = in[55] & in2[55];
    assign P[33] = in[55] ^ in2[55];
    assign G[34] = in[54] & in2[54];
    assign P[34] = in[54] ^ in2[54];
    assign G[35] = in[53] & in2[53];
    assign P[35] = in[53] ^ in2[53];
    assign G[36] = in[52] & in2[52];
    assign P[36] = in[52] ^ in2[52];
    assign G[37] = in[51] & in2[51];
    assign P[37] = in[51] ^ in2[51];
    assign G[38] = in[50] & in2[50];
    assign P[38] = in[50] ^ in2[50];
    assign G[39] = in[49] & in2[49];
    assign P[39] = in[49] ^ in2[49];
    assign G[40] = in[48] & in2[48];
    assign P[40] = in[48] ^ in2[48];
    assign G[41] = in[47] & in2[47];
    assign P[41] = in[47] ^ in2[47];
    assign G[42] = in[46] & in2[46];
    assign P[42] = in[46] ^ in2[46];
    assign G[43] = in[45] & in2[45];
    assign P[43] = in[45] ^ in2[45];
    assign G[44] = in[44] & in2[44];
    assign P[44] = in[44] ^ in2[44];
    assign G[45] = in[43] & in2[43];
    assign P[45] = in[43] ^ in2[43];
    assign G[46] = in[42] & in2[42];
    assign P[46] = in[42] ^ in2[42];
    assign G[47] = in[41] & in2[41];
    assign P[47] = in[41] ^ in2[41];
    assign G[48] = in[40] & in2[40];
    assign P[48] = in[40] ^ in2[40];
    assign G[49] = in[39] & in2[39];
    assign P[49] = in[39] ^ in2[39];
    assign G[50] = in[38] & in2[38];
    assign P[50] = in[38] ^ in2[38];
    assign G[51] = in[37] & in2[37];
    assign P[51] = in[37] ^ in2[37];
    assign G[52] = in[36] & in2[36];
    assign P[52] = in[36] ^ in2[36];
    assign G[53] = in[35] & in2[35];
    assign P[53] = in[35] ^ in2[35];
    assign G[54] = in[34] & in2[34];
    assign P[54] = in[34] ^ in2[34];
    assign G[55] = in[33] & in2[33];
    assign P[55] = in[33] ^ in2[33];
    assign G[56] = in[32] & in2[32];
    assign P[56] = in[32] ^ in2[32];
    assign G[57] = in[31] & in2[31];
    assign P[57] = in[31] ^ in2[31];
    assign G[58] = in[30] & in2[30];
    assign P[58] = in[30] ^ in2[30];
    assign G[59] = in[29] & in2[29];
    assign P[59] = in[29] ^ in2[29];
    assign G[60] = in[28] & in2[28];
    assign P[60] = in[28] ^ in2[28];
    assign G[61] = in[27] & in2[27];
    assign P[61] = in[27] ^ in2[27];
    assign G[62] = in[26] & in2[26];
    assign P[62] = in[26] ^ in2[26];
    assign G[63] = in[25] & in2[25];
    assign P[63] = in[25] ^ in2[25];
    assign G[64] = in[24] & in2[24];
    assign P[64] = in[24] ^ in2[24];
    assign G[65] = in[23] & in2[23];
    assign P[65] = in[23] ^ in2[23];
    assign G[66] = in[22] & in2[22];
    assign P[66] = in[22] ^ in2[22];
    assign G[67] = in[21] & in2[21];
    assign P[67] = in[21] ^ in2[21];
    assign G[68] = in[20] & in2[20];
    assign P[68] = in[20] ^ in2[20];
    assign G[69] = in[19] & in2[19];
    assign P[69] = in[19] ^ in2[19];
    assign G[70] = in[18] & in2[18];
    assign P[70] = in[18] ^ in2[18];
    assign G[71] = in[17] & in2[17];
    assign P[71] = in[17] ^ in2[17];
    assign G[72] = in[16] & in2[16];
    assign P[72] = in[16] ^ in2[16];
    assign G[73] = in[15] & in2[15];
    assign P[73] = in[15] ^ in2[15];
    assign G[74] = in[14] & in2[14];
    assign P[74] = in[14] ^ in2[14];
    assign G[75] = in[13] & in2[13];
    assign P[75] = in[13] ^ in2[13];
    assign G[76] = in[12] & in2[12];
    assign P[76] = in[12] ^ in2[12];
    assign G[77] = in[11] & in2[11];
    assign P[77] = in[11] ^ in2[11];
    assign G[78] = in[10] & in2[10];
    assign P[78] = in[10] ^ in2[10];
    assign G[79] = in[9] & in2[9];
    assign P[79] = in[9] ^ in2[9];
    assign G[80] = in[8] & in2[8];
    assign P[80] = in[8] ^ in2[8];
    assign G[81] = in[7] & in2[7];
    assign P[81] = in[7] ^ in2[7];
    assign G[82] = in[6] & in2[6];
    assign P[82] = in[6] ^ in2[6];
    assign G[83] = in[5] & in2[5];
    assign P[83] = in[5] ^ in2[5];
    assign G[84] = in[4] & in2[4];
    assign P[84] = in[4] ^ in2[4];
    assign G[85] = in[3] & in2[3];
    assign P[85] = in[3] ^ in2[3];
    assign G[86] = in[2] & in2[2];
    assign P[86] = in[2] ^ in2[2];
    assign G[87] = in[1] & in2[1];
    assign P[87] = in[1] ^ in2[1];
    assign G[88] = in[0] & in2[0];
    assign P[88] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign C[88] = G[87] | (P[87] & C[87]);
    assign cout = G[88] | (P[88] & C[88]);
    assign sum = P ^ C;
endmodule

module CLA88(output [87:0] sum, output cout, input [87:0] in1, input [87:0] in2;

    wire[87:0] G;
    wire[87:0] C;
    wire[87:0] P;

    assign G[0] = in[87] & in2[87];
    assign P[0] = in[87] ^ in2[87];
    assign G[1] = in[86] & in2[86];
    assign P[1] = in[86] ^ in2[86];
    assign G[2] = in[85] & in2[85];
    assign P[2] = in[85] ^ in2[85];
    assign G[3] = in[84] & in2[84];
    assign P[3] = in[84] ^ in2[84];
    assign G[4] = in[83] & in2[83];
    assign P[4] = in[83] ^ in2[83];
    assign G[5] = in[82] & in2[82];
    assign P[5] = in[82] ^ in2[82];
    assign G[6] = in[81] & in2[81];
    assign P[6] = in[81] ^ in2[81];
    assign G[7] = in[80] & in2[80];
    assign P[7] = in[80] ^ in2[80];
    assign G[8] = in[79] & in2[79];
    assign P[8] = in[79] ^ in2[79];
    assign G[9] = in[78] & in2[78];
    assign P[9] = in[78] ^ in2[78];
    assign G[10] = in[77] & in2[77];
    assign P[10] = in[77] ^ in2[77];
    assign G[11] = in[76] & in2[76];
    assign P[11] = in[76] ^ in2[76];
    assign G[12] = in[75] & in2[75];
    assign P[12] = in[75] ^ in2[75];
    assign G[13] = in[74] & in2[74];
    assign P[13] = in[74] ^ in2[74];
    assign G[14] = in[73] & in2[73];
    assign P[14] = in[73] ^ in2[73];
    assign G[15] = in[72] & in2[72];
    assign P[15] = in[72] ^ in2[72];
    assign G[16] = in[71] & in2[71];
    assign P[16] = in[71] ^ in2[71];
    assign G[17] = in[70] & in2[70];
    assign P[17] = in[70] ^ in2[70];
    assign G[18] = in[69] & in2[69];
    assign P[18] = in[69] ^ in2[69];
    assign G[19] = in[68] & in2[68];
    assign P[19] = in[68] ^ in2[68];
    assign G[20] = in[67] & in2[67];
    assign P[20] = in[67] ^ in2[67];
    assign G[21] = in[66] & in2[66];
    assign P[21] = in[66] ^ in2[66];
    assign G[22] = in[65] & in2[65];
    assign P[22] = in[65] ^ in2[65];
    assign G[23] = in[64] & in2[64];
    assign P[23] = in[64] ^ in2[64];
    assign G[24] = in[63] & in2[63];
    assign P[24] = in[63] ^ in2[63];
    assign G[25] = in[62] & in2[62];
    assign P[25] = in[62] ^ in2[62];
    assign G[26] = in[61] & in2[61];
    assign P[26] = in[61] ^ in2[61];
    assign G[27] = in[60] & in2[60];
    assign P[27] = in[60] ^ in2[60];
    assign G[28] = in[59] & in2[59];
    assign P[28] = in[59] ^ in2[59];
    assign G[29] = in[58] & in2[58];
    assign P[29] = in[58] ^ in2[58];
    assign G[30] = in[57] & in2[57];
    assign P[30] = in[57] ^ in2[57];
    assign G[31] = in[56] & in2[56];
    assign P[31] = in[56] ^ in2[56];
    assign G[32] = in[55] & in2[55];
    assign P[32] = in[55] ^ in2[55];
    assign G[33] = in[54] & in2[54];
    assign P[33] = in[54] ^ in2[54];
    assign G[34] = in[53] & in2[53];
    assign P[34] = in[53] ^ in2[53];
    assign G[35] = in[52] & in2[52];
    assign P[35] = in[52] ^ in2[52];
    assign G[36] = in[51] & in2[51];
    assign P[36] = in[51] ^ in2[51];
    assign G[37] = in[50] & in2[50];
    assign P[37] = in[50] ^ in2[50];
    assign G[38] = in[49] & in2[49];
    assign P[38] = in[49] ^ in2[49];
    assign G[39] = in[48] & in2[48];
    assign P[39] = in[48] ^ in2[48];
    assign G[40] = in[47] & in2[47];
    assign P[40] = in[47] ^ in2[47];
    assign G[41] = in[46] & in2[46];
    assign P[41] = in[46] ^ in2[46];
    assign G[42] = in[45] & in2[45];
    assign P[42] = in[45] ^ in2[45];
    assign G[43] = in[44] & in2[44];
    assign P[43] = in[44] ^ in2[44];
    assign G[44] = in[43] & in2[43];
    assign P[44] = in[43] ^ in2[43];
    assign G[45] = in[42] & in2[42];
    assign P[45] = in[42] ^ in2[42];
    assign G[46] = in[41] & in2[41];
    assign P[46] = in[41] ^ in2[41];
    assign G[47] = in[40] & in2[40];
    assign P[47] = in[40] ^ in2[40];
    assign G[48] = in[39] & in2[39];
    assign P[48] = in[39] ^ in2[39];
    assign G[49] = in[38] & in2[38];
    assign P[49] = in[38] ^ in2[38];
    assign G[50] = in[37] & in2[37];
    assign P[50] = in[37] ^ in2[37];
    assign G[51] = in[36] & in2[36];
    assign P[51] = in[36] ^ in2[36];
    assign G[52] = in[35] & in2[35];
    assign P[52] = in[35] ^ in2[35];
    assign G[53] = in[34] & in2[34];
    assign P[53] = in[34] ^ in2[34];
    assign G[54] = in[33] & in2[33];
    assign P[54] = in[33] ^ in2[33];
    assign G[55] = in[32] & in2[32];
    assign P[55] = in[32] ^ in2[32];
    assign G[56] = in[31] & in2[31];
    assign P[56] = in[31] ^ in2[31];
    assign G[57] = in[30] & in2[30];
    assign P[57] = in[30] ^ in2[30];
    assign G[58] = in[29] & in2[29];
    assign P[58] = in[29] ^ in2[29];
    assign G[59] = in[28] & in2[28];
    assign P[59] = in[28] ^ in2[28];
    assign G[60] = in[27] & in2[27];
    assign P[60] = in[27] ^ in2[27];
    assign G[61] = in[26] & in2[26];
    assign P[61] = in[26] ^ in2[26];
    assign G[62] = in[25] & in2[25];
    assign P[62] = in[25] ^ in2[25];
    assign G[63] = in[24] & in2[24];
    assign P[63] = in[24] ^ in2[24];
    assign G[64] = in[23] & in2[23];
    assign P[64] = in[23] ^ in2[23];
    assign G[65] = in[22] & in2[22];
    assign P[65] = in[22] ^ in2[22];
    assign G[66] = in[21] & in2[21];
    assign P[66] = in[21] ^ in2[21];
    assign G[67] = in[20] & in2[20];
    assign P[67] = in[20] ^ in2[20];
    assign G[68] = in[19] & in2[19];
    assign P[68] = in[19] ^ in2[19];
    assign G[69] = in[18] & in2[18];
    assign P[69] = in[18] ^ in2[18];
    assign G[70] = in[17] & in2[17];
    assign P[70] = in[17] ^ in2[17];
    assign G[71] = in[16] & in2[16];
    assign P[71] = in[16] ^ in2[16];
    assign G[72] = in[15] & in2[15];
    assign P[72] = in[15] ^ in2[15];
    assign G[73] = in[14] & in2[14];
    assign P[73] = in[14] ^ in2[14];
    assign G[74] = in[13] & in2[13];
    assign P[74] = in[13] ^ in2[13];
    assign G[75] = in[12] & in2[12];
    assign P[75] = in[12] ^ in2[12];
    assign G[76] = in[11] & in2[11];
    assign P[76] = in[11] ^ in2[11];
    assign G[77] = in[10] & in2[10];
    assign P[77] = in[10] ^ in2[10];
    assign G[78] = in[9] & in2[9];
    assign P[78] = in[9] ^ in2[9];
    assign G[79] = in[8] & in2[8];
    assign P[79] = in[8] ^ in2[8];
    assign G[80] = in[7] & in2[7];
    assign P[80] = in[7] ^ in2[7];
    assign G[81] = in[6] & in2[6];
    assign P[81] = in[6] ^ in2[6];
    assign G[82] = in[5] & in2[5];
    assign P[82] = in[5] ^ in2[5];
    assign G[83] = in[4] & in2[4];
    assign P[83] = in[4] ^ in2[4];
    assign G[84] = in[3] & in2[3];
    assign P[84] = in[3] ^ in2[3];
    assign G[85] = in[2] & in2[2];
    assign P[85] = in[2] ^ in2[2];
    assign G[86] = in[1] & in2[1];
    assign P[86] = in[1] ^ in2[1];
    assign G[87] = in[0] & in2[0];
    assign P[87] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign C[87] = G[86] | (P[86] & C[86]);
    assign cout = G[87] | (P[87] & C[87]);
    assign sum = P ^ C;
endmodule

module CLA87(output [86:0] sum, output cout, input [86:0] in1, input [86:0] in2;

    wire[86:0] G;
    wire[86:0] C;
    wire[86:0] P;

    assign G[0] = in[86] & in2[86];
    assign P[0] = in[86] ^ in2[86];
    assign G[1] = in[85] & in2[85];
    assign P[1] = in[85] ^ in2[85];
    assign G[2] = in[84] & in2[84];
    assign P[2] = in[84] ^ in2[84];
    assign G[3] = in[83] & in2[83];
    assign P[3] = in[83] ^ in2[83];
    assign G[4] = in[82] & in2[82];
    assign P[4] = in[82] ^ in2[82];
    assign G[5] = in[81] & in2[81];
    assign P[5] = in[81] ^ in2[81];
    assign G[6] = in[80] & in2[80];
    assign P[6] = in[80] ^ in2[80];
    assign G[7] = in[79] & in2[79];
    assign P[7] = in[79] ^ in2[79];
    assign G[8] = in[78] & in2[78];
    assign P[8] = in[78] ^ in2[78];
    assign G[9] = in[77] & in2[77];
    assign P[9] = in[77] ^ in2[77];
    assign G[10] = in[76] & in2[76];
    assign P[10] = in[76] ^ in2[76];
    assign G[11] = in[75] & in2[75];
    assign P[11] = in[75] ^ in2[75];
    assign G[12] = in[74] & in2[74];
    assign P[12] = in[74] ^ in2[74];
    assign G[13] = in[73] & in2[73];
    assign P[13] = in[73] ^ in2[73];
    assign G[14] = in[72] & in2[72];
    assign P[14] = in[72] ^ in2[72];
    assign G[15] = in[71] & in2[71];
    assign P[15] = in[71] ^ in2[71];
    assign G[16] = in[70] & in2[70];
    assign P[16] = in[70] ^ in2[70];
    assign G[17] = in[69] & in2[69];
    assign P[17] = in[69] ^ in2[69];
    assign G[18] = in[68] & in2[68];
    assign P[18] = in[68] ^ in2[68];
    assign G[19] = in[67] & in2[67];
    assign P[19] = in[67] ^ in2[67];
    assign G[20] = in[66] & in2[66];
    assign P[20] = in[66] ^ in2[66];
    assign G[21] = in[65] & in2[65];
    assign P[21] = in[65] ^ in2[65];
    assign G[22] = in[64] & in2[64];
    assign P[22] = in[64] ^ in2[64];
    assign G[23] = in[63] & in2[63];
    assign P[23] = in[63] ^ in2[63];
    assign G[24] = in[62] & in2[62];
    assign P[24] = in[62] ^ in2[62];
    assign G[25] = in[61] & in2[61];
    assign P[25] = in[61] ^ in2[61];
    assign G[26] = in[60] & in2[60];
    assign P[26] = in[60] ^ in2[60];
    assign G[27] = in[59] & in2[59];
    assign P[27] = in[59] ^ in2[59];
    assign G[28] = in[58] & in2[58];
    assign P[28] = in[58] ^ in2[58];
    assign G[29] = in[57] & in2[57];
    assign P[29] = in[57] ^ in2[57];
    assign G[30] = in[56] & in2[56];
    assign P[30] = in[56] ^ in2[56];
    assign G[31] = in[55] & in2[55];
    assign P[31] = in[55] ^ in2[55];
    assign G[32] = in[54] & in2[54];
    assign P[32] = in[54] ^ in2[54];
    assign G[33] = in[53] & in2[53];
    assign P[33] = in[53] ^ in2[53];
    assign G[34] = in[52] & in2[52];
    assign P[34] = in[52] ^ in2[52];
    assign G[35] = in[51] & in2[51];
    assign P[35] = in[51] ^ in2[51];
    assign G[36] = in[50] & in2[50];
    assign P[36] = in[50] ^ in2[50];
    assign G[37] = in[49] & in2[49];
    assign P[37] = in[49] ^ in2[49];
    assign G[38] = in[48] & in2[48];
    assign P[38] = in[48] ^ in2[48];
    assign G[39] = in[47] & in2[47];
    assign P[39] = in[47] ^ in2[47];
    assign G[40] = in[46] & in2[46];
    assign P[40] = in[46] ^ in2[46];
    assign G[41] = in[45] & in2[45];
    assign P[41] = in[45] ^ in2[45];
    assign G[42] = in[44] & in2[44];
    assign P[42] = in[44] ^ in2[44];
    assign G[43] = in[43] & in2[43];
    assign P[43] = in[43] ^ in2[43];
    assign G[44] = in[42] & in2[42];
    assign P[44] = in[42] ^ in2[42];
    assign G[45] = in[41] & in2[41];
    assign P[45] = in[41] ^ in2[41];
    assign G[46] = in[40] & in2[40];
    assign P[46] = in[40] ^ in2[40];
    assign G[47] = in[39] & in2[39];
    assign P[47] = in[39] ^ in2[39];
    assign G[48] = in[38] & in2[38];
    assign P[48] = in[38] ^ in2[38];
    assign G[49] = in[37] & in2[37];
    assign P[49] = in[37] ^ in2[37];
    assign G[50] = in[36] & in2[36];
    assign P[50] = in[36] ^ in2[36];
    assign G[51] = in[35] & in2[35];
    assign P[51] = in[35] ^ in2[35];
    assign G[52] = in[34] & in2[34];
    assign P[52] = in[34] ^ in2[34];
    assign G[53] = in[33] & in2[33];
    assign P[53] = in[33] ^ in2[33];
    assign G[54] = in[32] & in2[32];
    assign P[54] = in[32] ^ in2[32];
    assign G[55] = in[31] & in2[31];
    assign P[55] = in[31] ^ in2[31];
    assign G[56] = in[30] & in2[30];
    assign P[56] = in[30] ^ in2[30];
    assign G[57] = in[29] & in2[29];
    assign P[57] = in[29] ^ in2[29];
    assign G[58] = in[28] & in2[28];
    assign P[58] = in[28] ^ in2[28];
    assign G[59] = in[27] & in2[27];
    assign P[59] = in[27] ^ in2[27];
    assign G[60] = in[26] & in2[26];
    assign P[60] = in[26] ^ in2[26];
    assign G[61] = in[25] & in2[25];
    assign P[61] = in[25] ^ in2[25];
    assign G[62] = in[24] & in2[24];
    assign P[62] = in[24] ^ in2[24];
    assign G[63] = in[23] & in2[23];
    assign P[63] = in[23] ^ in2[23];
    assign G[64] = in[22] & in2[22];
    assign P[64] = in[22] ^ in2[22];
    assign G[65] = in[21] & in2[21];
    assign P[65] = in[21] ^ in2[21];
    assign G[66] = in[20] & in2[20];
    assign P[66] = in[20] ^ in2[20];
    assign G[67] = in[19] & in2[19];
    assign P[67] = in[19] ^ in2[19];
    assign G[68] = in[18] & in2[18];
    assign P[68] = in[18] ^ in2[18];
    assign G[69] = in[17] & in2[17];
    assign P[69] = in[17] ^ in2[17];
    assign G[70] = in[16] & in2[16];
    assign P[70] = in[16] ^ in2[16];
    assign G[71] = in[15] & in2[15];
    assign P[71] = in[15] ^ in2[15];
    assign G[72] = in[14] & in2[14];
    assign P[72] = in[14] ^ in2[14];
    assign G[73] = in[13] & in2[13];
    assign P[73] = in[13] ^ in2[13];
    assign G[74] = in[12] & in2[12];
    assign P[74] = in[12] ^ in2[12];
    assign G[75] = in[11] & in2[11];
    assign P[75] = in[11] ^ in2[11];
    assign G[76] = in[10] & in2[10];
    assign P[76] = in[10] ^ in2[10];
    assign G[77] = in[9] & in2[9];
    assign P[77] = in[9] ^ in2[9];
    assign G[78] = in[8] & in2[8];
    assign P[78] = in[8] ^ in2[8];
    assign G[79] = in[7] & in2[7];
    assign P[79] = in[7] ^ in2[7];
    assign G[80] = in[6] & in2[6];
    assign P[80] = in[6] ^ in2[6];
    assign G[81] = in[5] & in2[5];
    assign P[81] = in[5] ^ in2[5];
    assign G[82] = in[4] & in2[4];
    assign P[82] = in[4] ^ in2[4];
    assign G[83] = in[3] & in2[3];
    assign P[83] = in[3] ^ in2[3];
    assign G[84] = in[2] & in2[2];
    assign P[84] = in[2] ^ in2[2];
    assign G[85] = in[1] & in2[1];
    assign P[85] = in[1] ^ in2[1];
    assign G[86] = in[0] & in2[0];
    assign P[86] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign C[86] = G[85] | (P[85] & C[85]);
    assign cout = G[86] | (P[86] & C[86]);
    assign sum = P ^ C;
endmodule

module CLA86(output [85:0] sum, output cout, input [85:0] in1, input [85:0] in2;

    wire[85:0] G;
    wire[85:0] C;
    wire[85:0] P;

    assign G[0] = in[85] & in2[85];
    assign P[0] = in[85] ^ in2[85];
    assign G[1] = in[84] & in2[84];
    assign P[1] = in[84] ^ in2[84];
    assign G[2] = in[83] & in2[83];
    assign P[2] = in[83] ^ in2[83];
    assign G[3] = in[82] & in2[82];
    assign P[3] = in[82] ^ in2[82];
    assign G[4] = in[81] & in2[81];
    assign P[4] = in[81] ^ in2[81];
    assign G[5] = in[80] & in2[80];
    assign P[5] = in[80] ^ in2[80];
    assign G[6] = in[79] & in2[79];
    assign P[6] = in[79] ^ in2[79];
    assign G[7] = in[78] & in2[78];
    assign P[7] = in[78] ^ in2[78];
    assign G[8] = in[77] & in2[77];
    assign P[8] = in[77] ^ in2[77];
    assign G[9] = in[76] & in2[76];
    assign P[9] = in[76] ^ in2[76];
    assign G[10] = in[75] & in2[75];
    assign P[10] = in[75] ^ in2[75];
    assign G[11] = in[74] & in2[74];
    assign P[11] = in[74] ^ in2[74];
    assign G[12] = in[73] & in2[73];
    assign P[12] = in[73] ^ in2[73];
    assign G[13] = in[72] & in2[72];
    assign P[13] = in[72] ^ in2[72];
    assign G[14] = in[71] & in2[71];
    assign P[14] = in[71] ^ in2[71];
    assign G[15] = in[70] & in2[70];
    assign P[15] = in[70] ^ in2[70];
    assign G[16] = in[69] & in2[69];
    assign P[16] = in[69] ^ in2[69];
    assign G[17] = in[68] & in2[68];
    assign P[17] = in[68] ^ in2[68];
    assign G[18] = in[67] & in2[67];
    assign P[18] = in[67] ^ in2[67];
    assign G[19] = in[66] & in2[66];
    assign P[19] = in[66] ^ in2[66];
    assign G[20] = in[65] & in2[65];
    assign P[20] = in[65] ^ in2[65];
    assign G[21] = in[64] & in2[64];
    assign P[21] = in[64] ^ in2[64];
    assign G[22] = in[63] & in2[63];
    assign P[22] = in[63] ^ in2[63];
    assign G[23] = in[62] & in2[62];
    assign P[23] = in[62] ^ in2[62];
    assign G[24] = in[61] & in2[61];
    assign P[24] = in[61] ^ in2[61];
    assign G[25] = in[60] & in2[60];
    assign P[25] = in[60] ^ in2[60];
    assign G[26] = in[59] & in2[59];
    assign P[26] = in[59] ^ in2[59];
    assign G[27] = in[58] & in2[58];
    assign P[27] = in[58] ^ in2[58];
    assign G[28] = in[57] & in2[57];
    assign P[28] = in[57] ^ in2[57];
    assign G[29] = in[56] & in2[56];
    assign P[29] = in[56] ^ in2[56];
    assign G[30] = in[55] & in2[55];
    assign P[30] = in[55] ^ in2[55];
    assign G[31] = in[54] & in2[54];
    assign P[31] = in[54] ^ in2[54];
    assign G[32] = in[53] & in2[53];
    assign P[32] = in[53] ^ in2[53];
    assign G[33] = in[52] & in2[52];
    assign P[33] = in[52] ^ in2[52];
    assign G[34] = in[51] & in2[51];
    assign P[34] = in[51] ^ in2[51];
    assign G[35] = in[50] & in2[50];
    assign P[35] = in[50] ^ in2[50];
    assign G[36] = in[49] & in2[49];
    assign P[36] = in[49] ^ in2[49];
    assign G[37] = in[48] & in2[48];
    assign P[37] = in[48] ^ in2[48];
    assign G[38] = in[47] & in2[47];
    assign P[38] = in[47] ^ in2[47];
    assign G[39] = in[46] & in2[46];
    assign P[39] = in[46] ^ in2[46];
    assign G[40] = in[45] & in2[45];
    assign P[40] = in[45] ^ in2[45];
    assign G[41] = in[44] & in2[44];
    assign P[41] = in[44] ^ in2[44];
    assign G[42] = in[43] & in2[43];
    assign P[42] = in[43] ^ in2[43];
    assign G[43] = in[42] & in2[42];
    assign P[43] = in[42] ^ in2[42];
    assign G[44] = in[41] & in2[41];
    assign P[44] = in[41] ^ in2[41];
    assign G[45] = in[40] & in2[40];
    assign P[45] = in[40] ^ in2[40];
    assign G[46] = in[39] & in2[39];
    assign P[46] = in[39] ^ in2[39];
    assign G[47] = in[38] & in2[38];
    assign P[47] = in[38] ^ in2[38];
    assign G[48] = in[37] & in2[37];
    assign P[48] = in[37] ^ in2[37];
    assign G[49] = in[36] & in2[36];
    assign P[49] = in[36] ^ in2[36];
    assign G[50] = in[35] & in2[35];
    assign P[50] = in[35] ^ in2[35];
    assign G[51] = in[34] & in2[34];
    assign P[51] = in[34] ^ in2[34];
    assign G[52] = in[33] & in2[33];
    assign P[52] = in[33] ^ in2[33];
    assign G[53] = in[32] & in2[32];
    assign P[53] = in[32] ^ in2[32];
    assign G[54] = in[31] & in2[31];
    assign P[54] = in[31] ^ in2[31];
    assign G[55] = in[30] & in2[30];
    assign P[55] = in[30] ^ in2[30];
    assign G[56] = in[29] & in2[29];
    assign P[56] = in[29] ^ in2[29];
    assign G[57] = in[28] & in2[28];
    assign P[57] = in[28] ^ in2[28];
    assign G[58] = in[27] & in2[27];
    assign P[58] = in[27] ^ in2[27];
    assign G[59] = in[26] & in2[26];
    assign P[59] = in[26] ^ in2[26];
    assign G[60] = in[25] & in2[25];
    assign P[60] = in[25] ^ in2[25];
    assign G[61] = in[24] & in2[24];
    assign P[61] = in[24] ^ in2[24];
    assign G[62] = in[23] & in2[23];
    assign P[62] = in[23] ^ in2[23];
    assign G[63] = in[22] & in2[22];
    assign P[63] = in[22] ^ in2[22];
    assign G[64] = in[21] & in2[21];
    assign P[64] = in[21] ^ in2[21];
    assign G[65] = in[20] & in2[20];
    assign P[65] = in[20] ^ in2[20];
    assign G[66] = in[19] & in2[19];
    assign P[66] = in[19] ^ in2[19];
    assign G[67] = in[18] & in2[18];
    assign P[67] = in[18] ^ in2[18];
    assign G[68] = in[17] & in2[17];
    assign P[68] = in[17] ^ in2[17];
    assign G[69] = in[16] & in2[16];
    assign P[69] = in[16] ^ in2[16];
    assign G[70] = in[15] & in2[15];
    assign P[70] = in[15] ^ in2[15];
    assign G[71] = in[14] & in2[14];
    assign P[71] = in[14] ^ in2[14];
    assign G[72] = in[13] & in2[13];
    assign P[72] = in[13] ^ in2[13];
    assign G[73] = in[12] & in2[12];
    assign P[73] = in[12] ^ in2[12];
    assign G[74] = in[11] & in2[11];
    assign P[74] = in[11] ^ in2[11];
    assign G[75] = in[10] & in2[10];
    assign P[75] = in[10] ^ in2[10];
    assign G[76] = in[9] & in2[9];
    assign P[76] = in[9] ^ in2[9];
    assign G[77] = in[8] & in2[8];
    assign P[77] = in[8] ^ in2[8];
    assign G[78] = in[7] & in2[7];
    assign P[78] = in[7] ^ in2[7];
    assign G[79] = in[6] & in2[6];
    assign P[79] = in[6] ^ in2[6];
    assign G[80] = in[5] & in2[5];
    assign P[80] = in[5] ^ in2[5];
    assign G[81] = in[4] & in2[4];
    assign P[81] = in[4] ^ in2[4];
    assign G[82] = in[3] & in2[3];
    assign P[82] = in[3] ^ in2[3];
    assign G[83] = in[2] & in2[2];
    assign P[83] = in[2] ^ in2[2];
    assign G[84] = in[1] & in2[1];
    assign P[84] = in[1] ^ in2[1];
    assign G[85] = in[0] & in2[0];
    assign P[85] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign C[85] = G[84] | (P[84] & C[84]);
    assign cout = G[85] | (P[85] & C[85]);
    assign sum = P ^ C;
endmodule

module CLA85(output [84:0] sum, output cout, input [84:0] in1, input [84:0] in2;

    wire[84:0] G;
    wire[84:0] C;
    wire[84:0] P;

    assign G[0] = in[84] & in2[84];
    assign P[0] = in[84] ^ in2[84];
    assign G[1] = in[83] & in2[83];
    assign P[1] = in[83] ^ in2[83];
    assign G[2] = in[82] & in2[82];
    assign P[2] = in[82] ^ in2[82];
    assign G[3] = in[81] & in2[81];
    assign P[3] = in[81] ^ in2[81];
    assign G[4] = in[80] & in2[80];
    assign P[4] = in[80] ^ in2[80];
    assign G[5] = in[79] & in2[79];
    assign P[5] = in[79] ^ in2[79];
    assign G[6] = in[78] & in2[78];
    assign P[6] = in[78] ^ in2[78];
    assign G[7] = in[77] & in2[77];
    assign P[7] = in[77] ^ in2[77];
    assign G[8] = in[76] & in2[76];
    assign P[8] = in[76] ^ in2[76];
    assign G[9] = in[75] & in2[75];
    assign P[9] = in[75] ^ in2[75];
    assign G[10] = in[74] & in2[74];
    assign P[10] = in[74] ^ in2[74];
    assign G[11] = in[73] & in2[73];
    assign P[11] = in[73] ^ in2[73];
    assign G[12] = in[72] & in2[72];
    assign P[12] = in[72] ^ in2[72];
    assign G[13] = in[71] & in2[71];
    assign P[13] = in[71] ^ in2[71];
    assign G[14] = in[70] & in2[70];
    assign P[14] = in[70] ^ in2[70];
    assign G[15] = in[69] & in2[69];
    assign P[15] = in[69] ^ in2[69];
    assign G[16] = in[68] & in2[68];
    assign P[16] = in[68] ^ in2[68];
    assign G[17] = in[67] & in2[67];
    assign P[17] = in[67] ^ in2[67];
    assign G[18] = in[66] & in2[66];
    assign P[18] = in[66] ^ in2[66];
    assign G[19] = in[65] & in2[65];
    assign P[19] = in[65] ^ in2[65];
    assign G[20] = in[64] & in2[64];
    assign P[20] = in[64] ^ in2[64];
    assign G[21] = in[63] & in2[63];
    assign P[21] = in[63] ^ in2[63];
    assign G[22] = in[62] & in2[62];
    assign P[22] = in[62] ^ in2[62];
    assign G[23] = in[61] & in2[61];
    assign P[23] = in[61] ^ in2[61];
    assign G[24] = in[60] & in2[60];
    assign P[24] = in[60] ^ in2[60];
    assign G[25] = in[59] & in2[59];
    assign P[25] = in[59] ^ in2[59];
    assign G[26] = in[58] & in2[58];
    assign P[26] = in[58] ^ in2[58];
    assign G[27] = in[57] & in2[57];
    assign P[27] = in[57] ^ in2[57];
    assign G[28] = in[56] & in2[56];
    assign P[28] = in[56] ^ in2[56];
    assign G[29] = in[55] & in2[55];
    assign P[29] = in[55] ^ in2[55];
    assign G[30] = in[54] & in2[54];
    assign P[30] = in[54] ^ in2[54];
    assign G[31] = in[53] & in2[53];
    assign P[31] = in[53] ^ in2[53];
    assign G[32] = in[52] & in2[52];
    assign P[32] = in[52] ^ in2[52];
    assign G[33] = in[51] & in2[51];
    assign P[33] = in[51] ^ in2[51];
    assign G[34] = in[50] & in2[50];
    assign P[34] = in[50] ^ in2[50];
    assign G[35] = in[49] & in2[49];
    assign P[35] = in[49] ^ in2[49];
    assign G[36] = in[48] & in2[48];
    assign P[36] = in[48] ^ in2[48];
    assign G[37] = in[47] & in2[47];
    assign P[37] = in[47] ^ in2[47];
    assign G[38] = in[46] & in2[46];
    assign P[38] = in[46] ^ in2[46];
    assign G[39] = in[45] & in2[45];
    assign P[39] = in[45] ^ in2[45];
    assign G[40] = in[44] & in2[44];
    assign P[40] = in[44] ^ in2[44];
    assign G[41] = in[43] & in2[43];
    assign P[41] = in[43] ^ in2[43];
    assign G[42] = in[42] & in2[42];
    assign P[42] = in[42] ^ in2[42];
    assign G[43] = in[41] & in2[41];
    assign P[43] = in[41] ^ in2[41];
    assign G[44] = in[40] & in2[40];
    assign P[44] = in[40] ^ in2[40];
    assign G[45] = in[39] & in2[39];
    assign P[45] = in[39] ^ in2[39];
    assign G[46] = in[38] & in2[38];
    assign P[46] = in[38] ^ in2[38];
    assign G[47] = in[37] & in2[37];
    assign P[47] = in[37] ^ in2[37];
    assign G[48] = in[36] & in2[36];
    assign P[48] = in[36] ^ in2[36];
    assign G[49] = in[35] & in2[35];
    assign P[49] = in[35] ^ in2[35];
    assign G[50] = in[34] & in2[34];
    assign P[50] = in[34] ^ in2[34];
    assign G[51] = in[33] & in2[33];
    assign P[51] = in[33] ^ in2[33];
    assign G[52] = in[32] & in2[32];
    assign P[52] = in[32] ^ in2[32];
    assign G[53] = in[31] & in2[31];
    assign P[53] = in[31] ^ in2[31];
    assign G[54] = in[30] & in2[30];
    assign P[54] = in[30] ^ in2[30];
    assign G[55] = in[29] & in2[29];
    assign P[55] = in[29] ^ in2[29];
    assign G[56] = in[28] & in2[28];
    assign P[56] = in[28] ^ in2[28];
    assign G[57] = in[27] & in2[27];
    assign P[57] = in[27] ^ in2[27];
    assign G[58] = in[26] & in2[26];
    assign P[58] = in[26] ^ in2[26];
    assign G[59] = in[25] & in2[25];
    assign P[59] = in[25] ^ in2[25];
    assign G[60] = in[24] & in2[24];
    assign P[60] = in[24] ^ in2[24];
    assign G[61] = in[23] & in2[23];
    assign P[61] = in[23] ^ in2[23];
    assign G[62] = in[22] & in2[22];
    assign P[62] = in[22] ^ in2[22];
    assign G[63] = in[21] & in2[21];
    assign P[63] = in[21] ^ in2[21];
    assign G[64] = in[20] & in2[20];
    assign P[64] = in[20] ^ in2[20];
    assign G[65] = in[19] & in2[19];
    assign P[65] = in[19] ^ in2[19];
    assign G[66] = in[18] & in2[18];
    assign P[66] = in[18] ^ in2[18];
    assign G[67] = in[17] & in2[17];
    assign P[67] = in[17] ^ in2[17];
    assign G[68] = in[16] & in2[16];
    assign P[68] = in[16] ^ in2[16];
    assign G[69] = in[15] & in2[15];
    assign P[69] = in[15] ^ in2[15];
    assign G[70] = in[14] & in2[14];
    assign P[70] = in[14] ^ in2[14];
    assign G[71] = in[13] & in2[13];
    assign P[71] = in[13] ^ in2[13];
    assign G[72] = in[12] & in2[12];
    assign P[72] = in[12] ^ in2[12];
    assign G[73] = in[11] & in2[11];
    assign P[73] = in[11] ^ in2[11];
    assign G[74] = in[10] & in2[10];
    assign P[74] = in[10] ^ in2[10];
    assign G[75] = in[9] & in2[9];
    assign P[75] = in[9] ^ in2[9];
    assign G[76] = in[8] & in2[8];
    assign P[76] = in[8] ^ in2[8];
    assign G[77] = in[7] & in2[7];
    assign P[77] = in[7] ^ in2[7];
    assign G[78] = in[6] & in2[6];
    assign P[78] = in[6] ^ in2[6];
    assign G[79] = in[5] & in2[5];
    assign P[79] = in[5] ^ in2[5];
    assign G[80] = in[4] & in2[4];
    assign P[80] = in[4] ^ in2[4];
    assign G[81] = in[3] & in2[3];
    assign P[81] = in[3] ^ in2[3];
    assign G[82] = in[2] & in2[2];
    assign P[82] = in[2] ^ in2[2];
    assign G[83] = in[1] & in2[1];
    assign P[83] = in[1] ^ in2[1];
    assign G[84] = in[0] & in2[0];
    assign P[84] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign C[84] = G[83] | (P[83] & C[83]);
    assign cout = G[84] | (P[84] & C[84]);
    assign sum = P ^ C;
endmodule

module CLA84(output [83:0] sum, output cout, input [83:0] in1, input [83:0] in2;

    wire[83:0] G;
    wire[83:0] C;
    wire[83:0] P;

    assign G[0] = in[83] & in2[83];
    assign P[0] = in[83] ^ in2[83];
    assign G[1] = in[82] & in2[82];
    assign P[1] = in[82] ^ in2[82];
    assign G[2] = in[81] & in2[81];
    assign P[2] = in[81] ^ in2[81];
    assign G[3] = in[80] & in2[80];
    assign P[3] = in[80] ^ in2[80];
    assign G[4] = in[79] & in2[79];
    assign P[4] = in[79] ^ in2[79];
    assign G[5] = in[78] & in2[78];
    assign P[5] = in[78] ^ in2[78];
    assign G[6] = in[77] & in2[77];
    assign P[6] = in[77] ^ in2[77];
    assign G[7] = in[76] & in2[76];
    assign P[7] = in[76] ^ in2[76];
    assign G[8] = in[75] & in2[75];
    assign P[8] = in[75] ^ in2[75];
    assign G[9] = in[74] & in2[74];
    assign P[9] = in[74] ^ in2[74];
    assign G[10] = in[73] & in2[73];
    assign P[10] = in[73] ^ in2[73];
    assign G[11] = in[72] & in2[72];
    assign P[11] = in[72] ^ in2[72];
    assign G[12] = in[71] & in2[71];
    assign P[12] = in[71] ^ in2[71];
    assign G[13] = in[70] & in2[70];
    assign P[13] = in[70] ^ in2[70];
    assign G[14] = in[69] & in2[69];
    assign P[14] = in[69] ^ in2[69];
    assign G[15] = in[68] & in2[68];
    assign P[15] = in[68] ^ in2[68];
    assign G[16] = in[67] & in2[67];
    assign P[16] = in[67] ^ in2[67];
    assign G[17] = in[66] & in2[66];
    assign P[17] = in[66] ^ in2[66];
    assign G[18] = in[65] & in2[65];
    assign P[18] = in[65] ^ in2[65];
    assign G[19] = in[64] & in2[64];
    assign P[19] = in[64] ^ in2[64];
    assign G[20] = in[63] & in2[63];
    assign P[20] = in[63] ^ in2[63];
    assign G[21] = in[62] & in2[62];
    assign P[21] = in[62] ^ in2[62];
    assign G[22] = in[61] & in2[61];
    assign P[22] = in[61] ^ in2[61];
    assign G[23] = in[60] & in2[60];
    assign P[23] = in[60] ^ in2[60];
    assign G[24] = in[59] & in2[59];
    assign P[24] = in[59] ^ in2[59];
    assign G[25] = in[58] & in2[58];
    assign P[25] = in[58] ^ in2[58];
    assign G[26] = in[57] & in2[57];
    assign P[26] = in[57] ^ in2[57];
    assign G[27] = in[56] & in2[56];
    assign P[27] = in[56] ^ in2[56];
    assign G[28] = in[55] & in2[55];
    assign P[28] = in[55] ^ in2[55];
    assign G[29] = in[54] & in2[54];
    assign P[29] = in[54] ^ in2[54];
    assign G[30] = in[53] & in2[53];
    assign P[30] = in[53] ^ in2[53];
    assign G[31] = in[52] & in2[52];
    assign P[31] = in[52] ^ in2[52];
    assign G[32] = in[51] & in2[51];
    assign P[32] = in[51] ^ in2[51];
    assign G[33] = in[50] & in2[50];
    assign P[33] = in[50] ^ in2[50];
    assign G[34] = in[49] & in2[49];
    assign P[34] = in[49] ^ in2[49];
    assign G[35] = in[48] & in2[48];
    assign P[35] = in[48] ^ in2[48];
    assign G[36] = in[47] & in2[47];
    assign P[36] = in[47] ^ in2[47];
    assign G[37] = in[46] & in2[46];
    assign P[37] = in[46] ^ in2[46];
    assign G[38] = in[45] & in2[45];
    assign P[38] = in[45] ^ in2[45];
    assign G[39] = in[44] & in2[44];
    assign P[39] = in[44] ^ in2[44];
    assign G[40] = in[43] & in2[43];
    assign P[40] = in[43] ^ in2[43];
    assign G[41] = in[42] & in2[42];
    assign P[41] = in[42] ^ in2[42];
    assign G[42] = in[41] & in2[41];
    assign P[42] = in[41] ^ in2[41];
    assign G[43] = in[40] & in2[40];
    assign P[43] = in[40] ^ in2[40];
    assign G[44] = in[39] & in2[39];
    assign P[44] = in[39] ^ in2[39];
    assign G[45] = in[38] & in2[38];
    assign P[45] = in[38] ^ in2[38];
    assign G[46] = in[37] & in2[37];
    assign P[46] = in[37] ^ in2[37];
    assign G[47] = in[36] & in2[36];
    assign P[47] = in[36] ^ in2[36];
    assign G[48] = in[35] & in2[35];
    assign P[48] = in[35] ^ in2[35];
    assign G[49] = in[34] & in2[34];
    assign P[49] = in[34] ^ in2[34];
    assign G[50] = in[33] & in2[33];
    assign P[50] = in[33] ^ in2[33];
    assign G[51] = in[32] & in2[32];
    assign P[51] = in[32] ^ in2[32];
    assign G[52] = in[31] & in2[31];
    assign P[52] = in[31] ^ in2[31];
    assign G[53] = in[30] & in2[30];
    assign P[53] = in[30] ^ in2[30];
    assign G[54] = in[29] & in2[29];
    assign P[54] = in[29] ^ in2[29];
    assign G[55] = in[28] & in2[28];
    assign P[55] = in[28] ^ in2[28];
    assign G[56] = in[27] & in2[27];
    assign P[56] = in[27] ^ in2[27];
    assign G[57] = in[26] & in2[26];
    assign P[57] = in[26] ^ in2[26];
    assign G[58] = in[25] & in2[25];
    assign P[58] = in[25] ^ in2[25];
    assign G[59] = in[24] & in2[24];
    assign P[59] = in[24] ^ in2[24];
    assign G[60] = in[23] & in2[23];
    assign P[60] = in[23] ^ in2[23];
    assign G[61] = in[22] & in2[22];
    assign P[61] = in[22] ^ in2[22];
    assign G[62] = in[21] & in2[21];
    assign P[62] = in[21] ^ in2[21];
    assign G[63] = in[20] & in2[20];
    assign P[63] = in[20] ^ in2[20];
    assign G[64] = in[19] & in2[19];
    assign P[64] = in[19] ^ in2[19];
    assign G[65] = in[18] & in2[18];
    assign P[65] = in[18] ^ in2[18];
    assign G[66] = in[17] & in2[17];
    assign P[66] = in[17] ^ in2[17];
    assign G[67] = in[16] & in2[16];
    assign P[67] = in[16] ^ in2[16];
    assign G[68] = in[15] & in2[15];
    assign P[68] = in[15] ^ in2[15];
    assign G[69] = in[14] & in2[14];
    assign P[69] = in[14] ^ in2[14];
    assign G[70] = in[13] & in2[13];
    assign P[70] = in[13] ^ in2[13];
    assign G[71] = in[12] & in2[12];
    assign P[71] = in[12] ^ in2[12];
    assign G[72] = in[11] & in2[11];
    assign P[72] = in[11] ^ in2[11];
    assign G[73] = in[10] & in2[10];
    assign P[73] = in[10] ^ in2[10];
    assign G[74] = in[9] & in2[9];
    assign P[74] = in[9] ^ in2[9];
    assign G[75] = in[8] & in2[8];
    assign P[75] = in[8] ^ in2[8];
    assign G[76] = in[7] & in2[7];
    assign P[76] = in[7] ^ in2[7];
    assign G[77] = in[6] & in2[6];
    assign P[77] = in[6] ^ in2[6];
    assign G[78] = in[5] & in2[5];
    assign P[78] = in[5] ^ in2[5];
    assign G[79] = in[4] & in2[4];
    assign P[79] = in[4] ^ in2[4];
    assign G[80] = in[3] & in2[3];
    assign P[80] = in[3] ^ in2[3];
    assign G[81] = in[2] & in2[2];
    assign P[81] = in[2] ^ in2[2];
    assign G[82] = in[1] & in2[1];
    assign P[82] = in[1] ^ in2[1];
    assign G[83] = in[0] & in2[0];
    assign P[83] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign C[83] = G[82] | (P[82] & C[82]);
    assign cout = G[83] | (P[83] & C[83]);
    assign sum = P ^ C;
endmodule

module CLA83(output [82:0] sum, output cout, input [82:0] in1, input [82:0] in2;

    wire[82:0] G;
    wire[82:0] C;
    wire[82:0] P;

    assign G[0] = in[82] & in2[82];
    assign P[0] = in[82] ^ in2[82];
    assign G[1] = in[81] & in2[81];
    assign P[1] = in[81] ^ in2[81];
    assign G[2] = in[80] & in2[80];
    assign P[2] = in[80] ^ in2[80];
    assign G[3] = in[79] & in2[79];
    assign P[3] = in[79] ^ in2[79];
    assign G[4] = in[78] & in2[78];
    assign P[4] = in[78] ^ in2[78];
    assign G[5] = in[77] & in2[77];
    assign P[5] = in[77] ^ in2[77];
    assign G[6] = in[76] & in2[76];
    assign P[6] = in[76] ^ in2[76];
    assign G[7] = in[75] & in2[75];
    assign P[7] = in[75] ^ in2[75];
    assign G[8] = in[74] & in2[74];
    assign P[8] = in[74] ^ in2[74];
    assign G[9] = in[73] & in2[73];
    assign P[9] = in[73] ^ in2[73];
    assign G[10] = in[72] & in2[72];
    assign P[10] = in[72] ^ in2[72];
    assign G[11] = in[71] & in2[71];
    assign P[11] = in[71] ^ in2[71];
    assign G[12] = in[70] & in2[70];
    assign P[12] = in[70] ^ in2[70];
    assign G[13] = in[69] & in2[69];
    assign P[13] = in[69] ^ in2[69];
    assign G[14] = in[68] & in2[68];
    assign P[14] = in[68] ^ in2[68];
    assign G[15] = in[67] & in2[67];
    assign P[15] = in[67] ^ in2[67];
    assign G[16] = in[66] & in2[66];
    assign P[16] = in[66] ^ in2[66];
    assign G[17] = in[65] & in2[65];
    assign P[17] = in[65] ^ in2[65];
    assign G[18] = in[64] & in2[64];
    assign P[18] = in[64] ^ in2[64];
    assign G[19] = in[63] & in2[63];
    assign P[19] = in[63] ^ in2[63];
    assign G[20] = in[62] & in2[62];
    assign P[20] = in[62] ^ in2[62];
    assign G[21] = in[61] & in2[61];
    assign P[21] = in[61] ^ in2[61];
    assign G[22] = in[60] & in2[60];
    assign P[22] = in[60] ^ in2[60];
    assign G[23] = in[59] & in2[59];
    assign P[23] = in[59] ^ in2[59];
    assign G[24] = in[58] & in2[58];
    assign P[24] = in[58] ^ in2[58];
    assign G[25] = in[57] & in2[57];
    assign P[25] = in[57] ^ in2[57];
    assign G[26] = in[56] & in2[56];
    assign P[26] = in[56] ^ in2[56];
    assign G[27] = in[55] & in2[55];
    assign P[27] = in[55] ^ in2[55];
    assign G[28] = in[54] & in2[54];
    assign P[28] = in[54] ^ in2[54];
    assign G[29] = in[53] & in2[53];
    assign P[29] = in[53] ^ in2[53];
    assign G[30] = in[52] & in2[52];
    assign P[30] = in[52] ^ in2[52];
    assign G[31] = in[51] & in2[51];
    assign P[31] = in[51] ^ in2[51];
    assign G[32] = in[50] & in2[50];
    assign P[32] = in[50] ^ in2[50];
    assign G[33] = in[49] & in2[49];
    assign P[33] = in[49] ^ in2[49];
    assign G[34] = in[48] & in2[48];
    assign P[34] = in[48] ^ in2[48];
    assign G[35] = in[47] & in2[47];
    assign P[35] = in[47] ^ in2[47];
    assign G[36] = in[46] & in2[46];
    assign P[36] = in[46] ^ in2[46];
    assign G[37] = in[45] & in2[45];
    assign P[37] = in[45] ^ in2[45];
    assign G[38] = in[44] & in2[44];
    assign P[38] = in[44] ^ in2[44];
    assign G[39] = in[43] & in2[43];
    assign P[39] = in[43] ^ in2[43];
    assign G[40] = in[42] & in2[42];
    assign P[40] = in[42] ^ in2[42];
    assign G[41] = in[41] & in2[41];
    assign P[41] = in[41] ^ in2[41];
    assign G[42] = in[40] & in2[40];
    assign P[42] = in[40] ^ in2[40];
    assign G[43] = in[39] & in2[39];
    assign P[43] = in[39] ^ in2[39];
    assign G[44] = in[38] & in2[38];
    assign P[44] = in[38] ^ in2[38];
    assign G[45] = in[37] & in2[37];
    assign P[45] = in[37] ^ in2[37];
    assign G[46] = in[36] & in2[36];
    assign P[46] = in[36] ^ in2[36];
    assign G[47] = in[35] & in2[35];
    assign P[47] = in[35] ^ in2[35];
    assign G[48] = in[34] & in2[34];
    assign P[48] = in[34] ^ in2[34];
    assign G[49] = in[33] & in2[33];
    assign P[49] = in[33] ^ in2[33];
    assign G[50] = in[32] & in2[32];
    assign P[50] = in[32] ^ in2[32];
    assign G[51] = in[31] & in2[31];
    assign P[51] = in[31] ^ in2[31];
    assign G[52] = in[30] & in2[30];
    assign P[52] = in[30] ^ in2[30];
    assign G[53] = in[29] & in2[29];
    assign P[53] = in[29] ^ in2[29];
    assign G[54] = in[28] & in2[28];
    assign P[54] = in[28] ^ in2[28];
    assign G[55] = in[27] & in2[27];
    assign P[55] = in[27] ^ in2[27];
    assign G[56] = in[26] & in2[26];
    assign P[56] = in[26] ^ in2[26];
    assign G[57] = in[25] & in2[25];
    assign P[57] = in[25] ^ in2[25];
    assign G[58] = in[24] & in2[24];
    assign P[58] = in[24] ^ in2[24];
    assign G[59] = in[23] & in2[23];
    assign P[59] = in[23] ^ in2[23];
    assign G[60] = in[22] & in2[22];
    assign P[60] = in[22] ^ in2[22];
    assign G[61] = in[21] & in2[21];
    assign P[61] = in[21] ^ in2[21];
    assign G[62] = in[20] & in2[20];
    assign P[62] = in[20] ^ in2[20];
    assign G[63] = in[19] & in2[19];
    assign P[63] = in[19] ^ in2[19];
    assign G[64] = in[18] & in2[18];
    assign P[64] = in[18] ^ in2[18];
    assign G[65] = in[17] & in2[17];
    assign P[65] = in[17] ^ in2[17];
    assign G[66] = in[16] & in2[16];
    assign P[66] = in[16] ^ in2[16];
    assign G[67] = in[15] & in2[15];
    assign P[67] = in[15] ^ in2[15];
    assign G[68] = in[14] & in2[14];
    assign P[68] = in[14] ^ in2[14];
    assign G[69] = in[13] & in2[13];
    assign P[69] = in[13] ^ in2[13];
    assign G[70] = in[12] & in2[12];
    assign P[70] = in[12] ^ in2[12];
    assign G[71] = in[11] & in2[11];
    assign P[71] = in[11] ^ in2[11];
    assign G[72] = in[10] & in2[10];
    assign P[72] = in[10] ^ in2[10];
    assign G[73] = in[9] & in2[9];
    assign P[73] = in[9] ^ in2[9];
    assign G[74] = in[8] & in2[8];
    assign P[74] = in[8] ^ in2[8];
    assign G[75] = in[7] & in2[7];
    assign P[75] = in[7] ^ in2[7];
    assign G[76] = in[6] & in2[6];
    assign P[76] = in[6] ^ in2[6];
    assign G[77] = in[5] & in2[5];
    assign P[77] = in[5] ^ in2[5];
    assign G[78] = in[4] & in2[4];
    assign P[78] = in[4] ^ in2[4];
    assign G[79] = in[3] & in2[3];
    assign P[79] = in[3] ^ in2[3];
    assign G[80] = in[2] & in2[2];
    assign P[80] = in[2] ^ in2[2];
    assign G[81] = in[1] & in2[1];
    assign P[81] = in[1] ^ in2[1];
    assign G[82] = in[0] & in2[0];
    assign P[82] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign C[82] = G[81] | (P[81] & C[81]);
    assign cout = G[82] | (P[82] & C[82]);
    assign sum = P ^ C;
endmodule

module CLA82(output [81:0] sum, output cout, input [81:0] in1, input [81:0] in2;

    wire[81:0] G;
    wire[81:0] C;
    wire[81:0] P;

    assign G[0] = in[81] & in2[81];
    assign P[0] = in[81] ^ in2[81];
    assign G[1] = in[80] & in2[80];
    assign P[1] = in[80] ^ in2[80];
    assign G[2] = in[79] & in2[79];
    assign P[2] = in[79] ^ in2[79];
    assign G[3] = in[78] & in2[78];
    assign P[3] = in[78] ^ in2[78];
    assign G[4] = in[77] & in2[77];
    assign P[4] = in[77] ^ in2[77];
    assign G[5] = in[76] & in2[76];
    assign P[5] = in[76] ^ in2[76];
    assign G[6] = in[75] & in2[75];
    assign P[6] = in[75] ^ in2[75];
    assign G[7] = in[74] & in2[74];
    assign P[7] = in[74] ^ in2[74];
    assign G[8] = in[73] & in2[73];
    assign P[8] = in[73] ^ in2[73];
    assign G[9] = in[72] & in2[72];
    assign P[9] = in[72] ^ in2[72];
    assign G[10] = in[71] & in2[71];
    assign P[10] = in[71] ^ in2[71];
    assign G[11] = in[70] & in2[70];
    assign P[11] = in[70] ^ in2[70];
    assign G[12] = in[69] & in2[69];
    assign P[12] = in[69] ^ in2[69];
    assign G[13] = in[68] & in2[68];
    assign P[13] = in[68] ^ in2[68];
    assign G[14] = in[67] & in2[67];
    assign P[14] = in[67] ^ in2[67];
    assign G[15] = in[66] & in2[66];
    assign P[15] = in[66] ^ in2[66];
    assign G[16] = in[65] & in2[65];
    assign P[16] = in[65] ^ in2[65];
    assign G[17] = in[64] & in2[64];
    assign P[17] = in[64] ^ in2[64];
    assign G[18] = in[63] & in2[63];
    assign P[18] = in[63] ^ in2[63];
    assign G[19] = in[62] & in2[62];
    assign P[19] = in[62] ^ in2[62];
    assign G[20] = in[61] & in2[61];
    assign P[20] = in[61] ^ in2[61];
    assign G[21] = in[60] & in2[60];
    assign P[21] = in[60] ^ in2[60];
    assign G[22] = in[59] & in2[59];
    assign P[22] = in[59] ^ in2[59];
    assign G[23] = in[58] & in2[58];
    assign P[23] = in[58] ^ in2[58];
    assign G[24] = in[57] & in2[57];
    assign P[24] = in[57] ^ in2[57];
    assign G[25] = in[56] & in2[56];
    assign P[25] = in[56] ^ in2[56];
    assign G[26] = in[55] & in2[55];
    assign P[26] = in[55] ^ in2[55];
    assign G[27] = in[54] & in2[54];
    assign P[27] = in[54] ^ in2[54];
    assign G[28] = in[53] & in2[53];
    assign P[28] = in[53] ^ in2[53];
    assign G[29] = in[52] & in2[52];
    assign P[29] = in[52] ^ in2[52];
    assign G[30] = in[51] & in2[51];
    assign P[30] = in[51] ^ in2[51];
    assign G[31] = in[50] & in2[50];
    assign P[31] = in[50] ^ in2[50];
    assign G[32] = in[49] & in2[49];
    assign P[32] = in[49] ^ in2[49];
    assign G[33] = in[48] & in2[48];
    assign P[33] = in[48] ^ in2[48];
    assign G[34] = in[47] & in2[47];
    assign P[34] = in[47] ^ in2[47];
    assign G[35] = in[46] & in2[46];
    assign P[35] = in[46] ^ in2[46];
    assign G[36] = in[45] & in2[45];
    assign P[36] = in[45] ^ in2[45];
    assign G[37] = in[44] & in2[44];
    assign P[37] = in[44] ^ in2[44];
    assign G[38] = in[43] & in2[43];
    assign P[38] = in[43] ^ in2[43];
    assign G[39] = in[42] & in2[42];
    assign P[39] = in[42] ^ in2[42];
    assign G[40] = in[41] & in2[41];
    assign P[40] = in[41] ^ in2[41];
    assign G[41] = in[40] & in2[40];
    assign P[41] = in[40] ^ in2[40];
    assign G[42] = in[39] & in2[39];
    assign P[42] = in[39] ^ in2[39];
    assign G[43] = in[38] & in2[38];
    assign P[43] = in[38] ^ in2[38];
    assign G[44] = in[37] & in2[37];
    assign P[44] = in[37] ^ in2[37];
    assign G[45] = in[36] & in2[36];
    assign P[45] = in[36] ^ in2[36];
    assign G[46] = in[35] & in2[35];
    assign P[46] = in[35] ^ in2[35];
    assign G[47] = in[34] & in2[34];
    assign P[47] = in[34] ^ in2[34];
    assign G[48] = in[33] & in2[33];
    assign P[48] = in[33] ^ in2[33];
    assign G[49] = in[32] & in2[32];
    assign P[49] = in[32] ^ in2[32];
    assign G[50] = in[31] & in2[31];
    assign P[50] = in[31] ^ in2[31];
    assign G[51] = in[30] & in2[30];
    assign P[51] = in[30] ^ in2[30];
    assign G[52] = in[29] & in2[29];
    assign P[52] = in[29] ^ in2[29];
    assign G[53] = in[28] & in2[28];
    assign P[53] = in[28] ^ in2[28];
    assign G[54] = in[27] & in2[27];
    assign P[54] = in[27] ^ in2[27];
    assign G[55] = in[26] & in2[26];
    assign P[55] = in[26] ^ in2[26];
    assign G[56] = in[25] & in2[25];
    assign P[56] = in[25] ^ in2[25];
    assign G[57] = in[24] & in2[24];
    assign P[57] = in[24] ^ in2[24];
    assign G[58] = in[23] & in2[23];
    assign P[58] = in[23] ^ in2[23];
    assign G[59] = in[22] & in2[22];
    assign P[59] = in[22] ^ in2[22];
    assign G[60] = in[21] & in2[21];
    assign P[60] = in[21] ^ in2[21];
    assign G[61] = in[20] & in2[20];
    assign P[61] = in[20] ^ in2[20];
    assign G[62] = in[19] & in2[19];
    assign P[62] = in[19] ^ in2[19];
    assign G[63] = in[18] & in2[18];
    assign P[63] = in[18] ^ in2[18];
    assign G[64] = in[17] & in2[17];
    assign P[64] = in[17] ^ in2[17];
    assign G[65] = in[16] & in2[16];
    assign P[65] = in[16] ^ in2[16];
    assign G[66] = in[15] & in2[15];
    assign P[66] = in[15] ^ in2[15];
    assign G[67] = in[14] & in2[14];
    assign P[67] = in[14] ^ in2[14];
    assign G[68] = in[13] & in2[13];
    assign P[68] = in[13] ^ in2[13];
    assign G[69] = in[12] & in2[12];
    assign P[69] = in[12] ^ in2[12];
    assign G[70] = in[11] & in2[11];
    assign P[70] = in[11] ^ in2[11];
    assign G[71] = in[10] & in2[10];
    assign P[71] = in[10] ^ in2[10];
    assign G[72] = in[9] & in2[9];
    assign P[72] = in[9] ^ in2[9];
    assign G[73] = in[8] & in2[8];
    assign P[73] = in[8] ^ in2[8];
    assign G[74] = in[7] & in2[7];
    assign P[74] = in[7] ^ in2[7];
    assign G[75] = in[6] & in2[6];
    assign P[75] = in[6] ^ in2[6];
    assign G[76] = in[5] & in2[5];
    assign P[76] = in[5] ^ in2[5];
    assign G[77] = in[4] & in2[4];
    assign P[77] = in[4] ^ in2[4];
    assign G[78] = in[3] & in2[3];
    assign P[78] = in[3] ^ in2[3];
    assign G[79] = in[2] & in2[2];
    assign P[79] = in[2] ^ in2[2];
    assign G[80] = in[1] & in2[1];
    assign P[80] = in[1] ^ in2[1];
    assign G[81] = in[0] & in2[0];
    assign P[81] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign C[81] = G[80] | (P[80] & C[80]);
    assign cout = G[81] | (P[81] & C[81]);
    assign sum = P ^ C;
endmodule

module CLA81(output [80:0] sum, output cout, input [80:0] in1, input [80:0] in2;

    wire[80:0] G;
    wire[80:0] C;
    wire[80:0] P;

    assign G[0] = in[80] & in2[80];
    assign P[0] = in[80] ^ in2[80];
    assign G[1] = in[79] & in2[79];
    assign P[1] = in[79] ^ in2[79];
    assign G[2] = in[78] & in2[78];
    assign P[2] = in[78] ^ in2[78];
    assign G[3] = in[77] & in2[77];
    assign P[3] = in[77] ^ in2[77];
    assign G[4] = in[76] & in2[76];
    assign P[4] = in[76] ^ in2[76];
    assign G[5] = in[75] & in2[75];
    assign P[5] = in[75] ^ in2[75];
    assign G[6] = in[74] & in2[74];
    assign P[6] = in[74] ^ in2[74];
    assign G[7] = in[73] & in2[73];
    assign P[7] = in[73] ^ in2[73];
    assign G[8] = in[72] & in2[72];
    assign P[8] = in[72] ^ in2[72];
    assign G[9] = in[71] & in2[71];
    assign P[9] = in[71] ^ in2[71];
    assign G[10] = in[70] & in2[70];
    assign P[10] = in[70] ^ in2[70];
    assign G[11] = in[69] & in2[69];
    assign P[11] = in[69] ^ in2[69];
    assign G[12] = in[68] & in2[68];
    assign P[12] = in[68] ^ in2[68];
    assign G[13] = in[67] & in2[67];
    assign P[13] = in[67] ^ in2[67];
    assign G[14] = in[66] & in2[66];
    assign P[14] = in[66] ^ in2[66];
    assign G[15] = in[65] & in2[65];
    assign P[15] = in[65] ^ in2[65];
    assign G[16] = in[64] & in2[64];
    assign P[16] = in[64] ^ in2[64];
    assign G[17] = in[63] & in2[63];
    assign P[17] = in[63] ^ in2[63];
    assign G[18] = in[62] & in2[62];
    assign P[18] = in[62] ^ in2[62];
    assign G[19] = in[61] & in2[61];
    assign P[19] = in[61] ^ in2[61];
    assign G[20] = in[60] & in2[60];
    assign P[20] = in[60] ^ in2[60];
    assign G[21] = in[59] & in2[59];
    assign P[21] = in[59] ^ in2[59];
    assign G[22] = in[58] & in2[58];
    assign P[22] = in[58] ^ in2[58];
    assign G[23] = in[57] & in2[57];
    assign P[23] = in[57] ^ in2[57];
    assign G[24] = in[56] & in2[56];
    assign P[24] = in[56] ^ in2[56];
    assign G[25] = in[55] & in2[55];
    assign P[25] = in[55] ^ in2[55];
    assign G[26] = in[54] & in2[54];
    assign P[26] = in[54] ^ in2[54];
    assign G[27] = in[53] & in2[53];
    assign P[27] = in[53] ^ in2[53];
    assign G[28] = in[52] & in2[52];
    assign P[28] = in[52] ^ in2[52];
    assign G[29] = in[51] & in2[51];
    assign P[29] = in[51] ^ in2[51];
    assign G[30] = in[50] & in2[50];
    assign P[30] = in[50] ^ in2[50];
    assign G[31] = in[49] & in2[49];
    assign P[31] = in[49] ^ in2[49];
    assign G[32] = in[48] & in2[48];
    assign P[32] = in[48] ^ in2[48];
    assign G[33] = in[47] & in2[47];
    assign P[33] = in[47] ^ in2[47];
    assign G[34] = in[46] & in2[46];
    assign P[34] = in[46] ^ in2[46];
    assign G[35] = in[45] & in2[45];
    assign P[35] = in[45] ^ in2[45];
    assign G[36] = in[44] & in2[44];
    assign P[36] = in[44] ^ in2[44];
    assign G[37] = in[43] & in2[43];
    assign P[37] = in[43] ^ in2[43];
    assign G[38] = in[42] & in2[42];
    assign P[38] = in[42] ^ in2[42];
    assign G[39] = in[41] & in2[41];
    assign P[39] = in[41] ^ in2[41];
    assign G[40] = in[40] & in2[40];
    assign P[40] = in[40] ^ in2[40];
    assign G[41] = in[39] & in2[39];
    assign P[41] = in[39] ^ in2[39];
    assign G[42] = in[38] & in2[38];
    assign P[42] = in[38] ^ in2[38];
    assign G[43] = in[37] & in2[37];
    assign P[43] = in[37] ^ in2[37];
    assign G[44] = in[36] & in2[36];
    assign P[44] = in[36] ^ in2[36];
    assign G[45] = in[35] & in2[35];
    assign P[45] = in[35] ^ in2[35];
    assign G[46] = in[34] & in2[34];
    assign P[46] = in[34] ^ in2[34];
    assign G[47] = in[33] & in2[33];
    assign P[47] = in[33] ^ in2[33];
    assign G[48] = in[32] & in2[32];
    assign P[48] = in[32] ^ in2[32];
    assign G[49] = in[31] & in2[31];
    assign P[49] = in[31] ^ in2[31];
    assign G[50] = in[30] & in2[30];
    assign P[50] = in[30] ^ in2[30];
    assign G[51] = in[29] & in2[29];
    assign P[51] = in[29] ^ in2[29];
    assign G[52] = in[28] & in2[28];
    assign P[52] = in[28] ^ in2[28];
    assign G[53] = in[27] & in2[27];
    assign P[53] = in[27] ^ in2[27];
    assign G[54] = in[26] & in2[26];
    assign P[54] = in[26] ^ in2[26];
    assign G[55] = in[25] & in2[25];
    assign P[55] = in[25] ^ in2[25];
    assign G[56] = in[24] & in2[24];
    assign P[56] = in[24] ^ in2[24];
    assign G[57] = in[23] & in2[23];
    assign P[57] = in[23] ^ in2[23];
    assign G[58] = in[22] & in2[22];
    assign P[58] = in[22] ^ in2[22];
    assign G[59] = in[21] & in2[21];
    assign P[59] = in[21] ^ in2[21];
    assign G[60] = in[20] & in2[20];
    assign P[60] = in[20] ^ in2[20];
    assign G[61] = in[19] & in2[19];
    assign P[61] = in[19] ^ in2[19];
    assign G[62] = in[18] & in2[18];
    assign P[62] = in[18] ^ in2[18];
    assign G[63] = in[17] & in2[17];
    assign P[63] = in[17] ^ in2[17];
    assign G[64] = in[16] & in2[16];
    assign P[64] = in[16] ^ in2[16];
    assign G[65] = in[15] & in2[15];
    assign P[65] = in[15] ^ in2[15];
    assign G[66] = in[14] & in2[14];
    assign P[66] = in[14] ^ in2[14];
    assign G[67] = in[13] & in2[13];
    assign P[67] = in[13] ^ in2[13];
    assign G[68] = in[12] & in2[12];
    assign P[68] = in[12] ^ in2[12];
    assign G[69] = in[11] & in2[11];
    assign P[69] = in[11] ^ in2[11];
    assign G[70] = in[10] & in2[10];
    assign P[70] = in[10] ^ in2[10];
    assign G[71] = in[9] & in2[9];
    assign P[71] = in[9] ^ in2[9];
    assign G[72] = in[8] & in2[8];
    assign P[72] = in[8] ^ in2[8];
    assign G[73] = in[7] & in2[7];
    assign P[73] = in[7] ^ in2[7];
    assign G[74] = in[6] & in2[6];
    assign P[74] = in[6] ^ in2[6];
    assign G[75] = in[5] & in2[5];
    assign P[75] = in[5] ^ in2[5];
    assign G[76] = in[4] & in2[4];
    assign P[76] = in[4] ^ in2[4];
    assign G[77] = in[3] & in2[3];
    assign P[77] = in[3] ^ in2[3];
    assign G[78] = in[2] & in2[2];
    assign P[78] = in[2] ^ in2[2];
    assign G[79] = in[1] & in2[1];
    assign P[79] = in[1] ^ in2[1];
    assign G[80] = in[0] & in2[0];
    assign P[80] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign C[80] = G[79] | (P[79] & C[79]);
    assign cout = G[80] | (P[80] & C[80]);
    assign sum = P ^ C;
endmodule

module CLA80(output [79:0] sum, output cout, input [79:0] in1, input [79:0] in2;

    wire[79:0] G;
    wire[79:0] C;
    wire[79:0] P;

    assign G[0] = in[79] & in2[79];
    assign P[0] = in[79] ^ in2[79];
    assign G[1] = in[78] & in2[78];
    assign P[1] = in[78] ^ in2[78];
    assign G[2] = in[77] & in2[77];
    assign P[2] = in[77] ^ in2[77];
    assign G[3] = in[76] & in2[76];
    assign P[3] = in[76] ^ in2[76];
    assign G[4] = in[75] & in2[75];
    assign P[4] = in[75] ^ in2[75];
    assign G[5] = in[74] & in2[74];
    assign P[5] = in[74] ^ in2[74];
    assign G[6] = in[73] & in2[73];
    assign P[6] = in[73] ^ in2[73];
    assign G[7] = in[72] & in2[72];
    assign P[7] = in[72] ^ in2[72];
    assign G[8] = in[71] & in2[71];
    assign P[8] = in[71] ^ in2[71];
    assign G[9] = in[70] & in2[70];
    assign P[9] = in[70] ^ in2[70];
    assign G[10] = in[69] & in2[69];
    assign P[10] = in[69] ^ in2[69];
    assign G[11] = in[68] & in2[68];
    assign P[11] = in[68] ^ in2[68];
    assign G[12] = in[67] & in2[67];
    assign P[12] = in[67] ^ in2[67];
    assign G[13] = in[66] & in2[66];
    assign P[13] = in[66] ^ in2[66];
    assign G[14] = in[65] & in2[65];
    assign P[14] = in[65] ^ in2[65];
    assign G[15] = in[64] & in2[64];
    assign P[15] = in[64] ^ in2[64];
    assign G[16] = in[63] & in2[63];
    assign P[16] = in[63] ^ in2[63];
    assign G[17] = in[62] & in2[62];
    assign P[17] = in[62] ^ in2[62];
    assign G[18] = in[61] & in2[61];
    assign P[18] = in[61] ^ in2[61];
    assign G[19] = in[60] & in2[60];
    assign P[19] = in[60] ^ in2[60];
    assign G[20] = in[59] & in2[59];
    assign P[20] = in[59] ^ in2[59];
    assign G[21] = in[58] & in2[58];
    assign P[21] = in[58] ^ in2[58];
    assign G[22] = in[57] & in2[57];
    assign P[22] = in[57] ^ in2[57];
    assign G[23] = in[56] & in2[56];
    assign P[23] = in[56] ^ in2[56];
    assign G[24] = in[55] & in2[55];
    assign P[24] = in[55] ^ in2[55];
    assign G[25] = in[54] & in2[54];
    assign P[25] = in[54] ^ in2[54];
    assign G[26] = in[53] & in2[53];
    assign P[26] = in[53] ^ in2[53];
    assign G[27] = in[52] & in2[52];
    assign P[27] = in[52] ^ in2[52];
    assign G[28] = in[51] & in2[51];
    assign P[28] = in[51] ^ in2[51];
    assign G[29] = in[50] & in2[50];
    assign P[29] = in[50] ^ in2[50];
    assign G[30] = in[49] & in2[49];
    assign P[30] = in[49] ^ in2[49];
    assign G[31] = in[48] & in2[48];
    assign P[31] = in[48] ^ in2[48];
    assign G[32] = in[47] & in2[47];
    assign P[32] = in[47] ^ in2[47];
    assign G[33] = in[46] & in2[46];
    assign P[33] = in[46] ^ in2[46];
    assign G[34] = in[45] & in2[45];
    assign P[34] = in[45] ^ in2[45];
    assign G[35] = in[44] & in2[44];
    assign P[35] = in[44] ^ in2[44];
    assign G[36] = in[43] & in2[43];
    assign P[36] = in[43] ^ in2[43];
    assign G[37] = in[42] & in2[42];
    assign P[37] = in[42] ^ in2[42];
    assign G[38] = in[41] & in2[41];
    assign P[38] = in[41] ^ in2[41];
    assign G[39] = in[40] & in2[40];
    assign P[39] = in[40] ^ in2[40];
    assign G[40] = in[39] & in2[39];
    assign P[40] = in[39] ^ in2[39];
    assign G[41] = in[38] & in2[38];
    assign P[41] = in[38] ^ in2[38];
    assign G[42] = in[37] & in2[37];
    assign P[42] = in[37] ^ in2[37];
    assign G[43] = in[36] & in2[36];
    assign P[43] = in[36] ^ in2[36];
    assign G[44] = in[35] & in2[35];
    assign P[44] = in[35] ^ in2[35];
    assign G[45] = in[34] & in2[34];
    assign P[45] = in[34] ^ in2[34];
    assign G[46] = in[33] & in2[33];
    assign P[46] = in[33] ^ in2[33];
    assign G[47] = in[32] & in2[32];
    assign P[47] = in[32] ^ in2[32];
    assign G[48] = in[31] & in2[31];
    assign P[48] = in[31] ^ in2[31];
    assign G[49] = in[30] & in2[30];
    assign P[49] = in[30] ^ in2[30];
    assign G[50] = in[29] & in2[29];
    assign P[50] = in[29] ^ in2[29];
    assign G[51] = in[28] & in2[28];
    assign P[51] = in[28] ^ in2[28];
    assign G[52] = in[27] & in2[27];
    assign P[52] = in[27] ^ in2[27];
    assign G[53] = in[26] & in2[26];
    assign P[53] = in[26] ^ in2[26];
    assign G[54] = in[25] & in2[25];
    assign P[54] = in[25] ^ in2[25];
    assign G[55] = in[24] & in2[24];
    assign P[55] = in[24] ^ in2[24];
    assign G[56] = in[23] & in2[23];
    assign P[56] = in[23] ^ in2[23];
    assign G[57] = in[22] & in2[22];
    assign P[57] = in[22] ^ in2[22];
    assign G[58] = in[21] & in2[21];
    assign P[58] = in[21] ^ in2[21];
    assign G[59] = in[20] & in2[20];
    assign P[59] = in[20] ^ in2[20];
    assign G[60] = in[19] & in2[19];
    assign P[60] = in[19] ^ in2[19];
    assign G[61] = in[18] & in2[18];
    assign P[61] = in[18] ^ in2[18];
    assign G[62] = in[17] & in2[17];
    assign P[62] = in[17] ^ in2[17];
    assign G[63] = in[16] & in2[16];
    assign P[63] = in[16] ^ in2[16];
    assign G[64] = in[15] & in2[15];
    assign P[64] = in[15] ^ in2[15];
    assign G[65] = in[14] & in2[14];
    assign P[65] = in[14] ^ in2[14];
    assign G[66] = in[13] & in2[13];
    assign P[66] = in[13] ^ in2[13];
    assign G[67] = in[12] & in2[12];
    assign P[67] = in[12] ^ in2[12];
    assign G[68] = in[11] & in2[11];
    assign P[68] = in[11] ^ in2[11];
    assign G[69] = in[10] & in2[10];
    assign P[69] = in[10] ^ in2[10];
    assign G[70] = in[9] & in2[9];
    assign P[70] = in[9] ^ in2[9];
    assign G[71] = in[8] & in2[8];
    assign P[71] = in[8] ^ in2[8];
    assign G[72] = in[7] & in2[7];
    assign P[72] = in[7] ^ in2[7];
    assign G[73] = in[6] & in2[6];
    assign P[73] = in[6] ^ in2[6];
    assign G[74] = in[5] & in2[5];
    assign P[74] = in[5] ^ in2[5];
    assign G[75] = in[4] & in2[4];
    assign P[75] = in[4] ^ in2[4];
    assign G[76] = in[3] & in2[3];
    assign P[76] = in[3] ^ in2[3];
    assign G[77] = in[2] & in2[2];
    assign P[77] = in[2] ^ in2[2];
    assign G[78] = in[1] & in2[1];
    assign P[78] = in[1] ^ in2[1];
    assign G[79] = in[0] & in2[0];
    assign P[79] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign C[79] = G[78] | (P[78] & C[78]);
    assign cout = G[79] | (P[79] & C[79]);
    assign sum = P ^ C;
endmodule

module CLA79(output [78:0] sum, output cout, input [78:0] in1, input [78:0] in2;

    wire[78:0] G;
    wire[78:0] C;
    wire[78:0] P;

    assign G[0] = in[78] & in2[78];
    assign P[0] = in[78] ^ in2[78];
    assign G[1] = in[77] & in2[77];
    assign P[1] = in[77] ^ in2[77];
    assign G[2] = in[76] & in2[76];
    assign P[2] = in[76] ^ in2[76];
    assign G[3] = in[75] & in2[75];
    assign P[3] = in[75] ^ in2[75];
    assign G[4] = in[74] & in2[74];
    assign P[4] = in[74] ^ in2[74];
    assign G[5] = in[73] & in2[73];
    assign P[5] = in[73] ^ in2[73];
    assign G[6] = in[72] & in2[72];
    assign P[6] = in[72] ^ in2[72];
    assign G[7] = in[71] & in2[71];
    assign P[7] = in[71] ^ in2[71];
    assign G[8] = in[70] & in2[70];
    assign P[8] = in[70] ^ in2[70];
    assign G[9] = in[69] & in2[69];
    assign P[9] = in[69] ^ in2[69];
    assign G[10] = in[68] & in2[68];
    assign P[10] = in[68] ^ in2[68];
    assign G[11] = in[67] & in2[67];
    assign P[11] = in[67] ^ in2[67];
    assign G[12] = in[66] & in2[66];
    assign P[12] = in[66] ^ in2[66];
    assign G[13] = in[65] & in2[65];
    assign P[13] = in[65] ^ in2[65];
    assign G[14] = in[64] & in2[64];
    assign P[14] = in[64] ^ in2[64];
    assign G[15] = in[63] & in2[63];
    assign P[15] = in[63] ^ in2[63];
    assign G[16] = in[62] & in2[62];
    assign P[16] = in[62] ^ in2[62];
    assign G[17] = in[61] & in2[61];
    assign P[17] = in[61] ^ in2[61];
    assign G[18] = in[60] & in2[60];
    assign P[18] = in[60] ^ in2[60];
    assign G[19] = in[59] & in2[59];
    assign P[19] = in[59] ^ in2[59];
    assign G[20] = in[58] & in2[58];
    assign P[20] = in[58] ^ in2[58];
    assign G[21] = in[57] & in2[57];
    assign P[21] = in[57] ^ in2[57];
    assign G[22] = in[56] & in2[56];
    assign P[22] = in[56] ^ in2[56];
    assign G[23] = in[55] & in2[55];
    assign P[23] = in[55] ^ in2[55];
    assign G[24] = in[54] & in2[54];
    assign P[24] = in[54] ^ in2[54];
    assign G[25] = in[53] & in2[53];
    assign P[25] = in[53] ^ in2[53];
    assign G[26] = in[52] & in2[52];
    assign P[26] = in[52] ^ in2[52];
    assign G[27] = in[51] & in2[51];
    assign P[27] = in[51] ^ in2[51];
    assign G[28] = in[50] & in2[50];
    assign P[28] = in[50] ^ in2[50];
    assign G[29] = in[49] & in2[49];
    assign P[29] = in[49] ^ in2[49];
    assign G[30] = in[48] & in2[48];
    assign P[30] = in[48] ^ in2[48];
    assign G[31] = in[47] & in2[47];
    assign P[31] = in[47] ^ in2[47];
    assign G[32] = in[46] & in2[46];
    assign P[32] = in[46] ^ in2[46];
    assign G[33] = in[45] & in2[45];
    assign P[33] = in[45] ^ in2[45];
    assign G[34] = in[44] & in2[44];
    assign P[34] = in[44] ^ in2[44];
    assign G[35] = in[43] & in2[43];
    assign P[35] = in[43] ^ in2[43];
    assign G[36] = in[42] & in2[42];
    assign P[36] = in[42] ^ in2[42];
    assign G[37] = in[41] & in2[41];
    assign P[37] = in[41] ^ in2[41];
    assign G[38] = in[40] & in2[40];
    assign P[38] = in[40] ^ in2[40];
    assign G[39] = in[39] & in2[39];
    assign P[39] = in[39] ^ in2[39];
    assign G[40] = in[38] & in2[38];
    assign P[40] = in[38] ^ in2[38];
    assign G[41] = in[37] & in2[37];
    assign P[41] = in[37] ^ in2[37];
    assign G[42] = in[36] & in2[36];
    assign P[42] = in[36] ^ in2[36];
    assign G[43] = in[35] & in2[35];
    assign P[43] = in[35] ^ in2[35];
    assign G[44] = in[34] & in2[34];
    assign P[44] = in[34] ^ in2[34];
    assign G[45] = in[33] & in2[33];
    assign P[45] = in[33] ^ in2[33];
    assign G[46] = in[32] & in2[32];
    assign P[46] = in[32] ^ in2[32];
    assign G[47] = in[31] & in2[31];
    assign P[47] = in[31] ^ in2[31];
    assign G[48] = in[30] & in2[30];
    assign P[48] = in[30] ^ in2[30];
    assign G[49] = in[29] & in2[29];
    assign P[49] = in[29] ^ in2[29];
    assign G[50] = in[28] & in2[28];
    assign P[50] = in[28] ^ in2[28];
    assign G[51] = in[27] & in2[27];
    assign P[51] = in[27] ^ in2[27];
    assign G[52] = in[26] & in2[26];
    assign P[52] = in[26] ^ in2[26];
    assign G[53] = in[25] & in2[25];
    assign P[53] = in[25] ^ in2[25];
    assign G[54] = in[24] & in2[24];
    assign P[54] = in[24] ^ in2[24];
    assign G[55] = in[23] & in2[23];
    assign P[55] = in[23] ^ in2[23];
    assign G[56] = in[22] & in2[22];
    assign P[56] = in[22] ^ in2[22];
    assign G[57] = in[21] & in2[21];
    assign P[57] = in[21] ^ in2[21];
    assign G[58] = in[20] & in2[20];
    assign P[58] = in[20] ^ in2[20];
    assign G[59] = in[19] & in2[19];
    assign P[59] = in[19] ^ in2[19];
    assign G[60] = in[18] & in2[18];
    assign P[60] = in[18] ^ in2[18];
    assign G[61] = in[17] & in2[17];
    assign P[61] = in[17] ^ in2[17];
    assign G[62] = in[16] & in2[16];
    assign P[62] = in[16] ^ in2[16];
    assign G[63] = in[15] & in2[15];
    assign P[63] = in[15] ^ in2[15];
    assign G[64] = in[14] & in2[14];
    assign P[64] = in[14] ^ in2[14];
    assign G[65] = in[13] & in2[13];
    assign P[65] = in[13] ^ in2[13];
    assign G[66] = in[12] & in2[12];
    assign P[66] = in[12] ^ in2[12];
    assign G[67] = in[11] & in2[11];
    assign P[67] = in[11] ^ in2[11];
    assign G[68] = in[10] & in2[10];
    assign P[68] = in[10] ^ in2[10];
    assign G[69] = in[9] & in2[9];
    assign P[69] = in[9] ^ in2[9];
    assign G[70] = in[8] & in2[8];
    assign P[70] = in[8] ^ in2[8];
    assign G[71] = in[7] & in2[7];
    assign P[71] = in[7] ^ in2[7];
    assign G[72] = in[6] & in2[6];
    assign P[72] = in[6] ^ in2[6];
    assign G[73] = in[5] & in2[5];
    assign P[73] = in[5] ^ in2[5];
    assign G[74] = in[4] & in2[4];
    assign P[74] = in[4] ^ in2[4];
    assign G[75] = in[3] & in2[3];
    assign P[75] = in[3] ^ in2[3];
    assign G[76] = in[2] & in2[2];
    assign P[76] = in[2] ^ in2[2];
    assign G[77] = in[1] & in2[1];
    assign P[77] = in[1] ^ in2[1];
    assign G[78] = in[0] & in2[0];
    assign P[78] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign C[78] = G[77] | (P[77] & C[77]);
    assign cout = G[78] | (P[78] & C[78]);
    assign sum = P ^ C;
endmodule

module CLA78(output [77:0] sum, output cout, input [77:0] in1, input [77:0] in2;

    wire[77:0] G;
    wire[77:0] C;
    wire[77:0] P;

    assign G[0] = in[77] & in2[77];
    assign P[0] = in[77] ^ in2[77];
    assign G[1] = in[76] & in2[76];
    assign P[1] = in[76] ^ in2[76];
    assign G[2] = in[75] & in2[75];
    assign P[2] = in[75] ^ in2[75];
    assign G[3] = in[74] & in2[74];
    assign P[3] = in[74] ^ in2[74];
    assign G[4] = in[73] & in2[73];
    assign P[4] = in[73] ^ in2[73];
    assign G[5] = in[72] & in2[72];
    assign P[5] = in[72] ^ in2[72];
    assign G[6] = in[71] & in2[71];
    assign P[6] = in[71] ^ in2[71];
    assign G[7] = in[70] & in2[70];
    assign P[7] = in[70] ^ in2[70];
    assign G[8] = in[69] & in2[69];
    assign P[8] = in[69] ^ in2[69];
    assign G[9] = in[68] & in2[68];
    assign P[9] = in[68] ^ in2[68];
    assign G[10] = in[67] & in2[67];
    assign P[10] = in[67] ^ in2[67];
    assign G[11] = in[66] & in2[66];
    assign P[11] = in[66] ^ in2[66];
    assign G[12] = in[65] & in2[65];
    assign P[12] = in[65] ^ in2[65];
    assign G[13] = in[64] & in2[64];
    assign P[13] = in[64] ^ in2[64];
    assign G[14] = in[63] & in2[63];
    assign P[14] = in[63] ^ in2[63];
    assign G[15] = in[62] & in2[62];
    assign P[15] = in[62] ^ in2[62];
    assign G[16] = in[61] & in2[61];
    assign P[16] = in[61] ^ in2[61];
    assign G[17] = in[60] & in2[60];
    assign P[17] = in[60] ^ in2[60];
    assign G[18] = in[59] & in2[59];
    assign P[18] = in[59] ^ in2[59];
    assign G[19] = in[58] & in2[58];
    assign P[19] = in[58] ^ in2[58];
    assign G[20] = in[57] & in2[57];
    assign P[20] = in[57] ^ in2[57];
    assign G[21] = in[56] & in2[56];
    assign P[21] = in[56] ^ in2[56];
    assign G[22] = in[55] & in2[55];
    assign P[22] = in[55] ^ in2[55];
    assign G[23] = in[54] & in2[54];
    assign P[23] = in[54] ^ in2[54];
    assign G[24] = in[53] & in2[53];
    assign P[24] = in[53] ^ in2[53];
    assign G[25] = in[52] & in2[52];
    assign P[25] = in[52] ^ in2[52];
    assign G[26] = in[51] & in2[51];
    assign P[26] = in[51] ^ in2[51];
    assign G[27] = in[50] & in2[50];
    assign P[27] = in[50] ^ in2[50];
    assign G[28] = in[49] & in2[49];
    assign P[28] = in[49] ^ in2[49];
    assign G[29] = in[48] & in2[48];
    assign P[29] = in[48] ^ in2[48];
    assign G[30] = in[47] & in2[47];
    assign P[30] = in[47] ^ in2[47];
    assign G[31] = in[46] & in2[46];
    assign P[31] = in[46] ^ in2[46];
    assign G[32] = in[45] & in2[45];
    assign P[32] = in[45] ^ in2[45];
    assign G[33] = in[44] & in2[44];
    assign P[33] = in[44] ^ in2[44];
    assign G[34] = in[43] & in2[43];
    assign P[34] = in[43] ^ in2[43];
    assign G[35] = in[42] & in2[42];
    assign P[35] = in[42] ^ in2[42];
    assign G[36] = in[41] & in2[41];
    assign P[36] = in[41] ^ in2[41];
    assign G[37] = in[40] & in2[40];
    assign P[37] = in[40] ^ in2[40];
    assign G[38] = in[39] & in2[39];
    assign P[38] = in[39] ^ in2[39];
    assign G[39] = in[38] & in2[38];
    assign P[39] = in[38] ^ in2[38];
    assign G[40] = in[37] & in2[37];
    assign P[40] = in[37] ^ in2[37];
    assign G[41] = in[36] & in2[36];
    assign P[41] = in[36] ^ in2[36];
    assign G[42] = in[35] & in2[35];
    assign P[42] = in[35] ^ in2[35];
    assign G[43] = in[34] & in2[34];
    assign P[43] = in[34] ^ in2[34];
    assign G[44] = in[33] & in2[33];
    assign P[44] = in[33] ^ in2[33];
    assign G[45] = in[32] & in2[32];
    assign P[45] = in[32] ^ in2[32];
    assign G[46] = in[31] & in2[31];
    assign P[46] = in[31] ^ in2[31];
    assign G[47] = in[30] & in2[30];
    assign P[47] = in[30] ^ in2[30];
    assign G[48] = in[29] & in2[29];
    assign P[48] = in[29] ^ in2[29];
    assign G[49] = in[28] & in2[28];
    assign P[49] = in[28] ^ in2[28];
    assign G[50] = in[27] & in2[27];
    assign P[50] = in[27] ^ in2[27];
    assign G[51] = in[26] & in2[26];
    assign P[51] = in[26] ^ in2[26];
    assign G[52] = in[25] & in2[25];
    assign P[52] = in[25] ^ in2[25];
    assign G[53] = in[24] & in2[24];
    assign P[53] = in[24] ^ in2[24];
    assign G[54] = in[23] & in2[23];
    assign P[54] = in[23] ^ in2[23];
    assign G[55] = in[22] & in2[22];
    assign P[55] = in[22] ^ in2[22];
    assign G[56] = in[21] & in2[21];
    assign P[56] = in[21] ^ in2[21];
    assign G[57] = in[20] & in2[20];
    assign P[57] = in[20] ^ in2[20];
    assign G[58] = in[19] & in2[19];
    assign P[58] = in[19] ^ in2[19];
    assign G[59] = in[18] & in2[18];
    assign P[59] = in[18] ^ in2[18];
    assign G[60] = in[17] & in2[17];
    assign P[60] = in[17] ^ in2[17];
    assign G[61] = in[16] & in2[16];
    assign P[61] = in[16] ^ in2[16];
    assign G[62] = in[15] & in2[15];
    assign P[62] = in[15] ^ in2[15];
    assign G[63] = in[14] & in2[14];
    assign P[63] = in[14] ^ in2[14];
    assign G[64] = in[13] & in2[13];
    assign P[64] = in[13] ^ in2[13];
    assign G[65] = in[12] & in2[12];
    assign P[65] = in[12] ^ in2[12];
    assign G[66] = in[11] & in2[11];
    assign P[66] = in[11] ^ in2[11];
    assign G[67] = in[10] & in2[10];
    assign P[67] = in[10] ^ in2[10];
    assign G[68] = in[9] & in2[9];
    assign P[68] = in[9] ^ in2[9];
    assign G[69] = in[8] & in2[8];
    assign P[69] = in[8] ^ in2[8];
    assign G[70] = in[7] & in2[7];
    assign P[70] = in[7] ^ in2[7];
    assign G[71] = in[6] & in2[6];
    assign P[71] = in[6] ^ in2[6];
    assign G[72] = in[5] & in2[5];
    assign P[72] = in[5] ^ in2[5];
    assign G[73] = in[4] & in2[4];
    assign P[73] = in[4] ^ in2[4];
    assign G[74] = in[3] & in2[3];
    assign P[74] = in[3] ^ in2[3];
    assign G[75] = in[2] & in2[2];
    assign P[75] = in[2] ^ in2[2];
    assign G[76] = in[1] & in2[1];
    assign P[76] = in[1] ^ in2[1];
    assign G[77] = in[0] & in2[0];
    assign P[77] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign C[77] = G[76] | (P[76] & C[76]);
    assign cout = G[77] | (P[77] & C[77]);
    assign sum = P ^ C;
endmodule

module CLA77(output [76:0] sum, output cout, input [76:0] in1, input [76:0] in2;

    wire[76:0] G;
    wire[76:0] C;
    wire[76:0] P;

    assign G[0] = in[76] & in2[76];
    assign P[0] = in[76] ^ in2[76];
    assign G[1] = in[75] & in2[75];
    assign P[1] = in[75] ^ in2[75];
    assign G[2] = in[74] & in2[74];
    assign P[2] = in[74] ^ in2[74];
    assign G[3] = in[73] & in2[73];
    assign P[3] = in[73] ^ in2[73];
    assign G[4] = in[72] & in2[72];
    assign P[4] = in[72] ^ in2[72];
    assign G[5] = in[71] & in2[71];
    assign P[5] = in[71] ^ in2[71];
    assign G[6] = in[70] & in2[70];
    assign P[6] = in[70] ^ in2[70];
    assign G[7] = in[69] & in2[69];
    assign P[7] = in[69] ^ in2[69];
    assign G[8] = in[68] & in2[68];
    assign P[8] = in[68] ^ in2[68];
    assign G[9] = in[67] & in2[67];
    assign P[9] = in[67] ^ in2[67];
    assign G[10] = in[66] & in2[66];
    assign P[10] = in[66] ^ in2[66];
    assign G[11] = in[65] & in2[65];
    assign P[11] = in[65] ^ in2[65];
    assign G[12] = in[64] & in2[64];
    assign P[12] = in[64] ^ in2[64];
    assign G[13] = in[63] & in2[63];
    assign P[13] = in[63] ^ in2[63];
    assign G[14] = in[62] & in2[62];
    assign P[14] = in[62] ^ in2[62];
    assign G[15] = in[61] & in2[61];
    assign P[15] = in[61] ^ in2[61];
    assign G[16] = in[60] & in2[60];
    assign P[16] = in[60] ^ in2[60];
    assign G[17] = in[59] & in2[59];
    assign P[17] = in[59] ^ in2[59];
    assign G[18] = in[58] & in2[58];
    assign P[18] = in[58] ^ in2[58];
    assign G[19] = in[57] & in2[57];
    assign P[19] = in[57] ^ in2[57];
    assign G[20] = in[56] & in2[56];
    assign P[20] = in[56] ^ in2[56];
    assign G[21] = in[55] & in2[55];
    assign P[21] = in[55] ^ in2[55];
    assign G[22] = in[54] & in2[54];
    assign P[22] = in[54] ^ in2[54];
    assign G[23] = in[53] & in2[53];
    assign P[23] = in[53] ^ in2[53];
    assign G[24] = in[52] & in2[52];
    assign P[24] = in[52] ^ in2[52];
    assign G[25] = in[51] & in2[51];
    assign P[25] = in[51] ^ in2[51];
    assign G[26] = in[50] & in2[50];
    assign P[26] = in[50] ^ in2[50];
    assign G[27] = in[49] & in2[49];
    assign P[27] = in[49] ^ in2[49];
    assign G[28] = in[48] & in2[48];
    assign P[28] = in[48] ^ in2[48];
    assign G[29] = in[47] & in2[47];
    assign P[29] = in[47] ^ in2[47];
    assign G[30] = in[46] & in2[46];
    assign P[30] = in[46] ^ in2[46];
    assign G[31] = in[45] & in2[45];
    assign P[31] = in[45] ^ in2[45];
    assign G[32] = in[44] & in2[44];
    assign P[32] = in[44] ^ in2[44];
    assign G[33] = in[43] & in2[43];
    assign P[33] = in[43] ^ in2[43];
    assign G[34] = in[42] & in2[42];
    assign P[34] = in[42] ^ in2[42];
    assign G[35] = in[41] & in2[41];
    assign P[35] = in[41] ^ in2[41];
    assign G[36] = in[40] & in2[40];
    assign P[36] = in[40] ^ in2[40];
    assign G[37] = in[39] & in2[39];
    assign P[37] = in[39] ^ in2[39];
    assign G[38] = in[38] & in2[38];
    assign P[38] = in[38] ^ in2[38];
    assign G[39] = in[37] & in2[37];
    assign P[39] = in[37] ^ in2[37];
    assign G[40] = in[36] & in2[36];
    assign P[40] = in[36] ^ in2[36];
    assign G[41] = in[35] & in2[35];
    assign P[41] = in[35] ^ in2[35];
    assign G[42] = in[34] & in2[34];
    assign P[42] = in[34] ^ in2[34];
    assign G[43] = in[33] & in2[33];
    assign P[43] = in[33] ^ in2[33];
    assign G[44] = in[32] & in2[32];
    assign P[44] = in[32] ^ in2[32];
    assign G[45] = in[31] & in2[31];
    assign P[45] = in[31] ^ in2[31];
    assign G[46] = in[30] & in2[30];
    assign P[46] = in[30] ^ in2[30];
    assign G[47] = in[29] & in2[29];
    assign P[47] = in[29] ^ in2[29];
    assign G[48] = in[28] & in2[28];
    assign P[48] = in[28] ^ in2[28];
    assign G[49] = in[27] & in2[27];
    assign P[49] = in[27] ^ in2[27];
    assign G[50] = in[26] & in2[26];
    assign P[50] = in[26] ^ in2[26];
    assign G[51] = in[25] & in2[25];
    assign P[51] = in[25] ^ in2[25];
    assign G[52] = in[24] & in2[24];
    assign P[52] = in[24] ^ in2[24];
    assign G[53] = in[23] & in2[23];
    assign P[53] = in[23] ^ in2[23];
    assign G[54] = in[22] & in2[22];
    assign P[54] = in[22] ^ in2[22];
    assign G[55] = in[21] & in2[21];
    assign P[55] = in[21] ^ in2[21];
    assign G[56] = in[20] & in2[20];
    assign P[56] = in[20] ^ in2[20];
    assign G[57] = in[19] & in2[19];
    assign P[57] = in[19] ^ in2[19];
    assign G[58] = in[18] & in2[18];
    assign P[58] = in[18] ^ in2[18];
    assign G[59] = in[17] & in2[17];
    assign P[59] = in[17] ^ in2[17];
    assign G[60] = in[16] & in2[16];
    assign P[60] = in[16] ^ in2[16];
    assign G[61] = in[15] & in2[15];
    assign P[61] = in[15] ^ in2[15];
    assign G[62] = in[14] & in2[14];
    assign P[62] = in[14] ^ in2[14];
    assign G[63] = in[13] & in2[13];
    assign P[63] = in[13] ^ in2[13];
    assign G[64] = in[12] & in2[12];
    assign P[64] = in[12] ^ in2[12];
    assign G[65] = in[11] & in2[11];
    assign P[65] = in[11] ^ in2[11];
    assign G[66] = in[10] & in2[10];
    assign P[66] = in[10] ^ in2[10];
    assign G[67] = in[9] & in2[9];
    assign P[67] = in[9] ^ in2[9];
    assign G[68] = in[8] & in2[8];
    assign P[68] = in[8] ^ in2[8];
    assign G[69] = in[7] & in2[7];
    assign P[69] = in[7] ^ in2[7];
    assign G[70] = in[6] & in2[6];
    assign P[70] = in[6] ^ in2[6];
    assign G[71] = in[5] & in2[5];
    assign P[71] = in[5] ^ in2[5];
    assign G[72] = in[4] & in2[4];
    assign P[72] = in[4] ^ in2[4];
    assign G[73] = in[3] & in2[3];
    assign P[73] = in[3] ^ in2[3];
    assign G[74] = in[2] & in2[2];
    assign P[74] = in[2] ^ in2[2];
    assign G[75] = in[1] & in2[1];
    assign P[75] = in[1] ^ in2[1];
    assign G[76] = in[0] & in2[0];
    assign P[76] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign C[76] = G[75] | (P[75] & C[75]);
    assign cout = G[76] | (P[76] & C[76]);
    assign sum = P ^ C;
endmodule

module CLA76(output [75:0] sum, output cout, input [75:0] in1, input [75:0] in2;

    wire[75:0] G;
    wire[75:0] C;
    wire[75:0] P;

    assign G[0] = in[75] & in2[75];
    assign P[0] = in[75] ^ in2[75];
    assign G[1] = in[74] & in2[74];
    assign P[1] = in[74] ^ in2[74];
    assign G[2] = in[73] & in2[73];
    assign P[2] = in[73] ^ in2[73];
    assign G[3] = in[72] & in2[72];
    assign P[3] = in[72] ^ in2[72];
    assign G[4] = in[71] & in2[71];
    assign P[4] = in[71] ^ in2[71];
    assign G[5] = in[70] & in2[70];
    assign P[5] = in[70] ^ in2[70];
    assign G[6] = in[69] & in2[69];
    assign P[6] = in[69] ^ in2[69];
    assign G[7] = in[68] & in2[68];
    assign P[7] = in[68] ^ in2[68];
    assign G[8] = in[67] & in2[67];
    assign P[8] = in[67] ^ in2[67];
    assign G[9] = in[66] & in2[66];
    assign P[9] = in[66] ^ in2[66];
    assign G[10] = in[65] & in2[65];
    assign P[10] = in[65] ^ in2[65];
    assign G[11] = in[64] & in2[64];
    assign P[11] = in[64] ^ in2[64];
    assign G[12] = in[63] & in2[63];
    assign P[12] = in[63] ^ in2[63];
    assign G[13] = in[62] & in2[62];
    assign P[13] = in[62] ^ in2[62];
    assign G[14] = in[61] & in2[61];
    assign P[14] = in[61] ^ in2[61];
    assign G[15] = in[60] & in2[60];
    assign P[15] = in[60] ^ in2[60];
    assign G[16] = in[59] & in2[59];
    assign P[16] = in[59] ^ in2[59];
    assign G[17] = in[58] & in2[58];
    assign P[17] = in[58] ^ in2[58];
    assign G[18] = in[57] & in2[57];
    assign P[18] = in[57] ^ in2[57];
    assign G[19] = in[56] & in2[56];
    assign P[19] = in[56] ^ in2[56];
    assign G[20] = in[55] & in2[55];
    assign P[20] = in[55] ^ in2[55];
    assign G[21] = in[54] & in2[54];
    assign P[21] = in[54] ^ in2[54];
    assign G[22] = in[53] & in2[53];
    assign P[22] = in[53] ^ in2[53];
    assign G[23] = in[52] & in2[52];
    assign P[23] = in[52] ^ in2[52];
    assign G[24] = in[51] & in2[51];
    assign P[24] = in[51] ^ in2[51];
    assign G[25] = in[50] & in2[50];
    assign P[25] = in[50] ^ in2[50];
    assign G[26] = in[49] & in2[49];
    assign P[26] = in[49] ^ in2[49];
    assign G[27] = in[48] & in2[48];
    assign P[27] = in[48] ^ in2[48];
    assign G[28] = in[47] & in2[47];
    assign P[28] = in[47] ^ in2[47];
    assign G[29] = in[46] & in2[46];
    assign P[29] = in[46] ^ in2[46];
    assign G[30] = in[45] & in2[45];
    assign P[30] = in[45] ^ in2[45];
    assign G[31] = in[44] & in2[44];
    assign P[31] = in[44] ^ in2[44];
    assign G[32] = in[43] & in2[43];
    assign P[32] = in[43] ^ in2[43];
    assign G[33] = in[42] & in2[42];
    assign P[33] = in[42] ^ in2[42];
    assign G[34] = in[41] & in2[41];
    assign P[34] = in[41] ^ in2[41];
    assign G[35] = in[40] & in2[40];
    assign P[35] = in[40] ^ in2[40];
    assign G[36] = in[39] & in2[39];
    assign P[36] = in[39] ^ in2[39];
    assign G[37] = in[38] & in2[38];
    assign P[37] = in[38] ^ in2[38];
    assign G[38] = in[37] & in2[37];
    assign P[38] = in[37] ^ in2[37];
    assign G[39] = in[36] & in2[36];
    assign P[39] = in[36] ^ in2[36];
    assign G[40] = in[35] & in2[35];
    assign P[40] = in[35] ^ in2[35];
    assign G[41] = in[34] & in2[34];
    assign P[41] = in[34] ^ in2[34];
    assign G[42] = in[33] & in2[33];
    assign P[42] = in[33] ^ in2[33];
    assign G[43] = in[32] & in2[32];
    assign P[43] = in[32] ^ in2[32];
    assign G[44] = in[31] & in2[31];
    assign P[44] = in[31] ^ in2[31];
    assign G[45] = in[30] & in2[30];
    assign P[45] = in[30] ^ in2[30];
    assign G[46] = in[29] & in2[29];
    assign P[46] = in[29] ^ in2[29];
    assign G[47] = in[28] & in2[28];
    assign P[47] = in[28] ^ in2[28];
    assign G[48] = in[27] & in2[27];
    assign P[48] = in[27] ^ in2[27];
    assign G[49] = in[26] & in2[26];
    assign P[49] = in[26] ^ in2[26];
    assign G[50] = in[25] & in2[25];
    assign P[50] = in[25] ^ in2[25];
    assign G[51] = in[24] & in2[24];
    assign P[51] = in[24] ^ in2[24];
    assign G[52] = in[23] & in2[23];
    assign P[52] = in[23] ^ in2[23];
    assign G[53] = in[22] & in2[22];
    assign P[53] = in[22] ^ in2[22];
    assign G[54] = in[21] & in2[21];
    assign P[54] = in[21] ^ in2[21];
    assign G[55] = in[20] & in2[20];
    assign P[55] = in[20] ^ in2[20];
    assign G[56] = in[19] & in2[19];
    assign P[56] = in[19] ^ in2[19];
    assign G[57] = in[18] & in2[18];
    assign P[57] = in[18] ^ in2[18];
    assign G[58] = in[17] & in2[17];
    assign P[58] = in[17] ^ in2[17];
    assign G[59] = in[16] & in2[16];
    assign P[59] = in[16] ^ in2[16];
    assign G[60] = in[15] & in2[15];
    assign P[60] = in[15] ^ in2[15];
    assign G[61] = in[14] & in2[14];
    assign P[61] = in[14] ^ in2[14];
    assign G[62] = in[13] & in2[13];
    assign P[62] = in[13] ^ in2[13];
    assign G[63] = in[12] & in2[12];
    assign P[63] = in[12] ^ in2[12];
    assign G[64] = in[11] & in2[11];
    assign P[64] = in[11] ^ in2[11];
    assign G[65] = in[10] & in2[10];
    assign P[65] = in[10] ^ in2[10];
    assign G[66] = in[9] & in2[9];
    assign P[66] = in[9] ^ in2[9];
    assign G[67] = in[8] & in2[8];
    assign P[67] = in[8] ^ in2[8];
    assign G[68] = in[7] & in2[7];
    assign P[68] = in[7] ^ in2[7];
    assign G[69] = in[6] & in2[6];
    assign P[69] = in[6] ^ in2[6];
    assign G[70] = in[5] & in2[5];
    assign P[70] = in[5] ^ in2[5];
    assign G[71] = in[4] & in2[4];
    assign P[71] = in[4] ^ in2[4];
    assign G[72] = in[3] & in2[3];
    assign P[72] = in[3] ^ in2[3];
    assign G[73] = in[2] & in2[2];
    assign P[73] = in[2] ^ in2[2];
    assign G[74] = in[1] & in2[1];
    assign P[74] = in[1] ^ in2[1];
    assign G[75] = in[0] & in2[0];
    assign P[75] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign C[75] = G[74] | (P[74] & C[74]);
    assign cout = G[75] | (P[75] & C[75]);
    assign sum = P ^ C;
endmodule

module CLA75(output [74:0] sum, output cout, input [74:0] in1, input [74:0] in2;

    wire[74:0] G;
    wire[74:0] C;
    wire[74:0] P;

    assign G[0] = in[74] & in2[74];
    assign P[0] = in[74] ^ in2[74];
    assign G[1] = in[73] & in2[73];
    assign P[1] = in[73] ^ in2[73];
    assign G[2] = in[72] & in2[72];
    assign P[2] = in[72] ^ in2[72];
    assign G[3] = in[71] & in2[71];
    assign P[3] = in[71] ^ in2[71];
    assign G[4] = in[70] & in2[70];
    assign P[4] = in[70] ^ in2[70];
    assign G[5] = in[69] & in2[69];
    assign P[5] = in[69] ^ in2[69];
    assign G[6] = in[68] & in2[68];
    assign P[6] = in[68] ^ in2[68];
    assign G[7] = in[67] & in2[67];
    assign P[7] = in[67] ^ in2[67];
    assign G[8] = in[66] & in2[66];
    assign P[8] = in[66] ^ in2[66];
    assign G[9] = in[65] & in2[65];
    assign P[9] = in[65] ^ in2[65];
    assign G[10] = in[64] & in2[64];
    assign P[10] = in[64] ^ in2[64];
    assign G[11] = in[63] & in2[63];
    assign P[11] = in[63] ^ in2[63];
    assign G[12] = in[62] & in2[62];
    assign P[12] = in[62] ^ in2[62];
    assign G[13] = in[61] & in2[61];
    assign P[13] = in[61] ^ in2[61];
    assign G[14] = in[60] & in2[60];
    assign P[14] = in[60] ^ in2[60];
    assign G[15] = in[59] & in2[59];
    assign P[15] = in[59] ^ in2[59];
    assign G[16] = in[58] & in2[58];
    assign P[16] = in[58] ^ in2[58];
    assign G[17] = in[57] & in2[57];
    assign P[17] = in[57] ^ in2[57];
    assign G[18] = in[56] & in2[56];
    assign P[18] = in[56] ^ in2[56];
    assign G[19] = in[55] & in2[55];
    assign P[19] = in[55] ^ in2[55];
    assign G[20] = in[54] & in2[54];
    assign P[20] = in[54] ^ in2[54];
    assign G[21] = in[53] & in2[53];
    assign P[21] = in[53] ^ in2[53];
    assign G[22] = in[52] & in2[52];
    assign P[22] = in[52] ^ in2[52];
    assign G[23] = in[51] & in2[51];
    assign P[23] = in[51] ^ in2[51];
    assign G[24] = in[50] & in2[50];
    assign P[24] = in[50] ^ in2[50];
    assign G[25] = in[49] & in2[49];
    assign P[25] = in[49] ^ in2[49];
    assign G[26] = in[48] & in2[48];
    assign P[26] = in[48] ^ in2[48];
    assign G[27] = in[47] & in2[47];
    assign P[27] = in[47] ^ in2[47];
    assign G[28] = in[46] & in2[46];
    assign P[28] = in[46] ^ in2[46];
    assign G[29] = in[45] & in2[45];
    assign P[29] = in[45] ^ in2[45];
    assign G[30] = in[44] & in2[44];
    assign P[30] = in[44] ^ in2[44];
    assign G[31] = in[43] & in2[43];
    assign P[31] = in[43] ^ in2[43];
    assign G[32] = in[42] & in2[42];
    assign P[32] = in[42] ^ in2[42];
    assign G[33] = in[41] & in2[41];
    assign P[33] = in[41] ^ in2[41];
    assign G[34] = in[40] & in2[40];
    assign P[34] = in[40] ^ in2[40];
    assign G[35] = in[39] & in2[39];
    assign P[35] = in[39] ^ in2[39];
    assign G[36] = in[38] & in2[38];
    assign P[36] = in[38] ^ in2[38];
    assign G[37] = in[37] & in2[37];
    assign P[37] = in[37] ^ in2[37];
    assign G[38] = in[36] & in2[36];
    assign P[38] = in[36] ^ in2[36];
    assign G[39] = in[35] & in2[35];
    assign P[39] = in[35] ^ in2[35];
    assign G[40] = in[34] & in2[34];
    assign P[40] = in[34] ^ in2[34];
    assign G[41] = in[33] & in2[33];
    assign P[41] = in[33] ^ in2[33];
    assign G[42] = in[32] & in2[32];
    assign P[42] = in[32] ^ in2[32];
    assign G[43] = in[31] & in2[31];
    assign P[43] = in[31] ^ in2[31];
    assign G[44] = in[30] & in2[30];
    assign P[44] = in[30] ^ in2[30];
    assign G[45] = in[29] & in2[29];
    assign P[45] = in[29] ^ in2[29];
    assign G[46] = in[28] & in2[28];
    assign P[46] = in[28] ^ in2[28];
    assign G[47] = in[27] & in2[27];
    assign P[47] = in[27] ^ in2[27];
    assign G[48] = in[26] & in2[26];
    assign P[48] = in[26] ^ in2[26];
    assign G[49] = in[25] & in2[25];
    assign P[49] = in[25] ^ in2[25];
    assign G[50] = in[24] & in2[24];
    assign P[50] = in[24] ^ in2[24];
    assign G[51] = in[23] & in2[23];
    assign P[51] = in[23] ^ in2[23];
    assign G[52] = in[22] & in2[22];
    assign P[52] = in[22] ^ in2[22];
    assign G[53] = in[21] & in2[21];
    assign P[53] = in[21] ^ in2[21];
    assign G[54] = in[20] & in2[20];
    assign P[54] = in[20] ^ in2[20];
    assign G[55] = in[19] & in2[19];
    assign P[55] = in[19] ^ in2[19];
    assign G[56] = in[18] & in2[18];
    assign P[56] = in[18] ^ in2[18];
    assign G[57] = in[17] & in2[17];
    assign P[57] = in[17] ^ in2[17];
    assign G[58] = in[16] & in2[16];
    assign P[58] = in[16] ^ in2[16];
    assign G[59] = in[15] & in2[15];
    assign P[59] = in[15] ^ in2[15];
    assign G[60] = in[14] & in2[14];
    assign P[60] = in[14] ^ in2[14];
    assign G[61] = in[13] & in2[13];
    assign P[61] = in[13] ^ in2[13];
    assign G[62] = in[12] & in2[12];
    assign P[62] = in[12] ^ in2[12];
    assign G[63] = in[11] & in2[11];
    assign P[63] = in[11] ^ in2[11];
    assign G[64] = in[10] & in2[10];
    assign P[64] = in[10] ^ in2[10];
    assign G[65] = in[9] & in2[9];
    assign P[65] = in[9] ^ in2[9];
    assign G[66] = in[8] & in2[8];
    assign P[66] = in[8] ^ in2[8];
    assign G[67] = in[7] & in2[7];
    assign P[67] = in[7] ^ in2[7];
    assign G[68] = in[6] & in2[6];
    assign P[68] = in[6] ^ in2[6];
    assign G[69] = in[5] & in2[5];
    assign P[69] = in[5] ^ in2[5];
    assign G[70] = in[4] & in2[4];
    assign P[70] = in[4] ^ in2[4];
    assign G[71] = in[3] & in2[3];
    assign P[71] = in[3] ^ in2[3];
    assign G[72] = in[2] & in2[2];
    assign P[72] = in[2] ^ in2[2];
    assign G[73] = in[1] & in2[1];
    assign P[73] = in[1] ^ in2[1];
    assign G[74] = in[0] & in2[0];
    assign P[74] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign C[74] = G[73] | (P[73] & C[73]);
    assign cout = G[74] | (P[74] & C[74]);
    assign sum = P ^ C;
endmodule

module CLA74(output [73:0] sum, output cout, input [73:0] in1, input [73:0] in2;

    wire[73:0] G;
    wire[73:0] C;
    wire[73:0] P;

    assign G[0] = in[73] & in2[73];
    assign P[0] = in[73] ^ in2[73];
    assign G[1] = in[72] & in2[72];
    assign P[1] = in[72] ^ in2[72];
    assign G[2] = in[71] & in2[71];
    assign P[2] = in[71] ^ in2[71];
    assign G[3] = in[70] & in2[70];
    assign P[3] = in[70] ^ in2[70];
    assign G[4] = in[69] & in2[69];
    assign P[4] = in[69] ^ in2[69];
    assign G[5] = in[68] & in2[68];
    assign P[5] = in[68] ^ in2[68];
    assign G[6] = in[67] & in2[67];
    assign P[6] = in[67] ^ in2[67];
    assign G[7] = in[66] & in2[66];
    assign P[7] = in[66] ^ in2[66];
    assign G[8] = in[65] & in2[65];
    assign P[8] = in[65] ^ in2[65];
    assign G[9] = in[64] & in2[64];
    assign P[9] = in[64] ^ in2[64];
    assign G[10] = in[63] & in2[63];
    assign P[10] = in[63] ^ in2[63];
    assign G[11] = in[62] & in2[62];
    assign P[11] = in[62] ^ in2[62];
    assign G[12] = in[61] & in2[61];
    assign P[12] = in[61] ^ in2[61];
    assign G[13] = in[60] & in2[60];
    assign P[13] = in[60] ^ in2[60];
    assign G[14] = in[59] & in2[59];
    assign P[14] = in[59] ^ in2[59];
    assign G[15] = in[58] & in2[58];
    assign P[15] = in[58] ^ in2[58];
    assign G[16] = in[57] & in2[57];
    assign P[16] = in[57] ^ in2[57];
    assign G[17] = in[56] & in2[56];
    assign P[17] = in[56] ^ in2[56];
    assign G[18] = in[55] & in2[55];
    assign P[18] = in[55] ^ in2[55];
    assign G[19] = in[54] & in2[54];
    assign P[19] = in[54] ^ in2[54];
    assign G[20] = in[53] & in2[53];
    assign P[20] = in[53] ^ in2[53];
    assign G[21] = in[52] & in2[52];
    assign P[21] = in[52] ^ in2[52];
    assign G[22] = in[51] & in2[51];
    assign P[22] = in[51] ^ in2[51];
    assign G[23] = in[50] & in2[50];
    assign P[23] = in[50] ^ in2[50];
    assign G[24] = in[49] & in2[49];
    assign P[24] = in[49] ^ in2[49];
    assign G[25] = in[48] & in2[48];
    assign P[25] = in[48] ^ in2[48];
    assign G[26] = in[47] & in2[47];
    assign P[26] = in[47] ^ in2[47];
    assign G[27] = in[46] & in2[46];
    assign P[27] = in[46] ^ in2[46];
    assign G[28] = in[45] & in2[45];
    assign P[28] = in[45] ^ in2[45];
    assign G[29] = in[44] & in2[44];
    assign P[29] = in[44] ^ in2[44];
    assign G[30] = in[43] & in2[43];
    assign P[30] = in[43] ^ in2[43];
    assign G[31] = in[42] & in2[42];
    assign P[31] = in[42] ^ in2[42];
    assign G[32] = in[41] & in2[41];
    assign P[32] = in[41] ^ in2[41];
    assign G[33] = in[40] & in2[40];
    assign P[33] = in[40] ^ in2[40];
    assign G[34] = in[39] & in2[39];
    assign P[34] = in[39] ^ in2[39];
    assign G[35] = in[38] & in2[38];
    assign P[35] = in[38] ^ in2[38];
    assign G[36] = in[37] & in2[37];
    assign P[36] = in[37] ^ in2[37];
    assign G[37] = in[36] & in2[36];
    assign P[37] = in[36] ^ in2[36];
    assign G[38] = in[35] & in2[35];
    assign P[38] = in[35] ^ in2[35];
    assign G[39] = in[34] & in2[34];
    assign P[39] = in[34] ^ in2[34];
    assign G[40] = in[33] & in2[33];
    assign P[40] = in[33] ^ in2[33];
    assign G[41] = in[32] & in2[32];
    assign P[41] = in[32] ^ in2[32];
    assign G[42] = in[31] & in2[31];
    assign P[42] = in[31] ^ in2[31];
    assign G[43] = in[30] & in2[30];
    assign P[43] = in[30] ^ in2[30];
    assign G[44] = in[29] & in2[29];
    assign P[44] = in[29] ^ in2[29];
    assign G[45] = in[28] & in2[28];
    assign P[45] = in[28] ^ in2[28];
    assign G[46] = in[27] & in2[27];
    assign P[46] = in[27] ^ in2[27];
    assign G[47] = in[26] & in2[26];
    assign P[47] = in[26] ^ in2[26];
    assign G[48] = in[25] & in2[25];
    assign P[48] = in[25] ^ in2[25];
    assign G[49] = in[24] & in2[24];
    assign P[49] = in[24] ^ in2[24];
    assign G[50] = in[23] & in2[23];
    assign P[50] = in[23] ^ in2[23];
    assign G[51] = in[22] & in2[22];
    assign P[51] = in[22] ^ in2[22];
    assign G[52] = in[21] & in2[21];
    assign P[52] = in[21] ^ in2[21];
    assign G[53] = in[20] & in2[20];
    assign P[53] = in[20] ^ in2[20];
    assign G[54] = in[19] & in2[19];
    assign P[54] = in[19] ^ in2[19];
    assign G[55] = in[18] & in2[18];
    assign P[55] = in[18] ^ in2[18];
    assign G[56] = in[17] & in2[17];
    assign P[56] = in[17] ^ in2[17];
    assign G[57] = in[16] & in2[16];
    assign P[57] = in[16] ^ in2[16];
    assign G[58] = in[15] & in2[15];
    assign P[58] = in[15] ^ in2[15];
    assign G[59] = in[14] & in2[14];
    assign P[59] = in[14] ^ in2[14];
    assign G[60] = in[13] & in2[13];
    assign P[60] = in[13] ^ in2[13];
    assign G[61] = in[12] & in2[12];
    assign P[61] = in[12] ^ in2[12];
    assign G[62] = in[11] & in2[11];
    assign P[62] = in[11] ^ in2[11];
    assign G[63] = in[10] & in2[10];
    assign P[63] = in[10] ^ in2[10];
    assign G[64] = in[9] & in2[9];
    assign P[64] = in[9] ^ in2[9];
    assign G[65] = in[8] & in2[8];
    assign P[65] = in[8] ^ in2[8];
    assign G[66] = in[7] & in2[7];
    assign P[66] = in[7] ^ in2[7];
    assign G[67] = in[6] & in2[6];
    assign P[67] = in[6] ^ in2[6];
    assign G[68] = in[5] & in2[5];
    assign P[68] = in[5] ^ in2[5];
    assign G[69] = in[4] & in2[4];
    assign P[69] = in[4] ^ in2[4];
    assign G[70] = in[3] & in2[3];
    assign P[70] = in[3] ^ in2[3];
    assign G[71] = in[2] & in2[2];
    assign P[71] = in[2] ^ in2[2];
    assign G[72] = in[1] & in2[1];
    assign P[72] = in[1] ^ in2[1];
    assign G[73] = in[0] & in2[0];
    assign P[73] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign C[73] = G[72] | (P[72] & C[72]);
    assign cout = G[73] | (P[73] & C[73]);
    assign sum = P ^ C;
endmodule

module CLA73(output [72:0] sum, output cout, input [72:0] in1, input [72:0] in2;

    wire[72:0] G;
    wire[72:0] C;
    wire[72:0] P;

    assign G[0] = in[72] & in2[72];
    assign P[0] = in[72] ^ in2[72];
    assign G[1] = in[71] & in2[71];
    assign P[1] = in[71] ^ in2[71];
    assign G[2] = in[70] & in2[70];
    assign P[2] = in[70] ^ in2[70];
    assign G[3] = in[69] & in2[69];
    assign P[3] = in[69] ^ in2[69];
    assign G[4] = in[68] & in2[68];
    assign P[4] = in[68] ^ in2[68];
    assign G[5] = in[67] & in2[67];
    assign P[5] = in[67] ^ in2[67];
    assign G[6] = in[66] & in2[66];
    assign P[6] = in[66] ^ in2[66];
    assign G[7] = in[65] & in2[65];
    assign P[7] = in[65] ^ in2[65];
    assign G[8] = in[64] & in2[64];
    assign P[8] = in[64] ^ in2[64];
    assign G[9] = in[63] & in2[63];
    assign P[9] = in[63] ^ in2[63];
    assign G[10] = in[62] & in2[62];
    assign P[10] = in[62] ^ in2[62];
    assign G[11] = in[61] & in2[61];
    assign P[11] = in[61] ^ in2[61];
    assign G[12] = in[60] & in2[60];
    assign P[12] = in[60] ^ in2[60];
    assign G[13] = in[59] & in2[59];
    assign P[13] = in[59] ^ in2[59];
    assign G[14] = in[58] & in2[58];
    assign P[14] = in[58] ^ in2[58];
    assign G[15] = in[57] & in2[57];
    assign P[15] = in[57] ^ in2[57];
    assign G[16] = in[56] & in2[56];
    assign P[16] = in[56] ^ in2[56];
    assign G[17] = in[55] & in2[55];
    assign P[17] = in[55] ^ in2[55];
    assign G[18] = in[54] & in2[54];
    assign P[18] = in[54] ^ in2[54];
    assign G[19] = in[53] & in2[53];
    assign P[19] = in[53] ^ in2[53];
    assign G[20] = in[52] & in2[52];
    assign P[20] = in[52] ^ in2[52];
    assign G[21] = in[51] & in2[51];
    assign P[21] = in[51] ^ in2[51];
    assign G[22] = in[50] & in2[50];
    assign P[22] = in[50] ^ in2[50];
    assign G[23] = in[49] & in2[49];
    assign P[23] = in[49] ^ in2[49];
    assign G[24] = in[48] & in2[48];
    assign P[24] = in[48] ^ in2[48];
    assign G[25] = in[47] & in2[47];
    assign P[25] = in[47] ^ in2[47];
    assign G[26] = in[46] & in2[46];
    assign P[26] = in[46] ^ in2[46];
    assign G[27] = in[45] & in2[45];
    assign P[27] = in[45] ^ in2[45];
    assign G[28] = in[44] & in2[44];
    assign P[28] = in[44] ^ in2[44];
    assign G[29] = in[43] & in2[43];
    assign P[29] = in[43] ^ in2[43];
    assign G[30] = in[42] & in2[42];
    assign P[30] = in[42] ^ in2[42];
    assign G[31] = in[41] & in2[41];
    assign P[31] = in[41] ^ in2[41];
    assign G[32] = in[40] & in2[40];
    assign P[32] = in[40] ^ in2[40];
    assign G[33] = in[39] & in2[39];
    assign P[33] = in[39] ^ in2[39];
    assign G[34] = in[38] & in2[38];
    assign P[34] = in[38] ^ in2[38];
    assign G[35] = in[37] & in2[37];
    assign P[35] = in[37] ^ in2[37];
    assign G[36] = in[36] & in2[36];
    assign P[36] = in[36] ^ in2[36];
    assign G[37] = in[35] & in2[35];
    assign P[37] = in[35] ^ in2[35];
    assign G[38] = in[34] & in2[34];
    assign P[38] = in[34] ^ in2[34];
    assign G[39] = in[33] & in2[33];
    assign P[39] = in[33] ^ in2[33];
    assign G[40] = in[32] & in2[32];
    assign P[40] = in[32] ^ in2[32];
    assign G[41] = in[31] & in2[31];
    assign P[41] = in[31] ^ in2[31];
    assign G[42] = in[30] & in2[30];
    assign P[42] = in[30] ^ in2[30];
    assign G[43] = in[29] & in2[29];
    assign P[43] = in[29] ^ in2[29];
    assign G[44] = in[28] & in2[28];
    assign P[44] = in[28] ^ in2[28];
    assign G[45] = in[27] & in2[27];
    assign P[45] = in[27] ^ in2[27];
    assign G[46] = in[26] & in2[26];
    assign P[46] = in[26] ^ in2[26];
    assign G[47] = in[25] & in2[25];
    assign P[47] = in[25] ^ in2[25];
    assign G[48] = in[24] & in2[24];
    assign P[48] = in[24] ^ in2[24];
    assign G[49] = in[23] & in2[23];
    assign P[49] = in[23] ^ in2[23];
    assign G[50] = in[22] & in2[22];
    assign P[50] = in[22] ^ in2[22];
    assign G[51] = in[21] & in2[21];
    assign P[51] = in[21] ^ in2[21];
    assign G[52] = in[20] & in2[20];
    assign P[52] = in[20] ^ in2[20];
    assign G[53] = in[19] & in2[19];
    assign P[53] = in[19] ^ in2[19];
    assign G[54] = in[18] & in2[18];
    assign P[54] = in[18] ^ in2[18];
    assign G[55] = in[17] & in2[17];
    assign P[55] = in[17] ^ in2[17];
    assign G[56] = in[16] & in2[16];
    assign P[56] = in[16] ^ in2[16];
    assign G[57] = in[15] & in2[15];
    assign P[57] = in[15] ^ in2[15];
    assign G[58] = in[14] & in2[14];
    assign P[58] = in[14] ^ in2[14];
    assign G[59] = in[13] & in2[13];
    assign P[59] = in[13] ^ in2[13];
    assign G[60] = in[12] & in2[12];
    assign P[60] = in[12] ^ in2[12];
    assign G[61] = in[11] & in2[11];
    assign P[61] = in[11] ^ in2[11];
    assign G[62] = in[10] & in2[10];
    assign P[62] = in[10] ^ in2[10];
    assign G[63] = in[9] & in2[9];
    assign P[63] = in[9] ^ in2[9];
    assign G[64] = in[8] & in2[8];
    assign P[64] = in[8] ^ in2[8];
    assign G[65] = in[7] & in2[7];
    assign P[65] = in[7] ^ in2[7];
    assign G[66] = in[6] & in2[6];
    assign P[66] = in[6] ^ in2[6];
    assign G[67] = in[5] & in2[5];
    assign P[67] = in[5] ^ in2[5];
    assign G[68] = in[4] & in2[4];
    assign P[68] = in[4] ^ in2[4];
    assign G[69] = in[3] & in2[3];
    assign P[69] = in[3] ^ in2[3];
    assign G[70] = in[2] & in2[2];
    assign P[70] = in[2] ^ in2[2];
    assign G[71] = in[1] & in2[1];
    assign P[71] = in[1] ^ in2[1];
    assign G[72] = in[0] & in2[0];
    assign P[72] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign C[72] = G[71] | (P[71] & C[71]);
    assign cout = G[72] | (P[72] & C[72]);
    assign sum = P ^ C;
endmodule

module CLA72(output [71:0] sum, output cout, input [71:0] in1, input [71:0] in2;

    wire[71:0] G;
    wire[71:0] C;
    wire[71:0] P;

    assign G[0] = in[71] & in2[71];
    assign P[0] = in[71] ^ in2[71];
    assign G[1] = in[70] & in2[70];
    assign P[1] = in[70] ^ in2[70];
    assign G[2] = in[69] & in2[69];
    assign P[2] = in[69] ^ in2[69];
    assign G[3] = in[68] & in2[68];
    assign P[3] = in[68] ^ in2[68];
    assign G[4] = in[67] & in2[67];
    assign P[4] = in[67] ^ in2[67];
    assign G[5] = in[66] & in2[66];
    assign P[5] = in[66] ^ in2[66];
    assign G[6] = in[65] & in2[65];
    assign P[6] = in[65] ^ in2[65];
    assign G[7] = in[64] & in2[64];
    assign P[7] = in[64] ^ in2[64];
    assign G[8] = in[63] & in2[63];
    assign P[8] = in[63] ^ in2[63];
    assign G[9] = in[62] & in2[62];
    assign P[9] = in[62] ^ in2[62];
    assign G[10] = in[61] & in2[61];
    assign P[10] = in[61] ^ in2[61];
    assign G[11] = in[60] & in2[60];
    assign P[11] = in[60] ^ in2[60];
    assign G[12] = in[59] & in2[59];
    assign P[12] = in[59] ^ in2[59];
    assign G[13] = in[58] & in2[58];
    assign P[13] = in[58] ^ in2[58];
    assign G[14] = in[57] & in2[57];
    assign P[14] = in[57] ^ in2[57];
    assign G[15] = in[56] & in2[56];
    assign P[15] = in[56] ^ in2[56];
    assign G[16] = in[55] & in2[55];
    assign P[16] = in[55] ^ in2[55];
    assign G[17] = in[54] & in2[54];
    assign P[17] = in[54] ^ in2[54];
    assign G[18] = in[53] & in2[53];
    assign P[18] = in[53] ^ in2[53];
    assign G[19] = in[52] & in2[52];
    assign P[19] = in[52] ^ in2[52];
    assign G[20] = in[51] & in2[51];
    assign P[20] = in[51] ^ in2[51];
    assign G[21] = in[50] & in2[50];
    assign P[21] = in[50] ^ in2[50];
    assign G[22] = in[49] & in2[49];
    assign P[22] = in[49] ^ in2[49];
    assign G[23] = in[48] & in2[48];
    assign P[23] = in[48] ^ in2[48];
    assign G[24] = in[47] & in2[47];
    assign P[24] = in[47] ^ in2[47];
    assign G[25] = in[46] & in2[46];
    assign P[25] = in[46] ^ in2[46];
    assign G[26] = in[45] & in2[45];
    assign P[26] = in[45] ^ in2[45];
    assign G[27] = in[44] & in2[44];
    assign P[27] = in[44] ^ in2[44];
    assign G[28] = in[43] & in2[43];
    assign P[28] = in[43] ^ in2[43];
    assign G[29] = in[42] & in2[42];
    assign P[29] = in[42] ^ in2[42];
    assign G[30] = in[41] & in2[41];
    assign P[30] = in[41] ^ in2[41];
    assign G[31] = in[40] & in2[40];
    assign P[31] = in[40] ^ in2[40];
    assign G[32] = in[39] & in2[39];
    assign P[32] = in[39] ^ in2[39];
    assign G[33] = in[38] & in2[38];
    assign P[33] = in[38] ^ in2[38];
    assign G[34] = in[37] & in2[37];
    assign P[34] = in[37] ^ in2[37];
    assign G[35] = in[36] & in2[36];
    assign P[35] = in[36] ^ in2[36];
    assign G[36] = in[35] & in2[35];
    assign P[36] = in[35] ^ in2[35];
    assign G[37] = in[34] & in2[34];
    assign P[37] = in[34] ^ in2[34];
    assign G[38] = in[33] & in2[33];
    assign P[38] = in[33] ^ in2[33];
    assign G[39] = in[32] & in2[32];
    assign P[39] = in[32] ^ in2[32];
    assign G[40] = in[31] & in2[31];
    assign P[40] = in[31] ^ in2[31];
    assign G[41] = in[30] & in2[30];
    assign P[41] = in[30] ^ in2[30];
    assign G[42] = in[29] & in2[29];
    assign P[42] = in[29] ^ in2[29];
    assign G[43] = in[28] & in2[28];
    assign P[43] = in[28] ^ in2[28];
    assign G[44] = in[27] & in2[27];
    assign P[44] = in[27] ^ in2[27];
    assign G[45] = in[26] & in2[26];
    assign P[45] = in[26] ^ in2[26];
    assign G[46] = in[25] & in2[25];
    assign P[46] = in[25] ^ in2[25];
    assign G[47] = in[24] & in2[24];
    assign P[47] = in[24] ^ in2[24];
    assign G[48] = in[23] & in2[23];
    assign P[48] = in[23] ^ in2[23];
    assign G[49] = in[22] & in2[22];
    assign P[49] = in[22] ^ in2[22];
    assign G[50] = in[21] & in2[21];
    assign P[50] = in[21] ^ in2[21];
    assign G[51] = in[20] & in2[20];
    assign P[51] = in[20] ^ in2[20];
    assign G[52] = in[19] & in2[19];
    assign P[52] = in[19] ^ in2[19];
    assign G[53] = in[18] & in2[18];
    assign P[53] = in[18] ^ in2[18];
    assign G[54] = in[17] & in2[17];
    assign P[54] = in[17] ^ in2[17];
    assign G[55] = in[16] & in2[16];
    assign P[55] = in[16] ^ in2[16];
    assign G[56] = in[15] & in2[15];
    assign P[56] = in[15] ^ in2[15];
    assign G[57] = in[14] & in2[14];
    assign P[57] = in[14] ^ in2[14];
    assign G[58] = in[13] & in2[13];
    assign P[58] = in[13] ^ in2[13];
    assign G[59] = in[12] & in2[12];
    assign P[59] = in[12] ^ in2[12];
    assign G[60] = in[11] & in2[11];
    assign P[60] = in[11] ^ in2[11];
    assign G[61] = in[10] & in2[10];
    assign P[61] = in[10] ^ in2[10];
    assign G[62] = in[9] & in2[9];
    assign P[62] = in[9] ^ in2[9];
    assign G[63] = in[8] & in2[8];
    assign P[63] = in[8] ^ in2[8];
    assign G[64] = in[7] & in2[7];
    assign P[64] = in[7] ^ in2[7];
    assign G[65] = in[6] & in2[6];
    assign P[65] = in[6] ^ in2[6];
    assign G[66] = in[5] & in2[5];
    assign P[66] = in[5] ^ in2[5];
    assign G[67] = in[4] & in2[4];
    assign P[67] = in[4] ^ in2[4];
    assign G[68] = in[3] & in2[3];
    assign P[68] = in[3] ^ in2[3];
    assign G[69] = in[2] & in2[2];
    assign P[69] = in[2] ^ in2[2];
    assign G[70] = in[1] & in2[1];
    assign P[70] = in[1] ^ in2[1];
    assign G[71] = in[0] & in2[0];
    assign P[71] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign C[71] = G[70] | (P[70] & C[70]);
    assign cout = G[71] | (P[71] & C[71]);
    assign sum = P ^ C;
endmodule

module CLA71(output [70:0] sum, output cout, input [70:0] in1, input [70:0] in2;

    wire[70:0] G;
    wire[70:0] C;
    wire[70:0] P;

    assign G[0] = in[70] & in2[70];
    assign P[0] = in[70] ^ in2[70];
    assign G[1] = in[69] & in2[69];
    assign P[1] = in[69] ^ in2[69];
    assign G[2] = in[68] & in2[68];
    assign P[2] = in[68] ^ in2[68];
    assign G[3] = in[67] & in2[67];
    assign P[3] = in[67] ^ in2[67];
    assign G[4] = in[66] & in2[66];
    assign P[4] = in[66] ^ in2[66];
    assign G[5] = in[65] & in2[65];
    assign P[5] = in[65] ^ in2[65];
    assign G[6] = in[64] & in2[64];
    assign P[6] = in[64] ^ in2[64];
    assign G[7] = in[63] & in2[63];
    assign P[7] = in[63] ^ in2[63];
    assign G[8] = in[62] & in2[62];
    assign P[8] = in[62] ^ in2[62];
    assign G[9] = in[61] & in2[61];
    assign P[9] = in[61] ^ in2[61];
    assign G[10] = in[60] & in2[60];
    assign P[10] = in[60] ^ in2[60];
    assign G[11] = in[59] & in2[59];
    assign P[11] = in[59] ^ in2[59];
    assign G[12] = in[58] & in2[58];
    assign P[12] = in[58] ^ in2[58];
    assign G[13] = in[57] & in2[57];
    assign P[13] = in[57] ^ in2[57];
    assign G[14] = in[56] & in2[56];
    assign P[14] = in[56] ^ in2[56];
    assign G[15] = in[55] & in2[55];
    assign P[15] = in[55] ^ in2[55];
    assign G[16] = in[54] & in2[54];
    assign P[16] = in[54] ^ in2[54];
    assign G[17] = in[53] & in2[53];
    assign P[17] = in[53] ^ in2[53];
    assign G[18] = in[52] & in2[52];
    assign P[18] = in[52] ^ in2[52];
    assign G[19] = in[51] & in2[51];
    assign P[19] = in[51] ^ in2[51];
    assign G[20] = in[50] & in2[50];
    assign P[20] = in[50] ^ in2[50];
    assign G[21] = in[49] & in2[49];
    assign P[21] = in[49] ^ in2[49];
    assign G[22] = in[48] & in2[48];
    assign P[22] = in[48] ^ in2[48];
    assign G[23] = in[47] & in2[47];
    assign P[23] = in[47] ^ in2[47];
    assign G[24] = in[46] & in2[46];
    assign P[24] = in[46] ^ in2[46];
    assign G[25] = in[45] & in2[45];
    assign P[25] = in[45] ^ in2[45];
    assign G[26] = in[44] & in2[44];
    assign P[26] = in[44] ^ in2[44];
    assign G[27] = in[43] & in2[43];
    assign P[27] = in[43] ^ in2[43];
    assign G[28] = in[42] & in2[42];
    assign P[28] = in[42] ^ in2[42];
    assign G[29] = in[41] & in2[41];
    assign P[29] = in[41] ^ in2[41];
    assign G[30] = in[40] & in2[40];
    assign P[30] = in[40] ^ in2[40];
    assign G[31] = in[39] & in2[39];
    assign P[31] = in[39] ^ in2[39];
    assign G[32] = in[38] & in2[38];
    assign P[32] = in[38] ^ in2[38];
    assign G[33] = in[37] & in2[37];
    assign P[33] = in[37] ^ in2[37];
    assign G[34] = in[36] & in2[36];
    assign P[34] = in[36] ^ in2[36];
    assign G[35] = in[35] & in2[35];
    assign P[35] = in[35] ^ in2[35];
    assign G[36] = in[34] & in2[34];
    assign P[36] = in[34] ^ in2[34];
    assign G[37] = in[33] & in2[33];
    assign P[37] = in[33] ^ in2[33];
    assign G[38] = in[32] & in2[32];
    assign P[38] = in[32] ^ in2[32];
    assign G[39] = in[31] & in2[31];
    assign P[39] = in[31] ^ in2[31];
    assign G[40] = in[30] & in2[30];
    assign P[40] = in[30] ^ in2[30];
    assign G[41] = in[29] & in2[29];
    assign P[41] = in[29] ^ in2[29];
    assign G[42] = in[28] & in2[28];
    assign P[42] = in[28] ^ in2[28];
    assign G[43] = in[27] & in2[27];
    assign P[43] = in[27] ^ in2[27];
    assign G[44] = in[26] & in2[26];
    assign P[44] = in[26] ^ in2[26];
    assign G[45] = in[25] & in2[25];
    assign P[45] = in[25] ^ in2[25];
    assign G[46] = in[24] & in2[24];
    assign P[46] = in[24] ^ in2[24];
    assign G[47] = in[23] & in2[23];
    assign P[47] = in[23] ^ in2[23];
    assign G[48] = in[22] & in2[22];
    assign P[48] = in[22] ^ in2[22];
    assign G[49] = in[21] & in2[21];
    assign P[49] = in[21] ^ in2[21];
    assign G[50] = in[20] & in2[20];
    assign P[50] = in[20] ^ in2[20];
    assign G[51] = in[19] & in2[19];
    assign P[51] = in[19] ^ in2[19];
    assign G[52] = in[18] & in2[18];
    assign P[52] = in[18] ^ in2[18];
    assign G[53] = in[17] & in2[17];
    assign P[53] = in[17] ^ in2[17];
    assign G[54] = in[16] & in2[16];
    assign P[54] = in[16] ^ in2[16];
    assign G[55] = in[15] & in2[15];
    assign P[55] = in[15] ^ in2[15];
    assign G[56] = in[14] & in2[14];
    assign P[56] = in[14] ^ in2[14];
    assign G[57] = in[13] & in2[13];
    assign P[57] = in[13] ^ in2[13];
    assign G[58] = in[12] & in2[12];
    assign P[58] = in[12] ^ in2[12];
    assign G[59] = in[11] & in2[11];
    assign P[59] = in[11] ^ in2[11];
    assign G[60] = in[10] & in2[10];
    assign P[60] = in[10] ^ in2[10];
    assign G[61] = in[9] & in2[9];
    assign P[61] = in[9] ^ in2[9];
    assign G[62] = in[8] & in2[8];
    assign P[62] = in[8] ^ in2[8];
    assign G[63] = in[7] & in2[7];
    assign P[63] = in[7] ^ in2[7];
    assign G[64] = in[6] & in2[6];
    assign P[64] = in[6] ^ in2[6];
    assign G[65] = in[5] & in2[5];
    assign P[65] = in[5] ^ in2[5];
    assign G[66] = in[4] & in2[4];
    assign P[66] = in[4] ^ in2[4];
    assign G[67] = in[3] & in2[3];
    assign P[67] = in[3] ^ in2[3];
    assign G[68] = in[2] & in2[2];
    assign P[68] = in[2] ^ in2[2];
    assign G[69] = in[1] & in2[1];
    assign P[69] = in[1] ^ in2[1];
    assign G[70] = in[0] & in2[0];
    assign P[70] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign C[70] = G[69] | (P[69] & C[69]);
    assign cout = G[70] | (P[70] & C[70]);
    assign sum = P ^ C;
endmodule

module CLA70(output [69:0] sum, output cout, input [69:0] in1, input [69:0] in2;

    wire[69:0] G;
    wire[69:0] C;
    wire[69:0] P;

    assign G[0] = in[69] & in2[69];
    assign P[0] = in[69] ^ in2[69];
    assign G[1] = in[68] & in2[68];
    assign P[1] = in[68] ^ in2[68];
    assign G[2] = in[67] & in2[67];
    assign P[2] = in[67] ^ in2[67];
    assign G[3] = in[66] & in2[66];
    assign P[3] = in[66] ^ in2[66];
    assign G[4] = in[65] & in2[65];
    assign P[4] = in[65] ^ in2[65];
    assign G[5] = in[64] & in2[64];
    assign P[5] = in[64] ^ in2[64];
    assign G[6] = in[63] & in2[63];
    assign P[6] = in[63] ^ in2[63];
    assign G[7] = in[62] & in2[62];
    assign P[7] = in[62] ^ in2[62];
    assign G[8] = in[61] & in2[61];
    assign P[8] = in[61] ^ in2[61];
    assign G[9] = in[60] & in2[60];
    assign P[9] = in[60] ^ in2[60];
    assign G[10] = in[59] & in2[59];
    assign P[10] = in[59] ^ in2[59];
    assign G[11] = in[58] & in2[58];
    assign P[11] = in[58] ^ in2[58];
    assign G[12] = in[57] & in2[57];
    assign P[12] = in[57] ^ in2[57];
    assign G[13] = in[56] & in2[56];
    assign P[13] = in[56] ^ in2[56];
    assign G[14] = in[55] & in2[55];
    assign P[14] = in[55] ^ in2[55];
    assign G[15] = in[54] & in2[54];
    assign P[15] = in[54] ^ in2[54];
    assign G[16] = in[53] & in2[53];
    assign P[16] = in[53] ^ in2[53];
    assign G[17] = in[52] & in2[52];
    assign P[17] = in[52] ^ in2[52];
    assign G[18] = in[51] & in2[51];
    assign P[18] = in[51] ^ in2[51];
    assign G[19] = in[50] & in2[50];
    assign P[19] = in[50] ^ in2[50];
    assign G[20] = in[49] & in2[49];
    assign P[20] = in[49] ^ in2[49];
    assign G[21] = in[48] & in2[48];
    assign P[21] = in[48] ^ in2[48];
    assign G[22] = in[47] & in2[47];
    assign P[22] = in[47] ^ in2[47];
    assign G[23] = in[46] & in2[46];
    assign P[23] = in[46] ^ in2[46];
    assign G[24] = in[45] & in2[45];
    assign P[24] = in[45] ^ in2[45];
    assign G[25] = in[44] & in2[44];
    assign P[25] = in[44] ^ in2[44];
    assign G[26] = in[43] & in2[43];
    assign P[26] = in[43] ^ in2[43];
    assign G[27] = in[42] & in2[42];
    assign P[27] = in[42] ^ in2[42];
    assign G[28] = in[41] & in2[41];
    assign P[28] = in[41] ^ in2[41];
    assign G[29] = in[40] & in2[40];
    assign P[29] = in[40] ^ in2[40];
    assign G[30] = in[39] & in2[39];
    assign P[30] = in[39] ^ in2[39];
    assign G[31] = in[38] & in2[38];
    assign P[31] = in[38] ^ in2[38];
    assign G[32] = in[37] & in2[37];
    assign P[32] = in[37] ^ in2[37];
    assign G[33] = in[36] & in2[36];
    assign P[33] = in[36] ^ in2[36];
    assign G[34] = in[35] & in2[35];
    assign P[34] = in[35] ^ in2[35];
    assign G[35] = in[34] & in2[34];
    assign P[35] = in[34] ^ in2[34];
    assign G[36] = in[33] & in2[33];
    assign P[36] = in[33] ^ in2[33];
    assign G[37] = in[32] & in2[32];
    assign P[37] = in[32] ^ in2[32];
    assign G[38] = in[31] & in2[31];
    assign P[38] = in[31] ^ in2[31];
    assign G[39] = in[30] & in2[30];
    assign P[39] = in[30] ^ in2[30];
    assign G[40] = in[29] & in2[29];
    assign P[40] = in[29] ^ in2[29];
    assign G[41] = in[28] & in2[28];
    assign P[41] = in[28] ^ in2[28];
    assign G[42] = in[27] & in2[27];
    assign P[42] = in[27] ^ in2[27];
    assign G[43] = in[26] & in2[26];
    assign P[43] = in[26] ^ in2[26];
    assign G[44] = in[25] & in2[25];
    assign P[44] = in[25] ^ in2[25];
    assign G[45] = in[24] & in2[24];
    assign P[45] = in[24] ^ in2[24];
    assign G[46] = in[23] & in2[23];
    assign P[46] = in[23] ^ in2[23];
    assign G[47] = in[22] & in2[22];
    assign P[47] = in[22] ^ in2[22];
    assign G[48] = in[21] & in2[21];
    assign P[48] = in[21] ^ in2[21];
    assign G[49] = in[20] & in2[20];
    assign P[49] = in[20] ^ in2[20];
    assign G[50] = in[19] & in2[19];
    assign P[50] = in[19] ^ in2[19];
    assign G[51] = in[18] & in2[18];
    assign P[51] = in[18] ^ in2[18];
    assign G[52] = in[17] & in2[17];
    assign P[52] = in[17] ^ in2[17];
    assign G[53] = in[16] & in2[16];
    assign P[53] = in[16] ^ in2[16];
    assign G[54] = in[15] & in2[15];
    assign P[54] = in[15] ^ in2[15];
    assign G[55] = in[14] & in2[14];
    assign P[55] = in[14] ^ in2[14];
    assign G[56] = in[13] & in2[13];
    assign P[56] = in[13] ^ in2[13];
    assign G[57] = in[12] & in2[12];
    assign P[57] = in[12] ^ in2[12];
    assign G[58] = in[11] & in2[11];
    assign P[58] = in[11] ^ in2[11];
    assign G[59] = in[10] & in2[10];
    assign P[59] = in[10] ^ in2[10];
    assign G[60] = in[9] & in2[9];
    assign P[60] = in[9] ^ in2[9];
    assign G[61] = in[8] & in2[8];
    assign P[61] = in[8] ^ in2[8];
    assign G[62] = in[7] & in2[7];
    assign P[62] = in[7] ^ in2[7];
    assign G[63] = in[6] & in2[6];
    assign P[63] = in[6] ^ in2[6];
    assign G[64] = in[5] & in2[5];
    assign P[64] = in[5] ^ in2[5];
    assign G[65] = in[4] & in2[4];
    assign P[65] = in[4] ^ in2[4];
    assign G[66] = in[3] & in2[3];
    assign P[66] = in[3] ^ in2[3];
    assign G[67] = in[2] & in2[2];
    assign P[67] = in[2] ^ in2[2];
    assign G[68] = in[1] & in2[1];
    assign P[68] = in[1] ^ in2[1];
    assign G[69] = in[0] & in2[0];
    assign P[69] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign C[69] = G[68] | (P[68] & C[68]);
    assign cout = G[69] | (P[69] & C[69]);
    assign sum = P ^ C;
endmodule

module CLA69(output [68:0] sum, output cout, input [68:0] in1, input [68:0] in2;

    wire[68:0] G;
    wire[68:0] C;
    wire[68:0] P;

    assign G[0] = in[68] & in2[68];
    assign P[0] = in[68] ^ in2[68];
    assign G[1] = in[67] & in2[67];
    assign P[1] = in[67] ^ in2[67];
    assign G[2] = in[66] & in2[66];
    assign P[2] = in[66] ^ in2[66];
    assign G[3] = in[65] & in2[65];
    assign P[3] = in[65] ^ in2[65];
    assign G[4] = in[64] & in2[64];
    assign P[4] = in[64] ^ in2[64];
    assign G[5] = in[63] & in2[63];
    assign P[5] = in[63] ^ in2[63];
    assign G[6] = in[62] & in2[62];
    assign P[6] = in[62] ^ in2[62];
    assign G[7] = in[61] & in2[61];
    assign P[7] = in[61] ^ in2[61];
    assign G[8] = in[60] & in2[60];
    assign P[8] = in[60] ^ in2[60];
    assign G[9] = in[59] & in2[59];
    assign P[9] = in[59] ^ in2[59];
    assign G[10] = in[58] & in2[58];
    assign P[10] = in[58] ^ in2[58];
    assign G[11] = in[57] & in2[57];
    assign P[11] = in[57] ^ in2[57];
    assign G[12] = in[56] & in2[56];
    assign P[12] = in[56] ^ in2[56];
    assign G[13] = in[55] & in2[55];
    assign P[13] = in[55] ^ in2[55];
    assign G[14] = in[54] & in2[54];
    assign P[14] = in[54] ^ in2[54];
    assign G[15] = in[53] & in2[53];
    assign P[15] = in[53] ^ in2[53];
    assign G[16] = in[52] & in2[52];
    assign P[16] = in[52] ^ in2[52];
    assign G[17] = in[51] & in2[51];
    assign P[17] = in[51] ^ in2[51];
    assign G[18] = in[50] & in2[50];
    assign P[18] = in[50] ^ in2[50];
    assign G[19] = in[49] & in2[49];
    assign P[19] = in[49] ^ in2[49];
    assign G[20] = in[48] & in2[48];
    assign P[20] = in[48] ^ in2[48];
    assign G[21] = in[47] & in2[47];
    assign P[21] = in[47] ^ in2[47];
    assign G[22] = in[46] & in2[46];
    assign P[22] = in[46] ^ in2[46];
    assign G[23] = in[45] & in2[45];
    assign P[23] = in[45] ^ in2[45];
    assign G[24] = in[44] & in2[44];
    assign P[24] = in[44] ^ in2[44];
    assign G[25] = in[43] & in2[43];
    assign P[25] = in[43] ^ in2[43];
    assign G[26] = in[42] & in2[42];
    assign P[26] = in[42] ^ in2[42];
    assign G[27] = in[41] & in2[41];
    assign P[27] = in[41] ^ in2[41];
    assign G[28] = in[40] & in2[40];
    assign P[28] = in[40] ^ in2[40];
    assign G[29] = in[39] & in2[39];
    assign P[29] = in[39] ^ in2[39];
    assign G[30] = in[38] & in2[38];
    assign P[30] = in[38] ^ in2[38];
    assign G[31] = in[37] & in2[37];
    assign P[31] = in[37] ^ in2[37];
    assign G[32] = in[36] & in2[36];
    assign P[32] = in[36] ^ in2[36];
    assign G[33] = in[35] & in2[35];
    assign P[33] = in[35] ^ in2[35];
    assign G[34] = in[34] & in2[34];
    assign P[34] = in[34] ^ in2[34];
    assign G[35] = in[33] & in2[33];
    assign P[35] = in[33] ^ in2[33];
    assign G[36] = in[32] & in2[32];
    assign P[36] = in[32] ^ in2[32];
    assign G[37] = in[31] & in2[31];
    assign P[37] = in[31] ^ in2[31];
    assign G[38] = in[30] & in2[30];
    assign P[38] = in[30] ^ in2[30];
    assign G[39] = in[29] & in2[29];
    assign P[39] = in[29] ^ in2[29];
    assign G[40] = in[28] & in2[28];
    assign P[40] = in[28] ^ in2[28];
    assign G[41] = in[27] & in2[27];
    assign P[41] = in[27] ^ in2[27];
    assign G[42] = in[26] & in2[26];
    assign P[42] = in[26] ^ in2[26];
    assign G[43] = in[25] & in2[25];
    assign P[43] = in[25] ^ in2[25];
    assign G[44] = in[24] & in2[24];
    assign P[44] = in[24] ^ in2[24];
    assign G[45] = in[23] & in2[23];
    assign P[45] = in[23] ^ in2[23];
    assign G[46] = in[22] & in2[22];
    assign P[46] = in[22] ^ in2[22];
    assign G[47] = in[21] & in2[21];
    assign P[47] = in[21] ^ in2[21];
    assign G[48] = in[20] & in2[20];
    assign P[48] = in[20] ^ in2[20];
    assign G[49] = in[19] & in2[19];
    assign P[49] = in[19] ^ in2[19];
    assign G[50] = in[18] & in2[18];
    assign P[50] = in[18] ^ in2[18];
    assign G[51] = in[17] & in2[17];
    assign P[51] = in[17] ^ in2[17];
    assign G[52] = in[16] & in2[16];
    assign P[52] = in[16] ^ in2[16];
    assign G[53] = in[15] & in2[15];
    assign P[53] = in[15] ^ in2[15];
    assign G[54] = in[14] & in2[14];
    assign P[54] = in[14] ^ in2[14];
    assign G[55] = in[13] & in2[13];
    assign P[55] = in[13] ^ in2[13];
    assign G[56] = in[12] & in2[12];
    assign P[56] = in[12] ^ in2[12];
    assign G[57] = in[11] & in2[11];
    assign P[57] = in[11] ^ in2[11];
    assign G[58] = in[10] & in2[10];
    assign P[58] = in[10] ^ in2[10];
    assign G[59] = in[9] & in2[9];
    assign P[59] = in[9] ^ in2[9];
    assign G[60] = in[8] & in2[8];
    assign P[60] = in[8] ^ in2[8];
    assign G[61] = in[7] & in2[7];
    assign P[61] = in[7] ^ in2[7];
    assign G[62] = in[6] & in2[6];
    assign P[62] = in[6] ^ in2[6];
    assign G[63] = in[5] & in2[5];
    assign P[63] = in[5] ^ in2[5];
    assign G[64] = in[4] & in2[4];
    assign P[64] = in[4] ^ in2[4];
    assign G[65] = in[3] & in2[3];
    assign P[65] = in[3] ^ in2[3];
    assign G[66] = in[2] & in2[2];
    assign P[66] = in[2] ^ in2[2];
    assign G[67] = in[1] & in2[1];
    assign P[67] = in[1] ^ in2[1];
    assign G[68] = in[0] & in2[0];
    assign P[68] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign C[68] = G[67] | (P[67] & C[67]);
    assign cout = G[68] | (P[68] & C[68]);
    assign sum = P ^ C;
endmodule

module CLA68(output [67:0] sum, output cout, input [67:0] in1, input [67:0] in2;

    wire[67:0] G;
    wire[67:0] C;
    wire[67:0] P;

    assign G[0] = in[67] & in2[67];
    assign P[0] = in[67] ^ in2[67];
    assign G[1] = in[66] & in2[66];
    assign P[1] = in[66] ^ in2[66];
    assign G[2] = in[65] & in2[65];
    assign P[2] = in[65] ^ in2[65];
    assign G[3] = in[64] & in2[64];
    assign P[3] = in[64] ^ in2[64];
    assign G[4] = in[63] & in2[63];
    assign P[4] = in[63] ^ in2[63];
    assign G[5] = in[62] & in2[62];
    assign P[5] = in[62] ^ in2[62];
    assign G[6] = in[61] & in2[61];
    assign P[6] = in[61] ^ in2[61];
    assign G[7] = in[60] & in2[60];
    assign P[7] = in[60] ^ in2[60];
    assign G[8] = in[59] & in2[59];
    assign P[8] = in[59] ^ in2[59];
    assign G[9] = in[58] & in2[58];
    assign P[9] = in[58] ^ in2[58];
    assign G[10] = in[57] & in2[57];
    assign P[10] = in[57] ^ in2[57];
    assign G[11] = in[56] & in2[56];
    assign P[11] = in[56] ^ in2[56];
    assign G[12] = in[55] & in2[55];
    assign P[12] = in[55] ^ in2[55];
    assign G[13] = in[54] & in2[54];
    assign P[13] = in[54] ^ in2[54];
    assign G[14] = in[53] & in2[53];
    assign P[14] = in[53] ^ in2[53];
    assign G[15] = in[52] & in2[52];
    assign P[15] = in[52] ^ in2[52];
    assign G[16] = in[51] & in2[51];
    assign P[16] = in[51] ^ in2[51];
    assign G[17] = in[50] & in2[50];
    assign P[17] = in[50] ^ in2[50];
    assign G[18] = in[49] & in2[49];
    assign P[18] = in[49] ^ in2[49];
    assign G[19] = in[48] & in2[48];
    assign P[19] = in[48] ^ in2[48];
    assign G[20] = in[47] & in2[47];
    assign P[20] = in[47] ^ in2[47];
    assign G[21] = in[46] & in2[46];
    assign P[21] = in[46] ^ in2[46];
    assign G[22] = in[45] & in2[45];
    assign P[22] = in[45] ^ in2[45];
    assign G[23] = in[44] & in2[44];
    assign P[23] = in[44] ^ in2[44];
    assign G[24] = in[43] & in2[43];
    assign P[24] = in[43] ^ in2[43];
    assign G[25] = in[42] & in2[42];
    assign P[25] = in[42] ^ in2[42];
    assign G[26] = in[41] & in2[41];
    assign P[26] = in[41] ^ in2[41];
    assign G[27] = in[40] & in2[40];
    assign P[27] = in[40] ^ in2[40];
    assign G[28] = in[39] & in2[39];
    assign P[28] = in[39] ^ in2[39];
    assign G[29] = in[38] & in2[38];
    assign P[29] = in[38] ^ in2[38];
    assign G[30] = in[37] & in2[37];
    assign P[30] = in[37] ^ in2[37];
    assign G[31] = in[36] & in2[36];
    assign P[31] = in[36] ^ in2[36];
    assign G[32] = in[35] & in2[35];
    assign P[32] = in[35] ^ in2[35];
    assign G[33] = in[34] & in2[34];
    assign P[33] = in[34] ^ in2[34];
    assign G[34] = in[33] & in2[33];
    assign P[34] = in[33] ^ in2[33];
    assign G[35] = in[32] & in2[32];
    assign P[35] = in[32] ^ in2[32];
    assign G[36] = in[31] & in2[31];
    assign P[36] = in[31] ^ in2[31];
    assign G[37] = in[30] & in2[30];
    assign P[37] = in[30] ^ in2[30];
    assign G[38] = in[29] & in2[29];
    assign P[38] = in[29] ^ in2[29];
    assign G[39] = in[28] & in2[28];
    assign P[39] = in[28] ^ in2[28];
    assign G[40] = in[27] & in2[27];
    assign P[40] = in[27] ^ in2[27];
    assign G[41] = in[26] & in2[26];
    assign P[41] = in[26] ^ in2[26];
    assign G[42] = in[25] & in2[25];
    assign P[42] = in[25] ^ in2[25];
    assign G[43] = in[24] & in2[24];
    assign P[43] = in[24] ^ in2[24];
    assign G[44] = in[23] & in2[23];
    assign P[44] = in[23] ^ in2[23];
    assign G[45] = in[22] & in2[22];
    assign P[45] = in[22] ^ in2[22];
    assign G[46] = in[21] & in2[21];
    assign P[46] = in[21] ^ in2[21];
    assign G[47] = in[20] & in2[20];
    assign P[47] = in[20] ^ in2[20];
    assign G[48] = in[19] & in2[19];
    assign P[48] = in[19] ^ in2[19];
    assign G[49] = in[18] & in2[18];
    assign P[49] = in[18] ^ in2[18];
    assign G[50] = in[17] & in2[17];
    assign P[50] = in[17] ^ in2[17];
    assign G[51] = in[16] & in2[16];
    assign P[51] = in[16] ^ in2[16];
    assign G[52] = in[15] & in2[15];
    assign P[52] = in[15] ^ in2[15];
    assign G[53] = in[14] & in2[14];
    assign P[53] = in[14] ^ in2[14];
    assign G[54] = in[13] & in2[13];
    assign P[54] = in[13] ^ in2[13];
    assign G[55] = in[12] & in2[12];
    assign P[55] = in[12] ^ in2[12];
    assign G[56] = in[11] & in2[11];
    assign P[56] = in[11] ^ in2[11];
    assign G[57] = in[10] & in2[10];
    assign P[57] = in[10] ^ in2[10];
    assign G[58] = in[9] & in2[9];
    assign P[58] = in[9] ^ in2[9];
    assign G[59] = in[8] & in2[8];
    assign P[59] = in[8] ^ in2[8];
    assign G[60] = in[7] & in2[7];
    assign P[60] = in[7] ^ in2[7];
    assign G[61] = in[6] & in2[6];
    assign P[61] = in[6] ^ in2[6];
    assign G[62] = in[5] & in2[5];
    assign P[62] = in[5] ^ in2[5];
    assign G[63] = in[4] & in2[4];
    assign P[63] = in[4] ^ in2[4];
    assign G[64] = in[3] & in2[3];
    assign P[64] = in[3] ^ in2[3];
    assign G[65] = in[2] & in2[2];
    assign P[65] = in[2] ^ in2[2];
    assign G[66] = in[1] & in2[1];
    assign P[66] = in[1] ^ in2[1];
    assign G[67] = in[0] & in2[0];
    assign P[67] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign C[67] = G[66] | (P[66] & C[66]);
    assign cout = G[67] | (P[67] & C[67]);
    assign sum = P ^ C;
endmodule

module CLA67(output [66:0] sum, output cout, input [66:0] in1, input [66:0] in2;

    wire[66:0] G;
    wire[66:0] C;
    wire[66:0] P;

    assign G[0] = in[66] & in2[66];
    assign P[0] = in[66] ^ in2[66];
    assign G[1] = in[65] & in2[65];
    assign P[1] = in[65] ^ in2[65];
    assign G[2] = in[64] & in2[64];
    assign P[2] = in[64] ^ in2[64];
    assign G[3] = in[63] & in2[63];
    assign P[3] = in[63] ^ in2[63];
    assign G[4] = in[62] & in2[62];
    assign P[4] = in[62] ^ in2[62];
    assign G[5] = in[61] & in2[61];
    assign P[5] = in[61] ^ in2[61];
    assign G[6] = in[60] & in2[60];
    assign P[6] = in[60] ^ in2[60];
    assign G[7] = in[59] & in2[59];
    assign P[7] = in[59] ^ in2[59];
    assign G[8] = in[58] & in2[58];
    assign P[8] = in[58] ^ in2[58];
    assign G[9] = in[57] & in2[57];
    assign P[9] = in[57] ^ in2[57];
    assign G[10] = in[56] & in2[56];
    assign P[10] = in[56] ^ in2[56];
    assign G[11] = in[55] & in2[55];
    assign P[11] = in[55] ^ in2[55];
    assign G[12] = in[54] & in2[54];
    assign P[12] = in[54] ^ in2[54];
    assign G[13] = in[53] & in2[53];
    assign P[13] = in[53] ^ in2[53];
    assign G[14] = in[52] & in2[52];
    assign P[14] = in[52] ^ in2[52];
    assign G[15] = in[51] & in2[51];
    assign P[15] = in[51] ^ in2[51];
    assign G[16] = in[50] & in2[50];
    assign P[16] = in[50] ^ in2[50];
    assign G[17] = in[49] & in2[49];
    assign P[17] = in[49] ^ in2[49];
    assign G[18] = in[48] & in2[48];
    assign P[18] = in[48] ^ in2[48];
    assign G[19] = in[47] & in2[47];
    assign P[19] = in[47] ^ in2[47];
    assign G[20] = in[46] & in2[46];
    assign P[20] = in[46] ^ in2[46];
    assign G[21] = in[45] & in2[45];
    assign P[21] = in[45] ^ in2[45];
    assign G[22] = in[44] & in2[44];
    assign P[22] = in[44] ^ in2[44];
    assign G[23] = in[43] & in2[43];
    assign P[23] = in[43] ^ in2[43];
    assign G[24] = in[42] & in2[42];
    assign P[24] = in[42] ^ in2[42];
    assign G[25] = in[41] & in2[41];
    assign P[25] = in[41] ^ in2[41];
    assign G[26] = in[40] & in2[40];
    assign P[26] = in[40] ^ in2[40];
    assign G[27] = in[39] & in2[39];
    assign P[27] = in[39] ^ in2[39];
    assign G[28] = in[38] & in2[38];
    assign P[28] = in[38] ^ in2[38];
    assign G[29] = in[37] & in2[37];
    assign P[29] = in[37] ^ in2[37];
    assign G[30] = in[36] & in2[36];
    assign P[30] = in[36] ^ in2[36];
    assign G[31] = in[35] & in2[35];
    assign P[31] = in[35] ^ in2[35];
    assign G[32] = in[34] & in2[34];
    assign P[32] = in[34] ^ in2[34];
    assign G[33] = in[33] & in2[33];
    assign P[33] = in[33] ^ in2[33];
    assign G[34] = in[32] & in2[32];
    assign P[34] = in[32] ^ in2[32];
    assign G[35] = in[31] & in2[31];
    assign P[35] = in[31] ^ in2[31];
    assign G[36] = in[30] & in2[30];
    assign P[36] = in[30] ^ in2[30];
    assign G[37] = in[29] & in2[29];
    assign P[37] = in[29] ^ in2[29];
    assign G[38] = in[28] & in2[28];
    assign P[38] = in[28] ^ in2[28];
    assign G[39] = in[27] & in2[27];
    assign P[39] = in[27] ^ in2[27];
    assign G[40] = in[26] & in2[26];
    assign P[40] = in[26] ^ in2[26];
    assign G[41] = in[25] & in2[25];
    assign P[41] = in[25] ^ in2[25];
    assign G[42] = in[24] & in2[24];
    assign P[42] = in[24] ^ in2[24];
    assign G[43] = in[23] & in2[23];
    assign P[43] = in[23] ^ in2[23];
    assign G[44] = in[22] & in2[22];
    assign P[44] = in[22] ^ in2[22];
    assign G[45] = in[21] & in2[21];
    assign P[45] = in[21] ^ in2[21];
    assign G[46] = in[20] & in2[20];
    assign P[46] = in[20] ^ in2[20];
    assign G[47] = in[19] & in2[19];
    assign P[47] = in[19] ^ in2[19];
    assign G[48] = in[18] & in2[18];
    assign P[48] = in[18] ^ in2[18];
    assign G[49] = in[17] & in2[17];
    assign P[49] = in[17] ^ in2[17];
    assign G[50] = in[16] & in2[16];
    assign P[50] = in[16] ^ in2[16];
    assign G[51] = in[15] & in2[15];
    assign P[51] = in[15] ^ in2[15];
    assign G[52] = in[14] & in2[14];
    assign P[52] = in[14] ^ in2[14];
    assign G[53] = in[13] & in2[13];
    assign P[53] = in[13] ^ in2[13];
    assign G[54] = in[12] & in2[12];
    assign P[54] = in[12] ^ in2[12];
    assign G[55] = in[11] & in2[11];
    assign P[55] = in[11] ^ in2[11];
    assign G[56] = in[10] & in2[10];
    assign P[56] = in[10] ^ in2[10];
    assign G[57] = in[9] & in2[9];
    assign P[57] = in[9] ^ in2[9];
    assign G[58] = in[8] & in2[8];
    assign P[58] = in[8] ^ in2[8];
    assign G[59] = in[7] & in2[7];
    assign P[59] = in[7] ^ in2[7];
    assign G[60] = in[6] & in2[6];
    assign P[60] = in[6] ^ in2[6];
    assign G[61] = in[5] & in2[5];
    assign P[61] = in[5] ^ in2[5];
    assign G[62] = in[4] & in2[4];
    assign P[62] = in[4] ^ in2[4];
    assign G[63] = in[3] & in2[3];
    assign P[63] = in[3] ^ in2[3];
    assign G[64] = in[2] & in2[2];
    assign P[64] = in[2] ^ in2[2];
    assign G[65] = in[1] & in2[1];
    assign P[65] = in[1] ^ in2[1];
    assign G[66] = in[0] & in2[0];
    assign P[66] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign C[66] = G[65] | (P[65] & C[65]);
    assign cout = G[66] | (P[66] & C[66]);
    assign sum = P ^ C;
endmodule

module CLA66(output [65:0] sum, output cout, input [65:0] in1, input [65:0] in2;

    wire[65:0] G;
    wire[65:0] C;
    wire[65:0] P;

    assign G[0] = in[65] & in2[65];
    assign P[0] = in[65] ^ in2[65];
    assign G[1] = in[64] & in2[64];
    assign P[1] = in[64] ^ in2[64];
    assign G[2] = in[63] & in2[63];
    assign P[2] = in[63] ^ in2[63];
    assign G[3] = in[62] & in2[62];
    assign P[3] = in[62] ^ in2[62];
    assign G[4] = in[61] & in2[61];
    assign P[4] = in[61] ^ in2[61];
    assign G[5] = in[60] & in2[60];
    assign P[5] = in[60] ^ in2[60];
    assign G[6] = in[59] & in2[59];
    assign P[6] = in[59] ^ in2[59];
    assign G[7] = in[58] & in2[58];
    assign P[7] = in[58] ^ in2[58];
    assign G[8] = in[57] & in2[57];
    assign P[8] = in[57] ^ in2[57];
    assign G[9] = in[56] & in2[56];
    assign P[9] = in[56] ^ in2[56];
    assign G[10] = in[55] & in2[55];
    assign P[10] = in[55] ^ in2[55];
    assign G[11] = in[54] & in2[54];
    assign P[11] = in[54] ^ in2[54];
    assign G[12] = in[53] & in2[53];
    assign P[12] = in[53] ^ in2[53];
    assign G[13] = in[52] & in2[52];
    assign P[13] = in[52] ^ in2[52];
    assign G[14] = in[51] & in2[51];
    assign P[14] = in[51] ^ in2[51];
    assign G[15] = in[50] & in2[50];
    assign P[15] = in[50] ^ in2[50];
    assign G[16] = in[49] & in2[49];
    assign P[16] = in[49] ^ in2[49];
    assign G[17] = in[48] & in2[48];
    assign P[17] = in[48] ^ in2[48];
    assign G[18] = in[47] & in2[47];
    assign P[18] = in[47] ^ in2[47];
    assign G[19] = in[46] & in2[46];
    assign P[19] = in[46] ^ in2[46];
    assign G[20] = in[45] & in2[45];
    assign P[20] = in[45] ^ in2[45];
    assign G[21] = in[44] & in2[44];
    assign P[21] = in[44] ^ in2[44];
    assign G[22] = in[43] & in2[43];
    assign P[22] = in[43] ^ in2[43];
    assign G[23] = in[42] & in2[42];
    assign P[23] = in[42] ^ in2[42];
    assign G[24] = in[41] & in2[41];
    assign P[24] = in[41] ^ in2[41];
    assign G[25] = in[40] & in2[40];
    assign P[25] = in[40] ^ in2[40];
    assign G[26] = in[39] & in2[39];
    assign P[26] = in[39] ^ in2[39];
    assign G[27] = in[38] & in2[38];
    assign P[27] = in[38] ^ in2[38];
    assign G[28] = in[37] & in2[37];
    assign P[28] = in[37] ^ in2[37];
    assign G[29] = in[36] & in2[36];
    assign P[29] = in[36] ^ in2[36];
    assign G[30] = in[35] & in2[35];
    assign P[30] = in[35] ^ in2[35];
    assign G[31] = in[34] & in2[34];
    assign P[31] = in[34] ^ in2[34];
    assign G[32] = in[33] & in2[33];
    assign P[32] = in[33] ^ in2[33];
    assign G[33] = in[32] & in2[32];
    assign P[33] = in[32] ^ in2[32];
    assign G[34] = in[31] & in2[31];
    assign P[34] = in[31] ^ in2[31];
    assign G[35] = in[30] & in2[30];
    assign P[35] = in[30] ^ in2[30];
    assign G[36] = in[29] & in2[29];
    assign P[36] = in[29] ^ in2[29];
    assign G[37] = in[28] & in2[28];
    assign P[37] = in[28] ^ in2[28];
    assign G[38] = in[27] & in2[27];
    assign P[38] = in[27] ^ in2[27];
    assign G[39] = in[26] & in2[26];
    assign P[39] = in[26] ^ in2[26];
    assign G[40] = in[25] & in2[25];
    assign P[40] = in[25] ^ in2[25];
    assign G[41] = in[24] & in2[24];
    assign P[41] = in[24] ^ in2[24];
    assign G[42] = in[23] & in2[23];
    assign P[42] = in[23] ^ in2[23];
    assign G[43] = in[22] & in2[22];
    assign P[43] = in[22] ^ in2[22];
    assign G[44] = in[21] & in2[21];
    assign P[44] = in[21] ^ in2[21];
    assign G[45] = in[20] & in2[20];
    assign P[45] = in[20] ^ in2[20];
    assign G[46] = in[19] & in2[19];
    assign P[46] = in[19] ^ in2[19];
    assign G[47] = in[18] & in2[18];
    assign P[47] = in[18] ^ in2[18];
    assign G[48] = in[17] & in2[17];
    assign P[48] = in[17] ^ in2[17];
    assign G[49] = in[16] & in2[16];
    assign P[49] = in[16] ^ in2[16];
    assign G[50] = in[15] & in2[15];
    assign P[50] = in[15] ^ in2[15];
    assign G[51] = in[14] & in2[14];
    assign P[51] = in[14] ^ in2[14];
    assign G[52] = in[13] & in2[13];
    assign P[52] = in[13] ^ in2[13];
    assign G[53] = in[12] & in2[12];
    assign P[53] = in[12] ^ in2[12];
    assign G[54] = in[11] & in2[11];
    assign P[54] = in[11] ^ in2[11];
    assign G[55] = in[10] & in2[10];
    assign P[55] = in[10] ^ in2[10];
    assign G[56] = in[9] & in2[9];
    assign P[56] = in[9] ^ in2[9];
    assign G[57] = in[8] & in2[8];
    assign P[57] = in[8] ^ in2[8];
    assign G[58] = in[7] & in2[7];
    assign P[58] = in[7] ^ in2[7];
    assign G[59] = in[6] & in2[6];
    assign P[59] = in[6] ^ in2[6];
    assign G[60] = in[5] & in2[5];
    assign P[60] = in[5] ^ in2[5];
    assign G[61] = in[4] & in2[4];
    assign P[61] = in[4] ^ in2[4];
    assign G[62] = in[3] & in2[3];
    assign P[62] = in[3] ^ in2[3];
    assign G[63] = in[2] & in2[2];
    assign P[63] = in[2] ^ in2[2];
    assign G[64] = in[1] & in2[1];
    assign P[64] = in[1] ^ in2[1];
    assign G[65] = in[0] & in2[0];
    assign P[65] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign C[65] = G[64] | (P[64] & C[64]);
    assign cout = G[65] | (P[65] & C[65]);
    assign sum = P ^ C;
endmodule

module CLA65(output [64:0] sum, output cout, input [64:0] in1, input [64:0] in2;

    wire[64:0] G;
    wire[64:0] C;
    wire[64:0] P;

    assign G[0] = in[64] & in2[64];
    assign P[0] = in[64] ^ in2[64];
    assign G[1] = in[63] & in2[63];
    assign P[1] = in[63] ^ in2[63];
    assign G[2] = in[62] & in2[62];
    assign P[2] = in[62] ^ in2[62];
    assign G[3] = in[61] & in2[61];
    assign P[3] = in[61] ^ in2[61];
    assign G[4] = in[60] & in2[60];
    assign P[4] = in[60] ^ in2[60];
    assign G[5] = in[59] & in2[59];
    assign P[5] = in[59] ^ in2[59];
    assign G[6] = in[58] & in2[58];
    assign P[6] = in[58] ^ in2[58];
    assign G[7] = in[57] & in2[57];
    assign P[7] = in[57] ^ in2[57];
    assign G[8] = in[56] & in2[56];
    assign P[8] = in[56] ^ in2[56];
    assign G[9] = in[55] & in2[55];
    assign P[9] = in[55] ^ in2[55];
    assign G[10] = in[54] & in2[54];
    assign P[10] = in[54] ^ in2[54];
    assign G[11] = in[53] & in2[53];
    assign P[11] = in[53] ^ in2[53];
    assign G[12] = in[52] & in2[52];
    assign P[12] = in[52] ^ in2[52];
    assign G[13] = in[51] & in2[51];
    assign P[13] = in[51] ^ in2[51];
    assign G[14] = in[50] & in2[50];
    assign P[14] = in[50] ^ in2[50];
    assign G[15] = in[49] & in2[49];
    assign P[15] = in[49] ^ in2[49];
    assign G[16] = in[48] & in2[48];
    assign P[16] = in[48] ^ in2[48];
    assign G[17] = in[47] & in2[47];
    assign P[17] = in[47] ^ in2[47];
    assign G[18] = in[46] & in2[46];
    assign P[18] = in[46] ^ in2[46];
    assign G[19] = in[45] & in2[45];
    assign P[19] = in[45] ^ in2[45];
    assign G[20] = in[44] & in2[44];
    assign P[20] = in[44] ^ in2[44];
    assign G[21] = in[43] & in2[43];
    assign P[21] = in[43] ^ in2[43];
    assign G[22] = in[42] & in2[42];
    assign P[22] = in[42] ^ in2[42];
    assign G[23] = in[41] & in2[41];
    assign P[23] = in[41] ^ in2[41];
    assign G[24] = in[40] & in2[40];
    assign P[24] = in[40] ^ in2[40];
    assign G[25] = in[39] & in2[39];
    assign P[25] = in[39] ^ in2[39];
    assign G[26] = in[38] & in2[38];
    assign P[26] = in[38] ^ in2[38];
    assign G[27] = in[37] & in2[37];
    assign P[27] = in[37] ^ in2[37];
    assign G[28] = in[36] & in2[36];
    assign P[28] = in[36] ^ in2[36];
    assign G[29] = in[35] & in2[35];
    assign P[29] = in[35] ^ in2[35];
    assign G[30] = in[34] & in2[34];
    assign P[30] = in[34] ^ in2[34];
    assign G[31] = in[33] & in2[33];
    assign P[31] = in[33] ^ in2[33];
    assign G[32] = in[32] & in2[32];
    assign P[32] = in[32] ^ in2[32];
    assign G[33] = in[31] & in2[31];
    assign P[33] = in[31] ^ in2[31];
    assign G[34] = in[30] & in2[30];
    assign P[34] = in[30] ^ in2[30];
    assign G[35] = in[29] & in2[29];
    assign P[35] = in[29] ^ in2[29];
    assign G[36] = in[28] & in2[28];
    assign P[36] = in[28] ^ in2[28];
    assign G[37] = in[27] & in2[27];
    assign P[37] = in[27] ^ in2[27];
    assign G[38] = in[26] & in2[26];
    assign P[38] = in[26] ^ in2[26];
    assign G[39] = in[25] & in2[25];
    assign P[39] = in[25] ^ in2[25];
    assign G[40] = in[24] & in2[24];
    assign P[40] = in[24] ^ in2[24];
    assign G[41] = in[23] & in2[23];
    assign P[41] = in[23] ^ in2[23];
    assign G[42] = in[22] & in2[22];
    assign P[42] = in[22] ^ in2[22];
    assign G[43] = in[21] & in2[21];
    assign P[43] = in[21] ^ in2[21];
    assign G[44] = in[20] & in2[20];
    assign P[44] = in[20] ^ in2[20];
    assign G[45] = in[19] & in2[19];
    assign P[45] = in[19] ^ in2[19];
    assign G[46] = in[18] & in2[18];
    assign P[46] = in[18] ^ in2[18];
    assign G[47] = in[17] & in2[17];
    assign P[47] = in[17] ^ in2[17];
    assign G[48] = in[16] & in2[16];
    assign P[48] = in[16] ^ in2[16];
    assign G[49] = in[15] & in2[15];
    assign P[49] = in[15] ^ in2[15];
    assign G[50] = in[14] & in2[14];
    assign P[50] = in[14] ^ in2[14];
    assign G[51] = in[13] & in2[13];
    assign P[51] = in[13] ^ in2[13];
    assign G[52] = in[12] & in2[12];
    assign P[52] = in[12] ^ in2[12];
    assign G[53] = in[11] & in2[11];
    assign P[53] = in[11] ^ in2[11];
    assign G[54] = in[10] & in2[10];
    assign P[54] = in[10] ^ in2[10];
    assign G[55] = in[9] & in2[9];
    assign P[55] = in[9] ^ in2[9];
    assign G[56] = in[8] & in2[8];
    assign P[56] = in[8] ^ in2[8];
    assign G[57] = in[7] & in2[7];
    assign P[57] = in[7] ^ in2[7];
    assign G[58] = in[6] & in2[6];
    assign P[58] = in[6] ^ in2[6];
    assign G[59] = in[5] & in2[5];
    assign P[59] = in[5] ^ in2[5];
    assign G[60] = in[4] & in2[4];
    assign P[60] = in[4] ^ in2[4];
    assign G[61] = in[3] & in2[3];
    assign P[61] = in[3] ^ in2[3];
    assign G[62] = in[2] & in2[2];
    assign P[62] = in[2] ^ in2[2];
    assign G[63] = in[1] & in2[1];
    assign P[63] = in[1] ^ in2[1];
    assign G[64] = in[0] & in2[0];
    assign P[64] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign C[64] = G[63] | (P[63] & C[63]);
    assign cout = G[64] | (P[64] & C[64]);
    assign sum = P ^ C;
endmodule

module CLA64(output [63:0] sum, output cout, input [63:0] in1, input [63:0] in2;

    wire[63:0] G;
    wire[63:0] C;
    wire[63:0] P;

    assign G[0] = in[63] & in2[63];
    assign P[0] = in[63] ^ in2[63];
    assign G[1] = in[62] & in2[62];
    assign P[1] = in[62] ^ in2[62];
    assign G[2] = in[61] & in2[61];
    assign P[2] = in[61] ^ in2[61];
    assign G[3] = in[60] & in2[60];
    assign P[3] = in[60] ^ in2[60];
    assign G[4] = in[59] & in2[59];
    assign P[4] = in[59] ^ in2[59];
    assign G[5] = in[58] & in2[58];
    assign P[5] = in[58] ^ in2[58];
    assign G[6] = in[57] & in2[57];
    assign P[6] = in[57] ^ in2[57];
    assign G[7] = in[56] & in2[56];
    assign P[7] = in[56] ^ in2[56];
    assign G[8] = in[55] & in2[55];
    assign P[8] = in[55] ^ in2[55];
    assign G[9] = in[54] & in2[54];
    assign P[9] = in[54] ^ in2[54];
    assign G[10] = in[53] & in2[53];
    assign P[10] = in[53] ^ in2[53];
    assign G[11] = in[52] & in2[52];
    assign P[11] = in[52] ^ in2[52];
    assign G[12] = in[51] & in2[51];
    assign P[12] = in[51] ^ in2[51];
    assign G[13] = in[50] & in2[50];
    assign P[13] = in[50] ^ in2[50];
    assign G[14] = in[49] & in2[49];
    assign P[14] = in[49] ^ in2[49];
    assign G[15] = in[48] & in2[48];
    assign P[15] = in[48] ^ in2[48];
    assign G[16] = in[47] & in2[47];
    assign P[16] = in[47] ^ in2[47];
    assign G[17] = in[46] & in2[46];
    assign P[17] = in[46] ^ in2[46];
    assign G[18] = in[45] & in2[45];
    assign P[18] = in[45] ^ in2[45];
    assign G[19] = in[44] & in2[44];
    assign P[19] = in[44] ^ in2[44];
    assign G[20] = in[43] & in2[43];
    assign P[20] = in[43] ^ in2[43];
    assign G[21] = in[42] & in2[42];
    assign P[21] = in[42] ^ in2[42];
    assign G[22] = in[41] & in2[41];
    assign P[22] = in[41] ^ in2[41];
    assign G[23] = in[40] & in2[40];
    assign P[23] = in[40] ^ in2[40];
    assign G[24] = in[39] & in2[39];
    assign P[24] = in[39] ^ in2[39];
    assign G[25] = in[38] & in2[38];
    assign P[25] = in[38] ^ in2[38];
    assign G[26] = in[37] & in2[37];
    assign P[26] = in[37] ^ in2[37];
    assign G[27] = in[36] & in2[36];
    assign P[27] = in[36] ^ in2[36];
    assign G[28] = in[35] & in2[35];
    assign P[28] = in[35] ^ in2[35];
    assign G[29] = in[34] & in2[34];
    assign P[29] = in[34] ^ in2[34];
    assign G[30] = in[33] & in2[33];
    assign P[30] = in[33] ^ in2[33];
    assign G[31] = in[32] & in2[32];
    assign P[31] = in[32] ^ in2[32];
    assign G[32] = in[31] & in2[31];
    assign P[32] = in[31] ^ in2[31];
    assign G[33] = in[30] & in2[30];
    assign P[33] = in[30] ^ in2[30];
    assign G[34] = in[29] & in2[29];
    assign P[34] = in[29] ^ in2[29];
    assign G[35] = in[28] & in2[28];
    assign P[35] = in[28] ^ in2[28];
    assign G[36] = in[27] & in2[27];
    assign P[36] = in[27] ^ in2[27];
    assign G[37] = in[26] & in2[26];
    assign P[37] = in[26] ^ in2[26];
    assign G[38] = in[25] & in2[25];
    assign P[38] = in[25] ^ in2[25];
    assign G[39] = in[24] & in2[24];
    assign P[39] = in[24] ^ in2[24];
    assign G[40] = in[23] & in2[23];
    assign P[40] = in[23] ^ in2[23];
    assign G[41] = in[22] & in2[22];
    assign P[41] = in[22] ^ in2[22];
    assign G[42] = in[21] & in2[21];
    assign P[42] = in[21] ^ in2[21];
    assign G[43] = in[20] & in2[20];
    assign P[43] = in[20] ^ in2[20];
    assign G[44] = in[19] & in2[19];
    assign P[44] = in[19] ^ in2[19];
    assign G[45] = in[18] & in2[18];
    assign P[45] = in[18] ^ in2[18];
    assign G[46] = in[17] & in2[17];
    assign P[46] = in[17] ^ in2[17];
    assign G[47] = in[16] & in2[16];
    assign P[47] = in[16] ^ in2[16];
    assign G[48] = in[15] & in2[15];
    assign P[48] = in[15] ^ in2[15];
    assign G[49] = in[14] & in2[14];
    assign P[49] = in[14] ^ in2[14];
    assign G[50] = in[13] & in2[13];
    assign P[50] = in[13] ^ in2[13];
    assign G[51] = in[12] & in2[12];
    assign P[51] = in[12] ^ in2[12];
    assign G[52] = in[11] & in2[11];
    assign P[52] = in[11] ^ in2[11];
    assign G[53] = in[10] & in2[10];
    assign P[53] = in[10] ^ in2[10];
    assign G[54] = in[9] & in2[9];
    assign P[54] = in[9] ^ in2[9];
    assign G[55] = in[8] & in2[8];
    assign P[55] = in[8] ^ in2[8];
    assign G[56] = in[7] & in2[7];
    assign P[56] = in[7] ^ in2[7];
    assign G[57] = in[6] & in2[6];
    assign P[57] = in[6] ^ in2[6];
    assign G[58] = in[5] & in2[5];
    assign P[58] = in[5] ^ in2[5];
    assign G[59] = in[4] & in2[4];
    assign P[59] = in[4] ^ in2[4];
    assign G[60] = in[3] & in2[3];
    assign P[60] = in[3] ^ in2[3];
    assign G[61] = in[2] & in2[2];
    assign P[61] = in[2] ^ in2[2];
    assign G[62] = in[1] & in2[1];
    assign P[62] = in[1] ^ in2[1];
    assign G[63] = in[0] & in2[0];
    assign P[63] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign C[63] = G[62] | (P[62] & C[62]);
    assign cout = G[63] | (P[63] & C[63]);
    assign sum = P ^ C;
endmodule

module CLA63(output [62:0] sum, output cout, input [62:0] in1, input [62:0] in2;

    wire[62:0] G;
    wire[62:0] C;
    wire[62:0] P;

    assign G[0] = in[62] & in2[62];
    assign P[0] = in[62] ^ in2[62];
    assign G[1] = in[61] & in2[61];
    assign P[1] = in[61] ^ in2[61];
    assign G[2] = in[60] & in2[60];
    assign P[2] = in[60] ^ in2[60];
    assign G[3] = in[59] & in2[59];
    assign P[3] = in[59] ^ in2[59];
    assign G[4] = in[58] & in2[58];
    assign P[4] = in[58] ^ in2[58];
    assign G[5] = in[57] & in2[57];
    assign P[5] = in[57] ^ in2[57];
    assign G[6] = in[56] & in2[56];
    assign P[6] = in[56] ^ in2[56];
    assign G[7] = in[55] & in2[55];
    assign P[7] = in[55] ^ in2[55];
    assign G[8] = in[54] & in2[54];
    assign P[8] = in[54] ^ in2[54];
    assign G[9] = in[53] & in2[53];
    assign P[9] = in[53] ^ in2[53];
    assign G[10] = in[52] & in2[52];
    assign P[10] = in[52] ^ in2[52];
    assign G[11] = in[51] & in2[51];
    assign P[11] = in[51] ^ in2[51];
    assign G[12] = in[50] & in2[50];
    assign P[12] = in[50] ^ in2[50];
    assign G[13] = in[49] & in2[49];
    assign P[13] = in[49] ^ in2[49];
    assign G[14] = in[48] & in2[48];
    assign P[14] = in[48] ^ in2[48];
    assign G[15] = in[47] & in2[47];
    assign P[15] = in[47] ^ in2[47];
    assign G[16] = in[46] & in2[46];
    assign P[16] = in[46] ^ in2[46];
    assign G[17] = in[45] & in2[45];
    assign P[17] = in[45] ^ in2[45];
    assign G[18] = in[44] & in2[44];
    assign P[18] = in[44] ^ in2[44];
    assign G[19] = in[43] & in2[43];
    assign P[19] = in[43] ^ in2[43];
    assign G[20] = in[42] & in2[42];
    assign P[20] = in[42] ^ in2[42];
    assign G[21] = in[41] & in2[41];
    assign P[21] = in[41] ^ in2[41];
    assign G[22] = in[40] & in2[40];
    assign P[22] = in[40] ^ in2[40];
    assign G[23] = in[39] & in2[39];
    assign P[23] = in[39] ^ in2[39];
    assign G[24] = in[38] & in2[38];
    assign P[24] = in[38] ^ in2[38];
    assign G[25] = in[37] & in2[37];
    assign P[25] = in[37] ^ in2[37];
    assign G[26] = in[36] & in2[36];
    assign P[26] = in[36] ^ in2[36];
    assign G[27] = in[35] & in2[35];
    assign P[27] = in[35] ^ in2[35];
    assign G[28] = in[34] & in2[34];
    assign P[28] = in[34] ^ in2[34];
    assign G[29] = in[33] & in2[33];
    assign P[29] = in[33] ^ in2[33];
    assign G[30] = in[32] & in2[32];
    assign P[30] = in[32] ^ in2[32];
    assign G[31] = in[31] & in2[31];
    assign P[31] = in[31] ^ in2[31];
    assign G[32] = in[30] & in2[30];
    assign P[32] = in[30] ^ in2[30];
    assign G[33] = in[29] & in2[29];
    assign P[33] = in[29] ^ in2[29];
    assign G[34] = in[28] & in2[28];
    assign P[34] = in[28] ^ in2[28];
    assign G[35] = in[27] & in2[27];
    assign P[35] = in[27] ^ in2[27];
    assign G[36] = in[26] & in2[26];
    assign P[36] = in[26] ^ in2[26];
    assign G[37] = in[25] & in2[25];
    assign P[37] = in[25] ^ in2[25];
    assign G[38] = in[24] & in2[24];
    assign P[38] = in[24] ^ in2[24];
    assign G[39] = in[23] & in2[23];
    assign P[39] = in[23] ^ in2[23];
    assign G[40] = in[22] & in2[22];
    assign P[40] = in[22] ^ in2[22];
    assign G[41] = in[21] & in2[21];
    assign P[41] = in[21] ^ in2[21];
    assign G[42] = in[20] & in2[20];
    assign P[42] = in[20] ^ in2[20];
    assign G[43] = in[19] & in2[19];
    assign P[43] = in[19] ^ in2[19];
    assign G[44] = in[18] & in2[18];
    assign P[44] = in[18] ^ in2[18];
    assign G[45] = in[17] & in2[17];
    assign P[45] = in[17] ^ in2[17];
    assign G[46] = in[16] & in2[16];
    assign P[46] = in[16] ^ in2[16];
    assign G[47] = in[15] & in2[15];
    assign P[47] = in[15] ^ in2[15];
    assign G[48] = in[14] & in2[14];
    assign P[48] = in[14] ^ in2[14];
    assign G[49] = in[13] & in2[13];
    assign P[49] = in[13] ^ in2[13];
    assign G[50] = in[12] & in2[12];
    assign P[50] = in[12] ^ in2[12];
    assign G[51] = in[11] & in2[11];
    assign P[51] = in[11] ^ in2[11];
    assign G[52] = in[10] & in2[10];
    assign P[52] = in[10] ^ in2[10];
    assign G[53] = in[9] & in2[9];
    assign P[53] = in[9] ^ in2[9];
    assign G[54] = in[8] & in2[8];
    assign P[54] = in[8] ^ in2[8];
    assign G[55] = in[7] & in2[7];
    assign P[55] = in[7] ^ in2[7];
    assign G[56] = in[6] & in2[6];
    assign P[56] = in[6] ^ in2[6];
    assign G[57] = in[5] & in2[5];
    assign P[57] = in[5] ^ in2[5];
    assign G[58] = in[4] & in2[4];
    assign P[58] = in[4] ^ in2[4];
    assign G[59] = in[3] & in2[3];
    assign P[59] = in[3] ^ in2[3];
    assign G[60] = in[2] & in2[2];
    assign P[60] = in[2] ^ in2[2];
    assign G[61] = in[1] & in2[1];
    assign P[61] = in[1] ^ in2[1];
    assign G[62] = in[0] & in2[0];
    assign P[62] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign C[62] = G[61] | (P[61] & C[61]);
    assign cout = G[62] | (P[62] & C[62]);
    assign sum = P ^ C;
endmodule

module CLA62(output [61:0] sum, output cout, input [61:0] in1, input [61:0] in2;

    wire[61:0] G;
    wire[61:0] C;
    wire[61:0] P;

    assign G[0] = in[61] & in2[61];
    assign P[0] = in[61] ^ in2[61];
    assign G[1] = in[60] & in2[60];
    assign P[1] = in[60] ^ in2[60];
    assign G[2] = in[59] & in2[59];
    assign P[2] = in[59] ^ in2[59];
    assign G[3] = in[58] & in2[58];
    assign P[3] = in[58] ^ in2[58];
    assign G[4] = in[57] & in2[57];
    assign P[4] = in[57] ^ in2[57];
    assign G[5] = in[56] & in2[56];
    assign P[5] = in[56] ^ in2[56];
    assign G[6] = in[55] & in2[55];
    assign P[6] = in[55] ^ in2[55];
    assign G[7] = in[54] & in2[54];
    assign P[7] = in[54] ^ in2[54];
    assign G[8] = in[53] & in2[53];
    assign P[8] = in[53] ^ in2[53];
    assign G[9] = in[52] & in2[52];
    assign P[9] = in[52] ^ in2[52];
    assign G[10] = in[51] & in2[51];
    assign P[10] = in[51] ^ in2[51];
    assign G[11] = in[50] & in2[50];
    assign P[11] = in[50] ^ in2[50];
    assign G[12] = in[49] & in2[49];
    assign P[12] = in[49] ^ in2[49];
    assign G[13] = in[48] & in2[48];
    assign P[13] = in[48] ^ in2[48];
    assign G[14] = in[47] & in2[47];
    assign P[14] = in[47] ^ in2[47];
    assign G[15] = in[46] & in2[46];
    assign P[15] = in[46] ^ in2[46];
    assign G[16] = in[45] & in2[45];
    assign P[16] = in[45] ^ in2[45];
    assign G[17] = in[44] & in2[44];
    assign P[17] = in[44] ^ in2[44];
    assign G[18] = in[43] & in2[43];
    assign P[18] = in[43] ^ in2[43];
    assign G[19] = in[42] & in2[42];
    assign P[19] = in[42] ^ in2[42];
    assign G[20] = in[41] & in2[41];
    assign P[20] = in[41] ^ in2[41];
    assign G[21] = in[40] & in2[40];
    assign P[21] = in[40] ^ in2[40];
    assign G[22] = in[39] & in2[39];
    assign P[22] = in[39] ^ in2[39];
    assign G[23] = in[38] & in2[38];
    assign P[23] = in[38] ^ in2[38];
    assign G[24] = in[37] & in2[37];
    assign P[24] = in[37] ^ in2[37];
    assign G[25] = in[36] & in2[36];
    assign P[25] = in[36] ^ in2[36];
    assign G[26] = in[35] & in2[35];
    assign P[26] = in[35] ^ in2[35];
    assign G[27] = in[34] & in2[34];
    assign P[27] = in[34] ^ in2[34];
    assign G[28] = in[33] & in2[33];
    assign P[28] = in[33] ^ in2[33];
    assign G[29] = in[32] & in2[32];
    assign P[29] = in[32] ^ in2[32];
    assign G[30] = in[31] & in2[31];
    assign P[30] = in[31] ^ in2[31];
    assign G[31] = in[30] & in2[30];
    assign P[31] = in[30] ^ in2[30];
    assign G[32] = in[29] & in2[29];
    assign P[32] = in[29] ^ in2[29];
    assign G[33] = in[28] & in2[28];
    assign P[33] = in[28] ^ in2[28];
    assign G[34] = in[27] & in2[27];
    assign P[34] = in[27] ^ in2[27];
    assign G[35] = in[26] & in2[26];
    assign P[35] = in[26] ^ in2[26];
    assign G[36] = in[25] & in2[25];
    assign P[36] = in[25] ^ in2[25];
    assign G[37] = in[24] & in2[24];
    assign P[37] = in[24] ^ in2[24];
    assign G[38] = in[23] & in2[23];
    assign P[38] = in[23] ^ in2[23];
    assign G[39] = in[22] & in2[22];
    assign P[39] = in[22] ^ in2[22];
    assign G[40] = in[21] & in2[21];
    assign P[40] = in[21] ^ in2[21];
    assign G[41] = in[20] & in2[20];
    assign P[41] = in[20] ^ in2[20];
    assign G[42] = in[19] & in2[19];
    assign P[42] = in[19] ^ in2[19];
    assign G[43] = in[18] & in2[18];
    assign P[43] = in[18] ^ in2[18];
    assign G[44] = in[17] & in2[17];
    assign P[44] = in[17] ^ in2[17];
    assign G[45] = in[16] & in2[16];
    assign P[45] = in[16] ^ in2[16];
    assign G[46] = in[15] & in2[15];
    assign P[46] = in[15] ^ in2[15];
    assign G[47] = in[14] & in2[14];
    assign P[47] = in[14] ^ in2[14];
    assign G[48] = in[13] & in2[13];
    assign P[48] = in[13] ^ in2[13];
    assign G[49] = in[12] & in2[12];
    assign P[49] = in[12] ^ in2[12];
    assign G[50] = in[11] & in2[11];
    assign P[50] = in[11] ^ in2[11];
    assign G[51] = in[10] & in2[10];
    assign P[51] = in[10] ^ in2[10];
    assign G[52] = in[9] & in2[9];
    assign P[52] = in[9] ^ in2[9];
    assign G[53] = in[8] & in2[8];
    assign P[53] = in[8] ^ in2[8];
    assign G[54] = in[7] & in2[7];
    assign P[54] = in[7] ^ in2[7];
    assign G[55] = in[6] & in2[6];
    assign P[55] = in[6] ^ in2[6];
    assign G[56] = in[5] & in2[5];
    assign P[56] = in[5] ^ in2[5];
    assign G[57] = in[4] & in2[4];
    assign P[57] = in[4] ^ in2[4];
    assign G[58] = in[3] & in2[3];
    assign P[58] = in[3] ^ in2[3];
    assign G[59] = in[2] & in2[2];
    assign P[59] = in[2] ^ in2[2];
    assign G[60] = in[1] & in2[1];
    assign P[60] = in[1] ^ in2[1];
    assign G[61] = in[0] & in2[0];
    assign P[61] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign C[61] = G[60] | (P[60] & C[60]);
    assign cout = G[61] | (P[61] & C[61]);
    assign sum = P ^ C;
endmodule

module CLA61(output [60:0] sum, output cout, input [60:0] in1, input [60:0] in2;

    wire[60:0] G;
    wire[60:0] C;
    wire[60:0] P;

    assign G[0] = in[60] & in2[60];
    assign P[0] = in[60] ^ in2[60];
    assign G[1] = in[59] & in2[59];
    assign P[1] = in[59] ^ in2[59];
    assign G[2] = in[58] & in2[58];
    assign P[2] = in[58] ^ in2[58];
    assign G[3] = in[57] & in2[57];
    assign P[3] = in[57] ^ in2[57];
    assign G[4] = in[56] & in2[56];
    assign P[4] = in[56] ^ in2[56];
    assign G[5] = in[55] & in2[55];
    assign P[5] = in[55] ^ in2[55];
    assign G[6] = in[54] & in2[54];
    assign P[6] = in[54] ^ in2[54];
    assign G[7] = in[53] & in2[53];
    assign P[7] = in[53] ^ in2[53];
    assign G[8] = in[52] & in2[52];
    assign P[8] = in[52] ^ in2[52];
    assign G[9] = in[51] & in2[51];
    assign P[9] = in[51] ^ in2[51];
    assign G[10] = in[50] & in2[50];
    assign P[10] = in[50] ^ in2[50];
    assign G[11] = in[49] & in2[49];
    assign P[11] = in[49] ^ in2[49];
    assign G[12] = in[48] & in2[48];
    assign P[12] = in[48] ^ in2[48];
    assign G[13] = in[47] & in2[47];
    assign P[13] = in[47] ^ in2[47];
    assign G[14] = in[46] & in2[46];
    assign P[14] = in[46] ^ in2[46];
    assign G[15] = in[45] & in2[45];
    assign P[15] = in[45] ^ in2[45];
    assign G[16] = in[44] & in2[44];
    assign P[16] = in[44] ^ in2[44];
    assign G[17] = in[43] & in2[43];
    assign P[17] = in[43] ^ in2[43];
    assign G[18] = in[42] & in2[42];
    assign P[18] = in[42] ^ in2[42];
    assign G[19] = in[41] & in2[41];
    assign P[19] = in[41] ^ in2[41];
    assign G[20] = in[40] & in2[40];
    assign P[20] = in[40] ^ in2[40];
    assign G[21] = in[39] & in2[39];
    assign P[21] = in[39] ^ in2[39];
    assign G[22] = in[38] & in2[38];
    assign P[22] = in[38] ^ in2[38];
    assign G[23] = in[37] & in2[37];
    assign P[23] = in[37] ^ in2[37];
    assign G[24] = in[36] & in2[36];
    assign P[24] = in[36] ^ in2[36];
    assign G[25] = in[35] & in2[35];
    assign P[25] = in[35] ^ in2[35];
    assign G[26] = in[34] & in2[34];
    assign P[26] = in[34] ^ in2[34];
    assign G[27] = in[33] & in2[33];
    assign P[27] = in[33] ^ in2[33];
    assign G[28] = in[32] & in2[32];
    assign P[28] = in[32] ^ in2[32];
    assign G[29] = in[31] & in2[31];
    assign P[29] = in[31] ^ in2[31];
    assign G[30] = in[30] & in2[30];
    assign P[30] = in[30] ^ in2[30];
    assign G[31] = in[29] & in2[29];
    assign P[31] = in[29] ^ in2[29];
    assign G[32] = in[28] & in2[28];
    assign P[32] = in[28] ^ in2[28];
    assign G[33] = in[27] & in2[27];
    assign P[33] = in[27] ^ in2[27];
    assign G[34] = in[26] & in2[26];
    assign P[34] = in[26] ^ in2[26];
    assign G[35] = in[25] & in2[25];
    assign P[35] = in[25] ^ in2[25];
    assign G[36] = in[24] & in2[24];
    assign P[36] = in[24] ^ in2[24];
    assign G[37] = in[23] & in2[23];
    assign P[37] = in[23] ^ in2[23];
    assign G[38] = in[22] & in2[22];
    assign P[38] = in[22] ^ in2[22];
    assign G[39] = in[21] & in2[21];
    assign P[39] = in[21] ^ in2[21];
    assign G[40] = in[20] & in2[20];
    assign P[40] = in[20] ^ in2[20];
    assign G[41] = in[19] & in2[19];
    assign P[41] = in[19] ^ in2[19];
    assign G[42] = in[18] & in2[18];
    assign P[42] = in[18] ^ in2[18];
    assign G[43] = in[17] & in2[17];
    assign P[43] = in[17] ^ in2[17];
    assign G[44] = in[16] & in2[16];
    assign P[44] = in[16] ^ in2[16];
    assign G[45] = in[15] & in2[15];
    assign P[45] = in[15] ^ in2[15];
    assign G[46] = in[14] & in2[14];
    assign P[46] = in[14] ^ in2[14];
    assign G[47] = in[13] & in2[13];
    assign P[47] = in[13] ^ in2[13];
    assign G[48] = in[12] & in2[12];
    assign P[48] = in[12] ^ in2[12];
    assign G[49] = in[11] & in2[11];
    assign P[49] = in[11] ^ in2[11];
    assign G[50] = in[10] & in2[10];
    assign P[50] = in[10] ^ in2[10];
    assign G[51] = in[9] & in2[9];
    assign P[51] = in[9] ^ in2[9];
    assign G[52] = in[8] & in2[8];
    assign P[52] = in[8] ^ in2[8];
    assign G[53] = in[7] & in2[7];
    assign P[53] = in[7] ^ in2[7];
    assign G[54] = in[6] & in2[6];
    assign P[54] = in[6] ^ in2[6];
    assign G[55] = in[5] & in2[5];
    assign P[55] = in[5] ^ in2[5];
    assign G[56] = in[4] & in2[4];
    assign P[56] = in[4] ^ in2[4];
    assign G[57] = in[3] & in2[3];
    assign P[57] = in[3] ^ in2[3];
    assign G[58] = in[2] & in2[2];
    assign P[58] = in[2] ^ in2[2];
    assign G[59] = in[1] & in2[1];
    assign P[59] = in[1] ^ in2[1];
    assign G[60] = in[0] & in2[0];
    assign P[60] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign C[60] = G[59] | (P[59] & C[59]);
    assign cout = G[60] | (P[60] & C[60]);
    assign sum = P ^ C;
endmodule

module CLA60(output [59:0] sum, output cout, input [59:0] in1, input [59:0] in2;

    wire[59:0] G;
    wire[59:0] C;
    wire[59:0] P;

    assign G[0] = in[59] & in2[59];
    assign P[0] = in[59] ^ in2[59];
    assign G[1] = in[58] & in2[58];
    assign P[1] = in[58] ^ in2[58];
    assign G[2] = in[57] & in2[57];
    assign P[2] = in[57] ^ in2[57];
    assign G[3] = in[56] & in2[56];
    assign P[3] = in[56] ^ in2[56];
    assign G[4] = in[55] & in2[55];
    assign P[4] = in[55] ^ in2[55];
    assign G[5] = in[54] & in2[54];
    assign P[5] = in[54] ^ in2[54];
    assign G[6] = in[53] & in2[53];
    assign P[6] = in[53] ^ in2[53];
    assign G[7] = in[52] & in2[52];
    assign P[7] = in[52] ^ in2[52];
    assign G[8] = in[51] & in2[51];
    assign P[8] = in[51] ^ in2[51];
    assign G[9] = in[50] & in2[50];
    assign P[9] = in[50] ^ in2[50];
    assign G[10] = in[49] & in2[49];
    assign P[10] = in[49] ^ in2[49];
    assign G[11] = in[48] & in2[48];
    assign P[11] = in[48] ^ in2[48];
    assign G[12] = in[47] & in2[47];
    assign P[12] = in[47] ^ in2[47];
    assign G[13] = in[46] & in2[46];
    assign P[13] = in[46] ^ in2[46];
    assign G[14] = in[45] & in2[45];
    assign P[14] = in[45] ^ in2[45];
    assign G[15] = in[44] & in2[44];
    assign P[15] = in[44] ^ in2[44];
    assign G[16] = in[43] & in2[43];
    assign P[16] = in[43] ^ in2[43];
    assign G[17] = in[42] & in2[42];
    assign P[17] = in[42] ^ in2[42];
    assign G[18] = in[41] & in2[41];
    assign P[18] = in[41] ^ in2[41];
    assign G[19] = in[40] & in2[40];
    assign P[19] = in[40] ^ in2[40];
    assign G[20] = in[39] & in2[39];
    assign P[20] = in[39] ^ in2[39];
    assign G[21] = in[38] & in2[38];
    assign P[21] = in[38] ^ in2[38];
    assign G[22] = in[37] & in2[37];
    assign P[22] = in[37] ^ in2[37];
    assign G[23] = in[36] & in2[36];
    assign P[23] = in[36] ^ in2[36];
    assign G[24] = in[35] & in2[35];
    assign P[24] = in[35] ^ in2[35];
    assign G[25] = in[34] & in2[34];
    assign P[25] = in[34] ^ in2[34];
    assign G[26] = in[33] & in2[33];
    assign P[26] = in[33] ^ in2[33];
    assign G[27] = in[32] & in2[32];
    assign P[27] = in[32] ^ in2[32];
    assign G[28] = in[31] & in2[31];
    assign P[28] = in[31] ^ in2[31];
    assign G[29] = in[30] & in2[30];
    assign P[29] = in[30] ^ in2[30];
    assign G[30] = in[29] & in2[29];
    assign P[30] = in[29] ^ in2[29];
    assign G[31] = in[28] & in2[28];
    assign P[31] = in[28] ^ in2[28];
    assign G[32] = in[27] & in2[27];
    assign P[32] = in[27] ^ in2[27];
    assign G[33] = in[26] & in2[26];
    assign P[33] = in[26] ^ in2[26];
    assign G[34] = in[25] & in2[25];
    assign P[34] = in[25] ^ in2[25];
    assign G[35] = in[24] & in2[24];
    assign P[35] = in[24] ^ in2[24];
    assign G[36] = in[23] & in2[23];
    assign P[36] = in[23] ^ in2[23];
    assign G[37] = in[22] & in2[22];
    assign P[37] = in[22] ^ in2[22];
    assign G[38] = in[21] & in2[21];
    assign P[38] = in[21] ^ in2[21];
    assign G[39] = in[20] & in2[20];
    assign P[39] = in[20] ^ in2[20];
    assign G[40] = in[19] & in2[19];
    assign P[40] = in[19] ^ in2[19];
    assign G[41] = in[18] & in2[18];
    assign P[41] = in[18] ^ in2[18];
    assign G[42] = in[17] & in2[17];
    assign P[42] = in[17] ^ in2[17];
    assign G[43] = in[16] & in2[16];
    assign P[43] = in[16] ^ in2[16];
    assign G[44] = in[15] & in2[15];
    assign P[44] = in[15] ^ in2[15];
    assign G[45] = in[14] & in2[14];
    assign P[45] = in[14] ^ in2[14];
    assign G[46] = in[13] & in2[13];
    assign P[46] = in[13] ^ in2[13];
    assign G[47] = in[12] & in2[12];
    assign P[47] = in[12] ^ in2[12];
    assign G[48] = in[11] & in2[11];
    assign P[48] = in[11] ^ in2[11];
    assign G[49] = in[10] & in2[10];
    assign P[49] = in[10] ^ in2[10];
    assign G[50] = in[9] & in2[9];
    assign P[50] = in[9] ^ in2[9];
    assign G[51] = in[8] & in2[8];
    assign P[51] = in[8] ^ in2[8];
    assign G[52] = in[7] & in2[7];
    assign P[52] = in[7] ^ in2[7];
    assign G[53] = in[6] & in2[6];
    assign P[53] = in[6] ^ in2[6];
    assign G[54] = in[5] & in2[5];
    assign P[54] = in[5] ^ in2[5];
    assign G[55] = in[4] & in2[4];
    assign P[55] = in[4] ^ in2[4];
    assign G[56] = in[3] & in2[3];
    assign P[56] = in[3] ^ in2[3];
    assign G[57] = in[2] & in2[2];
    assign P[57] = in[2] ^ in2[2];
    assign G[58] = in[1] & in2[1];
    assign P[58] = in[1] ^ in2[1];
    assign G[59] = in[0] & in2[0];
    assign P[59] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign C[59] = G[58] | (P[58] & C[58]);
    assign cout = G[59] | (P[59] & C[59]);
    assign sum = P ^ C;
endmodule

module CLA59(output [58:0] sum, output cout, input [58:0] in1, input [58:0] in2;

    wire[58:0] G;
    wire[58:0] C;
    wire[58:0] P;

    assign G[0] = in[58] & in2[58];
    assign P[0] = in[58] ^ in2[58];
    assign G[1] = in[57] & in2[57];
    assign P[1] = in[57] ^ in2[57];
    assign G[2] = in[56] & in2[56];
    assign P[2] = in[56] ^ in2[56];
    assign G[3] = in[55] & in2[55];
    assign P[3] = in[55] ^ in2[55];
    assign G[4] = in[54] & in2[54];
    assign P[4] = in[54] ^ in2[54];
    assign G[5] = in[53] & in2[53];
    assign P[5] = in[53] ^ in2[53];
    assign G[6] = in[52] & in2[52];
    assign P[6] = in[52] ^ in2[52];
    assign G[7] = in[51] & in2[51];
    assign P[7] = in[51] ^ in2[51];
    assign G[8] = in[50] & in2[50];
    assign P[8] = in[50] ^ in2[50];
    assign G[9] = in[49] & in2[49];
    assign P[9] = in[49] ^ in2[49];
    assign G[10] = in[48] & in2[48];
    assign P[10] = in[48] ^ in2[48];
    assign G[11] = in[47] & in2[47];
    assign P[11] = in[47] ^ in2[47];
    assign G[12] = in[46] & in2[46];
    assign P[12] = in[46] ^ in2[46];
    assign G[13] = in[45] & in2[45];
    assign P[13] = in[45] ^ in2[45];
    assign G[14] = in[44] & in2[44];
    assign P[14] = in[44] ^ in2[44];
    assign G[15] = in[43] & in2[43];
    assign P[15] = in[43] ^ in2[43];
    assign G[16] = in[42] & in2[42];
    assign P[16] = in[42] ^ in2[42];
    assign G[17] = in[41] & in2[41];
    assign P[17] = in[41] ^ in2[41];
    assign G[18] = in[40] & in2[40];
    assign P[18] = in[40] ^ in2[40];
    assign G[19] = in[39] & in2[39];
    assign P[19] = in[39] ^ in2[39];
    assign G[20] = in[38] & in2[38];
    assign P[20] = in[38] ^ in2[38];
    assign G[21] = in[37] & in2[37];
    assign P[21] = in[37] ^ in2[37];
    assign G[22] = in[36] & in2[36];
    assign P[22] = in[36] ^ in2[36];
    assign G[23] = in[35] & in2[35];
    assign P[23] = in[35] ^ in2[35];
    assign G[24] = in[34] & in2[34];
    assign P[24] = in[34] ^ in2[34];
    assign G[25] = in[33] & in2[33];
    assign P[25] = in[33] ^ in2[33];
    assign G[26] = in[32] & in2[32];
    assign P[26] = in[32] ^ in2[32];
    assign G[27] = in[31] & in2[31];
    assign P[27] = in[31] ^ in2[31];
    assign G[28] = in[30] & in2[30];
    assign P[28] = in[30] ^ in2[30];
    assign G[29] = in[29] & in2[29];
    assign P[29] = in[29] ^ in2[29];
    assign G[30] = in[28] & in2[28];
    assign P[30] = in[28] ^ in2[28];
    assign G[31] = in[27] & in2[27];
    assign P[31] = in[27] ^ in2[27];
    assign G[32] = in[26] & in2[26];
    assign P[32] = in[26] ^ in2[26];
    assign G[33] = in[25] & in2[25];
    assign P[33] = in[25] ^ in2[25];
    assign G[34] = in[24] & in2[24];
    assign P[34] = in[24] ^ in2[24];
    assign G[35] = in[23] & in2[23];
    assign P[35] = in[23] ^ in2[23];
    assign G[36] = in[22] & in2[22];
    assign P[36] = in[22] ^ in2[22];
    assign G[37] = in[21] & in2[21];
    assign P[37] = in[21] ^ in2[21];
    assign G[38] = in[20] & in2[20];
    assign P[38] = in[20] ^ in2[20];
    assign G[39] = in[19] & in2[19];
    assign P[39] = in[19] ^ in2[19];
    assign G[40] = in[18] & in2[18];
    assign P[40] = in[18] ^ in2[18];
    assign G[41] = in[17] & in2[17];
    assign P[41] = in[17] ^ in2[17];
    assign G[42] = in[16] & in2[16];
    assign P[42] = in[16] ^ in2[16];
    assign G[43] = in[15] & in2[15];
    assign P[43] = in[15] ^ in2[15];
    assign G[44] = in[14] & in2[14];
    assign P[44] = in[14] ^ in2[14];
    assign G[45] = in[13] & in2[13];
    assign P[45] = in[13] ^ in2[13];
    assign G[46] = in[12] & in2[12];
    assign P[46] = in[12] ^ in2[12];
    assign G[47] = in[11] & in2[11];
    assign P[47] = in[11] ^ in2[11];
    assign G[48] = in[10] & in2[10];
    assign P[48] = in[10] ^ in2[10];
    assign G[49] = in[9] & in2[9];
    assign P[49] = in[9] ^ in2[9];
    assign G[50] = in[8] & in2[8];
    assign P[50] = in[8] ^ in2[8];
    assign G[51] = in[7] & in2[7];
    assign P[51] = in[7] ^ in2[7];
    assign G[52] = in[6] & in2[6];
    assign P[52] = in[6] ^ in2[6];
    assign G[53] = in[5] & in2[5];
    assign P[53] = in[5] ^ in2[5];
    assign G[54] = in[4] & in2[4];
    assign P[54] = in[4] ^ in2[4];
    assign G[55] = in[3] & in2[3];
    assign P[55] = in[3] ^ in2[3];
    assign G[56] = in[2] & in2[2];
    assign P[56] = in[2] ^ in2[2];
    assign G[57] = in[1] & in2[1];
    assign P[57] = in[1] ^ in2[1];
    assign G[58] = in[0] & in2[0];
    assign P[58] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign C[58] = G[57] | (P[57] & C[57]);
    assign cout = G[58] | (P[58] & C[58]);
    assign sum = P ^ C;
endmodule

module CLA58(output [57:0] sum, output cout, input [57:0] in1, input [57:0] in2;

    wire[57:0] G;
    wire[57:0] C;
    wire[57:0] P;

    assign G[0] = in[57] & in2[57];
    assign P[0] = in[57] ^ in2[57];
    assign G[1] = in[56] & in2[56];
    assign P[1] = in[56] ^ in2[56];
    assign G[2] = in[55] & in2[55];
    assign P[2] = in[55] ^ in2[55];
    assign G[3] = in[54] & in2[54];
    assign P[3] = in[54] ^ in2[54];
    assign G[4] = in[53] & in2[53];
    assign P[4] = in[53] ^ in2[53];
    assign G[5] = in[52] & in2[52];
    assign P[5] = in[52] ^ in2[52];
    assign G[6] = in[51] & in2[51];
    assign P[6] = in[51] ^ in2[51];
    assign G[7] = in[50] & in2[50];
    assign P[7] = in[50] ^ in2[50];
    assign G[8] = in[49] & in2[49];
    assign P[8] = in[49] ^ in2[49];
    assign G[9] = in[48] & in2[48];
    assign P[9] = in[48] ^ in2[48];
    assign G[10] = in[47] & in2[47];
    assign P[10] = in[47] ^ in2[47];
    assign G[11] = in[46] & in2[46];
    assign P[11] = in[46] ^ in2[46];
    assign G[12] = in[45] & in2[45];
    assign P[12] = in[45] ^ in2[45];
    assign G[13] = in[44] & in2[44];
    assign P[13] = in[44] ^ in2[44];
    assign G[14] = in[43] & in2[43];
    assign P[14] = in[43] ^ in2[43];
    assign G[15] = in[42] & in2[42];
    assign P[15] = in[42] ^ in2[42];
    assign G[16] = in[41] & in2[41];
    assign P[16] = in[41] ^ in2[41];
    assign G[17] = in[40] & in2[40];
    assign P[17] = in[40] ^ in2[40];
    assign G[18] = in[39] & in2[39];
    assign P[18] = in[39] ^ in2[39];
    assign G[19] = in[38] & in2[38];
    assign P[19] = in[38] ^ in2[38];
    assign G[20] = in[37] & in2[37];
    assign P[20] = in[37] ^ in2[37];
    assign G[21] = in[36] & in2[36];
    assign P[21] = in[36] ^ in2[36];
    assign G[22] = in[35] & in2[35];
    assign P[22] = in[35] ^ in2[35];
    assign G[23] = in[34] & in2[34];
    assign P[23] = in[34] ^ in2[34];
    assign G[24] = in[33] & in2[33];
    assign P[24] = in[33] ^ in2[33];
    assign G[25] = in[32] & in2[32];
    assign P[25] = in[32] ^ in2[32];
    assign G[26] = in[31] & in2[31];
    assign P[26] = in[31] ^ in2[31];
    assign G[27] = in[30] & in2[30];
    assign P[27] = in[30] ^ in2[30];
    assign G[28] = in[29] & in2[29];
    assign P[28] = in[29] ^ in2[29];
    assign G[29] = in[28] & in2[28];
    assign P[29] = in[28] ^ in2[28];
    assign G[30] = in[27] & in2[27];
    assign P[30] = in[27] ^ in2[27];
    assign G[31] = in[26] & in2[26];
    assign P[31] = in[26] ^ in2[26];
    assign G[32] = in[25] & in2[25];
    assign P[32] = in[25] ^ in2[25];
    assign G[33] = in[24] & in2[24];
    assign P[33] = in[24] ^ in2[24];
    assign G[34] = in[23] & in2[23];
    assign P[34] = in[23] ^ in2[23];
    assign G[35] = in[22] & in2[22];
    assign P[35] = in[22] ^ in2[22];
    assign G[36] = in[21] & in2[21];
    assign P[36] = in[21] ^ in2[21];
    assign G[37] = in[20] & in2[20];
    assign P[37] = in[20] ^ in2[20];
    assign G[38] = in[19] & in2[19];
    assign P[38] = in[19] ^ in2[19];
    assign G[39] = in[18] & in2[18];
    assign P[39] = in[18] ^ in2[18];
    assign G[40] = in[17] & in2[17];
    assign P[40] = in[17] ^ in2[17];
    assign G[41] = in[16] & in2[16];
    assign P[41] = in[16] ^ in2[16];
    assign G[42] = in[15] & in2[15];
    assign P[42] = in[15] ^ in2[15];
    assign G[43] = in[14] & in2[14];
    assign P[43] = in[14] ^ in2[14];
    assign G[44] = in[13] & in2[13];
    assign P[44] = in[13] ^ in2[13];
    assign G[45] = in[12] & in2[12];
    assign P[45] = in[12] ^ in2[12];
    assign G[46] = in[11] & in2[11];
    assign P[46] = in[11] ^ in2[11];
    assign G[47] = in[10] & in2[10];
    assign P[47] = in[10] ^ in2[10];
    assign G[48] = in[9] & in2[9];
    assign P[48] = in[9] ^ in2[9];
    assign G[49] = in[8] & in2[8];
    assign P[49] = in[8] ^ in2[8];
    assign G[50] = in[7] & in2[7];
    assign P[50] = in[7] ^ in2[7];
    assign G[51] = in[6] & in2[6];
    assign P[51] = in[6] ^ in2[6];
    assign G[52] = in[5] & in2[5];
    assign P[52] = in[5] ^ in2[5];
    assign G[53] = in[4] & in2[4];
    assign P[53] = in[4] ^ in2[4];
    assign G[54] = in[3] & in2[3];
    assign P[54] = in[3] ^ in2[3];
    assign G[55] = in[2] & in2[2];
    assign P[55] = in[2] ^ in2[2];
    assign G[56] = in[1] & in2[1];
    assign P[56] = in[1] ^ in2[1];
    assign G[57] = in[0] & in2[0];
    assign P[57] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign C[57] = G[56] | (P[56] & C[56]);
    assign cout = G[57] | (P[57] & C[57]);
    assign sum = P ^ C;
endmodule

module CLA57(output [56:0] sum, output cout, input [56:0] in1, input [56:0] in2;

    wire[56:0] G;
    wire[56:0] C;
    wire[56:0] P;

    assign G[0] = in[56] & in2[56];
    assign P[0] = in[56] ^ in2[56];
    assign G[1] = in[55] & in2[55];
    assign P[1] = in[55] ^ in2[55];
    assign G[2] = in[54] & in2[54];
    assign P[2] = in[54] ^ in2[54];
    assign G[3] = in[53] & in2[53];
    assign P[3] = in[53] ^ in2[53];
    assign G[4] = in[52] & in2[52];
    assign P[4] = in[52] ^ in2[52];
    assign G[5] = in[51] & in2[51];
    assign P[5] = in[51] ^ in2[51];
    assign G[6] = in[50] & in2[50];
    assign P[6] = in[50] ^ in2[50];
    assign G[7] = in[49] & in2[49];
    assign P[7] = in[49] ^ in2[49];
    assign G[8] = in[48] & in2[48];
    assign P[8] = in[48] ^ in2[48];
    assign G[9] = in[47] & in2[47];
    assign P[9] = in[47] ^ in2[47];
    assign G[10] = in[46] & in2[46];
    assign P[10] = in[46] ^ in2[46];
    assign G[11] = in[45] & in2[45];
    assign P[11] = in[45] ^ in2[45];
    assign G[12] = in[44] & in2[44];
    assign P[12] = in[44] ^ in2[44];
    assign G[13] = in[43] & in2[43];
    assign P[13] = in[43] ^ in2[43];
    assign G[14] = in[42] & in2[42];
    assign P[14] = in[42] ^ in2[42];
    assign G[15] = in[41] & in2[41];
    assign P[15] = in[41] ^ in2[41];
    assign G[16] = in[40] & in2[40];
    assign P[16] = in[40] ^ in2[40];
    assign G[17] = in[39] & in2[39];
    assign P[17] = in[39] ^ in2[39];
    assign G[18] = in[38] & in2[38];
    assign P[18] = in[38] ^ in2[38];
    assign G[19] = in[37] & in2[37];
    assign P[19] = in[37] ^ in2[37];
    assign G[20] = in[36] & in2[36];
    assign P[20] = in[36] ^ in2[36];
    assign G[21] = in[35] & in2[35];
    assign P[21] = in[35] ^ in2[35];
    assign G[22] = in[34] & in2[34];
    assign P[22] = in[34] ^ in2[34];
    assign G[23] = in[33] & in2[33];
    assign P[23] = in[33] ^ in2[33];
    assign G[24] = in[32] & in2[32];
    assign P[24] = in[32] ^ in2[32];
    assign G[25] = in[31] & in2[31];
    assign P[25] = in[31] ^ in2[31];
    assign G[26] = in[30] & in2[30];
    assign P[26] = in[30] ^ in2[30];
    assign G[27] = in[29] & in2[29];
    assign P[27] = in[29] ^ in2[29];
    assign G[28] = in[28] & in2[28];
    assign P[28] = in[28] ^ in2[28];
    assign G[29] = in[27] & in2[27];
    assign P[29] = in[27] ^ in2[27];
    assign G[30] = in[26] & in2[26];
    assign P[30] = in[26] ^ in2[26];
    assign G[31] = in[25] & in2[25];
    assign P[31] = in[25] ^ in2[25];
    assign G[32] = in[24] & in2[24];
    assign P[32] = in[24] ^ in2[24];
    assign G[33] = in[23] & in2[23];
    assign P[33] = in[23] ^ in2[23];
    assign G[34] = in[22] & in2[22];
    assign P[34] = in[22] ^ in2[22];
    assign G[35] = in[21] & in2[21];
    assign P[35] = in[21] ^ in2[21];
    assign G[36] = in[20] & in2[20];
    assign P[36] = in[20] ^ in2[20];
    assign G[37] = in[19] & in2[19];
    assign P[37] = in[19] ^ in2[19];
    assign G[38] = in[18] & in2[18];
    assign P[38] = in[18] ^ in2[18];
    assign G[39] = in[17] & in2[17];
    assign P[39] = in[17] ^ in2[17];
    assign G[40] = in[16] & in2[16];
    assign P[40] = in[16] ^ in2[16];
    assign G[41] = in[15] & in2[15];
    assign P[41] = in[15] ^ in2[15];
    assign G[42] = in[14] & in2[14];
    assign P[42] = in[14] ^ in2[14];
    assign G[43] = in[13] & in2[13];
    assign P[43] = in[13] ^ in2[13];
    assign G[44] = in[12] & in2[12];
    assign P[44] = in[12] ^ in2[12];
    assign G[45] = in[11] & in2[11];
    assign P[45] = in[11] ^ in2[11];
    assign G[46] = in[10] & in2[10];
    assign P[46] = in[10] ^ in2[10];
    assign G[47] = in[9] & in2[9];
    assign P[47] = in[9] ^ in2[9];
    assign G[48] = in[8] & in2[8];
    assign P[48] = in[8] ^ in2[8];
    assign G[49] = in[7] & in2[7];
    assign P[49] = in[7] ^ in2[7];
    assign G[50] = in[6] & in2[6];
    assign P[50] = in[6] ^ in2[6];
    assign G[51] = in[5] & in2[5];
    assign P[51] = in[5] ^ in2[5];
    assign G[52] = in[4] & in2[4];
    assign P[52] = in[4] ^ in2[4];
    assign G[53] = in[3] & in2[3];
    assign P[53] = in[3] ^ in2[3];
    assign G[54] = in[2] & in2[2];
    assign P[54] = in[2] ^ in2[2];
    assign G[55] = in[1] & in2[1];
    assign P[55] = in[1] ^ in2[1];
    assign G[56] = in[0] & in2[0];
    assign P[56] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign C[56] = G[55] | (P[55] & C[55]);
    assign cout = G[56] | (P[56] & C[56]);
    assign sum = P ^ C;
endmodule

module CLA56(output [55:0] sum, output cout, input [55:0] in1, input [55:0] in2;

    wire[55:0] G;
    wire[55:0] C;
    wire[55:0] P;

    assign G[0] = in[55] & in2[55];
    assign P[0] = in[55] ^ in2[55];
    assign G[1] = in[54] & in2[54];
    assign P[1] = in[54] ^ in2[54];
    assign G[2] = in[53] & in2[53];
    assign P[2] = in[53] ^ in2[53];
    assign G[3] = in[52] & in2[52];
    assign P[3] = in[52] ^ in2[52];
    assign G[4] = in[51] & in2[51];
    assign P[4] = in[51] ^ in2[51];
    assign G[5] = in[50] & in2[50];
    assign P[5] = in[50] ^ in2[50];
    assign G[6] = in[49] & in2[49];
    assign P[6] = in[49] ^ in2[49];
    assign G[7] = in[48] & in2[48];
    assign P[7] = in[48] ^ in2[48];
    assign G[8] = in[47] & in2[47];
    assign P[8] = in[47] ^ in2[47];
    assign G[9] = in[46] & in2[46];
    assign P[9] = in[46] ^ in2[46];
    assign G[10] = in[45] & in2[45];
    assign P[10] = in[45] ^ in2[45];
    assign G[11] = in[44] & in2[44];
    assign P[11] = in[44] ^ in2[44];
    assign G[12] = in[43] & in2[43];
    assign P[12] = in[43] ^ in2[43];
    assign G[13] = in[42] & in2[42];
    assign P[13] = in[42] ^ in2[42];
    assign G[14] = in[41] & in2[41];
    assign P[14] = in[41] ^ in2[41];
    assign G[15] = in[40] & in2[40];
    assign P[15] = in[40] ^ in2[40];
    assign G[16] = in[39] & in2[39];
    assign P[16] = in[39] ^ in2[39];
    assign G[17] = in[38] & in2[38];
    assign P[17] = in[38] ^ in2[38];
    assign G[18] = in[37] & in2[37];
    assign P[18] = in[37] ^ in2[37];
    assign G[19] = in[36] & in2[36];
    assign P[19] = in[36] ^ in2[36];
    assign G[20] = in[35] & in2[35];
    assign P[20] = in[35] ^ in2[35];
    assign G[21] = in[34] & in2[34];
    assign P[21] = in[34] ^ in2[34];
    assign G[22] = in[33] & in2[33];
    assign P[22] = in[33] ^ in2[33];
    assign G[23] = in[32] & in2[32];
    assign P[23] = in[32] ^ in2[32];
    assign G[24] = in[31] & in2[31];
    assign P[24] = in[31] ^ in2[31];
    assign G[25] = in[30] & in2[30];
    assign P[25] = in[30] ^ in2[30];
    assign G[26] = in[29] & in2[29];
    assign P[26] = in[29] ^ in2[29];
    assign G[27] = in[28] & in2[28];
    assign P[27] = in[28] ^ in2[28];
    assign G[28] = in[27] & in2[27];
    assign P[28] = in[27] ^ in2[27];
    assign G[29] = in[26] & in2[26];
    assign P[29] = in[26] ^ in2[26];
    assign G[30] = in[25] & in2[25];
    assign P[30] = in[25] ^ in2[25];
    assign G[31] = in[24] & in2[24];
    assign P[31] = in[24] ^ in2[24];
    assign G[32] = in[23] & in2[23];
    assign P[32] = in[23] ^ in2[23];
    assign G[33] = in[22] & in2[22];
    assign P[33] = in[22] ^ in2[22];
    assign G[34] = in[21] & in2[21];
    assign P[34] = in[21] ^ in2[21];
    assign G[35] = in[20] & in2[20];
    assign P[35] = in[20] ^ in2[20];
    assign G[36] = in[19] & in2[19];
    assign P[36] = in[19] ^ in2[19];
    assign G[37] = in[18] & in2[18];
    assign P[37] = in[18] ^ in2[18];
    assign G[38] = in[17] & in2[17];
    assign P[38] = in[17] ^ in2[17];
    assign G[39] = in[16] & in2[16];
    assign P[39] = in[16] ^ in2[16];
    assign G[40] = in[15] & in2[15];
    assign P[40] = in[15] ^ in2[15];
    assign G[41] = in[14] & in2[14];
    assign P[41] = in[14] ^ in2[14];
    assign G[42] = in[13] & in2[13];
    assign P[42] = in[13] ^ in2[13];
    assign G[43] = in[12] & in2[12];
    assign P[43] = in[12] ^ in2[12];
    assign G[44] = in[11] & in2[11];
    assign P[44] = in[11] ^ in2[11];
    assign G[45] = in[10] & in2[10];
    assign P[45] = in[10] ^ in2[10];
    assign G[46] = in[9] & in2[9];
    assign P[46] = in[9] ^ in2[9];
    assign G[47] = in[8] & in2[8];
    assign P[47] = in[8] ^ in2[8];
    assign G[48] = in[7] & in2[7];
    assign P[48] = in[7] ^ in2[7];
    assign G[49] = in[6] & in2[6];
    assign P[49] = in[6] ^ in2[6];
    assign G[50] = in[5] & in2[5];
    assign P[50] = in[5] ^ in2[5];
    assign G[51] = in[4] & in2[4];
    assign P[51] = in[4] ^ in2[4];
    assign G[52] = in[3] & in2[3];
    assign P[52] = in[3] ^ in2[3];
    assign G[53] = in[2] & in2[2];
    assign P[53] = in[2] ^ in2[2];
    assign G[54] = in[1] & in2[1];
    assign P[54] = in[1] ^ in2[1];
    assign G[55] = in[0] & in2[0];
    assign P[55] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign C[55] = G[54] | (P[54] & C[54]);
    assign cout = G[55] | (P[55] & C[55]);
    assign sum = P ^ C;
endmodule

module CLA55(output [54:0] sum, output cout, input [54:0] in1, input [54:0] in2;

    wire[54:0] G;
    wire[54:0] C;
    wire[54:0] P;

    assign G[0] = in[54] & in2[54];
    assign P[0] = in[54] ^ in2[54];
    assign G[1] = in[53] & in2[53];
    assign P[1] = in[53] ^ in2[53];
    assign G[2] = in[52] & in2[52];
    assign P[2] = in[52] ^ in2[52];
    assign G[3] = in[51] & in2[51];
    assign P[3] = in[51] ^ in2[51];
    assign G[4] = in[50] & in2[50];
    assign P[4] = in[50] ^ in2[50];
    assign G[5] = in[49] & in2[49];
    assign P[5] = in[49] ^ in2[49];
    assign G[6] = in[48] & in2[48];
    assign P[6] = in[48] ^ in2[48];
    assign G[7] = in[47] & in2[47];
    assign P[7] = in[47] ^ in2[47];
    assign G[8] = in[46] & in2[46];
    assign P[8] = in[46] ^ in2[46];
    assign G[9] = in[45] & in2[45];
    assign P[9] = in[45] ^ in2[45];
    assign G[10] = in[44] & in2[44];
    assign P[10] = in[44] ^ in2[44];
    assign G[11] = in[43] & in2[43];
    assign P[11] = in[43] ^ in2[43];
    assign G[12] = in[42] & in2[42];
    assign P[12] = in[42] ^ in2[42];
    assign G[13] = in[41] & in2[41];
    assign P[13] = in[41] ^ in2[41];
    assign G[14] = in[40] & in2[40];
    assign P[14] = in[40] ^ in2[40];
    assign G[15] = in[39] & in2[39];
    assign P[15] = in[39] ^ in2[39];
    assign G[16] = in[38] & in2[38];
    assign P[16] = in[38] ^ in2[38];
    assign G[17] = in[37] & in2[37];
    assign P[17] = in[37] ^ in2[37];
    assign G[18] = in[36] & in2[36];
    assign P[18] = in[36] ^ in2[36];
    assign G[19] = in[35] & in2[35];
    assign P[19] = in[35] ^ in2[35];
    assign G[20] = in[34] & in2[34];
    assign P[20] = in[34] ^ in2[34];
    assign G[21] = in[33] & in2[33];
    assign P[21] = in[33] ^ in2[33];
    assign G[22] = in[32] & in2[32];
    assign P[22] = in[32] ^ in2[32];
    assign G[23] = in[31] & in2[31];
    assign P[23] = in[31] ^ in2[31];
    assign G[24] = in[30] & in2[30];
    assign P[24] = in[30] ^ in2[30];
    assign G[25] = in[29] & in2[29];
    assign P[25] = in[29] ^ in2[29];
    assign G[26] = in[28] & in2[28];
    assign P[26] = in[28] ^ in2[28];
    assign G[27] = in[27] & in2[27];
    assign P[27] = in[27] ^ in2[27];
    assign G[28] = in[26] & in2[26];
    assign P[28] = in[26] ^ in2[26];
    assign G[29] = in[25] & in2[25];
    assign P[29] = in[25] ^ in2[25];
    assign G[30] = in[24] & in2[24];
    assign P[30] = in[24] ^ in2[24];
    assign G[31] = in[23] & in2[23];
    assign P[31] = in[23] ^ in2[23];
    assign G[32] = in[22] & in2[22];
    assign P[32] = in[22] ^ in2[22];
    assign G[33] = in[21] & in2[21];
    assign P[33] = in[21] ^ in2[21];
    assign G[34] = in[20] & in2[20];
    assign P[34] = in[20] ^ in2[20];
    assign G[35] = in[19] & in2[19];
    assign P[35] = in[19] ^ in2[19];
    assign G[36] = in[18] & in2[18];
    assign P[36] = in[18] ^ in2[18];
    assign G[37] = in[17] & in2[17];
    assign P[37] = in[17] ^ in2[17];
    assign G[38] = in[16] & in2[16];
    assign P[38] = in[16] ^ in2[16];
    assign G[39] = in[15] & in2[15];
    assign P[39] = in[15] ^ in2[15];
    assign G[40] = in[14] & in2[14];
    assign P[40] = in[14] ^ in2[14];
    assign G[41] = in[13] & in2[13];
    assign P[41] = in[13] ^ in2[13];
    assign G[42] = in[12] & in2[12];
    assign P[42] = in[12] ^ in2[12];
    assign G[43] = in[11] & in2[11];
    assign P[43] = in[11] ^ in2[11];
    assign G[44] = in[10] & in2[10];
    assign P[44] = in[10] ^ in2[10];
    assign G[45] = in[9] & in2[9];
    assign P[45] = in[9] ^ in2[9];
    assign G[46] = in[8] & in2[8];
    assign P[46] = in[8] ^ in2[8];
    assign G[47] = in[7] & in2[7];
    assign P[47] = in[7] ^ in2[7];
    assign G[48] = in[6] & in2[6];
    assign P[48] = in[6] ^ in2[6];
    assign G[49] = in[5] & in2[5];
    assign P[49] = in[5] ^ in2[5];
    assign G[50] = in[4] & in2[4];
    assign P[50] = in[4] ^ in2[4];
    assign G[51] = in[3] & in2[3];
    assign P[51] = in[3] ^ in2[3];
    assign G[52] = in[2] & in2[2];
    assign P[52] = in[2] ^ in2[2];
    assign G[53] = in[1] & in2[1];
    assign P[53] = in[1] ^ in2[1];
    assign G[54] = in[0] & in2[0];
    assign P[54] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign C[54] = G[53] | (P[53] & C[53]);
    assign cout = G[54] | (P[54] & C[54]);
    assign sum = P ^ C;
endmodule

module CLA54(output [53:0] sum, output cout, input [53:0] in1, input [53:0] in2;

    wire[53:0] G;
    wire[53:0] C;
    wire[53:0] P;

    assign G[0] = in[53] & in2[53];
    assign P[0] = in[53] ^ in2[53];
    assign G[1] = in[52] & in2[52];
    assign P[1] = in[52] ^ in2[52];
    assign G[2] = in[51] & in2[51];
    assign P[2] = in[51] ^ in2[51];
    assign G[3] = in[50] & in2[50];
    assign P[3] = in[50] ^ in2[50];
    assign G[4] = in[49] & in2[49];
    assign P[4] = in[49] ^ in2[49];
    assign G[5] = in[48] & in2[48];
    assign P[5] = in[48] ^ in2[48];
    assign G[6] = in[47] & in2[47];
    assign P[6] = in[47] ^ in2[47];
    assign G[7] = in[46] & in2[46];
    assign P[7] = in[46] ^ in2[46];
    assign G[8] = in[45] & in2[45];
    assign P[8] = in[45] ^ in2[45];
    assign G[9] = in[44] & in2[44];
    assign P[9] = in[44] ^ in2[44];
    assign G[10] = in[43] & in2[43];
    assign P[10] = in[43] ^ in2[43];
    assign G[11] = in[42] & in2[42];
    assign P[11] = in[42] ^ in2[42];
    assign G[12] = in[41] & in2[41];
    assign P[12] = in[41] ^ in2[41];
    assign G[13] = in[40] & in2[40];
    assign P[13] = in[40] ^ in2[40];
    assign G[14] = in[39] & in2[39];
    assign P[14] = in[39] ^ in2[39];
    assign G[15] = in[38] & in2[38];
    assign P[15] = in[38] ^ in2[38];
    assign G[16] = in[37] & in2[37];
    assign P[16] = in[37] ^ in2[37];
    assign G[17] = in[36] & in2[36];
    assign P[17] = in[36] ^ in2[36];
    assign G[18] = in[35] & in2[35];
    assign P[18] = in[35] ^ in2[35];
    assign G[19] = in[34] & in2[34];
    assign P[19] = in[34] ^ in2[34];
    assign G[20] = in[33] & in2[33];
    assign P[20] = in[33] ^ in2[33];
    assign G[21] = in[32] & in2[32];
    assign P[21] = in[32] ^ in2[32];
    assign G[22] = in[31] & in2[31];
    assign P[22] = in[31] ^ in2[31];
    assign G[23] = in[30] & in2[30];
    assign P[23] = in[30] ^ in2[30];
    assign G[24] = in[29] & in2[29];
    assign P[24] = in[29] ^ in2[29];
    assign G[25] = in[28] & in2[28];
    assign P[25] = in[28] ^ in2[28];
    assign G[26] = in[27] & in2[27];
    assign P[26] = in[27] ^ in2[27];
    assign G[27] = in[26] & in2[26];
    assign P[27] = in[26] ^ in2[26];
    assign G[28] = in[25] & in2[25];
    assign P[28] = in[25] ^ in2[25];
    assign G[29] = in[24] & in2[24];
    assign P[29] = in[24] ^ in2[24];
    assign G[30] = in[23] & in2[23];
    assign P[30] = in[23] ^ in2[23];
    assign G[31] = in[22] & in2[22];
    assign P[31] = in[22] ^ in2[22];
    assign G[32] = in[21] & in2[21];
    assign P[32] = in[21] ^ in2[21];
    assign G[33] = in[20] & in2[20];
    assign P[33] = in[20] ^ in2[20];
    assign G[34] = in[19] & in2[19];
    assign P[34] = in[19] ^ in2[19];
    assign G[35] = in[18] & in2[18];
    assign P[35] = in[18] ^ in2[18];
    assign G[36] = in[17] & in2[17];
    assign P[36] = in[17] ^ in2[17];
    assign G[37] = in[16] & in2[16];
    assign P[37] = in[16] ^ in2[16];
    assign G[38] = in[15] & in2[15];
    assign P[38] = in[15] ^ in2[15];
    assign G[39] = in[14] & in2[14];
    assign P[39] = in[14] ^ in2[14];
    assign G[40] = in[13] & in2[13];
    assign P[40] = in[13] ^ in2[13];
    assign G[41] = in[12] & in2[12];
    assign P[41] = in[12] ^ in2[12];
    assign G[42] = in[11] & in2[11];
    assign P[42] = in[11] ^ in2[11];
    assign G[43] = in[10] & in2[10];
    assign P[43] = in[10] ^ in2[10];
    assign G[44] = in[9] & in2[9];
    assign P[44] = in[9] ^ in2[9];
    assign G[45] = in[8] & in2[8];
    assign P[45] = in[8] ^ in2[8];
    assign G[46] = in[7] & in2[7];
    assign P[46] = in[7] ^ in2[7];
    assign G[47] = in[6] & in2[6];
    assign P[47] = in[6] ^ in2[6];
    assign G[48] = in[5] & in2[5];
    assign P[48] = in[5] ^ in2[5];
    assign G[49] = in[4] & in2[4];
    assign P[49] = in[4] ^ in2[4];
    assign G[50] = in[3] & in2[3];
    assign P[50] = in[3] ^ in2[3];
    assign G[51] = in[2] & in2[2];
    assign P[51] = in[2] ^ in2[2];
    assign G[52] = in[1] & in2[1];
    assign P[52] = in[1] ^ in2[1];
    assign G[53] = in[0] & in2[0];
    assign P[53] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign C[53] = G[52] | (P[52] & C[52]);
    assign cout = G[53] | (P[53] & C[53]);
    assign sum = P ^ C;
endmodule

module CLA53(output [52:0] sum, output cout, input [52:0] in1, input [52:0] in2;

    wire[52:0] G;
    wire[52:0] C;
    wire[52:0] P;

    assign G[0] = in[52] & in2[52];
    assign P[0] = in[52] ^ in2[52];
    assign G[1] = in[51] & in2[51];
    assign P[1] = in[51] ^ in2[51];
    assign G[2] = in[50] & in2[50];
    assign P[2] = in[50] ^ in2[50];
    assign G[3] = in[49] & in2[49];
    assign P[3] = in[49] ^ in2[49];
    assign G[4] = in[48] & in2[48];
    assign P[4] = in[48] ^ in2[48];
    assign G[5] = in[47] & in2[47];
    assign P[5] = in[47] ^ in2[47];
    assign G[6] = in[46] & in2[46];
    assign P[6] = in[46] ^ in2[46];
    assign G[7] = in[45] & in2[45];
    assign P[7] = in[45] ^ in2[45];
    assign G[8] = in[44] & in2[44];
    assign P[8] = in[44] ^ in2[44];
    assign G[9] = in[43] & in2[43];
    assign P[9] = in[43] ^ in2[43];
    assign G[10] = in[42] & in2[42];
    assign P[10] = in[42] ^ in2[42];
    assign G[11] = in[41] & in2[41];
    assign P[11] = in[41] ^ in2[41];
    assign G[12] = in[40] & in2[40];
    assign P[12] = in[40] ^ in2[40];
    assign G[13] = in[39] & in2[39];
    assign P[13] = in[39] ^ in2[39];
    assign G[14] = in[38] & in2[38];
    assign P[14] = in[38] ^ in2[38];
    assign G[15] = in[37] & in2[37];
    assign P[15] = in[37] ^ in2[37];
    assign G[16] = in[36] & in2[36];
    assign P[16] = in[36] ^ in2[36];
    assign G[17] = in[35] & in2[35];
    assign P[17] = in[35] ^ in2[35];
    assign G[18] = in[34] & in2[34];
    assign P[18] = in[34] ^ in2[34];
    assign G[19] = in[33] & in2[33];
    assign P[19] = in[33] ^ in2[33];
    assign G[20] = in[32] & in2[32];
    assign P[20] = in[32] ^ in2[32];
    assign G[21] = in[31] & in2[31];
    assign P[21] = in[31] ^ in2[31];
    assign G[22] = in[30] & in2[30];
    assign P[22] = in[30] ^ in2[30];
    assign G[23] = in[29] & in2[29];
    assign P[23] = in[29] ^ in2[29];
    assign G[24] = in[28] & in2[28];
    assign P[24] = in[28] ^ in2[28];
    assign G[25] = in[27] & in2[27];
    assign P[25] = in[27] ^ in2[27];
    assign G[26] = in[26] & in2[26];
    assign P[26] = in[26] ^ in2[26];
    assign G[27] = in[25] & in2[25];
    assign P[27] = in[25] ^ in2[25];
    assign G[28] = in[24] & in2[24];
    assign P[28] = in[24] ^ in2[24];
    assign G[29] = in[23] & in2[23];
    assign P[29] = in[23] ^ in2[23];
    assign G[30] = in[22] & in2[22];
    assign P[30] = in[22] ^ in2[22];
    assign G[31] = in[21] & in2[21];
    assign P[31] = in[21] ^ in2[21];
    assign G[32] = in[20] & in2[20];
    assign P[32] = in[20] ^ in2[20];
    assign G[33] = in[19] & in2[19];
    assign P[33] = in[19] ^ in2[19];
    assign G[34] = in[18] & in2[18];
    assign P[34] = in[18] ^ in2[18];
    assign G[35] = in[17] & in2[17];
    assign P[35] = in[17] ^ in2[17];
    assign G[36] = in[16] & in2[16];
    assign P[36] = in[16] ^ in2[16];
    assign G[37] = in[15] & in2[15];
    assign P[37] = in[15] ^ in2[15];
    assign G[38] = in[14] & in2[14];
    assign P[38] = in[14] ^ in2[14];
    assign G[39] = in[13] & in2[13];
    assign P[39] = in[13] ^ in2[13];
    assign G[40] = in[12] & in2[12];
    assign P[40] = in[12] ^ in2[12];
    assign G[41] = in[11] & in2[11];
    assign P[41] = in[11] ^ in2[11];
    assign G[42] = in[10] & in2[10];
    assign P[42] = in[10] ^ in2[10];
    assign G[43] = in[9] & in2[9];
    assign P[43] = in[9] ^ in2[9];
    assign G[44] = in[8] & in2[8];
    assign P[44] = in[8] ^ in2[8];
    assign G[45] = in[7] & in2[7];
    assign P[45] = in[7] ^ in2[7];
    assign G[46] = in[6] & in2[6];
    assign P[46] = in[6] ^ in2[6];
    assign G[47] = in[5] & in2[5];
    assign P[47] = in[5] ^ in2[5];
    assign G[48] = in[4] & in2[4];
    assign P[48] = in[4] ^ in2[4];
    assign G[49] = in[3] & in2[3];
    assign P[49] = in[3] ^ in2[3];
    assign G[50] = in[2] & in2[2];
    assign P[50] = in[2] ^ in2[2];
    assign G[51] = in[1] & in2[1];
    assign P[51] = in[1] ^ in2[1];
    assign G[52] = in[0] & in2[0];
    assign P[52] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign C[52] = G[51] | (P[51] & C[51]);
    assign cout = G[52] | (P[52] & C[52]);
    assign sum = P ^ C;
endmodule

module CLA52(output [51:0] sum, output cout, input [51:0] in1, input [51:0] in2;

    wire[51:0] G;
    wire[51:0] C;
    wire[51:0] P;

    assign G[0] = in[51] & in2[51];
    assign P[0] = in[51] ^ in2[51];
    assign G[1] = in[50] & in2[50];
    assign P[1] = in[50] ^ in2[50];
    assign G[2] = in[49] & in2[49];
    assign P[2] = in[49] ^ in2[49];
    assign G[3] = in[48] & in2[48];
    assign P[3] = in[48] ^ in2[48];
    assign G[4] = in[47] & in2[47];
    assign P[4] = in[47] ^ in2[47];
    assign G[5] = in[46] & in2[46];
    assign P[5] = in[46] ^ in2[46];
    assign G[6] = in[45] & in2[45];
    assign P[6] = in[45] ^ in2[45];
    assign G[7] = in[44] & in2[44];
    assign P[7] = in[44] ^ in2[44];
    assign G[8] = in[43] & in2[43];
    assign P[8] = in[43] ^ in2[43];
    assign G[9] = in[42] & in2[42];
    assign P[9] = in[42] ^ in2[42];
    assign G[10] = in[41] & in2[41];
    assign P[10] = in[41] ^ in2[41];
    assign G[11] = in[40] & in2[40];
    assign P[11] = in[40] ^ in2[40];
    assign G[12] = in[39] & in2[39];
    assign P[12] = in[39] ^ in2[39];
    assign G[13] = in[38] & in2[38];
    assign P[13] = in[38] ^ in2[38];
    assign G[14] = in[37] & in2[37];
    assign P[14] = in[37] ^ in2[37];
    assign G[15] = in[36] & in2[36];
    assign P[15] = in[36] ^ in2[36];
    assign G[16] = in[35] & in2[35];
    assign P[16] = in[35] ^ in2[35];
    assign G[17] = in[34] & in2[34];
    assign P[17] = in[34] ^ in2[34];
    assign G[18] = in[33] & in2[33];
    assign P[18] = in[33] ^ in2[33];
    assign G[19] = in[32] & in2[32];
    assign P[19] = in[32] ^ in2[32];
    assign G[20] = in[31] & in2[31];
    assign P[20] = in[31] ^ in2[31];
    assign G[21] = in[30] & in2[30];
    assign P[21] = in[30] ^ in2[30];
    assign G[22] = in[29] & in2[29];
    assign P[22] = in[29] ^ in2[29];
    assign G[23] = in[28] & in2[28];
    assign P[23] = in[28] ^ in2[28];
    assign G[24] = in[27] & in2[27];
    assign P[24] = in[27] ^ in2[27];
    assign G[25] = in[26] & in2[26];
    assign P[25] = in[26] ^ in2[26];
    assign G[26] = in[25] & in2[25];
    assign P[26] = in[25] ^ in2[25];
    assign G[27] = in[24] & in2[24];
    assign P[27] = in[24] ^ in2[24];
    assign G[28] = in[23] & in2[23];
    assign P[28] = in[23] ^ in2[23];
    assign G[29] = in[22] & in2[22];
    assign P[29] = in[22] ^ in2[22];
    assign G[30] = in[21] & in2[21];
    assign P[30] = in[21] ^ in2[21];
    assign G[31] = in[20] & in2[20];
    assign P[31] = in[20] ^ in2[20];
    assign G[32] = in[19] & in2[19];
    assign P[32] = in[19] ^ in2[19];
    assign G[33] = in[18] & in2[18];
    assign P[33] = in[18] ^ in2[18];
    assign G[34] = in[17] & in2[17];
    assign P[34] = in[17] ^ in2[17];
    assign G[35] = in[16] & in2[16];
    assign P[35] = in[16] ^ in2[16];
    assign G[36] = in[15] & in2[15];
    assign P[36] = in[15] ^ in2[15];
    assign G[37] = in[14] & in2[14];
    assign P[37] = in[14] ^ in2[14];
    assign G[38] = in[13] & in2[13];
    assign P[38] = in[13] ^ in2[13];
    assign G[39] = in[12] & in2[12];
    assign P[39] = in[12] ^ in2[12];
    assign G[40] = in[11] & in2[11];
    assign P[40] = in[11] ^ in2[11];
    assign G[41] = in[10] & in2[10];
    assign P[41] = in[10] ^ in2[10];
    assign G[42] = in[9] & in2[9];
    assign P[42] = in[9] ^ in2[9];
    assign G[43] = in[8] & in2[8];
    assign P[43] = in[8] ^ in2[8];
    assign G[44] = in[7] & in2[7];
    assign P[44] = in[7] ^ in2[7];
    assign G[45] = in[6] & in2[6];
    assign P[45] = in[6] ^ in2[6];
    assign G[46] = in[5] & in2[5];
    assign P[46] = in[5] ^ in2[5];
    assign G[47] = in[4] & in2[4];
    assign P[47] = in[4] ^ in2[4];
    assign G[48] = in[3] & in2[3];
    assign P[48] = in[3] ^ in2[3];
    assign G[49] = in[2] & in2[2];
    assign P[49] = in[2] ^ in2[2];
    assign G[50] = in[1] & in2[1];
    assign P[50] = in[1] ^ in2[1];
    assign G[51] = in[0] & in2[0];
    assign P[51] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign C[51] = G[50] | (P[50] & C[50]);
    assign cout = G[51] | (P[51] & C[51]);
    assign sum = P ^ C;
endmodule

module CLA51(output [50:0] sum, output cout, input [50:0] in1, input [50:0] in2;

    wire[50:0] G;
    wire[50:0] C;
    wire[50:0] P;

    assign G[0] = in[50] & in2[50];
    assign P[0] = in[50] ^ in2[50];
    assign G[1] = in[49] & in2[49];
    assign P[1] = in[49] ^ in2[49];
    assign G[2] = in[48] & in2[48];
    assign P[2] = in[48] ^ in2[48];
    assign G[3] = in[47] & in2[47];
    assign P[3] = in[47] ^ in2[47];
    assign G[4] = in[46] & in2[46];
    assign P[4] = in[46] ^ in2[46];
    assign G[5] = in[45] & in2[45];
    assign P[5] = in[45] ^ in2[45];
    assign G[6] = in[44] & in2[44];
    assign P[6] = in[44] ^ in2[44];
    assign G[7] = in[43] & in2[43];
    assign P[7] = in[43] ^ in2[43];
    assign G[8] = in[42] & in2[42];
    assign P[8] = in[42] ^ in2[42];
    assign G[9] = in[41] & in2[41];
    assign P[9] = in[41] ^ in2[41];
    assign G[10] = in[40] & in2[40];
    assign P[10] = in[40] ^ in2[40];
    assign G[11] = in[39] & in2[39];
    assign P[11] = in[39] ^ in2[39];
    assign G[12] = in[38] & in2[38];
    assign P[12] = in[38] ^ in2[38];
    assign G[13] = in[37] & in2[37];
    assign P[13] = in[37] ^ in2[37];
    assign G[14] = in[36] & in2[36];
    assign P[14] = in[36] ^ in2[36];
    assign G[15] = in[35] & in2[35];
    assign P[15] = in[35] ^ in2[35];
    assign G[16] = in[34] & in2[34];
    assign P[16] = in[34] ^ in2[34];
    assign G[17] = in[33] & in2[33];
    assign P[17] = in[33] ^ in2[33];
    assign G[18] = in[32] & in2[32];
    assign P[18] = in[32] ^ in2[32];
    assign G[19] = in[31] & in2[31];
    assign P[19] = in[31] ^ in2[31];
    assign G[20] = in[30] & in2[30];
    assign P[20] = in[30] ^ in2[30];
    assign G[21] = in[29] & in2[29];
    assign P[21] = in[29] ^ in2[29];
    assign G[22] = in[28] & in2[28];
    assign P[22] = in[28] ^ in2[28];
    assign G[23] = in[27] & in2[27];
    assign P[23] = in[27] ^ in2[27];
    assign G[24] = in[26] & in2[26];
    assign P[24] = in[26] ^ in2[26];
    assign G[25] = in[25] & in2[25];
    assign P[25] = in[25] ^ in2[25];
    assign G[26] = in[24] & in2[24];
    assign P[26] = in[24] ^ in2[24];
    assign G[27] = in[23] & in2[23];
    assign P[27] = in[23] ^ in2[23];
    assign G[28] = in[22] & in2[22];
    assign P[28] = in[22] ^ in2[22];
    assign G[29] = in[21] & in2[21];
    assign P[29] = in[21] ^ in2[21];
    assign G[30] = in[20] & in2[20];
    assign P[30] = in[20] ^ in2[20];
    assign G[31] = in[19] & in2[19];
    assign P[31] = in[19] ^ in2[19];
    assign G[32] = in[18] & in2[18];
    assign P[32] = in[18] ^ in2[18];
    assign G[33] = in[17] & in2[17];
    assign P[33] = in[17] ^ in2[17];
    assign G[34] = in[16] & in2[16];
    assign P[34] = in[16] ^ in2[16];
    assign G[35] = in[15] & in2[15];
    assign P[35] = in[15] ^ in2[15];
    assign G[36] = in[14] & in2[14];
    assign P[36] = in[14] ^ in2[14];
    assign G[37] = in[13] & in2[13];
    assign P[37] = in[13] ^ in2[13];
    assign G[38] = in[12] & in2[12];
    assign P[38] = in[12] ^ in2[12];
    assign G[39] = in[11] & in2[11];
    assign P[39] = in[11] ^ in2[11];
    assign G[40] = in[10] & in2[10];
    assign P[40] = in[10] ^ in2[10];
    assign G[41] = in[9] & in2[9];
    assign P[41] = in[9] ^ in2[9];
    assign G[42] = in[8] & in2[8];
    assign P[42] = in[8] ^ in2[8];
    assign G[43] = in[7] & in2[7];
    assign P[43] = in[7] ^ in2[7];
    assign G[44] = in[6] & in2[6];
    assign P[44] = in[6] ^ in2[6];
    assign G[45] = in[5] & in2[5];
    assign P[45] = in[5] ^ in2[5];
    assign G[46] = in[4] & in2[4];
    assign P[46] = in[4] ^ in2[4];
    assign G[47] = in[3] & in2[3];
    assign P[47] = in[3] ^ in2[3];
    assign G[48] = in[2] & in2[2];
    assign P[48] = in[2] ^ in2[2];
    assign G[49] = in[1] & in2[1];
    assign P[49] = in[1] ^ in2[1];
    assign G[50] = in[0] & in2[0];
    assign P[50] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign C[50] = G[49] | (P[49] & C[49]);
    assign cout = G[50] | (P[50] & C[50]);
    assign sum = P ^ C;
endmodule

module CLA50(output [49:0] sum, output cout, input [49:0] in1, input [49:0] in2;

    wire[49:0] G;
    wire[49:0] C;
    wire[49:0] P;

    assign G[0] = in[49] & in2[49];
    assign P[0] = in[49] ^ in2[49];
    assign G[1] = in[48] & in2[48];
    assign P[1] = in[48] ^ in2[48];
    assign G[2] = in[47] & in2[47];
    assign P[2] = in[47] ^ in2[47];
    assign G[3] = in[46] & in2[46];
    assign P[3] = in[46] ^ in2[46];
    assign G[4] = in[45] & in2[45];
    assign P[4] = in[45] ^ in2[45];
    assign G[5] = in[44] & in2[44];
    assign P[5] = in[44] ^ in2[44];
    assign G[6] = in[43] & in2[43];
    assign P[6] = in[43] ^ in2[43];
    assign G[7] = in[42] & in2[42];
    assign P[7] = in[42] ^ in2[42];
    assign G[8] = in[41] & in2[41];
    assign P[8] = in[41] ^ in2[41];
    assign G[9] = in[40] & in2[40];
    assign P[9] = in[40] ^ in2[40];
    assign G[10] = in[39] & in2[39];
    assign P[10] = in[39] ^ in2[39];
    assign G[11] = in[38] & in2[38];
    assign P[11] = in[38] ^ in2[38];
    assign G[12] = in[37] & in2[37];
    assign P[12] = in[37] ^ in2[37];
    assign G[13] = in[36] & in2[36];
    assign P[13] = in[36] ^ in2[36];
    assign G[14] = in[35] & in2[35];
    assign P[14] = in[35] ^ in2[35];
    assign G[15] = in[34] & in2[34];
    assign P[15] = in[34] ^ in2[34];
    assign G[16] = in[33] & in2[33];
    assign P[16] = in[33] ^ in2[33];
    assign G[17] = in[32] & in2[32];
    assign P[17] = in[32] ^ in2[32];
    assign G[18] = in[31] & in2[31];
    assign P[18] = in[31] ^ in2[31];
    assign G[19] = in[30] & in2[30];
    assign P[19] = in[30] ^ in2[30];
    assign G[20] = in[29] & in2[29];
    assign P[20] = in[29] ^ in2[29];
    assign G[21] = in[28] & in2[28];
    assign P[21] = in[28] ^ in2[28];
    assign G[22] = in[27] & in2[27];
    assign P[22] = in[27] ^ in2[27];
    assign G[23] = in[26] & in2[26];
    assign P[23] = in[26] ^ in2[26];
    assign G[24] = in[25] & in2[25];
    assign P[24] = in[25] ^ in2[25];
    assign G[25] = in[24] & in2[24];
    assign P[25] = in[24] ^ in2[24];
    assign G[26] = in[23] & in2[23];
    assign P[26] = in[23] ^ in2[23];
    assign G[27] = in[22] & in2[22];
    assign P[27] = in[22] ^ in2[22];
    assign G[28] = in[21] & in2[21];
    assign P[28] = in[21] ^ in2[21];
    assign G[29] = in[20] & in2[20];
    assign P[29] = in[20] ^ in2[20];
    assign G[30] = in[19] & in2[19];
    assign P[30] = in[19] ^ in2[19];
    assign G[31] = in[18] & in2[18];
    assign P[31] = in[18] ^ in2[18];
    assign G[32] = in[17] & in2[17];
    assign P[32] = in[17] ^ in2[17];
    assign G[33] = in[16] & in2[16];
    assign P[33] = in[16] ^ in2[16];
    assign G[34] = in[15] & in2[15];
    assign P[34] = in[15] ^ in2[15];
    assign G[35] = in[14] & in2[14];
    assign P[35] = in[14] ^ in2[14];
    assign G[36] = in[13] & in2[13];
    assign P[36] = in[13] ^ in2[13];
    assign G[37] = in[12] & in2[12];
    assign P[37] = in[12] ^ in2[12];
    assign G[38] = in[11] & in2[11];
    assign P[38] = in[11] ^ in2[11];
    assign G[39] = in[10] & in2[10];
    assign P[39] = in[10] ^ in2[10];
    assign G[40] = in[9] & in2[9];
    assign P[40] = in[9] ^ in2[9];
    assign G[41] = in[8] & in2[8];
    assign P[41] = in[8] ^ in2[8];
    assign G[42] = in[7] & in2[7];
    assign P[42] = in[7] ^ in2[7];
    assign G[43] = in[6] & in2[6];
    assign P[43] = in[6] ^ in2[6];
    assign G[44] = in[5] & in2[5];
    assign P[44] = in[5] ^ in2[5];
    assign G[45] = in[4] & in2[4];
    assign P[45] = in[4] ^ in2[4];
    assign G[46] = in[3] & in2[3];
    assign P[46] = in[3] ^ in2[3];
    assign G[47] = in[2] & in2[2];
    assign P[47] = in[2] ^ in2[2];
    assign G[48] = in[1] & in2[1];
    assign P[48] = in[1] ^ in2[1];
    assign G[49] = in[0] & in2[0];
    assign P[49] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign C[49] = G[48] | (P[48] & C[48]);
    assign cout = G[49] | (P[49] & C[49]);
    assign sum = P ^ C;
endmodule

module CLA49(output [48:0] sum, output cout, input [48:0] in1, input [48:0] in2;

    wire[48:0] G;
    wire[48:0] C;
    wire[48:0] P;

    assign G[0] = in[48] & in2[48];
    assign P[0] = in[48] ^ in2[48];
    assign G[1] = in[47] & in2[47];
    assign P[1] = in[47] ^ in2[47];
    assign G[2] = in[46] & in2[46];
    assign P[2] = in[46] ^ in2[46];
    assign G[3] = in[45] & in2[45];
    assign P[3] = in[45] ^ in2[45];
    assign G[4] = in[44] & in2[44];
    assign P[4] = in[44] ^ in2[44];
    assign G[5] = in[43] & in2[43];
    assign P[5] = in[43] ^ in2[43];
    assign G[6] = in[42] & in2[42];
    assign P[6] = in[42] ^ in2[42];
    assign G[7] = in[41] & in2[41];
    assign P[7] = in[41] ^ in2[41];
    assign G[8] = in[40] & in2[40];
    assign P[8] = in[40] ^ in2[40];
    assign G[9] = in[39] & in2[39];
    assign P[9] = in[39] ^ in2[39];
    assign G[10] = in[38] & in2[38];
    assign P[10] = in[38] ^ in2[38];
    assign G[11] = in[37] & in2[37];
    assign P[11] = in[37] ^ in2[37];
    assign G[12] = in[36] & in2[36];
    assign P[12] = in[36] ^ in2[36];
    assign G[13] = in[35] & in2[35];
    assign P[13] = in[35] ^ in2[35];
    assign G[14] = in[34] & in2[34];
    assign P[14] = in[34] ^ in2[34];
    assign G[15] = in[33] & in2[33];
    assign P[15] = in[33] ^ in2[33];
    assign G[16] = in[32] & in2[32];
    assign P[16] = in[32] ^ in2[32];
    assign G[17] = in[31] & in2[31];
    assign P[17] = in[31] ^ in2[31];
    assign G[18] = in[30] & in2[30];
    assign P[18] = in[30] ^ in2[30];
    assign G[19] = in[29] & in2[29];
    assign P[19] = in[29] ^ in2[29];
    assign G[20] = in[28] & in2[28];
    assign P[20] = in[28] ^ in2[28];
    assign G[21] = in[27] & in2[27];
    assign P[21] = in[27] ^ in2[27];
    assign G[22] = in[26] & in2[26];
    assign P[22] = in[26] ^ in2[26];
    assign G[23] = in[25] & in2[25];
    assign P[23] = in[25] ^ in2[25];
    assign G[24] = in[24] & in2[24];
    assign P[24] = in[24] ^ in2[24];
    assign G[25] = in[23] & in2[23];
    assign P[25] = in[23] ^ in2[23];
    assign G[26] = in[22] & in2[22];
    assign P[26] = in[22] ^ in2[22];
    assign G[27] = in[21] & in2[21];
    assign P[27] = in[21] ^ in2[21];
    assign G[28] = in[20] & in2[20];
    assign P[28] = in[20] ^ in2[20];
    assign G[29] = in[19] & in2[19];
    assign P[29] = in[19] ^ in2[19];
    assign G[30] = in[18] & in2[18];
    assign P[30] = in[18] ^ in2[18];
    assign G[31] = in[17] & in2[17];
    assign P[31] = in[17] ^ in2[17];
    assign G[32] = in[16] & in2[16];
    assign P[32] = in[16] ^ in2[16];
    assign G[33] = in[15] & in2[15];
    assign P[33] = in[15] ^ in2[15];
    assign G[34] = in[14] & in2[14];
    assign P[34] = in[14] ^ in2[14];
    assign G[35] = in[13] & in2[13];
    assign P[35] = in[13] ^ in2[13];
    assign G[36] = in[12] & in2[12];
    assign P[36] = in[12] ^ in2[12];
    assign G[37] = in[11] & in2[11];
    assign P[37] = in[11] ^ in2[11];
    assign G[38] = in[10] & in2[10];
    assign P[38] = in[10] ^ in2[10];
    assign G[39] = in[9] & in2[9];
    assign P[39] = in[9] ^ in2[9];
    assign G[40] = in[8] & in2[8];
    assign P[40] = in[8] ^ in2[8];
    assign G[41] = in[7] & in2[7];
    assign P[41] = in[7] ^ in2[7];
    assign G[42] = in[6] & in2[6];
    assign P[42] = in[6] ^ in2[6];
    assign G[43] = in[5] & in2[5];
    assign P[43] = in[5] ^ in2[5];
    assign G[44] = in[4] & in2[4];
    assign P[44] = in[4] ^ in2[4];
    assign G[45] = in[3] & in2[3];
    assign P[45] = in[3] ^ in2[3];
    assign G[46] = in[2] & in2[2];
    assign P[46] = in[2] ^ in2[2];
    assign G[47] = in[1] & in2[1];
    assign P[47] = in[1] ^ in2[1];
    assign G[48] = in[0] & in2[0];
    assign P[48] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign C[48] = G[47] | (P[47] & C[47]);
    assign cout = G[48] | (P[48] & C[48]);
    assign sum = P ^ C;
endmodule

module CLA48(output [47:0] sum, output cout, input [47:0] in1, input [47:0] in2;

    wire[47:0] G;
    wire[47:0] C;
    wire[47:0] P;

    assign G[0] = in[47] & in2[47];
    assign P[0] = in[47] ^ in2[47];
    assign G[1] = in[46] & in2[46];
    assign P[1] = in[46] ^ in2[46];
    assign G[2] = in[45] & in2[45];
    assign P[2] = in[45] ^ in2[45];
    assign G[3] = in[44] & in2[44];
    assign P[3] = in[44] ^ in2[44];
    assign G[4] = in[43] & in2[43];
    assign P[4] = in[43] ^ in2[43];
    assign G[5] = in[42] & in2[42];
    assign P[5] = in[42] ^ in2[42];
    assign G[6] = in[41] & in2[41];
    assign P[6] = in[41] ^ in2[41];
    assign G[7] = in[40] & in2[40];
    assign P[7] = in[40] ^ in2[40];
    assign G[8] = in[39] & in2[39];
    assign P[8] = in[39] ^ in2[39];
    assign G[9] = in[38] & in2[38];
    assign P[9] = in[38] ^ in2[38];
    assign G[10] = in[37] & in2[37];
    assign P[10] = in[37] ^ in2[37];
    assign G[11] = in[36] & in2[36];
    assign P[11] = in[36] ^ in2[36];
    assign G[12] = in[35] & in2[35];
    assign P[12] = in[35] ^ in2[35];
    assign G[13] = in[34] & in2[34];
    assign P[13] = in[34] ^ in2[34];
    assign G[14] = in[33] & in2[33];
    assign P[14] = in[33] ^ in2[33];
    assign G[15] = in[32] & in2[32];
    assign P[15] = in[32] ^ in2[32];
    assign G[16] = in[31] & in2[31];
    assign P[16] = in[31] ^ in2[31];
    assign G[17] = in[30] & in2[30];
    assign P[17] = in[30] ^ in2[30];
    assign G[18] = in[29] & in2[29];
    assign P[18] = in[29] ^ in2[29];
    assign G[19] = in[28] & in2[28];
    assign P[19] = in[28] ^ in2[28];
    assign G[20] = in[27] & in2[27];
    assign P[20] = in[27] ^ in2[27];
    assign G[21] = in[26] & in2[26];
    assign P[21] = in[26] ^ in2[26];
    assign G[22] = in[25] & in2[25];
    assign P[22] = in[25] ^ in2[25];
    assign G[23] = in[24] & in2[24];
    assign P[23] = in[24] ^ in2[24];
    assign G[24] = in[23] & in2[23];
    assign P[24] = in[23] ^ in2[23];
    assign G[25] = in[22] & in2[22];
    assign P[25] = in[22] ^ in2[22];
    assign G[26] = in[21] & in2[21];
    assign P[26] = in[21] ^ in2[21];
    assign G[27] = in[20] & in2[20];
    assign P[27] = in[20] ^ in2[20];
    assign G[28] = in[19] & in2[19];
    assign P[28] = in[19] ^ in2[19];
    assign G[29] = in[18] & in2[18];
    assign P[29] = in[18] ^ in2[18];
    assign G[30] = in[17] & in2[17];
    assign P[30] = in[17] ^ in2[17];
    assign G[31] = in[16] & in2[16];
    assign P[31] = in[16] ^ in2[16];
    assign G[32] = in[15] & in2[15];
    assign P[32] = in[15] ^ in2[15];
    assign G[33] = in[14] & in2[14];
    assign P[33] = in[14] ^ in2[14];
    assign G[34] = in[13] & in2[13];
    assign P[34] = in[13] ^ in2[13];
    assign G[35] = in[12] & in2[12];
    assign P[35] = in[12] ^ in2[12];
    assign G[36] = in[11] & in2[11];
    assign P[36] = in[11] ^ in2[11];
    assign G[37] = in[10] & in2[10];
    assign P[37] = in[10] ^ in2[10];
    assign G[38] = in[9] & in2[9];
    assign P[38] = in[9] ^ in2[9];
    assign G[39] = in[8] & in2[8];
    assign P[39] = in[8] ^ in2[8];
    assign G[40] = in[7] & in2[7];
    assign P[40] = in[7] ^ in2[7];
    assign G[41] = in[6] & in2[6];
    assign P[41] = in[6] ^ in2[6];
    assign G[42] = in[5] & in2[5];
    assign P[42] = in[5] ^ in2[5];
    assign G[43] = in[4] & in2[4];
    assign P[43] = in[4] ^ in2[4];
    assign G[44] = in[3] & in2[3];
    assign P[44] = in[3] ^ in2[3];
    assign G[45] = in[2] & in2[2];
    assign P[45] = in[2] ^ in2[2];
    assign G[46] = in[1] & in2[1];
    assign P[46] = in[1] ^ in2[1];
    assign G[47] = in[0] & in2[0];
    assign P[47] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign C[47] = G[46] | (P[46] & C[46]);
    assign cout = G[47] | (P[47] & C[47]);
    assign sum = P ^ C;
endmodule

module CLA47(output [46:0] sum, output cout, input [46:0] in1, input [46:0] in2;

    wire[46:0] G;
    wire[46:0] C;
    wire[46:0] P;

    assign G[0] = in[46] & in2[46];
    assign P[0] = in[46] ^ in2[46];
    assign G[1] = in[45] & in2[45];
    assign P[1] = in[45] ^ in2[45];
    assign G[2] = in[44] & in2[44];
    assign P[2] = in[44] ^ in2[44];
    assign G[3] = in[43] & in2[43];
    assign P[3] = in[43] ^ in2[43];
    assign G[4] = in[42] & in2[42];
    assign P[4] = in[42] ^ in2[42];
    assign G[5] = in[41] & in2[41];
    assign P[5] = in[41] ^ in2[41];
    assign G[6] = in[40] & in2[40];
    assign P[6] = in[40] ^ in2[40];
    assign G[7] = in[39] & in2[39];
    assign P[7] = in[39] ^ in2[39];
    assign G[8] = in[38] & in2[38];
    assign P[8] = in[38] ^ in2[38];
    assign G[9] = in[37] & in2[37];
    assign P[9] = in[37] ^ in2[37];
    assign G[10] = in[36] & in2[36];
    assign P[10] = in[36] ^ in2[36];
    assign G[11] = in[35] & in2[35];
    assign P[11] = in[35] ^ in2[35];
    assign G[12] = in[34] & in2[34];
    assign P[12] = in[34] ^ in2[34];
    assign G[13] = in[33] & in2[33];
    assign P[13] = in[33] ^ in2[33];
    assign G[14] = in[32] & in2[32];
    assign P[14] = in[32] ^ in2[32];
    assign G[15] = in[31] & in2[31];
    assign P[15] = in[31] ^ in2[31];
    assign G[16] = in[30] & in2[30];
    assign P[16] = in[30] ^ in2[30];
    assign G[17] = in[29] & in2[29];
    assign P[17] = in[29] ^ in2[29];
    assign G[18] = in[28] & in2[28];
    assign P[18] = in[28] ^ in2[28];
    assign G[19] = in[27] & in2[27];
    assign P[19] = in[27] ^ in2[27];
    assign G[20] = in[26] & in2[26];
    assign P[20] = in[26] ^ in2[26];
    assign G[21] = in[25] & in2[25];
    assign P[21] = in[25] ^ in2[25];
    assign G[22] = in[24] & in2[24];
    assign P[22] = in[24] ^ in2[24];
    assign G[23] = in[23] & in2[23];
    assign P[23] = in[23] ^ in2[23];
    assign G[24] = in[22] & in2[22];
    assign P[24] = in[22] ^ in2[22];
    assign G[25] = in[21] & in2[21];
    assign P[25] = in[21] ^ in2[21];
    assign G[26] = in[20] & in2[20];
    assign P[26] = in[20] ^ in2[20];
    assign G[27] = in[19] & in2[19];
    assign P[27] = in[19] ^ in2[19];
    assign G[28] = in[18] & in2[18];
    assign P[28] = in[18] ^ in2[18];
    assign G[29] = in[17] & in2[17];
    assign P[29] = in[17] ^ in2[17];
    assign G[30] = in[16] & in2[16];
    assign P[30] = in[16] ^ in2[16];
    assign G[31] = in[15] & in2[15];
    assign P[31] = in[15] ^ in2[15];
    assign G[32] = in[14] & in2[14];
    assign P[32] = in[14] ^ in2[14];
    assign G[33] = in[13] & in2[13];
    assign P[33] = in[13] ^ in2[13];
    assign G[34] = in[12] & in2[12];
    assign P[34] = in[12] ^ in2[12];
    assign G[35] = in[11] & in2[11];
    assign P[35] = in[11] ^ in2[11];
    assign G[36] = in[10] & in2[10];
    assign P[36] = in[10] ^ in2[10];
    assign G[37] = in[9] & in2[9];
    assign P[37] = in[9] ^ in2[9];
    assign G[38] = in[8] & in2[8];
    assign P[38] = in[8] ^ in2[8];
    assign G[39] = in[7] & in2[7];
    assign P[39] = in[7] ^ in2[7];
    assign G[40] = in[6] & in2[6];
    assign P[40] = in[6] ^ in2[6];
    assign G[41] = in[5] & in2[5];
    assign P[41] = in[5] ^ in2[5];
    assign G[42] = in[4] & in2[4];
    assign P[42] = in[4] ^ in2[4];
    assign G[43] = in[3] & in2[3];
    assign P[43] = in[3] ^ in2[3];
    assign G[44] = in[2] & in2[2];
    assign P[44] = in[2] ^ in2[2];
    assign G[45] = in[1] & in2[1];
    assign P[45] = in[1] ^ in2[1];
    assign G[46] = in[0] & in2[0];
    assign P[46] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign C[46] = G[45] | (P[45] & C[45]);
    assign cout = G[46] | (P[46] & C[46]);
    assign sum = P ^ C;
endmodule

module CLA46(output [45:0] sum, output cout, input [45:0] in1, input [45:0] in2;

    wire[45:0] G;
    wire[45:0] C;
    wire[45:0] P;

    assign G[0] = in[45] & in2[45];
    assign P[0] = in[45] ^ in2[45];
    assign G[1] = in[44] & in2[44];
    assign P[1] = in[44] ^ in2[44];
    assign G[2] = in[43] & in2[43];
    assign P[2] = in[43] ^ in2[43];
    assign G[3] = in[42] & in2[42];
    assign P[3] = in[42] ^ in2[42];
    assign G[4] = in[41] & in2[41];
    assign P[4] = in[41] ^ in2[41];
    assign G[5] = in[40] & in2[40];
    assign P[5] = in[40] ^ in2[40];
    assign G[6] = in[39] & in2[39];
    assign P[6] = in[39] ^ in2[39];
    assign G[7] = in[38] & in2[38];
    assign P[7] = in[38] ^ in2[38];
    assign G[8] = in[37] & in2[37];
    assign P[8] = in[37] ^ in2[37];
    assign G[9] = in[36] & in2[36];
    assign P[9] = in[36] ^ in2[36];
    assign G[10] = in[35] & in2[35];
    assign P[10] = in[35] ^ in2[35];
    assign G[11] = in[34] & in2[34];
    assign P[11] = in[34] ^ in2[34];
    assign G[12] = in[33] & in2[33];
    assign P[12] = in[33] ^ in2[33];
    assign G[13] = in[32] & in2[32];
    assign P[13] = in[32] ^ in2[32];
    assign G[14] = in[31] & in2[31];
    assign P[14] = in[31] ^ in2[31];
    assign G[15] = in[30] & in2[30];
    assign P[15] = in[30] ^ in2[30];
    assign G[16] = in[29] & in2[29];
    assign P[16] = in[29] ^ in2[29];
    assign G[17] = in[28] & in2[28];
    assign P[17] = in[28] ^ in2[28];
    assign G[18] = in[27] & in2[27];
    assign P[18] = in[27] ^ in2[27];
    assign G[19] = in[26] & in2[26];
    assign P[19] = in[26] ^ in2[26];
    assign G[20] = in[25] & in2[25];
    assign P[20] = in[25] ^ in2[25];
    assign G[21] = in[24] & in2[24];
    assign P[21] = in[24] ^ in2[24];
    assign G[22] = in[23] & in2[23];
    assign P[22] = in[23] ^ in2[23];
    assign G[23] = in[22] & in2[22];
    assign P[23] = in[22] ^ in2[22];
    assign G[24] = in[21] & in2[21];
    assign P[24] = in[21] ^ in2[21];
    assign G[25] = in[20] & in2[20];
    assign P[25] = in[20] ^ in2[20];
    assign G[26] = in[19] & in2[19];
    assign P[26] = in[19] ^ in2[19];
    assign G[27] = in[18] & in2[18];
    assign P[27] = in[18] ^ in2[18];
    assign G[28] = in[17] & in2[17];
    assign P[28] = in[17] ^ in2[17];
    assign G[29] = in[16] & in2[16];
    assign P[29] = in[16] ^ in2[16];
    assign G[30] = in[15] & in2[15];
    assign P[30] = in[15] ^ in2[15];
    assign G[31] = in[14] & in2[14];
    assign P[31] = in[14] ^ in2[14];
    assign G[32] = in[13] & in2[13];
    assign P[32] = in[13] ^ in2[13];
    assign G[33] = in[12] & in2[12];
    assign P[33] = in[12] ^ in2[12];
    assign G[34] = in[11] & in2[11];
    assign P[34] = in[11] ^ in2[11];
    assign G[35] = in[10] & in2[10];
    assign P[35] = in[10] ^ in2[10];
    assign G[36] = in[9] & in2[9];
    assign P[36] = in[9] ^ in2[9];
    assign G[37] = in[8] & in2[8];
    assign P[37] = in[8] ^ in2[8];
    assign G[38] = in[7] & in2[7];
    assign P[38] = in[7] ^ in2[7];
    assign G[39] = in[6] & in2[6];
    assign P[39] = in[6] ^ in2[6];
    assign G[40] = in[5] & in2[5];
    assign P[40] = in[5] ^ in2[5];
    assign G[41] = in[4] & in2[4];
    assign P[41] = in[4] ^ in2[4];
    assign G[42] = in[3] & in2[3];
    assign P[42] = in[3] ^ in2[3];
    assign G[43] = in[2] & in2[2];
    assign P[43] = in[2] ^ in2[2];
    assign G[44] = in[1] & in2[1];
    assign P[44] = in[1] ^ in2[1];
    assign G[45] = in[0] & in2[0];
    assign P[45] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign C[45] = G[44] | (P[44] & C[44]);
    assign cout = G[45] | (P[45] & C[45]);
    assign sum = P ^ C;
endmodule

module CLA45(output [44:0] sum, output cout, input [44:0] in1, input [44:0] in2;

    wire[44:0] G;
    wire[44:0] C;
    wire[44:0] P;

    assign G[0] = in[44] & in2[44];
    assign P[0] = in[44] ^ in2[44];
    assign G[1] = in[43] & in2[43];
    assign P[1] = in[43] ^ in2[43];
    assign G[2] = in[42] & in2[42];
    assign P[2] = in[42] ^ in2[42];
    assign G[3] = in[41] & in2[41];
    assign P[3] = in[41] ^ in2[41];
    assign G[4] = in[40] & in2[40];
    assign P[4] = in[40] ^ in2[40];
    assign G[5] = in[39] & in2[39];
    assign P[5] = in[39] ^ in2[39];
    assign G[6] = in[38] & in2[38];
    assign P[6] = in[38] ^ in2[38];
    assign G[7] = in[37] & in2[37];
    assign P[7] = in[37] ^ in2[37];
    assign G[8] = in[36] & in2[36];
    assign P[8] = in[36] ^ in2[36];
    assign G[9] = in[35] & in2[35];
    assign P[9] = in[35] ^ in2[35];
    assign G[10] = in[34] & in2[34];
    assign P[10] = in[34] ^ in2[34];
    assign G[11] = in[33] & in2[33];
    assign P[11] = in[33] ^ in2[33];
    assign G[12] = in[32] & in2[32];
    assign P[12] = in[32] ^ in2[32];
    assign G[13] = in[31] & in2[31];
    assign P[13] = in[31] ^ in2[31];
    assign G[14] = in[30] & in2[30];
    assign P[14] = in[30] ^ in2[30];
    assign G[15] = in[29] & in2[29];
    assign P[15] = in[29] ^ in2[29];
    assign G[16] = in[28] & in2[28];
    assign P[16] = in[28] ^ in2[28];
    assign G[17] = in[27] & in2[27];
    assign P[17] = in[27] ^ in2[27];
    assign G[18] = in[26] & in2[26];
    assign P[18] = in[26] ^ in2[26];
    assign G[19] = in[25] & in2[25];
    assign P[19] = in[25] ^ in2[25];
    assign G[20] = in[24] & in2[24];
    assign P[20] = in[24] ^ in2[24];
    assign G[21] = in[23] & in2[23];
    assign P[21] = in[23] ^ in2[23];
    assign G[22] = in[22] & in2[22];
    assign P[22] = in[22] ^ in2[22];
    assign G[23] = in[21] & in2[21];
    assign P[23] = in[21] ^ in2[21];
    assign G[24] = in[20] & in2[20];
    assign P[24] = in[20] ^ in2[20];
    assign G[25] = in[19] & in2[19];
    assign P[25] = in[19] ^ in2[19];
    assign G[26] = in[18] & in2[18];
    assign P[26] = in[18] ^ in2[18];
    assign G[27] = in[17] & in2[17];
    assign P[27] = in[17] ^ in2[17];
    assign G[28] = in[16] & in2[16];
    assign P[28] = in[16] ^ in2[16];
    assign G[29] = in[15] & in2[15];
    assign P[29] = in[15] ^ in2[15];
    assign G[30] = in[14] & in2[14];
    assign P[30] = in[14] ^ in2[14];
    assign G[31] = in[13] & in2[13];
    assign P[31] = in[13] ^ in2[13];
    assign G[32] = in[12] & in2[12];
    assign P[32] = in[12] ^ in2[12];
    assign G[33] = in[11] & in2[11];
    assign P[33] = in[11] ^ in2[11];
    assign G[34] = in[10] & in2[10];
    assign P[34] = in[10] ^ in2[10];
    assign G[35] = in[9] & in2[9];
    assign P[35] = in[9] ^ in2[9];
    assign G[36] = in[8] & in2[8];
    assign P[36] = in[8] ^ in2[8];
    assign G[37] = in[7] & in2[7];
    assign P[37] = in[7] ^ in2[7];
    assign G[38] = in[6] & in2[6];
    assign P[38] = in[6] ^ in2[6];
    assign G[39] = in[5] & in2[5];
    assign P[39] = in[5] ^ in2[5];
    assign G[40] = in[4] & in2[4];
    assign P[40] = in[4] ^ in2[4];
    assign G[41] = in[3] & in2[3];
    assign P[41] = in[3] ^ in2[3];
    assign G[42] = in[2] & in2[2];
    assign P[42] = in[2] ^ in2[2];
    assign G[43] = in[1] & in2[1];
    assign P[43] = in[1] ^ in2[1];
    assign G[44] = in[0] & in2[0];
    assign P[44] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign C[44] = G[43] | (P[43] & C[43]);
    assign cout = G[44] | (P[44] & C[44]);
    assign sum = P ^ C;
endmodule

module CLA44(output [43:0] sum, output cout, input [43:0] in1, input [43:0] in2;

    wire[43:0] G;
    wire[43:0] C;
    wire[43:0] P;

    assign G[0] = in[43] & in2[43];
    assign P[0] = in[43] ^ in2[43];
    assign G[1] = in[42] & in2[42];
    assign P[1] = in[42] ^ in2[42];
    assign G[2] = in[41] & in2[41];
    assign P[2] = in[41] ^ in2[41];
    assign G[3] = in[40] & in2[40];
    assign P[3] = in[40] ^ in2[40];
    assign G[4] = in[39] & in2[39];
    assign P[4] = in[39] ^ in2[39];
    assign G[5] = in[38] & in2[38];
    assign P[5] = in[38] ^ in2[38];
    assign G[6] = in[37] & in2[37];
    assign P[6] = in[37] ^ in2[37];
    assign G[7] = in[36] & in2[36];
    assign P[7] = in[36] ^ in2[36];
    assign G[8] = in[35] & in2[35];
    assign P[8] = in[35] ^ in2[35];
    assign G[9] = in[34] & in2[34];
    assign P[9] = in[34] ^ in2[34];
    assign G[10] = in[33] & in2[33];
    assign P[10] = in[33] ^ in2[33];
    assign G[11] = in[32] & in2[32];
    assign P[11] = in[32] ^ in2[32];
    assign G[12] = in[31] & in2[31];
    assign P[12] = in[31] ^ in2[31];
    assign G[13] = in[30] & in2[30];
    assign P[13] = in[30] ^ in2[30];
    assign G[14] = in[29] & in2[29];
    assign P[14] = in[29] ^ in2[29];
    assign G[15] = in[28] & in2[28];
    assign P[15] = in[28] ^ in2[28];
    assign G[16] = in[27] & in2[27];
    assign P[16] = in[27] ^ in2[27];
    assign G[17] = in[26] & in2[26];
    assign P[17] = in[26] ^ in2[26];
    assign G[18] = in[25] & in2[25];
    assign P[18] = in[25] ^ in2[25];
    assign G[19] = in[24] & in2[24];
    assign P[19] = in[24] ^ in2[24];
    assign G[20] = in[23] & in2[23];
    assign P[20] = in[23] ^ in2[23];
    assign G[21] = in[22] & in2[22];
    assign P[21] = in[22] ^ in2[22];
    assign G[22] = in[21] & in2[21];
    assign P[22] = in[21] ^ in2[21];
    assign G[23] = in[20] & in2[20];
    assign P[23] = in[20] ^ in2[20];
    assign G[24] = in[19] & in2[19];
    assign P[24] = in[19] ^ in2[19];
    assign G[25] = in[18] & in2[18];
    assign P[25] = in[18] ^ in2[18];
    assign G[26] = in[17] & in2[17];
    assign P[26] = in[17] ^ in2[17];
    assign G[27] = in[16] & in2[16];
    assign P[27] = in[16] ^ in2[16];
    assign G[28] = in[15] & in2[15];
    assign P[28] = in[15] ^ in2[15];
    assign G[29] = in[14] & in2[14];
    assign P[29] = in[14] ^ in2[14];
    assign G[30] = in[13] & in2[13];
    assign P[30] = in[13] ^ in2[13];
    assign G[31] = in[12] & in2[12];
    assign P[31] = in[12] ^ in2[12];
    assign G[32] = in[11] & in2[11];
    assign P[32] = in[11] ^ in2[11];
    assign G[33] = in[10] & in2[10];
    assign P[33] = in[10] ^ in2[10];
    assign G[34] = in[9] & in2[9];
    assign P[34] = in[9] ^ in2[9];
    assign G[35] = in[8] & in2[8];
    assign P[35] = in[8] ^ in2[8];
    assign G[36] = in[7] & in2[7];
    assign P[36] = in[7] ^ in2[7];
    assign G[37] = in[6] & in2[6];
    assign P[37] = in[6] ^ in2[6];
    assign G[38] = in[5] & in2[5];
    assign P[38] = in[5] ^ in2[5];
    assign G[39] = in[4] & in2[4];
    assign P[39] = in[4] ^ in2[4];
    assign G[40] = in[3] & in2[3];
    assign P[40] = in[3] ^ in2[3];
    assign G[41] = in[2] & in2[2];
    assign P[41] = in[2] ^ in2[2];
    assign G[42] = in[1] & in2[1];
    assign P[42] = in[1] ^ in2[1];
    assign G[43] = in[0] & in2[0];
    assign P[43] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign C[43] = G[42] | (P[42] & C[42]);
    assign cout = G[43] | (P[43] & C[43]);
    assign sum = P ^ C;
endmodule

module CLA43(output [42:0] sum, output cout, input [42:0] in1, input [42:0] in2;

    wire[42:0] G;
    wire[42:0] C;
    wire[42:0] P;

    assign G[0] = in[42] & in2[42];
    assign P[0] = in[42] ^ in2[42];
    assign G[1] = in[41] & in2[41];
    assign P[1] = in[41] ^ in2[41];
    assign G[2] = in[40] & in2[40];
    assign P[2] = in[40] ^ in2[40];
    assign G[3] = in[39] & in2[39];
    assign P[3] = in[39] ^ in2[39];
    assign G[4] = in[38] & in2[38];
    assign P[4] = in[38] ^ in2[38];
    assign G[5] = in[37] & in2[37];
    assign P[5] = in[37] ^ in2[37];
    assign G[6] = in[36] & in2[36];
    assign P[6] = in[36] ^ in2[36];
    assign G[7] = in[35] & in2[35];
    assign P[7] = in[35] ^ in2[35];
    assign G[8] = in[34] & in2[34];
    assign P[8] = in[34] ^ in2[34];
    assign G[9] = in[33] & in2[33];
    assign P[9] = in[33] ^ in2[33];
    assign G[10] = in[32] & in2[32];
    assign P[10] = in[32] ^ in2[32];
    assign G[11] = in[31] & in2[31];
    assign P[11] = in[31] ^ in2[31];
    assign G[12] = in[30] & in2[30];
    assign P[12] = in[30] ^ in2[30];
    assign G[13] = in[29] & in2[29];
    assign P[13] = in[29] ^ in2[29];
    assign G[14] = in[28] & in2[28];
    assign P[14] = in[28] ^ in2[28];
    assign G[15] = in[27] & in2[27];
    assign P[15] = in[27] ^ in2[27];
    assign G[16] = in[26] & in2[26];
    assign P[16] = in[26] ^ in2[26];
    assign G[17] = in[25] & in2[25];
    assign P[17] = in[25] ^ in2[25];
    assign G[18] = in[24] & in2[24];
    assign P[18] = in[24] ^ in2[24];
    assign G[19] = in[23] & in2[23];
    assign P[19] = in[23] ^ in2[23];
    assign G[20] = in[22] & in2[22];
    assign P[20] = in[22] ^ in2[22];
    assign G[21] = in[21] & in2[21];
    assign P[21] = in[21] ^ in2[21];
    assign G[22] = in[20] & in2[20];
    assign P[22] = in[20] ^ in2[20];
    assign G[23] = in[19] & in2[19];
    assign P[23] = in[19] ^ in2[19];
    assign G[24] = in[18] & in2[18];
    assign P[24] = in[18] ^ in2[18];
    assign G[25] = in[17] & in2[17];
    assign P[25] = in[17] ^ in2[17];
    assign G[26] = in[16] & in2[16];
    assign P[26] = in[16] ^ in2[16];
    assign G[27] = in[15] & in2[15];
    assign P[27] = in[15] ^ in2[15];
    assign G[28] = in[14] & in2[14];
    assign P[28] = in[14] ^ in2[14];
    assign G[29] = in[13] & in2[13];
    assign P[29] = in[13] ^ in2[13];
    assign G[30] = in[12] & in2[12];
    assign P[30] = in[12] ^ in2[12];
    assign G[31] = in[11] & in2[11];
    assign P[31] = in[11] ^ in2[11];
    assign G[32] = in[10] & in2[10];
    assign P[32] = in[10] ^ in2[10];
    assign G[33] = in[9] & in2[9];
    assign P[33] = in[9] ^ in2[9];
    assign G[34] = in[8] & in2[8];
    assign P[34] = in[8] ^ in2[8];
    assign G[35] = in[7] & in2[7];
    assign P[35] = in[7] ^ in2[7];
    assign G[36] = in[6] & in2[6];
    assign P[36] = in[6] ^ in2[6];
    assign G[37] = in[5] & in2[5];
    assign P[37] = in[5] ^ in2[5];
    assign G[38] = in[4] & in2[4];
    assign P[38] = in[4] ^ in2[4];
    assign G[39] = in[3] & in2[3];
    assign P[39] = in[3] ^ in2[3];
    assign G[40] = in[2] & in2[2];
    assign P[40] = in[2] ^ in2[2];
    assign G[41] = in[1] & in2[1];
    assign P[41] = in[1] ^ in2[1];
    assign G[42] = in[0] & in2[0];
    assign P[42] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign C[42] = G[41] | (P[41] & C[41]);
    assign cout = G[42] | (P[42] & C[42]);
    assign sum = P ^ C;
endmodule

module CLA42(output [41:0] sum, output cout, input [41:0] in1, input [41:0] in2;

    wire[41:0] G;
    wire[41:0] C;
    wire[41:0] P;

    assign G[0] = in[41] & in2[41];
    assign P[0] = in[41] ^ in2[41];
    assign G[1] = in[40] & in2[40];
    assign P[1] = in[40] ^ in2[40];
    assign G[2] = in[39] & in2[39];
    assign P[2] = in[39] ^ in2[39];
    assign G[3] = in[38] & in2[38];
    assign P[3] = in[38] ^ in2[38];
    assign G[4] = in[37] & in2[37];
    assign P[4] = in[37] ^ in2[37];
    assign G[5] = in[36] & in2[36];
    assign P[5] = in[36] ^ in2[36];
    assign G[6] = in[35] & in2[35];
    assign P[6] = in[35] ^ in2[35];
    assign G[7] = in[34] & in2[34];
    assign P[7] = in[34] ^ in2[34];
    assign G[8] = in[33] & in2[33];
    assign P[8] = in[33] ^ in2[33];
    assign G[9] = in[32] & in2[32];
    assign P[9] = in[32] ^ in2[32];
    assign G[10] = in[31] & in2[31];
    assign P[10] = in[31] ^ in2[31];
    assign G[11] = in[30] & in2[30];
    assign P[11] = in[30] ^ in2[30];
    assign G[12] = in[29] & in2[29];
    assign P[12] = in[29] ^ in2[29];
    assign G[13] = in[28] & in2[28];
    assign P[13] = in[28] ^ in2[28];
    assign G[14] = in[27] & in2[27];
    assign P[14] = in[27] ^ in2[27];
    assign G[15] = in[26] & in2[26];
    assign P[15] = in[26] ^ in2[26];
    assign G[16] = in[25] & in2[25];
    assign P[16] = in[25] ^ in2[25];
    assign G[17] = in[24] & in2[24];
    assign P[17] = in[24] ^ in2[24];
    assign G[18] = in[23] & in2[23];
    assign P[18] = in[23] ^ in2[23];
    assign G[19] = in[22] & in2[22];
    assign P[19] = in[22] ^ in2[22];
    assign G[20] = in[21] & in2[21];
    assign P[20] = in[21] ^ in2[21];
    assign G[21] = in[20] & in2[20];
    assign P[21] = in[20] ^ in2[20];
    assign G[22] = in[19] & in2[19];
    assign P[22] = in[19] ^ in2[19];
    assign G[23] = in[18] & in2[18];
    assign P[23] = in[18] ^ in2[18];
    assign G[24] = in[17] & in2[17];
    assign P[24] = in[17] ^ in2[17];
    assign G[25] = in[16] & in2[16];
    assign P[25] = in[16] ^ in2[16];
    assign G[26] = in[15] & in2[15];
    assign P[26] = in[15] ^ in2[15];
    assign G[27] = in[14] & in2[14];
    assign P[27] = in[14] ^ in2[14];
    assign G[28] = in[13] & in2[13];
    assign P[28] = in[13] ^ in2[13];
    assign G[29] = in[12] & in2[12];
    assign P[29] = in[12] ^ in2[12];
    assign G[30] = in[11] & in2[11];
    assign P[30] = in[11] ^ in2[11];
    assign G[31] = in[10] & in2[10];
    assign P[31] = in[10] ^ in2[10];
    assign G[32] = in[9] & in2[9];
    assign P[32] = in[9] ^ in2[9];
    assign G[33] = in[8] & in2[8];
    assign P[33] = in[8] ^ in2[8];
    assign G[34] = in[7] & in2[7];
    assign P[34] = in[7] ^ in2[7];
    assign G[35] = in[6] & in2[6];
    assign P[35] = in[6] ^ in2[6];
    assign G[36] = in[5] & in2[5];
    assign P[36] = in[5] ^ in2[5];
    assign G[37] = in[4] & in2[4];
    assign P[37] = in[4] ^ in2[4];
    assign G[38] = in[3] & in2[3];
    assign P[38] = in[3] ^ in2[3];
    assign G[39] = in[2] & in2[2];
    assign P[39] = in[2] ^ in2[2];
    assign G[40] = in[1] & in2[1];
    assign P[40] = in[1] ^ in2[1];
    assign G[41] = in[0] & in2[0];
    assign P[41] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign C[41] = G[40] | (P[40] & C[40]);
    assign cout = G[41] | (P[41] & C[41]);
    assign sum = P ^ C;
endmodule

module CLA41(output [40:0] sum, output cout, input [40:0] in1, input [40:0] in2;

    wire[40:0] G;
    wire[40:0] C;
    wire[40:0] P;

    assign G[0] = in[40] & in2[40];
    assign P[0] = in[40] ^ in2[40];
    assign G[1] = in[39] & in2[39];
    assign P[1] = in[39] ^ in2[39];
    assign G[2] = in[38] & in2[38];
    assign P[2] = in[38] ^ in2[38];
    assign G[3] = in[37] & in2[37];
    assign P[3] = in[37] ^ in2[37];
    assign G[4] = in[36] & in2[36];
    assign P[4] = in[36] ^ in2[36];
    assign G[5] = in[35] & in2[35];
    assign P[5] = in[35] ^ in2[35];
    assign G[6] = in[34] & in2[34];
    assign P[6] = in[34] ^ in2[34];
    assign G[7] = in[33] & in2[33];
    assign P[7] = in[33] ^ in2[33];
    assign G[8] = in[32] & in2[32];
    assign P[8] = in[32] ^ in2[32];
    assign G[9] = in[31] & in2[31];
    assign P[9] = in[31] ^ in2[31];
    assign G[10] = in[30] & in2[30];
    assign P[10] = in[30] ^ in2[30];
    assign G[11] = in[29] & in2[29];
    assign P[11] = in[29] ^ in2[29];
    assign G[12] = in[28] & in2[28];
    assign P[12] = in[28] ^ in2[28];
    assign G[13] = in[27] & in2[27];
    assign P[13] = in[27] ^ in2[27];
    assign G[14] = in[26] & in2[26];
    assign P[14] = in[26] ^ in2[26];
    assign G[15] = in[25] & in2[25];
    assign P[15] = in[25] ^ in2[25];
    assign G[16] = in[24] & in2[24];
    assign P[16] = in[24] ^ in2[24];
    assign G[17] = in[23] & in2[23];
    assign P[17] = in[23] ^ in2[23];
    assign G[18] = in[22] & in2[22];
    assign P[18] = in[22] ^ in2[22];
    assign G[19] = in[21] & in2[21];
    assign P[19] = in[21] ^ in2[21];
    assign G[20] = in[20] & in2[20];
    assign P[20] = in[20] ^ in2[20];
    assign G[21] = in[19] & in2[19];
    assign P[21] = in[19] ^ in2[19];
    assign G[22] = in[18] & in2[18];
    assign P[22] = in[18] ^ in2[18];
    assign G[23] = in[17] & in2[17];
    assign P[23] = in[17] ^ in2[17];
    assign G[24] = in[16] & in2[16];
    assign P[24] = in[16] ^ in2[16];
    assign G[25] = in[15] & in2[15];
    assign P[25] = in[15] ^ in2[15];
    assign G[26] = in[14] & in2[14];
    assign P[26] = in[14] ^ in2[14];
    assign G[27] = in[13] & in2[13];
    assign P[27] = in[13] ^ in2[13];
    assign G[28] = in[12] & in2[12];
    assign P[28] = in[12] ^ in2[12];
    assign G[29] = in[11] & in2[11];
    assign P[29] = in[11] ^ in2[11];
    assign G[30] = in[10] & in2[10];
    assign P[30] = in[10] ^ in2[10];
    assign G[31] = in[9] & in2[9];
    assign P[31] = in[9] ^ in2[9];
    assign G[32] = in[8] & in2[8];
    assign P[32] = in[8] ^ in2[8];
    assign G[33] = in[7] & in2[7];
    assign P[33] = in[7] ^ in2[7];
    assign G[34] = in[6] & in2[6];
    assign P[34] = in[6] ^ in2[6];
    assign G[35] = in[5] & in2[5];
    assign P[35] = in[5] ^ in2[5];
    assign G[36] = in[4] & in2[4];
    assign P[36] = in[4] ^ in2[4];
    assign G[37] = in[3] & in2[3];
    assign P[37] = in[3] ^ in2[3];
    assign G[38] = in[2] & in2[2];
    assign P[38] = in[2] ^ in2[2];
    assign G[39] = in[1] & in2[1];
    assign P[39] = in[1] ^ in2[1];
    assign G[40] = in[0] & in2[0];
    assign P[40] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign C[40] = G[39] | (P[39] & C[39]);
    assign cout = G[40] | (P[40] & C[40]);
    assign sum = P ^ C;
endmodule

module CLA40(output [39:0] sum, output cout, input [39:0] in1, input [39:0] in2;

    wire[39:0] G;
    wire[39:0] C;
    wire[39:0] P;

    assign G[0] = in[39] & in2[39];
    assign P[0] = in[39] ^ in2[39];
    assign G[1] = in[38] & in2[38];
    assign P[1] = in[38] ^ in2[38];
    assign G[2] = in[37] & in2[37];
    assign P[2] = in[37] ^ in2[37];
    assign G[3] = in[36] & in2[36];
    assign P[3] = in[36] ^ in2[36];
    assign G[4] = in[35] & in2[35];
    assign P[4] = in[35] ^ in2[35];
    assign G[5] = in[34] & in2[34];
    assign P[5] = in[34] ^ in2[34];
    assign G[6] = in[33] & in2[33];
    assign P[6] = in[33] ^ in2[33];
    assign G[7] = in[32] & in2[32];
    assign P[7] = in[32] ^ in2[32];
    assign G[8] = in[31] & in2[31];
    assign P[8] = in[31] ^ in2[31];
    assign G[9] = in[30] & in2[30];
    assign P[9] = in[30] ^ in2[30];
    assign G[10] = in[29] & in2[29];
    assign P[10] = in[29] ^ in2[29];
    assign G[11] = in[28] & in2[28];
    assign P[11] = in[28] ^ in2[28];
    assign G[12] = in[27] & in2[27];
    assign P[12] = in[27] ^ in2[27];
    assign G[13] = in[26] & in2[26];
    assign P[13] = in[26] ^ in2[26];
    assign G[14] = in[25] & in2[25];
    assign P[14] = in[25] ^ in2[25];
    assign G[15] = in[24] & in2[24];
    assign P[15] = in[24] ^ in2[24];
    assign G[16] = in[23] & in2[23];
    assign P[16] = in[23] ^ in2[23];
    assign G[17] = in[22] & in2[22];
    assign P[17] = in[22] ^ in2[22];
    assign G[18] = in[21] & in2[21];
    assign P[18] = in[21] ^ in2[21];
    assign G[19] = in[20] & in2[20];
    assign P[19] = in[20] ^ in2[20];
    assign G[20] = in[19] & in2[19];
    assign P[20] = in[19] ^ in2[19];
    assign G[21] = in[18] & in2[18];
    assign P[21] = in[18] ^ in2[18];
    assign G[22] = in[17] & in2[17];
    assign P[22] = in[17] ^ in2[17];
    assign G[23] = in[16] & in2[16];
    assign P[23] = in[16] ^ in2[16];
    assign G[24] = in[15] & in2[15];
    assign P[24] = in[15] ^ in2[15];
    assign G[25] = in[14] & in2[14];
    assign P[25] = in[14] ^ in2[14];
    assign G[26] = in[13] & in2[13];
    assign P[26] = in[13] ^ in2[13];
    assign G[27] = in[12] & in2[12];
    assign P[27] = in[12] ^ in2[12];
    assign G[28] = in[11] & in2[11];
    assign P[28] = in[11] ^ in2[11];
    assign G[29] = in[10] & in2[10];
    assign P[29] = in[10] ^ in2[10];
    assign G[30] = in[9] & in2[9];
    assign P[30] = in[9] ^ in2[9];
    assign G[31] = in[8] & in2[8];
    assign P[31] = in[8] ^ in2[8];
    assign G[32] = in[7] & in2[7];
    assign P[32] = in[7] ^ in2[7];
    assign G[33] = in[6] & in2[6];
    assign P[33] = in[6] ^ in2[6];
    assign G[34] = in[5] & in2[5];
    assign P[34] = in[5] ^ in2[5];
    assign G[35] = in[4] & in2[4];
    assign P[35] = in[4] ^ in2[4];
    assign G[36] = in[3] & in2[3];
    assign P[36] = in[3] ^ in2[3];
    assign G[37] = in[2] & in2[2];
    assign P[37] = in[2] ^ in2[2];
    assign G[38] = in[1] & in2[1];
    assign P[38] = in[1] ^ in2[1];
    assign G[39] = in[0] & in2[0];
    assign P[39] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign C[39] = G[38] | (P[38] & C[38]);
    assign cout = G[39] | (P[39] & C[39]);
    assign sum = P ^ C;
endmodule

module CLA39(output [38:0] sum, output cout, input [38:0] in1, input [38:0] in2;

    wire[38:0] G;
    wire[38:0] C;
    wire[38:0] P;

    assign G[0] = in[38] & in2[38];
    assign P[0] = in[38] ^ in2[38];
    assign G[1] = in[37] & in2[37];
    assign P[1] = in[37] ^ in2[37];
    assign G[2] = in[36] & in2[36];
    assign P[2] = in[36] ^ in2[36];
    assign G[3] = in[35] & in2[35];
    assign P[3] = in[35] ^ in2[35];
    assign G[4] = in[34] & in2[34];
    assign P[4] = in[34] ^ in2[34];
    assign G[5] = in[33] & in2[33];
    assign P[5] = in[33] ^ in2[33];
    assign G[6] = in[32] & in2[32];
    assign P[6] = in[32] ^ in2[32];
    assign G[7] = in[31] & in2[31];
    assign P[7] = in[31] ^ in2[31];
    assign G[8] = in[30] & in2[30];
    assign P[8] = in[30] ^ in2[30];
    assign G[9] = in[29] & in2[29];
    assign P[9] = in[29] ^ in2[29];
    assign G[10] = in[28] & in2[28];
    assign P[10] = in[28] ^ in2[28];
    assign G[11] = in[27] & in2[27];
    assign P[11] = in[27] ^ in2[27];
    assign G[12] = in[26] & in2[26];
    assign P[12] = in[26] ^ in2[26];
    assign G[13] = in[25] & in2[25];
    assign P[13] = in[25] ^ in2[25];
    assign G[14] = in[24] & in2[24];
    assign P[14] = in[24] ^ in2[24];
    assign G[15] = in[23] & in2[23];
    assign P[15] = in[23] ^ in2[23];
    assign G[16] = in[22] & in2[22];
    assign P[16] = in[22] ^ in2[22];
    assign G[17] = in[21] & in2[21];
    assign P[17] = in[21] ^ in2[21];
    assign G[18] = in[20] & in2[20];
    assign P[18] = in[20] ^ in2[20];
    assign G[19] = in[19] & in2[19];
    assign P[19] = in[19] ^ in2[19];
    assign G[20] = in[18] & in2[18];
    assign P[20] = in[18] ^ in2[18];
    assign G[21] = in[17] & in2[17];
    assign P[21] = in[17] ^ in2[17];
    assign G[22] = in[16] & in2[16];
    assign P[22] = in[16] ^ in2[16];
    assign G[23] = in[15] & in2[15];
    assign P[23] = in[15] ^ in2[15];
    assign G[24] = in[14] & in2[14];
    assign P[24] = in[14] ^ in2[14];
    assign G[25] = in[13] & in2[13];
    assign P[25] = in[13] ^ in2[13];
    assign G[26] = in[12] & in2[12];
    assign P[26] = in[12] ^ in2[12];
    assign G[27] = in[11] & in2[11];
    assign P[27] = in[11] ^ in2[11];
    assign G[28] = in[10] & in2[10];
    assign P[28] = in[10] ^ in2[10];
    assign G[29] = in[9] & in2[9];
    assign P[29] = in[9] ^ in2[9];
    assign G[30] = in[8] & in2[8];
    assign P[30] = in[8] ^ in2[8];
    assign G[31] = in[7] & in2[7];
    assign P[31] = in[7] ^ in2[7];
    assign G[32] = in[6] & in2[6];
    assign P[32] = in[6] ^ in2[6];
    assign G[33] = in[5] & in2[5];
    assign P[33] = in[5] ^ in2[5];
    assign G[34] = in[4] & in2[4];
    assign P[34] = in[4] ^ in2[4];
    assign G[35] = in[3] & in2[3];
    assign P[35] = in[3] ^ in2[3];
    assign G[36] = in[2] & in2[2];
    assign P[36] = in[2] ^ in2[2];
    assign G[37] = in[1] & in2[1];
    assign P[37] = in[1] ^ in2[1];
    assign G[38] = in[0] & in2[0];
    assign P[38] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign C[38] = G[37] | (P[37] & C[37]);
    assign cout = G[38] | (P[38] & C[38]);
    assign sum = P ^ C;
endmodule

module CLA38(output [37:0] sum, output cout, input [37:0] in1, input [37:0] in2;

    wire[37:0] G;
    wire[37:0] C;
    wire[37:0] P;

    assign G[0] = in[37] & in2[37];
    assign P[0] = in[37] ^ in2[37];
    assign G[1] = in[36] & in2[36];
    assign P[1] = in[36] ^ in2[36];
    assign G[2] = in[35] & in2[35];
    assign P[2] = in[35] ^ in2[35];
    assign G[3] = in[34] & in2[34];
    assign P[3] = in[34] ^ in2[34];
    assign G[4] = in[33] & in2[33];
    assign P[4] = in[33] ^ in2[33];
    assign G[5] = in[32] & in2[32];
    assign P[5] = in[32] ^ in2[32];
    assign G[6] = in[31] & in2[31];
    assign P[6] = in[31] ^ in2[31];
    assign G[7] = in[30] & in2[30];
    assign P[7] = in[30] ^ in2[30];
    assign G[8] = in[29] & in2[29];
    assign P[8] = in[29] ^ in2[29];
    assign G[9] = in[28] & in2[28];
    assign P[9] = in[28] ^ in2[28];
    assign G[10] = in[27] & in2[27];
    assign P[10] = in[27] ^ in2[27];
    assign G[11] = in[26] & in2[26];
    assign P[11] = in[26] ^ in2[26];
    assign G[12] = in[25] & in2[25];
    assign P[12] = in[25] ^ in2[25];
    assign G[13] = in[24] & in2[24];
    assign P[13] = in[24] ^ in2[24];
    assign G[14] = in[23] & in2[23];
    assign P[14] = in[23] ^ in2[23];
    assign G[15] = in[22] & in2[22];
    assign P[15] = in[22] ^ in2[22];
    assign G[16] = in[21] & in2[21];
    assign P[16] = in[21] ^ in2[21];
    assign G[17] = in[20] & in2[20];
    assign P[17] = in[20] ^ in2[20];
    assign G[18] = in[19] & in2[19];
    assign P[18] = in[19] ^ in2[19];
    assign G[19] = in[18] & in2[18];
    assign P[19] = in[18] ^ in2[18];
    assign G[20] = in[17] & in2[17];
    assign P[20] = in[17] ^ in2[17];
    assign G[21] = in[16] & in2[16];
    assign P[21] = in[16] ^ in2[16];
    assign G[22] = in[15] & in2[15];
    assign P[22] = in[15] ^ in2[15];
    assign G[23] = in[14] & in2[14];
    assign P[23] = in[14] ^ in2[14];
    assign G[24] = in[13] & in2[13];
    assign P[24] = in[13] ^ in2[13];
    assign G[25] = in[12] & in2[12];
    assign P[25] = in[12] ^ in2[12];
    assign G[26] = in[11] & in2[11];
    assign P[26] = in[11] ^ in2[11];
    assign G[27] = in[10] & in2[10];
    assign P[27] = in[10] ^ in2[10];
    assign G[28] = in[9] & in2[9];
    assign P[28] = in[9] ^ in2[9];
    assign G[29] = in[8] & in2[8];
    assign P[29] = in[8] ^ in2[8];
    assign G[30] = in[7] & in2[7];
    assign P[30] = in[7] ^ in2[7];
    assign G[31] = in[6] & in2[6];
    assign P[31] = in[6] ^ in2[6];
    assign G[32] = in[5] & in2[5];
    assign P[32] = in[5] ^ in2[5];
    assign G[33] = in[4] & in2[4];
    assign P[33] = in[4] ^ in2[4];
    assign G[34] = in[3] & in2[3];
    assign P[34] = in[3] ^ in2[3];
    assign G[35] = in[2] & in2[2];
    assign P[35] = in[2] ^ in2[2];
    assign G[36] = in[1] & in2[1];
    assign P[36] = in[1] ^ in2[1];
    assign G[37] = in[0] & in2[0];
    assign P[37] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign C[37] = G[36] | (P[36] & C[36]);
    assign cout = G[37] | (P[37] & C[37]);
    assign sum = P ^ C;
endmodule

module CLA37(output [36:0] sum, output cout, input [36:0] in1, input [36:0] in2;

    wire[36:0] G;
    wire[36:0] C;
    wire[36:0] P;

    assign G[0] = in[36] & in2[36];
    assign P[0] = in[36] ^ in2[36];
    assign G[1] = in[35] & in2[35];
    assign P[1] = in[35] ^ in2[35];
    assign G[2] = in[34] & in2[34];
    assign P[2] = in[34] ^ in2[34];
    assign G[3] = in[33] & in2[33];
    assign P[3] = in[33] ^ in2[33];
    assign G[4] = in[32] & in2[32];
    assign P[4] = in[32] ^ in2[32];
    assign G[5] = in[31] & in2[31];
    assign P[5] = in[31] ^ in2[31];
    assign G[6] = in[30] & in2[30];
    assign P[6] = in[30] ^ in2[30];
    assign G[7] = in[29] & in2[29];
    assign P[7] = in[29] ^ in2[29];
    assign G[8] = in[28] & in2[28];
    assign P[8] = in[28] ^ in2[28];
    assign G[9] = in[27] & in2[27];
    assign P[9] = in[27] ^ in2[27];
    assign G[10] = in[26] & in2[26];
    assign P[10] = in[26] ^ in2[26];
    assign G[11] = in[25] & in2[25];
    assign P[11] = in[25] ^ in2[25];
    assign G[12] = in[24] & in2[24];
    assign P[12] = in[24] ^ in2[24];
    assign G[13] = in[23] & in2[23];
    assign P[13] = in[23] ^ in2[23];
    assign G[14] = in[22] & in2[22];
    assign P[14] = in[22] ^ in2[22];
    assign G[15] = in[21] & in2[21];
    assign P[15] = in[21] ^ in2[21];
    assign G[16] = in[20] & in2[20];
    assign P[16] = in[20] ^ in2[20];
    assign G[17] = in[19] & in2[19];
    assign P[17] = in[19] ^ in2[19];
    assign G[18] = in[18] & in2[18];
    assign P[18] = in[18] ^ in2[18];
    assign G[19] = in[17] & in2[17];
    assign P[19] = in[17] ^ in2[17];
    assign G[20] = in[16] & in2[16];
    assign P[20] = in[16] ^ in2[16];
    assign G[21] = in[15] & in2[15];
    assign P[21] = in[15] ^ in2[15];
    assign G[22] = in[14] & in2[14];
    assign P[22] = in[14] ^ in2[14];
    assign G[23] = in[13] & in2[13];
    assign P[23] = in[13] ^ in2[13];
    assign G[24] = in[12] & in2[12];
    assign P[24] = in[12] ^ in2[12];
    assign G[25] = in[11] & in2[11];
    assign P[25] = in[11] ^ in2[11];
    assign G[26] = in[10] & in2[10];
    assign P[26] = in[10] ^ in2[10];
    assign G[27] = in[9] & in2[9];
    assign P[27] = in[9] ^ in2[9];
    assign G[28] = in[8] & in2[8];
    assign P[28] = in[8] ^ in2[8];
    assign G[29] = in[7] & in2[7];
    assign P[29] = in[7] ^ in2[7];
    assign G[30] = in[6] & in2[6];
    assign P[30] = in[6] ^ in2[6];
    assign G[31] = in[5] & in2[5];
    assign P[31] = in[5] ^ in2[5];
    assign G[32] = in[4] & in2[4];
    assign P[32] = in[4] ^ in2[4];
    assign G[33] = in[3] & in2[3];
    assign P[33] = in[3] ^ in2[3];
    assign G[34] = in[2] & in2[2];
    assign P[34] = in[2] ^ in2[2];
    assign G[35] = in[1] & in2[1];
    assign P[35] = in[1] ^ in2[1];
    assign G[36] = in[0] & in2[0];
    assign P[36] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign C[36] = G[35] | (P[35] & C[35]);
    assign cout = G[36] | (P[36] & C[36]);
    assign sum = P ^ C;
endmodule

module CLA36(output [35:0] sum, output cout, input [35:0] in1, input [35:0] in2;

    wire[35:0] G;
    wire[35:0] C;
    wire[35:0] P;

    assign G[0] = in[35] & in2[35];
    assign P[0] = in[35] ^ in2[35];
    assign G[1] = in[34] & in2[34];
    assign P[1] = in[34] ^ in2[34];
    assign G[2] = in[33] & in2[33];
    assign P[2] = in[33] ^ in2[33];
    assign G[3] = in[32] & in2[32];
    assign P[3] = in[32] ^ in2[32];
    assign G[4] = in[31] & in2[31];
    assign P[4] = in[31] ^ in2[31];
    assign G[5] = in[30] & in2[30];
    assign P[5] = in[30] ^ in2[30];
    assign G[6] = in[29] & in2[29];
    assign P[6] = in[29] ^ in2[29];
    assign G[7] = in[28] & in2[28];
    assign P[7] = in[28] ^ in2[28];
    assign G[8] = in[27] & in2[27];
    assign P[8] = in[27] ^ in2[27];
    assign G[9] = in[26] & in2[26];
    assign P[9] = in[26] ^ in2[26];
    assign G[10] = in[25] & in2[25];
    assign P[10] = in[25] ^ in2[25];
    assign G[11] = in[24] & in2[24];
    assign P[11] = in[24] ^ in2[24];
    assign G[12] = in[23] & in2[23];
    assign P[12] = in[23] ^ in2[23];
    assign G[13] = in[22] & in2[22];
    assign P[13] = in[22] ^ in2[22];
    assign G[14] = in[21] & in2[21];
    assign P[14] = in[21] ^ in2[21];
    assign G[15] = in[20] & in2[20];
    assign P[15] = in[20] ^ in2[20];
    assign G[16] = in[19] & in2[19];
    assign P[16] = in[19] ^ in2[19];
    assign G[17] = in[18] & in2[18];
    assign P[17] = in[18] ^ in2[18];
    assign G[18] = in[17] & in2[17];
    assign P[18] = in[17] ^ in2[17];
    assign G[19] = in[16] & in2[16];
    assign P[19] = in[16] ^ in2[16];
    assign G[20] = in[15] & in2[15];
    assign P[20] = in[15] ^ in2[15];
    assign G[21] = in[14] & in2[14];
    assign P[21] = in[14] ^ in2[14];
    assign G[22] = in[13] & in2[13];
    assign P[22] = in[13] ^ in2[13];
    assign G[23] = in[12] & in2[12];
    assign P[23] = in[12] ^ in2[12];
    assign G[24] = in[11] & in2[11];
    assign P[24] = in[11] ^ in2[11];
    assign G[25] = in[10] & in2[10];
    assign P[25] = in[10] ^ in2[10];
    assign G[26] = in[9] & in2[9];
    assign P[26] = in[9] ^ in2[9];
    assign G[27] = in[8] & in2[8];
    assign P[27] = in[8] ^ in2[8];
    assign G[28] = in[7] & in2[7];
    assign P[28] = in[7] ^ in2[7];
    assign G[29] = in[6] & in2[6];
    assign P[29] = in[6] ^ in2[6];
    assign G[30] = in[5] & in2[5];
    assign P[30] = in[5] ^ in2[5];
    assign G[31] = in[4] & in2[4];
    assign P[31] = in[4] ^ in2[4];
    assign G[32] = in[3] & in2[3];
    assign P[32] = in[3] ^ in2[3];
    assign G[33] = in[2] & in2[2];
    assign P[33] = in[2] ^ in2[2];
    assign G[34] = in[1] & in2[1];
    assign P[34] = in[1] ^ in2[1];
    assign G[35] = in[0] & in2[0];
    assign P[35] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign C[35] = G[34] | (P[34] & C[34]);
    assign cout = G[35] | (P[35] & C[35]);
    assign sum = P ^ C;
endmodule

module CLA35(output [34:0] sum, output cout, input [34:0] in1, input [34:0] in2;

    wire[34:0] G;
    wire[34:0] C;
    wire[34:0] P;

    assign G[0] = in[34] & in2[34];
    assign P[0] = in[34] ^ in2[34];
    assign G[1] = in[33] & in2[33];
    assign P[1] = in[33] ^ in2[33];
    assign G[2] = in[32] & in2[32];
    assign P[2] = in[32] ^ in2[32];
    assign G[3] = in[31] & in2[31];
    assign P[3] = in[31] ^ in2[31];
    assign G[4] = in[30] & in2[30];
    assign P[4] = in[30] ^ in2[30];
    assign G[5] = in[29] & in2[29];
    assign P[5] = in[29] ^ in2[29];
    assign G[6] = in[28] & in2[28];
    assign P[6] = in[28] ^ in2[28];
    assign G[7] = in[27] & in2[27];
    assign P[7] = in[27] ^ in2[27];
    assign G[8] = in[26] & in2[26];
    assign P[8] = in[26] ^ in2[26];
    assign G[9] = in[25] & in2[25];
    assign P[9] = in[25] ^ in2[25];
    assign G[10] = in[24] & in2[24];
    assign P[10] = in[24] ^ in2[24];
    assign G[11] = in[23] & in2[23];
    assign P[11] = in[23] ^ in2[23];
    assign G[12] = in[22] & in2[22];
    assign P[12] = in[22] ^ in2[22];
    assign G[13] = in[21] & in2[21];
    assign P[13] = in[21] ^ in2[21];
    assign G[14] = in[20] & in2[20];
    assign P[14] = in[20] ^ in2[20];
    assign G[15] = in[19] & in2[19];
    assign P[15] = in[19] ^ in2[19];
    assign G[16] = in[18] & in2[18];
    assign P[16] = in[18] ^ in2[18];
    assign G[17] = in[17] & in2[17];
    assign P[17] = in[17] ^ in2[17];
    assign G[18] = in[16] & in2[16];
    assign P[18] = in[16] ^ in2[16];
    assign G[19] = in[15] & in2[15];
    assign P[19] = in[15] ^ in2[15];
    assign G[20] = in[14] & in2[14];
    assign P[20] = in[14] ^ in2[14];
    assign G[21] = in[13] & in2[13];
    assign P[21] = in[13] ^ in2[13];
    assign G[22] = in[12] & in2[12];
    assign P[22] = in[12] ^ in2[12];
    assign G[23] = in[11] & in2[11];
    assign P[23] = in[11] ^ in2[11];
    assign G[24] = in[10] & in2[10];
    assign P[24] = in[10] ^ in2[10];
    assign G[25] = in[9] & in2[9];
    assign P[25] = in[9] ^ in2[9];
    assign G[26] = in[8] & in2[8];
    assign P[26] = in[8] ^ in2[8];
    assign G[27] = in[7] & in2[7];
    assign P[27] = in[7] ^ in2[7];
    assign G[28] = in[6] & in2[6];
    assign P[28] = in[6] ^ in2[6];
    assign G[29] = in[5] & in2[5];
    assign P[29] = in[5] ^ in2[5];
    assign G[30] = in[4] & in2[4];
    assign P[30] = in[4] ^ in2[4];
    assign G[31] = in[3] & in2[3];
    assign P[31] = in[3] ^ in2[3];
    assign G[32] = in[2] & in2[2];
    assign P[32] = in[2] ^ in2[2];
    assign G[33] = in[1] & in2[1];
    assign P[33] = in[1] ^ in2[1];
    assign G[34] = in[0] & in2[0];
    assign P[34] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign C[34] = G[33] | (P[33] & C[33]);
    assign cout = G[34] | (P[34] & C[34]);
    assign sum = P ^ C;
endmodule

module CLA34(output [33:0] sum, output cout, input [33:0] in1, input [33:0] in2;

    wire[33:0] G;
    wire[33:0] C;
    wire[33:0] P;

    assign G[0] = in[33] & in2[33];
    assign P[0] = in[33] ^ in2[33];
    assign G[1] = in[32] & in2[32];
    assign P[1] = in[32] ^ in2[32];
    assign G[2] = in[31] & in2[31];
    assign P[2] = in[31] ^ in2[31];
    assign G[3] = in[30] & in2[30];
    assign P[3] = in[30] ^ in2[30];
    assign G[4] = in[29] & in2[29];
    assign P[4] = in[29] ^ in2[29];
    assign G[5] = in[28] & in2[28];
    assign P[5] = in[28] ^ in2[28];
    assign G[6] = in[27] & in2[27];
    assign P[6] = in[27] ^ in2[27];
    assign G[7] = in[26] & in2[26];
    assign P[7] = in[26] ^ in2[26];
    assign G[8] = in[25] & in2[25];
    assign P[8] = in[25] ^ in2[25];
    assign G[9] = in[24] & in2[24];
    assign P[9] = in[24] ^ in2[24];
    assign G[10] = in[23] & in2[23];
    assign P[10] = in[23] ^ in2[23];
    assign G[11] = in[22] & in2[22];
    assign P[11] = in[22] ^ in2[22];
    assign G[12] = in[21] & in2[21];
    assign P[12] = in[21] ^ in2[21];
    assign G[13] = in[20] & in2[20];
    assign P[13] = in[20] ^ in2[20];
    assign G[14] = in[19] & in2[19];
    assign P[14] = in[19] ^ in2[19];
    assign G[15] = in[18] & in2[18];
    assign P[15] = in[18] ^ in2[18];
    assign G[16] = in[17] & in2[17];
    assign P[16] = in[17] ^ in2[17];
    assign G[17] = in[16] & in2[16];
    assign P[17] = in[16] ^ in2[16];
    assign G[18] = in[15] & in2[15];
    assign P[18] = in[15] ^ in2[15];
    assign G[19] = in[14] & in2[14];
    assign P[19] = in[14] ^ in2[14];
    assign G[20] = in[13] & in2[13];
    assign P[20] = in[13] ^ in2[13];
    assign G[21] = in[12] & in2[12];
    assign P[21] = in[12] ^ in2[12];
    assign G[22] = in[11] & in2[11];
    assign P[22] = in[11] ^ in2[11];
    assign G[23] = in[10] & in2[10];
    assign P[23] = in[10] ^ in2[10];
    assign G[24] = in[9] & in2[9];
    assign P[24] = in[9] ^ in2[9];
    assign G[25] = in[8] & in2[8];
    assign P[25] = in[8] ^ in2[8];
    assign G[26] = in[7] & in2[7];
    assign P[26] = in[7] ^ in2[7];
    assign G[27] = in[6] & in2[6];
    assign P[27] = in[6] ^ in2[6];
    assign G[28] = in[5] & in2[5];
    assign P[28] = in[5] ^ in2[5];
    assign G[29] = in[4] & in2[4];
    assign P[29] = in[4] ^ in2[4];
    assign G[30] = in[3] & in2[3];
    assign P[30] = in[3] ^ in2[3];
    assign G[31] = in[2] & in2[2];
    assign P[31] = in[2] ^ in2[2];
    assign G[32] = in[1] & in2[1];
    assign P[32] = in[1] ^ in2[1];
    assign G[33] = in[0] & in2[0];
    assign P[33] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign C[33] = G[32] | (P[32] & C[32]);
    assign cout = G[33] | (P[33] & C[33]);
    assign sum = P ^ C;
endmodule

module CLA33(output [32:0] sum, output cout, input [32:0] in1, input [32:0] in2;

    wire[32:0] G;
    wire[32:0] C;
    wire[32:0] P;

    assign G[0] = in[32] & in2[32];
    assign P[0] = in[32] ^ in2[32];
    assign G[1] = in[31] & in2[31];
    assign P[1] = in[31] ^ in2[31];
    assign G[2] = in[30] & in2[30];
    assign P[2] = in[30] ^ in2[30];
    assign G[3] = in[29] & in2[29];
    assign P[3] = in[29] ^ in2[29];
    assign G[4] = in[28] & in2[28];
    assign P[4] = in[28] ^ in2[28];
    assign G[5] = in[27] & in2[27];
    assign P[5] = in[27] ^ in2[27];
    assign G[6] = in[26] & in2[26];
    assign P[6] = in[26] ^ in2[26];
    assign G[7] = in[25] & in2[25];
    assign P[7] = in[25] ^ in2[25];
    assign G[8] = in[24] & in2[24];
    assign P[8] = in[24] ^ in2[24];
    assign G[9] = in[23] & in2[23];
    assign P[9] = in[23] ^ in2[23];
    assign G[10] = in[22] & in2[22];
    assign P[10] = in[22] ^ in2[22];
    assign G[11] = in[21] & in2[21];
    assign P[11] = in[21] ^ in2[21];
    assign G[12] = in[20] & in2[20];
    assign P[12] = in[20] ^ in2[20];
    assign G[13] = in[19] & in2[19];
    assign P[13] = in[19] ^ in2[19];
    assign G[14] = in[18] & in2[18];
    assign P[14] = in[18] ^ in2[18];
    assign G[15] = in[17] & in2[17];
    assign P[15] = in[17] ^ in2[17];
    assign G[16] = in[16] & in2[16];
    assign P[16] = in[16] ^ in2[16];
    assign G[17] = in[15] & in2[15];
    assign P[17] = in[15] ^ in2[15];
    assign G[18] = in[14] & in2[14];
    assign P[18] = in[14] ^ in2[14];
    assign G[19] = in[13] & in2[13];
    assign P[19] = in[13] ^ in2[13];
    assign G[20] = in[12] & in2[12];
    assign P[20] = in[12] ^ in2[12];
    assign G[21] = in[11] & in2[11];
    assign P[21] = in[11] ^ in2[11];
    assign G[22] = in[10] & in2[10];
    assign P[22] = in[10] ^ in2[10];
    assign G[23] = in[9] & in2[9];
    assign P[23] = in[9] ^ in2[9];
    assign G[24] = in[8] & in2[8];
    assign P[24] = in[8] ^ in2[8];
    assign G[25] = in[7] & in2[7];
    assign P[25] = in[7] ^ in2[7];
    assign G[26] = in[6] & in2[6];
    assign P[26] = in[6] ^ in2[6];
    assign G[27] = in[5] & in2[5];
    assign P[27] = in[5] ^ in2[5];
    assign G[28] = in[4] & in2[4];
    assign P[28] = in[4] ^ in2[4];
    assign G[29] = in[3] & in2[3];
    assign P[29] = in[3] ^ in2[3];
    assign G[30] = in[2] & in2[2];
    assign P[30] = in[2] ^ in2[2];
    assign G[31] = in[1] & in2[1];
    assign P[31] = in[1] ^ in2[1];
    assign G[32] = in[0] & in2[0];
    assign P[32] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign C[32] = G[31] | (P[31] & C[31]);
    assign cout = G[32] | (P[32] & C[32]);
    assign sum = P ^ C;
endmodule

module CLA32(output [31:0] sum, output cout, input [31:0] in1, input [31:0] in2;

    wire[31:0] G;
    wire[31:0] C;
    wire[31:0] P;

    assign G[0] = in[31] & in2[31];
    assign P[0] = in[31] ^ in2[31];
    assign G[1] = in[30] & in2[30];
    assign P[1] = in[30] ^ in2[30];
    assign G[2] = in[29] & in2[29];
    assign P[2] = in[29] ^ in2[29];
    assign G[3] = in[28] & in2[28];
    assign P[3] = in[28] ^ in2[28];
    assign G[4] = in[27] & in2[27];
    assign P[4] = in[27] ^ in2[27];
    assign G[5] = in[26] & in2[26];
    assign P[5] = in[26] ^ in2[26];
    assign G[6] = in[25] & in2[25];
    assign P[6] = in[25] ^ in2[25];
    assign G[7] = in[24] & in2[24];
    assign P[7] = in[24] ^ in2[24];
    assign G[8] = in[23] & in2[23];
    assign P[8] = in[23] ^ in2[23];
    assign G[9] = in[22] & in2[22];
    assign P[9] = in[22] ^ in2[22];
    assign G[10] = in[21] & in2[21];
    assign P[10] = in[21] ^ in2[21];
    assign G[11] = in[20] & in2[20];
    assign P[11] = in[20] ^ in2[20];
    assign G[12] = in[19] & in2[19];
    assign P[12] = in[19] ^ in2[19];
    assign G[13] = in[18] & in2[18];
    assign P[13] = in[18] ^ in2[18];
    assign G[14] = in[17] & in2[17];
    assign P[14] = in[17] ^ in2[17];
    assign G[15] = in[16] & in2[16];
    assign P[15] = in[16] ^ in2[16];
    assign G[16] = in[15] & in2[15];
    assign P[16] = in[15] ^ in2[15];
    assign G[17] = in[14] & in2[14];
    assign P[17] = in[14] ^ in2[14];
    assign G[18] = in[13] & in2[13];
    assign P[18] = in[13] ^ in2[13];
    assign G[19] = in[12] & in2[12];
    assign P[19] = in[12] ^ in2[12];
    assign G[20] = in[11] & in2[11];
    assign P[20] = in[11] ^ in2[11];
    assign G[21] = in[10] & in2[10];
    assign P[21] = in[10] ^ in2[10];
    assign G[22] = in[9] & in2[9];
    assign P[22] = in[9] ^ in2[9];
    assign G[23] = in[8] & in2[8];
    assign P[23] = in[8] ^ in2[8];
    assign G[24] = in[7] & in2[7];
    assign P[24] = in[7] ^ in2[7];
    assign G[25] = in[6] & in2[6];
    assign P[25] = in[6] ^ in2[6];
    assign G[26] = in[5] & in2[5];
    assign P[26] = in[5] ^ in2[5];
    assign G[27] = in[4] & in2[4];
    assign P[27] = in[4] ^ in2[4];
    assign G[28] = in[3] & in2[3];
    assign P[28] = in[3] ^ in2[3];
    assign G[29] = in[2] & in2[2];
    assign P[29] = in[2] ^ in2[2];
    assign G[30] = in[1] & in2[1];
    assign P[30] = in[1] ^ in2[1];
    assign G[31] = in[0] & in2[0];
    assign P[31] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign C[31] = G[30] | (P[30] & C[30]);
    assign cout = G[31] | (P[31] & C[31]);
    assign sum = P ^ C;
endmodule

module CLA31(output [30:0] sum, output cout, input [30:0] in1, input [30:0] in2;

    wire[30:0] G;
    wire[30:0] C;
    wire[30:0] P;

    assign G[0] = in[30] & in2[30];
    assign P[0] = in[30] ^ in2[30];
    assign G[1] = in[29] & in2[29];
    assign P[1] = in[29] ^ in2[29];
    assign G[2] = in[28] & in2[28];
    assign P[2] = in[28] ^ in2[28];
    assign G[3] = in[27] & in2[27];
    assign P[3] = in[27] ^ in2[27];
    assign G[4] = in[26] & in2[26];
    assign P[4] = in[26] ^ in2[26];
    assign G[5] = in[25] & in2[25];
    assign P[5] = in[25] ^ in2[25];
    assign G[6] = in[24] & in2[24];
    assign P[6] = in[24] ^ in2[24];
    assign G[7] = in[23] & in2[23];
    assign P[7] = in[23] ^ in2[23];
    assign G[8] = in[22] & in2[22];
    assign P[8] = in[22] ^ in2[22];
    assign G[9] = in[21] & in2[21];
    assign P[9] = in[21] ^ in2[21];
    assign G[10] = in[20] & in2[20];
    assign P[10] = in[20] ^ in2[20];
    assign G[11] = in[19] & in2[19];
    assign P[11] = in[19] ^ in2[19];
    assign G[12] = in[18] & in2[18];
    assign P[12] = in[18] ^ in2[18];
    assign G[13] = in[17] & in2[17];
    assign P[13] = in[17] ^ in2[17];
    assign G[14] = in[16] & in2[16];
    assign P[14] = in[16] ^ in2[16];
    assign G[15] = in[15] & in2[15];
    assign P[15] = in[15] ^ in2[15];
    assign G[16] = in[14] & in2[14];
    assign P[16] = in[14] ^ in2[14];
    assign G[17] = in[13] & in2[13];
    assign P[17] = in[13] ^ in2[13];
    assign G[18] = in[12] & in2[12];
    assign P[18] = in[12] ^ in2[12];
    assign G[19] = in[11] & in2[11];
    assign P[19] = in[11] ^ in2[11];
    assign G[20] = in[10] & in2[10];
    assign P[20] = in[10] ^ in2[10];
    assign G[21] = in[9] & in2[9];
    assign P[21] = in[9] ^ in2[9];
    assign G[22] = in[8] & in2[8];
    assign P[22] = in[8] ^ in2[8];
    assign G[23] = in[7] & in2[7];
    assign P[23] = in[7] ^ in2[7];
    assign G[24] = in[6] & in2[6];
    assign P[24] = in[6] ^ in2[6];
    assign G[25] = in[5] & in2[5];
    assign P[25] = in[5] ^ in2[5];
    assign G[26] = in[4] & in2[4];
    assign P[26] = in[4] ^ in2[4];
    assign G[27] = in[3] & in2[3];
    assign P[27] = in[3] ^ in2[3];
    assign G[28] = in[2] & in2[2];
    assign P[28] = in[2] ^ in2[2];
    assign G[29] = in[1] & in2[1];
    assign P[29] = in[1] ^ in2[1];
    assign G[30] = in[0] & in2[0];
    assign P[30] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign C[30] = G[29] | (P[29] & C[29]);
    assign cout = G[30] | (P[30] & C[30]);
    assign sum = P ^ C;
endmodule

module CLA30(output [29:0] sum, output cout, input [29:0] in1, input [29:0] in2;

    wire[29:0] G;
    wire[29:0] C;
    wire[29:0] P;

    assign G[0] = in[29] & in2[29];
    assign P[0] = in[29] ^ in2[29];
    assign G[1] = in[28] & in2[28];
    assign P[1] = in[28] ^ in2[28];
    assign G[2] = in[27] & in2[27];
    assign P[2] = in[27] ^ in2[27];
    assign G[3] = in[26] & in2[26];
    assign P[3] = in[26] ^ in2[26];
    assign G[4] = in[25] & in2[25];
    assign P[4] = in[25] ^ in2[25];
    assign G[5] = in[24] & in2[24];
    assign P[5] = in[24] ^ in2[24];
    assign G[6] = in[23] & in2[23];
    assign P[6] = in[23] ^ in2[23];
    assign G[7] = in[22] & in2[22];
    assign P[7] = in[22] ^ in2[22];
    assign G[8] = in[21] & in2[21];
    assign P[8] = in[21] ^ in2[21];
    assign G[9] = in[20] & in2[20];
    assign P[9] = in[20] ^ in2[20];
    assign G[10] = in[19] & in2[19];
    assign P[10] = in[19] ^ in2[19];
    assign G[11] = in[18] & in2[18];
    assign P[11] = in[18] ^ in2[18];
    assign G[12] = in[17] & in2[17];
    assign P[12] = in[17] ^ in2[17];
    assign G[13] = in[16] & in2[16];
    assign P[13] = in[16] ^ in2[16];
    assign G[14] = in[15] & in2[15];
    assign P[14] = in[15] ^ in2[15];
    assign G[15] = in[14] & in2[14];
    assign P[15] = in[14] ^ in2[14];
    assign G[16] = in[13] & in2[13];
    assign P[16] = in[13] ^ in2[13];
    assign G[17] = in[12] & in2[12];
    assign P[17] = in[12] ^ in2[12];
    assign G[18] = in[11] & in2[11];
    assign P[18] = in[11] ^ in2[11];
    assign G[19] = in[10] & in2[10];
    assign P[19] = in[10] ^ in2[10];
    assign G[20] = in[9] & in2[9];
    assign P[20] = in[9] ^ in2[9];
    assign G[21] = in[8] & in2[8];
    assign P[21] = in[8] ^ in2[8];
    assign G[22] = in[7] & in2[7];
    assign P[22] = in[7] ^ in2[7];
    assign G[23] = in[6] & in2[6];
    assign P[23] = in[6] ^ in2[6];
    assign G[24] = in[5] & in2[5];
    assign P[24] = in[5] ^ in2[5];
    assign G[25] = in[4] & in2[4];
    assign P[25] = in[4] ^ in2[4];
    assign G[26] = in[3] & in2[3];
    assign P[26] = in[3] ^ in2[3];
    assign G[27] = in[2] & in2[2];
    assign P[27] = in[2] ^ in2[2];
    assign G[28] = in[1] & in2[1];
    assign P[28] = in[1] ^ in2[1];
    assign G[29] = in[0] & in2[0];
    assign P[29] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign C[29] = G[28] | (P[28] & C[28]);
    assign cout = G[29] | (P[29] & C[29]);
    assign sum = P ^ C;
endmodule

module CLA29(output [28:0] sum, output cout, input [28:0] in1, input [28:0] in2;

    wire[28:0] G;
    wire[28:0] C;
    wire[28:0] P;

    assign G[0] = in[28] & in2[28];
    assign P[0] = in[28] ^ in2[28];
    assign G[1] = in[27] & in2[27];
    assign P[1] = in[27] ^ in2[27];
    assign G[2] = in[26] & in2[26];
    assign P[2] = in[26] ^ in2[26];
    assign G[3] = in[25] & in2[25];
    assign P[3] = in[25] ^ in2[25];
    assign G[4] = in[24] & in2[24];
    assign P[4] = in[24] ^ in2[24];
    assign G[5] = in[23] & in2[23];
    assign P[5] = in[23] ^ in2[23];
    assign G[6] = in[22] & in2[22];
    assign P[6] = in[22] ^ in2[22];
    assign G[7] = in[21] & in2[21];
    assign P[7] = in[21] ^ in2[21];
    assign G[8] = in[20] & in2[20];
    assign P[8] = in[20] ^ in2[20];
    assign G[9] = in[19] & in2[19];
    assign P[9] = in[19] ^ in2[19];
    assign G[10] = in[18] & in2[18];
    assign P[10] = in[18] ^ in2[18];
    assign G[11] = in[17] & in2[17];
    assign P[11] = in[17] ^ in2[17];
    assign G[12] = in[16] & in2[16];
    assign P[12] = in[16] ^ in2[16];
    assign G[13] = in[15] & in2[15];
    assign P[13] = in[15] ^ in2[15];
    assign G[14] = in[14] & in2[14];
    assign P[14] = in[14] ^ in2[14];
    assign G[15] = in[13] & in2[13];
    assign P[15] = in[13] ^ in2[13];
    assign G[16] = in[12] & in2[12];
    assign P[16] = in[12] ^ in2[12];
    assign G[17] = in[11] & in2[11];
    assign P[17] = in[11] ^ in2[11];
    assign G[18] = in[10] & in2[10];
    assign P[18] = in[10] ^ in2[10];
    assign G[19] = in[9] & in2[9];
    assign P[19] = in[9] ^ in2[9];
    assign G[20] = in[8] & in2[8];
    assign P[20] = in[8] ^ in2[8];
    assign G[21] = in[7] & in2[7];
    assign P[21] = in[7] ^ in2[7];
    assign G[22] = in[6] & in2[6];
    assign P[22] = in[6] ^ in2[6];
    assign G[23] = in[5] & in2[5];
    assign P[23] = in[5] ^ in2[5];
    assign G[24] = in[4] & in2[4];
    assign P[24] = in[4] ^ in2[4];
    assign G[25] = in[3] & in2[3];
    assign P[25] = in[3] ^ in2[3];
    assign G[26] = in[2] & in2[2];
    assign P[26] = in[2] ^ in2[2];
    assign G[27] = in[1] & in2[1];
    assign P[27] = in[1] ^ in2[1];
    assign G[28] = in[0] & in2[0];
    assign P[28] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign C[28] = G[27] | (P[27] & C[27]);
    assign cout = G[28] | (P[28] & C[28]);
    assign sum = P ^ C;
endmodule

module CLA28(output [27:0] sum, output cout, input [27:0] in1, input [27:0] in2;

    wire[27:0] G;
    wire[27:0] C;
    wire[27:0] P;

    assign G[0] = in[27] & in2[27];
    assign P[0] = in[27] ^ in2[27];
    assign G[1] = in[26] & in2[26];
    assign P[1] = in[26] ^ in2[26];
    assign G[2] = in[25] & in2[25];
    assign P[2] = in[25] ^ in2[25];
    assign G[3] = in[24] & in2[24];
    assign P[3] = in[24] ^ in2[24];
    assign G[4] = in[23] & in2[23];
    assign P[4] = in[23] ^ in2[23];
    assign G[5] = in[22] & in2[22];
    assign P[5] = in[22] ^ in2[22];
    assign G[6] = in[21] & in2[21];
    assign P[6] = in[21] ^ in2[21];
    assign G[7] = in[20] & in2[20];
    assign P[7] = in[20] ^ in2[20];
    assign G[8] = in[19] & in2[19];
    assign P[8] = in[19] ^ in2[19];
    assign G[9] = in[18] & in2[18];
    assign P[9] = in[18] ^ in2[18];
    assign G[10] = in[17] & in2[17];
    assign P[10] = in[17] ^ in2[17];
    assign G[11] = in[16] & in2[16];
    assign P[11] = in[16] ^ in2[16];
    assign G[12] = in[15] & in2[15];
    assign P[12] = in[15] ^ in2[15];
    assign G[13] = in[14] & in2[14];
    assign P[13] = in[14] ^ in2[14];
    assign G[14] = in[13] & in2[13];
    assign P[14] = in[13] ^ in2[13];
    assign G[15] = in[12] & in2[12];
    assign P[15] = in[12] ^ in2[12];
    assign G[16] = in[11] & in2[11];
    assign P[16] = in[11] ^ in2[11];
    assign G[17] = in[10] & in2[10];
    assign P[17] = in[10] ^ in2[10];
    assign G[18] = in[9] & in2[9];
    assign P[18] = in[9] ^ in2[9];
    assign G[19] = in[8] & in2[8];
    assign P[19] = in[8] ^ in2[8];
    assign G[20] = in[7] & in2[7];
    assign P[20] = in[7] ^ in2[7];
    assign G[21] = in[6] & in2[6];
    assign P[21] = in[6] ^ in2[6];
    assign G[22] = in[5] & in2[5];
    assign P[22] = in[5] ^ in2[5];
    assign G[23] = in[4] & in2[4];
    assign P[23] = in[4] ^ in2[4];
    assign G[24] = in[3] & in2[3];
    assign P[24] = in[3] ^ in2[3];
    assign G[25] = in[2] & in2[2];
    assign P[25] = in[2] ^ in2[2];
    assign G[26] = in[1] & in2[1];
    assign P[26] = in[1] ^ in2[1];
    assign G[27] = in[0] & in2[0];
    assign P[27] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign C[27] = G[26] | (P[26] & C[26]);
    assign cout = G[27] | (P[27] & C[27]);
    assign sum = P ^ C;
endmodule

module CLA27(output [26:0] sum, output cout, input [26:0] in1, input [26:0] in2;

    wire[26:0] G;
    wire[26:0] C;
    wire[26:0] P;

    assign G[0] = in[26] & in2[26];
    assign P[0] = in[26] ^ in2[26];
    assign G[1] = in[25] & in2[25];
    assign P[1] = in[25] ^ in2[25];
    assign G[2] = in[24] & in2[24];
    assign P[2] = in[24] ^ in2[24];
    assign G[3] = in[23] & in2[23];
    assign P[3] = in[23] ^ in2[23];
    assign G[4] = in[22] & in2[22];
    assign P[4] = in[22] ^ in2[22];
    assign G[5] = in[21] & in2[21];
    assign P[5] = in[21] ^ in2[21];
    assign G[6] = in[20] & in2[20];
    assign P[6] = in[20] ^ in2[20];
    assign G[7] = in[19] & in2[19];
    assign P[7] = in[19] ^ in2[19];
    assign G[8] = in[18] & in2[18];
    assign P[8] = in[18] ^ in2[18];
    assign G[9] = in[17] & in2[17];
    assign P[9] = in[17] ^ in2[17];
    assign G[10] = in[16] & in2[16];
    assign P[10] = in[16] ^ in2[16];
    assign G[11] = in[15] & in2[15];
    assign P[11] = in[15] ^ in2[15];
    assign G[12] = in[14] & in2[14];
    assign P[12] = in[14] ^ in2[14];
    assign G[13] = in[13] & in2[13];
    assign P[13] = in[13] ^ in2[13];
    assign G[14] = in[12] & in2[12];
    assign P[14] = in[12] ^ in2[12];
    assign G[15] = in[11] & in2[11];
    assign P[15] = in[11] ^ in2[11];
    assign G[16] = in[10] & in2[10];
    assign P[16] = in[10] ^ in2[10];
    assign G[17] = in[9] & in2[9];
    assign P[17] = in[9] ^ in2[9];
    assign G[18] = in[8] & in2[8];
    assign P[18] = in[8] ^ in2[8];
    assign G[19] = in[7] & in2[7];
    assign P[19] = in[7] ^ in2[7];
    assign G[20] = in[6] & in2[6];
    assign P[20] = in[6] ^ in2[6];
    assign G[21] = in[5] & in2[5];
    assign P[21] = in[5] ^ in2[5];
    assign G[22] = in[4] & in2[4];
    assign P[22] = in[4] ^ in2[4];
    assign G[23] = in[3] & in2[3];
    assign P[23] = in[3] ^ in2[3];
    assign G[24] = in[2] & in2[2];
    assign P[24] = in[2] ^ in2[2];
    assign G[25] = in[1] & in2[1];
    assign P[25] = in[1] ^ in2[1];
    assign G[26] = in[0] & in2[0];
    assign P[26] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign C[26] = G[25] | (P[25] & C[25]);
    assign cout = G[26] | (P[26] & C[26]);
    assign sum = P ^ C;
endmodule

module CLA26(output [25:0] sum, output cout, input [25:0] in1, input [25:0] in2;

    wire[25:0] G;
    wire[25:0] C;
    wire[25:0] P;

    assign G[0] = in[25] & in2[25];
    assign P[0] = in[25] ^ in2[25];
    assign G[1] = in[24] & in2[24];
    assign P[1] = in[24] ^ in2[24];
    assign G[2] = in[23] & in2[23];
    assign P[2] = in[23] ^ in2[23];
    assign G[3] = in[22] & in2[22];
    assign P[3] = in[22] ^ in2[22];
    assign G[4] = in[21] & in2[21];
    assign P[4] = in[21] ^ in2[21];
    assign G[5] = in[20] & in2[20];
    assign P[5] = in[20] ^ in2[20];
    assign G[6] = in[19] & in2[19];
    assign P[6] = in[19] ^ in2[19];
    assign G[7] = in[18] & in2[18];
    assign P[7] = in[18] ^ in2[18];
    assign G[8] = in[17] & in2[17];
    assign P[8] = in[17] ^ in2[17];
    assign G[9] = in[16] & in2[16];
    assign P[9] = in[16] ^ in2[16];
    assign G[10] = in[15] & in2[15];
    assign P[10] = in[15] ^ in2[15];
    assign G[11] = in[14] & in2[14];
    assign P[11] = in[14] ^ in2[14];
    assign G[12] = in[13] & in2[13];
    assign P[12] = in[13] ^ in2[13];
    assign G[13] = in[12] & in2[12];
    assign P[13] = in[12] ^ in2[12];
    assign G[14] = in[11] & in2[11];
    assign P[14] = in[11] ^ in2[11];
    assign G[15] = in[10] & in2[10];
    assign P[15] = in[10] ^ in2[10];
    assign G[16] = in[9] & in2[9];
    assign P[16] = in[9] ^ in2[9];
    assign G[17] = in[8] & in2[8];
    assign P[17] = in[8] ^ in2[8];
    assign G[18] = in[7] & in2[7];
    assign P[18] = in[7] ^ in2[7];
    assign G[19] = in[6] & in2[6];
    assign P[19] = in[6] ^ in2[6];
    assign G[20] = in[5] & in2[5];
    assign P[20] = in[5] ^ in2[5];
    assign G[21] = in[4] & in2[4];
    assign P[21] = in[4] ^ in2[4];
    assign G[22] = in[3] & in2[3];
    assign P[22] = in[3] ^ in2[3];
    assign G[23] = in[2] & in2[2];
    assign P[23] = in[2] ^ in2[2];
    assign G[24] = in[1] & in2[1];
    assign P[24] = in[1] ^ in2[1];
    assign G[25] = in[0] & in2[0];
    assign P[25] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign C[25] = G[24] | (P[24] & C[24]);
    assign cout = G[25] | (P[25] & C[25]);
    assign sum = P ^ C;
endmodule

module CLA25(output [24:0] sum, output cout, input [24:0] in1, input [24:0] in2;

    wire[24:0] G;
    wire[24:0] C;
    wire[24:0] P;

    assign G[0] = in[24] & in2[24];
    assign P[0] = in[24] ^ in2[24];
    assign G[1] = in[23] & in2[23];
    assign P[1] = in[23] ^ in2[23];
    assign G[2] = in[22] & in2[22];
    assign P[2] = in[22] ^ in2[22];
    assign G[3] = in[21] & in2[21];
    assign P[3] = in[21] ^ in2[21];
    assign G[4] = in[20] & in2[20];
    assign P[4] = in[20] ^ in2[20];
    assign G[5] = in[19] & in2[19];
    assign P[5] = in[19] ^ in2[19];
    assign G[6] = in[18] & in2[18];
    assign P[6] = in[18] ^ in2[18];
    assign G[7] = in[17] & in2[17];
    assign P[7] = in[17] ^ in2[17];
    assign G[8] = in[16] & in2[16];
    assign P[8] = in[16] ^ in2[16];
    assign G[9] = in[15] & in2[15];
    assign P[9] = in[15] ^ in2[15];
    assign G[10] = in[14] & in2[14];
    assign P[10] = in[14] ^ in2[14];
    assign G[11] = in[13] & in2[13];
    assign P[11] = in[13] ^ in2[13];
    assign G[12] = in[12] & in2[12];
    assign P[12] = in[12] ^ in2[12];
    assign G[13] = in[11] & in2[11];
    assign P[13] = in[11] ^ in2[11];
    assign G[14] = in[10] & in2[10];
    assign P[14] = in[10] ^ in2[10];
    assign G[15] = in[9] & in2[9];
    assign P[15] = in[9] ^ in2[9];
    assign G[16] = in[8] & in2[8];
    assign P[16] = in[8] ^ in2[8];
    assign G[17] = in[7] & in2[7];
    assign P[17] = in[7] ^ in2[7];
    assign G[18] = in[6] & in2[6];
    assign P[18] = in[6] ^ in2[6];
    assign G[19] = in[5] & in2[5];
    assign P[19] = in[5] ^ in2[5];
    assign G[20] = in[4] & in2[4];
    assign P[20] = in[4] ^ in2[4];
    assign G[21] = in[3] & in2[3];
    assign P[21] = in[3] ^ in2[3];
    assign G[22] = in[2] & in2[2];
    assign P[22] = in[2] ^ in2[2];
    assign G[23] = in[1] & in2[1];
    assign P[23] = in[1] ^ in2[1];
    assign G[24] = in[0] & in2[0];
    assign P[24] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign C[24] = G[23] | (P[23] & C[23]);
    assign cout = G[24] | (P[24] & C[24]);
    assign sum = P ^ C;
endmodule

module CLA24(output [23:0] sum, output cout, input [23:0] in1, input [23:0] in2;

    wire[23:0] G;
    wire[23:0] C;
    wire[23:0] P;

    assign G[0] = in[23] & in2[23];
    assign P[0] = in[23] ^ in2[23];
    assign G[1] = in[22] & in2[22];
    assign P[1] = in[22] ^ in2[22];
    assign G[2] = in[21] & in2[21];
    assign P[2] = in[21] ^ in2[21];
    assign G[3] = in[20] & in2[20];
    assign P[3] = in[20] ^ in2[20];
    assign G[4] = in[19] & in2[19];
    assign P[4] = in[19] ^ in2[19];
    assign G[5] = in[18] & in2[18];
    assign P[5] = in[18] ^ in2[18];
    assign G[6] = in[17] & in2[17];
    assign P[6] = in[17] ^ in2[17];
    assign G[7] = in[16] & in2[16];
    assign P[7] = in[16] ^ in2[16];
    assign G[8] = in[15] & in2[15];
    assign P[8] = in[15] ^ in2[15];
    assign G[9] = in[14] & in2[14];
    assign P[9] = in[14] ^ in2[14];
    assign G[10] = in[13] & in2[13];
    assign P[10] = in[13] ^ in2[13];
    assign G[11] = in[12] & in2[12];
    assign P[11] = in[12] ^ in2[12];
    assign G[12] = in[11] & in2[11];
    assign P[12] = in[11] ^ in2[11];
    assign G[13] = in[10] & in2[10];
    assign P[13] = in[10] ^ in2[10];
    assign G[14] = in[9] & in2[9];
    assign P[14] = in[9] ^ in2[9];
    assign G[15] = in[8] & in2[8];
    assign P[15] = in[8] ^ in2[8];
    assign G[16] = in[7] & in2[7];
    assign P[16] = in[7] ^ in2[7];
    assign G[17] = in[6] & in2[6];
    assign P[17] = in[6] ^ in2[6];
    assign G[18] = in[5] & in2[5];
    assign P[18] = in[5] ^ in2[5];
    assign G[19] = in[4] & in2[4];
    assign P[19] = in[4] ^ in2[4];
    assign G[20] = in[3] & in2[3];
    assign P[20] = in[3] ^ in2[3];
    assign G[21] = in[2] & in2[2];
    assign P[21] = in[2] ^ in2[2];
    assign G[22] = in[1] & in2[1];
    assign P[22] = in[1] ^ in2[1];
    assign G[23] = in[0] & in2[0];
    assign P[23] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign C[23] = G[22] | (P[22] & C[22]);
    assign cout = G[23] | (P[23] & C[23]);
    assign sum = P ^ C;
endmodule

module CLA23(output [22:0] sum, output cout, input [22:0] in1, input [22:0] in2;

    wire[22:0] G;
    wire[22:0] C;
    wire[22:0] P;

    assign G[0] = in[22] & in2[22];
    assign P[0] = in[22] ^ in2[22];
    assign G[1] = in[21] & in2[21];
    assign P[1] = in[21] ^ in2[21];
    assign G[2] = in[20] & in2[20];
    assign P[2] = in[20] ^ in2[20];
    assign G[3] = in[19] & in2[19];
    assign P[3] = in[19] ^ in2[19];
    assign G[4] = in[18] & in2[18];
    assign P[4] = in[18] ^ in2[18];
    assign G[5] = in[17] & in2[17];
    assign P[5] = in[17] ^ in2[17];
    assign G[6] = in[16] & in2[16];
    assign P[6] = in[16] ^ in2[16];
    assign G[7] = in[15] & in2[15];
    assign P[7] = in[15] ^ in2[15];
    assign G[8] = in[14] & in2[14];
    assign P[8] = in[14] ^ in2[14];
    assign G[9] = in[13] & in2[13];
    assign P[9] = in[13] ^ in2[13];
    assign G[10] = in[12] & in2[12];
    assign P[10] = in[12] ^ in2[12];
    assign G[11] = in[11] & in2[11];
    assign P[11] = in[11] ^ in2[11];
    assign G[12] = in[10] & in2[10];
    assign P[12] = in[10] ^ in2[10];
    assign G[13] = in[9] & in2[9];
    assign P[13] = in[9] ^ in2[9];
    assign G[14] = in[8] & in2[8];
    assign P[14] = in[8] ^ in2[8];
    assign G[15] = in[7] & in2[7];
    assign P[15] = in[7] ^ in2[7];
    assign G[16] = in[6] & in2[6];
    assign P[16] = in[6] ^ in2[6];
    assign G[17] = in[5] & in2[5];
    assign P[17] = in[5] ^ in2[5];
    assign G[18] = in[4] & in2[4];
    assign P[18] = in[4] ^ in2[4];
    assign G[19] = in[3] & in2[3];
    assign P[19] = in[3] ^ in2[3];
    assign G[20] = in[2] & in2[2];
    assign P[20] = in[2] ^ in2[2];
    assign G[21] = in[1] & in2[1];
    assign P[21] = in[1] ^ in2[1];
    assign G[22] = in[0] & in2[0];
    assign P[22] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign C[22] = G[21] | (P[21] & C[21]);
    assign cout = G[22] | (P[22] & C[22]);
    assign sum = P ^ C;
endmodule

module CLA22(output [21:0] sum, output cout, input [21:0] in1, input [21:0] in2;

    wire[21:0] G;
    wire[21:0] C;
    wire[21:0] P;

    assign G[0] = in[21] & in2[21];
    assign P[0] = in[21] ^ in2[21];
    assign G[1] = in[20] & in2[20];
    assign P[1] = in[20] ^ in2[20];
    assign G[2] = in[19] & in2[19];
    assign P[2] = in[19] ^ in2[19];
    assign G[3] = in[18] & in2[18];
    assign P[3] = in[18] ^ in2[18];
    assign G[4] = in[17] & in2[17];
    assign P[4] = in[17] ^ in2[17];
    assign G[5] = in[16] & in2[16];
    assign P[5] = in[16] ^ in2[16];
    assign G[6] = in[15] & in2[15];
    assign P[6] = in[15] ^ in2[15];
    assign G[7] = in[14] & in2[14];
    assign P[7] = in[14] ^ in2[14];
    assign G[8] = in[13] & in2[13];
    assign P[8] = in[13] ^ in2[13];
    assign G[9] = in[12] & in2[12];
    assign P[9] = in[12] ^ in2[12];
    assign G[10] = in[11] & in2[11];
    assign P[10] = in[11] ^ in2[11];
    assign G[11] = in[10] & in2[10];
    assign P[11] = in[10] ^ in2[10];
    assign G[12] = in[9] & in2[9];
    assign P[12] = in[9] ^ in2[9];
    assign G[13] = in[8] & in2[8];
    assign P[13] = in[8] ^ in2[8];
    assign G[14] = in[7] & in2[7];
    assign P[14] = in[7] ^ in2[7];
    assign G[15] = in[6] & in2[6];
    assign P[15] = in[6] ^ in2[6];
    assign G[16] = in[5] & in2[5];
    assign P[16] = in[5] ^ in2[5];
    assign G[17] = in[4] & in2[4];
    assign P[17] = in[4] ^ in2[4];
    assign G[18] = in[3] & in2[3];
    assign P[18] = in[3] ^ in2[3];
    assign G[19] = in[2] & in2[2];
    assign P[19] = in[2] ^ in2[2];
    assign G[20] = in[1] & in2[1];
    assign P[20] = in[1] ^ in2[1];
    assign G[21] = in[0] & in2[0];
    assign P[21] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign C[21] = G[20] | (P[20] & C[20]);
    assign cout = G[21] | (P[21] & C[21]);
    assign sum = P ^ C;
endmodule

module CLA21(output [20:0] sum, output cout, input [20:0] in1, input [20:0] in2;

    wire[20:0] G;
    wire[20:0] C;
    wire[20:0] P;

    assign G[0] = in[20] & in2[20];
    assign P[0] = in[20] ^ in2[20];
    assign G[1] = in[19] & in2[19];
    assign P[1] = in[19] ^ in2[19];
    assign G[2] = in[18] & in2[18];
    assign P[2] = in[18] ^ in2[18];
    assign G[3] = in[17] & in2[17];
    assign P[3] = in[17] ^ in2[17];
    assign G[4] = in[16] & in2[16];
    assign P[4] = in[16] ^ in2[16];
    assign G[5] = in[15] & in2[15];
    assign P[5] = in[15] ^ in2[15];
    assign G[6] = in[14] & in2[14];
    assign P[6] = in[14] ^ in2[14];
    assign G[7] = in[13] & in2[13];
    assign P[7] = in[13] ^ in2[13];
    assign G[8] = in[12] & in2[12];
    assign P[8] = in[12] ^ in2[12];
    assign G[9] = in[11] & in2[11];
    assign P[9] = in[11] ^ in2[11];
    assign G[10] = in[10] & in2[10];
    assign P[10] = in[10] ^ in2[10];
    assign G[11] = in[9] & in2[9];
    assign P[11] = in[9] ^ in2[9];
    assign G[12] = in[8] & in2[8];
    assign P[12] = in[8] ^ in2[8];
    assign G[13] = in[7] & in2[7];
    assign P[13] = in[7] ^ in2[7];
    assign G[14] = in[6] & in2[6];
    assign P[14] = in[6] ^ in2[6];
    assign G[15] = in[5] & in2[5];
    assign P[15] = in[5] ^ in2[5];
    assign G[16] = in[4] & in2[4];
    assign P[16] = in[4] ^ in2[4];
    assign G[17] = in[3] & in2[3];
    assign P[17] = in[3] ^ in2[3];
    assign G[18] = in[2] & in2[2];
    assign P[18] = in[2] ^ in2[2];
    assign G[19] = in[1] & in2[1];
    assign P[19] = in[1] ^ in2[1];
    assign G[20] = in[0] & in2[0];
    assign P[20] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign C[20] = G[19] | (P[19] & C[19]);
    assign cout = G[20] | (P[20] & C[20]);
    assign sum = P ^ C;
endmodule

module CLA20(output [19:0] sum, output cout, input [19:0] in1, input [19:0] in2;

    wire[19:0] G;
    wire[19:0] C;
    wire[19:0] P;

    assign G[0] = in[19] & in2[19];
    assign P[0] = in[19] ^ in2[19];
    assign G[1] = in[18] & in2[18];
    assign P[1] = in[18] ^ in2[18];
    assign G[2] = in[17] & in2[17];
    assign P[2] = in[17] ^ in2[17];
    assign G[3] = in[16] & in2[16];
    assign P[3] = in[16] ^ in2[16];
    assign G[4] = in[15] & in2[15];
    assign P[4] = in[15] ^ in2[15];
    assign G[5] = in[14] & in2[14];
    assign P[5] = in[14] ^ in2[14];
    assign G[6] = in[13] & in2[13];
    assign P[6] = in[13] ^ in2[13];
    assign G[7] = in[12] & in2[12];
    assign P[7] = in[12] ^ in2[12];
    assign G[8] = in[11] & in2[11];
    assign P[8] = in[11] ^ in2[11];
    assign G[9] = in[10] & in2[10];
    assign P[9] = in[10] ^ in2[10];
    assign G[10] = in[9] & in2[9];
    assign P[10] = in[9] ^ in2[9];
    assign G[11] = in[8] & in2[8];
    assign P[11] = in[8] ^ in2[8];
    assign G[12] = in[7] & in2[7];
    assign P[12] = in[7] ^ in2[7];
    assign G[13] = in[6] & in2[6];
    assign P[13] = in[6] ^ in2[6];
    assign G[14] = in[5] & in2[5];
    assign P[14] = in[5] ^ in2[5];
    assign G[15] = in[4] & in2[4];
    assign P[15] = in[4] ^ in2[4];
    assign G[16] = in[3] & in2[3];
    assign P[16] = in[3] ^ in2[3];
    assign G[17] = in[2] & in2[2];
    assign P[17] = in[2] ^ in2[2];
    assign G[18] = in[1] & in2[1];
    assign P[18] = in[1] ^ in2[1];
    assign G[19] = in[0] & in2[0];
    assign P[19] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign C[19] = G[18] | (P[18] & C[18]);
    assign cout = G[19] | (P[19] & C[19]);
    assign sum = P ^ C;
endmodule

module CLA19(output [18:0] sum, output cout, input [18:0] in1, input [18:0] in2;

    wire[18:0] G;
    wire[18:0] C;
    wire[18:0] P;

    assign G[0] = in[18] & in2[18];
    assign P[0] = in[18] ^ in2[18];
    assign G[1] = in[17] & in2[17];
    assign P[1] = in[17] ^ in2[17];
    assign G[2] = in[16] & in2[16];
    assign P[2] = in[16] ^ in2[16];
    assign G[3] = in[15] & in2[15];
    assign P[3] = in[15] ^ in2[15];
    assign G[4] = in[14] & in2[14];
    assign P[4] = in[14] ^ in2[14];
    assign G[5] = in[13] & in2[13];
    assign P[5] = in[13] ^ in2[13];
    assign G[6] = in[12] & in2[12];
    assign P[6] = in[12] ^ in2[12];
    assign G[7] = in[11] & in2[11];
    assign P[7] = in[11] ^ in2[11];
    assign G[8] = in[10] & in2[10];
    assign P[8] = in[10] ^ in2[10];
    assign G[9] = in[9] & in2[9];
    assign P[9] = in[9] ^ in2[9];
    assign G[10] = in[8] & in2[8];
    assign P[10] = in[8] ^ in2[8];
    assign G[11] = in[7] & in2[7];
    assign P[11] = in[7] ^ in2[7];
    assign G[12] = in[6] & in2[6];
    assign P[12] = in[6] ^ in2[6];
    assign G[13] = in[5] & in2[5];
    assign P[13] = in[5] ^ in2[5];
    assign G[14] = in[4] & in2[4];
    assign P[14] = in[4] ^ in2[4];
    assign G[15] = in[3] & in2[3];
    assign P[15] = in[3] ^ in2[3];
    assign G[16] = in[2] & in2[2];
    assign P[16] = in[2] ^ in2[2];
    assign G[17] = in[1] & in2[1];
    assign P[17] = in[1] ^ in2[1];
    assign G[18] = in[0] & in2[0];
    assign P[18] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign C[18] = G[17] | (P[17] & C[17]);
    assign cout = G[18] | (P[18] & C[18]);
    assign sum = P ^ C;
endmodule

module CLA18(output [17:0] sum, output cout, input [17:0] in1, input [17:0] in2;

    wire[17:0] G;
    wire[17:0] C;
    wire[17:0] P;

    assign G[0] = in[17] & in2[17];
    assign P[0] = in[17] ^ in2[17];
    assign G[1] = in[16] & in2[16];
    assign P[1] = in[16] ^ in2[16];
    assign G[2] = in[15] & in2[15];
    assign P[2] = in[15] ^ in2[15];
    assign G[3] = in[14] & in2[14];
    assign P[3] = in[14] ^ in2[14];
    assign G[4] = in[13] & in2[13];
    assign P[4] = in[13] ^ in2[13];
    assign G[5] = in[12] & in2[12];
    assign P[5] = in[12] ^ in2[12];
    assign G[6] = in[11] & in2[11];
    assign P[6] = in[11] ^ in2[11];
    assign G[7] = in[10] & in2[10];
    assign P[7] = in[10] ^ in2[10];
    assign G[8] = in[9] & in2[9];
    assign P[8] = in[9] ^ in2[9];
    assign G[9] = in[8] & in2[8];
    assign P[9] = in[8] ^ in2[8];
    assign G[10] = in[7] & in2[7];
    assign P[10] = in[7] ^ in2[7];
    assign G[11] = in[6] & in2[6];
    assign P[11] = in[6] ^ in2[6];
    assign G[12] = in[5] & in2[5];
    assign P[12] = in[5] ^ in2[5];
    assign G[13] = in[4] & in2[4];
    assign P[13] = in[4] ^ in2[4];
    assign G[14] = in[3] & in2[3];
    assign P[14] = in[3] ^ in2[3];
    assign G[15] = in[2] & in2[2];
    assign P[15] = in[2] ^ in2[2];
    assign G[16] = in[1] & in2[1];
    assign P[16] = in[1] ^ in2[1];
    assign G[17] = in[0] & in2[0];
    assign P[17] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign C[17] = G[16] | (P[16] & C[16]);
    assign cout = G[17] | (P[17] & C[17]);
    assign sum = P ^ C;
endmodule

module CLA17(output [16:0] sum, output cout, input [16:0] in1, input [16:0] in2;

    wire[16:0] G;
    wire[16:0] C;
    wire[16:0] P;

    assign G[0] = in[16] & in2[16];
    assign P[0] = in[16] ^ in2[16];
    assign G[1] = in[15] & in2[15];
    assign P[1] = in[15] ^ in2[15];
    assign G[2] = in[14] & in2[14];
    assign P[2] = in[14] ^ in2[14];
    assign G[3] = in[13] & in2[13];
    assign P[3] = in[13] ^ in2[13];
    assign G[4] = in[12] & in2[12];
    assign P[4] = in[12] ^ in2[12];
    assign G[5] = in[11] & in2[11];
    assign P[5] = in[11] ^ in2[11];
    assign G[6] = in[10] & in2[10];
    assign P[6] = in[10] ^ in2[10];
    assign G[7] = in[9] & in2[9];
    assign P[7] = in[9] ^ in2[9];
    assign G[8] = in[8] & in2[8];
    assign P[8] = in[8] ^ in2[8];
    assign G[9] = in[7] & in2[7];
    assign P[9] = in[7] ^ in2[7];
    assign G[10] = in[6] & in2[6];
    assign P[10] = in[6] ^ in2[6];
    assign G[11] = in[5] & in2[5];
    assign P[11] = in[5] ^ in2[5];
    assign G[12] = in[4] & in2[4];
    assign P[12] = in[4] ^ in2[4];
    assign G[13] = in[3] & in2[3];
    assign P[13] = in[3] ^ in2[3];
    assign G[14] = in[2] & in2[2];
    assign P[14] = in[2] ^ in2[2];
    assign G[15] = in[1] & in2[1];
    assign P[15] = in[1] ^ in2[1];
    assign G[16] = in[0] & in2[0];
    assign P[16] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign C[16] = G[15] | (P[15] & C[15]);
    assign cout = G[16] | (P[16] & C[16]);
    assign sum = P ^ C;
endmodule

module CLA16(output [15:0] sum, output cout, input [15:0] in1, input [15:0] in2;

    wire[15:0] G;
    wire[15:0] C;
    wire[15:0] P;

    assign G[0] = in[15] & in2[15];
    assign P[0] = in[15] ^ in2[15];
    assign G[1] = in[14] & in2[14];
    assign P[1] = in[14] ^ in2[14];
    assign G[2] = in[13] & in2[13];
    assign P[2] = in[13] ^ in2[13];
    assign G[3] = in[12] & in2[12];
    assign P[3] = in[12] ^ in2[12];
    assign G[4] = in[11] & in2[11];
    assign P[4] = in[11] ^ in2[11];
    assign G[5] = in[10] & in2[10];
    assign P[5] = in[10] ^ in2[10];
    assign G[6] = in[9] & in2[9];
    assign P[6] = in[9] ^ in2[9];
    assign G[7] = in[8] & in2[8];
    assign P[7] = in[8] ^ in2[8];
    assign G[8] = in[7] & in2[7];
    assign P[8] = in[7] ^ in2[7];
    assign G[9] = in[6] & in2[6];
    assign P[9] = in[6] ^ in2[6];
    assign G[10] = in[5] & in2[5];
    assign P[10] = in[5] ^ in2[5];
    assign G[11] = in[4] & in2[4];
    assign P[11] = in[4] ^ in2[4];
    assign G[12] = in[3] & in2[3];
    assign P[12] = in[3] ^ in2[3];
    assign G[13] = in[2] & in2[2];
    assign P[13] = in[2] ^ in2[2];
    assign G[14] = in[1] & in2[1];
    assign P[14] = in[1] ^ in2[1];
    assign G[15] = in[0] & in2[0];
    assign P[15] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign C[15] = G[14] | (P[14] & C[14]);
    assign cout = G[15] | (P[15] & C[15]);
    assign sum = P ^ C;
endmodule

module CLA15(output [14:0] sum, output cout, input [14:0] in1, input [14:0] in2;

    wire[14:0] G;
    wire[14:0] C;
    wire[14:0] P;

    assign G[0] = in[14] & in2[14];
    assign P[0] = in[14] ^ in2[14];
    assign G[1] = in[13] & in2[13];
    assign P[1] = in[13] ^ in2[13];
    assign G[2] = in[12] & in2[12];
    assign P[2] = in[12] ^ in2[12];
    assign G[3] = in[11] & in2[11];
    assign P[3] = in[11] ^ in2[11];
    assign G[4] = in[10] & in2[10];
    assign P[4] = in[10] ^ in2[10];
    assign G[5] = in[9] & in2[9];
    assign P[5] = in[9] ^ in2[9];
    assign G[6] = in[8] & in2[8];
    assign P[6] = in[8] ^ in2[8];
    assign G[7] = in[7] & in2[7];
    assign P[7] = in[7] ^ in2[7];
    assign G[8] = in[6] & in2[6];
    assign P[8] = in[6] ^ in2[6];
    assign G[9] = in[5] & in2[5];
    assign P[9] = in[5] ^ in2[5];
    assign G[10] = in[4] & in2[4];
    assign P[10] = in[4] ^ in2[4];
    assign G[11] = in[3] & in2[3];
    assign P[11] = in[3] ^ in2[3];
    assign G[12] = in[2] & in2[2];
    assign P[12] = in[2] ^ in2[2];
    assign G[13] = in[1] & in2[1];
    assign P[13] = in[1] ^ in2[1];
    assign G[14] = in[0] & in2[0];
    assign P[14] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign C[14] = G[13] | (P[13] & C[13]);
    assign cout = G[14] | (P[14] & C[14]);
    assign sum = P ^ C;
endmodule

module CLA14(output [13:0] sum, output cout, input [13:0] in1, input [13:0] in2;

    wire[13:0] G;
    wire[13:0] C;
    wire[13:0] P;

    assign G[0] = in[13] & in2[13];
    assign P[0] = in[13] ^ in2[13];
    assign G[1] = in[12] & in2[12];
    assign P[1] = in[12] ^ in2[12];
    assign G[2] = in[11] & in2[11];
    assign P[2] = in[11] ^ in2[11];
    assign G[3] = in[10] & in2[10];
    assign P[3] = in[10] ^ in2[10];
    assign G[4] = in[9] & in2[9];
    assign P[4] = in[9] ^ in2[9];
    assign G[5] = in[8] & in2[8];
    assign P[5] = in[8] ^ in2[8];
    assign G[6] = in[7] & in2[7];
    assign P[6] = in[7] ^ in2[7];
    assign G[7] = in[6] & in2[6];
    assign P[7] = in[6] ^ in2[6];
    assign G[8] = in[5] & in2[5];
    assign P[8] = in[5] ^ in2[5];
    assign G[9] = in[4] & in2[4];
    assign P[9] = in[4] ^ in2[4];
    assign G[10] = in[3] & in2[3];
    assign P[10] = in[3] ^ in2[3];
    assign G[11] = in[2] & in2[2];
    assign P[11] = in[2] ^ in2[2];
    assign G[12] = in[1] & in2[1];
    assign P[12] = in[1] ^ in2[1];
    assign G[13] = in[0] & in2[0];
    assign P[13] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign C[13] = G[12] | (P[12] & C[12]);
    assign cout = G[13] | (P[13] & C[13]);
    assign sum = P ^ C;
endmodule

module CLA13(output [12:0] sum, output cout, input [12:0] in1, input [12:0] in2;

    wire[12:0] G;
    wire[12:0] C;
    wire[12:0] P;

    assign G[0] = in[12] & in2[12];
    assign P[0] = in[12] ^ in2[12];
    assign G[1] = in[11] & in2[11];
    assign P[1] = in[11] ^ in2[11];
    assign G[2] = in[10] & in2[10];
    assign P[2] = in[10] ^ in2[10];
    assign G[3] = in[9] & in2[9];
    assign P[3] = in[9] ^ in2[9];
    assign G[4] = in[8] & in2[8];
    assign P[4] = in[8] ^ in2[8];
    assign G[5] = in[7] & in2[7];
    assign P[5] = in[7] ^ in2[7];
    assign G[6] = in[6] & in2[6];
    assign P[6] = in[6] ^ in2[6];
    assign G[7] = in[5] & in2[5];
    assign P[7] = in[5] ^ in2[5];
    assign G[8] = in[4] & in2[4];
    assign P[8] = in[4] ^ in2[4];
    assign G[9] = in[3] & in2[3];
    assign P[9] = in[3] ^ in2[3];
    assign G[10] = in[2] & in2[2];
    assign P[10] = in[2] ^ in2[2];
    assign G[11] = in[1] & in2[1];
    assign P[11] = in[1] ^ in2[1];
    assign G[12] = in[0] & in2[0];
    assign P[12] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign C[12] = G[11] | (P[11] & C[11]);
    assign cout = G[12] | (P[12] & C[12]);
    assign sum = P ^ C;
endmodule

module CLA12(output [11:0] sum, output cout, input [11:0] in1, input [11:0] in2;

    wire[11:0] G;
    wire[11:0] C;
    wire[11:0] P;

    assign G[0] = in[11] & in2[11];
    assign P[0] = in[11] ^ in2[11];
    assign G[1] = in[10] & in2[10];
    assign P[1] = in[10] ^ in2[10];
    assign G[2] = in[9] & in2[9];
    assign P[2] = in[9] ^ in2[9];
    assign G[3] = in[8] & in2[8];
    assign P[3] = in[8] ^ in2[8];
    assign G[4] = in[7] & in2[7];
    assign P[4] = in[7] ^ in2[7];
    assign G[5] = in[6] & in2[6];
    assign P[5] = in[6] ^ in2[6];
    assign G[6] = in[5] & in2[5];
    assign P[6] = in[5] ^ in2[5];
    assign G[7] = in[4] & in2[4];
    assign P[7] = in[4] ^ in2[4];
    assign G[8] = in[3] & in2[3];
    assign P[8] = in[3] ^ in2[3];
    assign G[9] = in[2] & in2[2];
    assign P[9] = in[2] ^ in2[2];
    assign G[10] = in[1] & in2[1];
    assign P[10] = in[1] ^ in2[1];
    assign G[11] = in[0] & in2[0];
    assign P[11] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign C[11] = G[10] | (P[10] & C[10]);
    assign cout = G[11] | (P[11] & C[11]);
    assign sum = P ^ C;
endmodule

module CLA11(output [10:0] sum, output cout, input [10:0] in1, input [10:0] in2;

    wire[10:0] G;
    wire[10:0] C;
    wire[10:0] P;

    assign G[0] = in[10] & in2[10];
    assign P[0] = in[10] ^ in2[10];
    assign G[1] = in[9] & in2[9];
    assign P[1] = in[9] ^ in2[9];
    assign G[2] = in[8] & in2[8];
    assign P[2] = in[8] ^ in2[8];
    assign G[3] = in[7] & in2[7];
    assign P[3] = in[7] ^ in2[7];
    assign G[4] = in[6] & in2[6];
    assign P[4] = in[6] ^ in2[6];
    assign G[5] = in[5] & in2[5];
    assign P[5] = in[5] ^ in2[5];
    assign G[6] = in[4] & in2[4];
    assign P[6] = in[4] ^ in2[4];
    assign G[7] = in[3] & in2[3];
    assign P[7] = in[3] ^ in2[3];
    assign G[8] = in[2] & in2[2];
    assign P[8] = in[2] ^ in2[2];
    assign G[9] = in[1] & in2[1];
    assign P[9] = in[1] ^ in2[1];
    assign G[10] = in[0] & in2[0];
    assign P[10] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign C[10] = G[9] | (P[9] & C[9]);
    assign cout = G[10] | (P[10] & C[10]);
    assign sum = P ^ C;
endmodule

module CLA10(output [9:0] sum, output cout, input [9:0] in1, input [9:0] in2;

    wire[9:0] G;
    wire[9:0] C;
    wire[9:0] P;

    assign G[0] = in[9] & in2[9];
    assign P[0] = in[9] ^ in2[9];
    assign G[1] = in[8] & in2[8];
    assign P[1] = in[8] ^ in2[8];
    assign G[2] = in[7] & in2[7];
    assign P[2] = in[7] ^ in2[7];
    assign G[3] = in[6] & in2[6];
    assign P[3] = in[6] ^ in2[6];
    assign G[4] = in[5] & in2[5];
    assign P[4] = in[5] ^ in2[5];
    assign G[5] = in[4] & in2[4];
    assign P[5] = in[4] ^ in2[4];
    assign G[6] = in[3] & in2[3];
    assign P[6] = in[3] ^ in2[3];
    assign G[7] = in[2] & in2[2];
    assign P[7] = in[2] ^ in2[2];
    assign G[8] = in[1] & in2[1];
    assign P[8] = in[1] ^ in2[1];
    assign G[9] = in[0] & in2[0];
    assign P[9] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign C[9] = G[8] | (P[8] & C[8]);
    assign cout = G[9] | (P[9] & C[9]);
    assign sum = P ^ C;
endmodule

module CLA9(output [8:0] sum, output cout, input [8:0] in1, input [8:0] in2;

    wire[8:0] G;
    wire[8:0] C;
    wire[8:0] P;

    assign G[0] = in[8] & in2[8];
    assign P[0] = in[8] ^ in2[8];
    assign G[1] = in[7] & in2[7];
    assign P[1] = in[7] ^ in2[7];
    assign G[2] = in[6] & in2[6];
    assign P[2] = in[6] ^ in2[6];
    assign G[3] = in[5] & in2[5];
    assign P[3] = in[5] ^ in2[5];
    assign G[4] = in[4] & in2[4];
    assign P[4] = in[4] ^ in2[4];
    assign G[5] = in[3] & in2[3];
    assign P[5] = in[3] ^ in2[3];
    assign G[6] = in[2] & in2[2];
    assign P[6] = in[2] ^ in2[2];
    assign G[7] = in[1] & in2[1];
    assign P[7] = in[1] ^ in2[1];
    assign G[8] = in[0] & in2[0];
    assign P[8] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign C[8] = G[7] | (P[7] & C[7]);
    assign cout = G[8] | (P[8] & C[8]);
    assign sum = P ^ C;
endmodule

module CLA8(output [7:0] sum, output cout, input [7:0] in1, input [7:0] in2;

    wire[7:0] G;
    wire[7:0] C;
    wire[7:0] P;

    assign G[0] = in[7] & in2[7];
    assign P[0] = in[7] ^ in2[7];
    assign G[1] = in[6] & in2[6];
    assign P[1] = in[6] ^ in2[6];
    assign G[2] = in[5] & in2[5];
    assign P[2] = in[5] ^ in2[5];
    assign G[3] = in[4] & in2[4];
    assign P[3] = in[4] ^ in2[4];
    assign G[4] = in[3] & in2[3];
    assign P[4] = in[3] ^ in2[3];
    assign G[5] = in[2] & in2[2];
    assign P[5] = in[2] ^ in2[2];
    assign G[6] = in[1] & in2[1];
    assign P[6] = in[1] ^ in2[1];
    assign G[7] = in[0] & in2[0];
    assign P[7] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign C[7] = G[6] | (P[6] & C[6]);
    assign cout = G[7] | (P[7] & C[7]);
    assign sum = P ^ C;
endmodule

module CLA7(output [6:0] sum, output cout, input [6:0] in1, input [6:0] in2;

    wire[6:0] G;
    wire[6:0] C;
    wire[6:0] P;

    assign G[0] = in[6] & in2[6];
    assign P[0] = in[6] ^ in2[6];
    assign G[1] = in[5] & in2[5];
    assign P[1] = in[5] ^ in2[5];
    assign G[2] = in[4] & in2[4];
    assign P[2] = in[4] ^ in2[4];
    assign G[3] = in[3] & in2[3];
    assign P[3] = in[3] ^ in2[3];
    assign G[4] = in[2] & in2[2];
    assign P[4] = in[2] ^ in2[2];
    assign G[5] = in[1] & in2[1];
    assign P[5] = in[1] ^ in2[1];
    assign G[6] = in[0] & in2[0];
    assign P[6] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign C[6] = G[5] | (P[5] & C[5]);
    assign cout = G[6] | (P[6] & C[6]);
    assign sum = P ^ C;
endmodule

module CLA6(output [5:0] sum, output cout, input [5:0] in1, input [5:0] in2;

    wire[5:0] G;
    wire[5:0] C;
    wire[5:0] P;

    assign G[0] = in[5] & in2[5];
    assign P[0] = in[5] ^ in2[5];
    assign G[1] = in[4] & in2[4];
    assign P[1] = in[4] ^ in2[4];
    assign G[2] = in[3] & in2[3];
    assign P[2] = in[3] ^ in2[3];
    assign G[3] = in[2] & in2[2];
    assign P[3] = in[2] ^ in2[2];
    assign G[4] = in[1] & in2[1];
    assign P[4] = in[1] ^ in2[1];
    assign G[5] = in[0] & in2[0];
    assign P[5] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign C[5] = G[4] | (P[4] & C[4]);
    assign cout = G[5] | (P[5] & C[5]);
    assign sum = P ^ C;
endmodule

module CLA5(output [4:0] sum, output cout, input [4:0] in1, input [4:0] in2;

    wire[4:0] G;
    wire[4:0] C;
    wire[4:0] P;

    assign G[0] = in[4] & in2[4];
    assign P[0] = in[4] ^ in2[4];
    assign G[1] = in[3] & in2[3];
    assign P[1] = in[3] ^ in2[3];
    assign G[2] = in[2] & in2[2];
    assign P[2] = in[2] ^ in2[2];
    assign G[3] = in[1] & in2[1];
    assign P[3] = in[1] ^ in2[1];
    assign G[4] = in[0] & in2[0];
    assign P[4] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign C[4] = G[3] | (P[3] & C[3]);
    assign cout = G[4] | (P[4] & C[4]);
    assign sum = P ^ C;
endmodule

module CLA4(output [3:0] sum, output cout, input [3:0] in1, input [3:0] in2;

    wire[3:0] G;
    wire[3:0] C;
    wire[3:0] P;

    assign G[0] = in[3] & in2[3];
    assign P[0] = in[3] ^ in2[3];
    assign G[1] = in[2] & in2[2];
    assign P[1] = in[2] ^ in2[2];
    assign G[2] = in[1] & in2[1];
    assign P[2] = in[1] ^ in2[1];
    assign G[3] = in[0] & in2[0];
    assign P[3] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign C[3] = G[2] | (P[2] & C[2]);
    assign cout = G[3] | (P[3] & C[3]);
    assign sum = P ^ C;
endmodule

module CLA3(output [2:0] sum, output cout, input [2:0] in1, input [2:0] in2;

    wire[2:0] G;
    wire[2:0] C;
    wire[2:0] P;

    assign G[0] = in[2] & in2[2];
    assign P[0] = in[2] ^ in2[2];
    assign G[1] = in[1] & in2[1];
    assign P[1] = in[1] ^ in2[1];
    assign G[2] = in[0] & in2[0];
    assign P[2] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign C[2] = G[1] | (P[1] & C[1]);
    assign cout = G[2] | (P[2] & C[2]);
    assign sum = P ^ C;
endmodule

module CLA2(output [1:0] sum, output cout, input [1:0] in1, input [1:0] in2;

    wire[1:0] G;
    wire[1:0] C;
    wire[1:0] P;

    assign G[0] = in[1] & in2[1];
    assign P[0] = in[1] ^ in2[1];
    assign G[1] = in[0] & in2[0];
    assign P[1] = in[0] ^ in2[0];


    assign C[0] = 0;  /* Carry_out = Ci+1 = Gi + Pi*Ci */;
    assign C[1] = G[0] | (P[0] & C[0]);
    assign cout = G[1] | (P[1] & C[1]);
    assign sum = P ^ C;
endmodule

