module wallace_unsigned_multiplier_RCA_32(product, A, B);
    input [31:0] A, B;
    output [63:0] product;

wire [31:0] pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10, pp11, pp12, pp13, pp14, pp15;
wire [31:0] pp16, pp17, pp18, pp19, pp20, pp21, pp22, pp23, pp24, pp25, pp26, pp27, pp28, pp29, pp30, pp31;

assign P[0][0] = x[0] & y[0];
assign P[0][1] = x[0] & y[1];
assign P[0][2] = x[0] & y[2];
assign P[0][3] = x[0] & y[3];
assign P[0][4] = x[0] & y[4];
assign P[0][5] = x[0] & y[5];
assign P[0][6] = x[0] & y[6];
assign P[0][7] = x[0] & y[7];
assign P[0][8] = x[0] & y[8];
assign P[0][9] = x[0] & y[9];
assign P[0][10] = x[0] & y[10];
assign P[0][11] = x[0] & y[11];
assign P[0][12] = x[0] & y[12];
assign P[0][13] = x[0] & y[13];
assign P[0][14] = x[0] & y[14];
assign P[0][15] = x[0] & y[15];
assign P[0][16] = x[0] & y[16];
assign P[0][17] = x[0] & y[17];
assign P[0][18] = x[0] & y[18];
assign P[0][19] = x[0] & y[19];
assign P[0][20] = x[0] & y[20];
assign P[0][21] = x[0] & y[21];
assign P[0][22] = x[0] & y[22];
assign P[0][23] = x[0] & y[23];
assign P[0][24] = x[0] & y[24];
assign P[0][25] = x[0] & y[25];
assign P[0][26] = x[0] & y[26];
assign P[0][27] = x[0] & y[27];
assign P[0][28] = x[0] & y[28];
assign P[0][29] = x[0] & y[29];
assign P[0][30] = x[0] & y[30];
assign P[0][31] = x[0] & y[31];
assign P[1][0] = x[1] & y[0];
assign P[1][1] = x[1] & y[1];
assign P[1][2] = x[1] & y[2];
assign P[1][3] = x[1] & y[3];
assign P[1][4] = x[1] & y[4];
assign P[1][5] = x[1] & y[5];
assign P[1][6] = x[1] & y[6];
assign P[1][7] = x[1] & y[7];
assign P[1][8] = x[1] & y[8];
assign P[1][9] = x[1] & y[9];
assign P[1][10] = x[1] & y[10];
assign P[1][11] = x[1] & y[11];
assign P[1][12] = x[1] & y[12];
assign P[1][13] = x[1] & y[13];
assign P[1][14] = x[1] & y[14];
assign P[1][15] = x[1] & y[15];
assign P[1][16] = x[1] & y[16];
assign P[1][17] = x[1] & y[17];
assign P[1][18] = x[1] & y[18];
assign P[1][19] = x[1] & y[19];
assign P[1][20] = x[1] & y[20];
assign P[1][21] = x[1] & y[21];
assign P[1][22] = x[1] & y[22];
assign P[1][23] = x[1] & y[23];
assign P[1][24] = x[1] & y[24];
assign P[1][25] = x[1] & y[25];
assign P[1][26] = x[1] & y[26];
assign P[1][27] = x[1] & y[27];
assign P[1][28] = x[1] & y[28];
assign P[1][29] = x[1] & y[29];
assign P[1][30] = x[1] & y[30];
assign P[1][31] = x[1] & y[31];
assign P[2][0] = x[2] & y[0];
assign P[2][1] = x[2] & y[1];
assign P[2][2] = x[2] & y[2];
assign P[2][3] = x[2] & y[3];
assign P[2][4] = x[2] & y[4];
assign P[2][5] = x[2] & y[5];
assign P[2][6] = x[2] & y[6];
assign P[2][7] = x[2] & y[7];
assign P[2][8] = x[2] & y[8];
assign P[2][9] = x[2] & y[9];
assign P[2][10] = x[2] & y[10];
assign P[2][11] = x[2] & y[11];
assign P[2][12] = x[2] & y[12];
assign P[2][13] = x[2] & y[13];
assign P[2][14] = x[2] & y[14];
assign P[2][15] = x[2] & y[15];
assign P[2][16] = x[2] & y[16];
assign P[2][17] = x[2] & y[17];
assign P[2][18] = x[2] & y[18];
assign P[2][19] = x[2] & y[19];
assign P[2][20] = x[2] & y[20];
assign P[2][21] = x[2] & y[21];
assign P[2][22] = x[2] & y[22];
assign P[2][23] = x[2] & y[23];
assign P[2][24] = x[2] & y[24];
assign P[2][25] = x[2] & y[25];
assign P[2][26] = x[2] & y[26];
assign P[2][27] = x[2] & y[27];
assign P[2][28] = x[2] & y[28];
assign P[2][29] = x[2] & y[29];
assign P[2][30] = x[2] & y[30];
assign P[2][31] = x[2] & y[31];
assign P[3][0] = x[3] & y[0];
assign P[3][1] = x[3] & y[1];
assign P[3][2] = x[3] & y[2];
assign P[3][3] = x[3] & y[3];
assign P[3][4] = x[3] & y[4];
assign P[3][5] = x[3] & y[5];
assign P[3][6] = x[3] & y[6];
assign P[3][7] = x[3] & y[7];
assign P[3][8] = x[3] & y[8];
assign P[3][9] = x[3] & y[9];
assign P[3][10] = x[3] & y[10];
assign P[3][11] = x[3] & y[11];
assign P[3][12] = x[3] & y[12];
assign P[3][13] = x[3] & y[13];
assign P[3][14] = x[3] & y[14];
assign P[3][15] = x[3] & y[15];
assign P[3][16] = x[3] & y[16];
assign P[3][17] = x[3] & y[17];
assign P[3][18] = x[3] & y[18];
assign P[3][19] = x[3] & y[19];
assign P[3][20] = x[3] & y[20];
assign P[3][21] = x[3] & y[21];
assign P[3][22] = x[3] & y[22];
assign P[3][23] = x[3] & y[23];
assign P[3][24] = x[3] & y[24];
assign P[3][25] = x[3] & y[25];
assign P[3][26] = x[3] & y[26];
assign P[3][27] = x[3] & y[27];
assign P[3][28] = x[3] & y[28];
assign P[3][29] = x[3] & y[29];
assign P[3][30] = x[3] & y[30];
assign P[3][31] = x[3] & y[31];
assign P[4][0] = x[4] & y[0];
assign P[4][1] = x[4] & y[1];
assign P[4][2] = x[4] & y[2];
assign P[4][3] = x[4] & y[3];
assign P[4][4] = x[4] & y[4];
assign P[4][5] = x[4] & y[5];
assign P[4][6] = x[4] & y[6];
assign P[4][7] = x[4] & y[7];
assign P[4][8] = x[4] & y[8];
assign P[4][9] = x[4] & y[9];
assign P[4][10] = x[4] & y[10];
assign P[4][11] = x[4] & y[11];
assign P[4][12] = x[4] & y[12];
assign P[4][13] = x[4] & y[13];
assign P[4][14] = x[4] & y[14];
assign P[4][15] = x[4] & y[15];
assign P[4][16] = x[4] & y[16];
assign P[4][17] = x[4] & y[17];
assign P[4][18] = x[4] & y[18];
assign P[4][19] = x[4] & y[19];
assign P[4][20] = x[4] & y[20];
assign P[4][21] = x[4] & y[21];
assign P[4][22] = x[4] & y[22];
assign P[4][23] = x[4] & y[23];
assign P[4][24] = x[4] & y[24];
assign P[4][25] = x[4] & y[25];
assign P[4][26] = x[4] & y[26];
assign P[4][27] = x[4] & y[27];
assign P[4][28] = x[4] & y[28];
assign P[4][29] = x[4] & y[29];
assign P[4][30] = x[4] & y[30];
assign P[4][31] = x[4] & y[31];
assign P[5][0] = x[5] & y[0];
assign P[5][1] = x[5] & y[1];
assign P[5][2] = x[5] & y[2];
assign P[5][3] = x[5] & y[3];
assign P[5][4] = x[5] & y[4];
assign P[5][5] = x[5] & y[5];
assign P[5][6] = x[5] & y[6];
assign P[5][7] = x[5] & y[7];
assign P[5][8] = x[5] & y[8];
assign P[5][9] = x[5] & y[9];
assign P[5][10] = x[5] & y[10];
assign P[5][11] = x[5] & y[11];
assign P[5][12] = x[5] & y[12];
assign P[5][13] = x[5] & y[13];
assign P[5][14] = x[5] & y[14];
assign P[5][15] = x[5] & y[15];
assign P[5][16] = x[5] & y[16];
assign P[5][17] = x[5] & y[17];
assign P[5][18] = x[5] & y[18];
assign P[5][19] = x[5] & y[19];
assign P[5][20] = x[5] & y[20];
assign P[5][21] = x[5] & y[21];
assign P[5][22] = x[5] & y[22];
assign P[5][23] = x[5] & y[23];
assign P[5][24] = x[5] & y[24];
assign P[5][25] = x[5] & y[25];
assign P[5][26] = x[5] & y[26];
assign P[5][27] = x[5] & y[27];
assign P[5][28] = x[5] & y[28];
assign P[5][29] = x[5] & y[29];
assign P[5][30] = x[5] & y[30];
assign P[5][31] = x[5] & y[31];
assign P[6][0] = x[6] & y[0];
assign P[6][1] = x[6] & y[1];
assign P[6][2] = x[6] & y[2];
assign P[6][3] = x[6] & y[3];
assign P[6][4] = x[6] & y[4];
assign P[6][5] = x[6] & y[5];
assign P[6][6] = x[6] & y[6];
assign P[6][7] = x[6] & y[7];
assign P[6][8] = x[6] & y[8];
assign P[6][9] = x[6] & y[9];
assign P[6][10] = x[6] & y[10];
assign P[6][11] = x[6] & y[11];
assign P[6][12] = x[6] & y[12];
assign P[6][13] = x[6] & y[13];
assign P[6][14] = x[6] & y[14];
assign P[6][15] = x[6] & y[15];
assign P[6][16] = x[6] & y[16];
assign P[6][17] = x[6] & y[17];
assign P[6][18] = x[6] & y[18];
assign P[6][19] = x[6] & y[19];
assign P[6][20] = x[6] & y[20];
assign P[6][21] = x[6] & y[21];
assign P[6][22] = x[6] & y[22];
assign P[6][23] = x[6] & y[23];
assign P[6][24] = x[6] & y[24];
assign P[6][25] = x[6] & y[25];
assign P[6][26] = x[6] & y[26];
assign P[6][27] = x[6] & y[27];
assign P[6][28] = x[6] & y[28];
assign P[6][29] = x[6] & y[29];
assign P[6][30] = x[6] & y[30];
assign P[6][31] = x[6] & y[31];
assign P[7][0] = x[7] & y[0];
assign P[7][1] = x[7] & y[1];
assign P[7][2] = x[7] & y[2];
assign P[7][3] = x[7] & y[3];
assign P[7][4] = x[7] & y[4];
assign P[7][5] = x[7] & y[5];
assign P[7][6] = x[7] & y[6];
assign P[7][7] = x[7] & y[7];
assign P[7][8] = x[7] & y[8];
assign P[7][9] = x[7] & y[9];
assign P[7][10] = x[7] & y[10];
assign P[7][11] = x[7] & y[11];
assign P[7][12] = x[7] & y[12];
assign P[7][13] = x[7] & y[13];
assign P[7][14] = x[7] & y[14];
assign P[7][15] = x[7] & y[15];
assign P[7][16] = x[7] & y[16];
assign P[7][17] = x[7] & y[17];
assign P[7][18] = x[7] & y[18];
assign P[7][19] = x[7] & y[19];
assign P[7][20] = x[7] & y[20];
assign P[7][21] = x[7] & y[21];
assign P[7][22] = x[7] & y[22];
assign P[7][23] = x[7] & y[23];
assign P[7][24] = x[7] & y[24];
assign P[7][25] = x[7] & y[25];
assign P[7][26] = x[7] & y[26];
assign P[7][27] = x[7] & y[27];
assign P[7][28] = x[7] & y[28];
assign P[7][29] = x[7] & y[29];
assign P[7][30] = x[7] & y[30];
assign P[7][31] = x[7] & y[31];
assign P[8][0] = x[8] & y[0];
assign P[8][1] = x[8] & y[1];
assign P[8][2] = x[8] & y[2];
assign P[8][3] = x[8] & y[3];
assign P[8][4] = x[8] & y[4];
assign P[8][5] = x[8] & y[5];
assign P[8][6] = x[8] & y[6];
assign P[8][7] = x[8] & y[7];
assign P[8][8] = x[8] & y[8];
assign P[8][9] = x[8] & y[9];
assign P[8][10] = x[8] & y[10];
assign P[8][11] = x[8] & y[11];
assign P[8][12] = x[8] & y[12];
assign P[8][13] = x[8] & y[13];
assign P[8][14] = x[8] & y[14];
assign P[8][15] = x[8] & y[15];
assign P[8][16] = x[8] & y[16];
assign P[8][17] = x[8] & y[17];
assign P[8][18] = x[8] & y[18];
assign P[8][19] = x[8] & y[19];
assign P[8][20] = x[8] & y[20];
assign P[8][21] = x[8] & y[21];
assign P[8][22] = x[8] & y[22];
assign P[8][23] = x[8] & y[23];
assign P[8][24] = x[8] & y[24];
assign P[8][25] = x[8] & y[25];
assign P[8][26] = x[8] & y[26];
assign P[8][27] = x[8] & y[27];
assign P[8][28] = x[8] & y[28];
assign P[8][29] = x[8] & y[29];
assign P[8][30] = x[8] & y[30];
assign P[8][31] = x[8] & y[31];
assign P[9][0] = x[9] & y[0];
assign P[9][1] = x[9] & y[1];
assign P[9][2] = x[9] & y[2];
assign P[9][3] = x[9] & y[3];
assign P[9][4] = x[9] & y[4];
assign P[9][5] = x[9] & y[5];
assign P[9][6] = x[9] & y[6];
assign P[9][7] = x[9] & y[7];
assign P[9][8] = x[9] & y[8];
assign P[9][9] = x[9] & y[9];
assign P[9][10] = x[9] & y[10];
assign P[9][11] = x[9] & y[11];
assign P[9][12] = x[9] & y[12];
assign P[9][13] = x[9] & y[13];
assign P[9][14] = x[9] & y[14];
assign P[9][15] = x[9] & y[15];
assign P[9][16] = x[9] & y[16];
assign P[9][17] = x[9] & y[17];
assign P[9][18] = x[9] & y[18];
assign P[9][19] = x[9] & y[19];
assign P[9][20] = x[9] & y[20];
assign P[9][21] = x[9] & y[21];
assign P[9][22] = x[9] & y[22];
assign P[9][23] = x[9] & y[23];
assign P[9][24] = x[9] & y[24];
assign P[9][25] = x[9] & y[25];
assign P[9][26] = x[9] & y[26];
assign P[9][27] = x[9] & y[27];
assign P[9][28] = x[9] & y[28];
assign P[9][29] = x[9] & y[29];
assign P[9][30] = x[9] & y[30];
assign P[9][31] = x[9] & y[31];
assign P[10][0] = x[10] & y[0];
assign P[10][1] = x[10] & y[1];
assign P[10][2] = x[10] & y[2];
assign P[10][3] = x[10] & y[3];
assign P[10][4] = x[10] & y[4];
assign P[10][5] = x[10] & y[5];
assign P[10][6] = x[10] & y[6];
assign P[10][7] = x[10] & y[7];
assign P[10][8] = x[10] & y[8];
assign P[10][9] = x[10] & y[9];
assign P[10][10] = x[10] & y[10];
assign P[10][11] = x[10] & y[11];
assign P[10][12] = x[10] & y[12];
assign P[10][13] = x[10] & y[13];
assign P[10][14] = x[10] & y[14];
assign P[10][15] = x[10] & y[15];
assign P[10][16] = x[10] & y[16];
assign P[10][17] = x[10] & y[17];
assign P[10][18] = x[10] & y[18];
assign P[10][19] = x[10] & y[19];
assign P[10][20] = x[10] & y[20];
assign P[10][21] = x[10] & y[21];
assign P[10][22] = x[10] & y[22];
assign P[10][23] = x[10] & y[23];
assign P[10][24] = x[10] & y[24];
assign P[10][25] = x[10] & y[25];
assign P[10][26] = x[10] & y[26];
assign P[10][27] = x[10] & y[27];
assign P[10][28] = x[10] & y[28];
assign P[10][29] = x[10] & y[29];
assign P[10][30] = x[10] & y[30];
assign P[10][31] = x[10] & y[31];
assign P[11][0] = x[11] & y[0];
assign P[11][1] = x[11] & y[1];
assign P[11][2] = x[11] & y[2];
assign P[11][3] = x[11] & y[3];
assign P[11][4] = x[11] & y[4];
assign P[11][5] = x[11] & y[5];
assign P[11][6] = x[11] & y[6];
assign P[11][7] = x[11] & y[7];
assign P[11][8] = x[11] & y[8];
assign P[11][9] = x[11] & y[9];
assign P[11][10] = x[11] & y[10];
assign P[11][11] = x[11] & y[11];
assign P[11][12] = x[11] & y[12];
assign P[11][13] = x[11] & y[13];
assign P[11][14] = x[11] & y[14];
assign P[11][15] = x[11] & y[15];
assign P[11][16] = x[11] & y[16];
assign P[11][17] = x[11] & y[17];
assign P[11][18] = x[11] & y[18];
assign P[11][19] = x[11] & y[19];
assign P[11][20] = x[11] & y[20];
assign P[11][21] = x[11] & y[21];
assign P[11][22] = x[11] & y[22];
assign P[11][23] = x[11] & y[23];
assign P[11][24] = x[11] & y[24];
assign P[11][25] = x[11] & y[25];
assign P[11][26] = x[11] & y[26];
assign P[11][27] = x[11] & y[27];
assign P[11][28] = x[11] & y[28];
assign P[11][29] = x[11] & y[29];
assign P[11][30] = x[11] & y[30];
assign P[11][31] = x[11] & y[31];
assign P[12][0] = x[12] & y[0];
assign P[12][1] = x[12] & y[1];
assign P[12][2] = x[12] & y[2];
assign P[12][3] = x[12] & y[3];
assign P[12][4] = x[12] & y[4];
assign P[12][5] = x[12] & y[5];
assign P[12][6] = x[12] & y[6];
assign P[12][7] = x[12] & y[7];
assign P[12][8] = x[12] & y[8];
assign P[12][9] = x[12] & y[9];
assign P[12][10] = x[12] & y[10];
assign P[12][11] = x[12] & y[11];
assign P[12][12] = x[12] & y[12];
assign P[12][13] = x[12] & y[13];
assign P[12][14] = x[12] & y[14];
assign P[12][15] = x[12] & y[15];
assign P[12][16] = x[12] & y[16];
assign P[12][17] = x[12] & y[17];
assign P[12][18] = x[12] & y[18];
assign P[12][19] = x[12] & y[19];
assign P[12][20] = x[12] & y[20];
assign P[12][21] = x[12] & y[21];
assign P[12][22] = x[12] & y[22];
assign P[12][23] = x[12] & y[23];
assign P[12][24] = x[12] & y[24];
assign P[12][25] = x[12] & y[25];
assign P[12][26] = x[12] & y[26];
assign P[12][27] = x[12] & y[27];
assign P[12][28] = x[12] & y[28];
assign P[12][29] = x[12] & y[29];
assign P[12][30] = x[12] & y[30];
assign P[12][31] = x[12] & y[31];
assign P[13][0] = x[13] & y[0];
assign P[13][1] = x[13] & y[1];
assign P[13][2] = x[13] & y[2];
assign P[13][3] = x[13] & y[3];
assign P[13][4] = x[13] & y[4];
assign P[13][5] = x[13] & y[5];
assign P[13][6] = x[13] & y[6];
assign P[13][7] = x[13] & y[7];
assign P[13][8] = x[13] & y[8];
assign P[13][9] = x[13] & y[9];
assign P[13][10] = x[13] & y[10];
assign P[13][11] = x[13] & y[11];
assign P[13][12] = x[13] & y[12];
assign P[13][13] = x[13] & y[13];
assign P[13][14] = x[13] & y[14];
assign P[13][15] = x[13] & y[15];
assign P[13][16] = x[13] & y[16];
assign P[13][17] = x[13] & y[17];
assign P[13][18] = x[13] & y[18];
assign P[13][19] = x[13] & y[19];
assign P[13][20] = x[13] & y[20];
assign P[13][21] = x[13] & y[21];
assign P[13][22] = x[13] & y[22];
assign P[13][23] = x[13] & y[23];
assign P[13][24] = x[13] & y[24];
assign P[13][25] = x[13] & y[25];
assign P[13][26] = x[13] & y[26];
assign P[13][27] = x[13] & y[27];
assign P[13][28] = x[13] & y[28];
assign P[13][29] = x[13] & y[29];
assign P[13][30] = x[13] & y[30];
assign P[13][31] = x[13] & y[31];
assign P[14][0] = x[14] & y[0];
assign P[14][1] = x[14] & y[1];
assign P[14][2] = x[14] & y[2];
assign P[14][3] = x[14] & y[3];
assign P[14][4] = x[14] & y[4];
assign P[14][5] = x[14] & y[5];
assign P[14][6] = x[14] & y[6];
assign P[14][7] = x[14] & y[7];
assign P[14][8] = x[14] & y[8];
assign P[14][9] = x[14] & y[9];
assign P[14][10] = x[14] & y[10];
assign P[14][11] = x[14] & y[11];
assign P[14][12] = x[14] & y[12];
assign P[14][13] = x[14] & y[13];
assign P[14][14] = x[14] & y[14];
assign P[14][15] = x[14] & y[15];
assign P[14][16] = x[14] & y[16];
assign P[14][17] = x[14] & y[17];
assign P[14][18] = x[14] & y[18];
assign P[14][19] = x[14] & y[19];
assign P[14][20] = x[14] & y[20];
assign P[14][21] = x[14] & y[21];
assign P[14][22] = x[14] & y[22];
assign P[14][23] = x[14] & y[23];
assign P[14][24] = x[14] & y[24];
assign P[14][25] = x[14] & y[25];
assign P[14][26] = x[14] & y[26];
assign P[14][27] = x[14] & y[27];
assign P[14][28] = x[14] & y[28];
assign P[14][29] = x[14] & y[29];
assign P[14][30] = x[14] & y[30];
assign P[14][31] = x[14] & y[31];
assign P[15][0] = x[15] & y[0];
assign P[15][1] = x[15] & y[1];
assign P[15][2] = x[15] & y[2];
assign P[15][3] = x[15] & y[3];
assign P[15][4] = x[15] & y[4];
assign P[15][5] = x[15] & y[5];
assign P[15][6] = x[15] & y[6];
assign P[15][7] = x[15] & y[7];
assign P[15][8] = x[15] & y[8];
assign P[15][9] = x[15] & y[9];
assign P[15][10] = x[15] & y[10];
assign P[15][11] = x[15] & y[11];
assign P[15][12] = x[15] & y[12];
assign P[15][13] = x[15] & y[13];
assign P[15][14] = x[15] & y[14];
assign P[15][15] = x[15] & y[15];
assign P[15][16] = x[15] & y[16];
assign P[15][17] = x[15] & y[17];
assign P[15][18] = x[15] & y[18];
assign P[15][19] = x[15] & y[19];
assign P[15][20] = x[15] & y[20];
assign P[15][21] = x[15] & y[21];
assign P[15][22] = x[15] & y[22];
assign P[15][23] = x[15] & y[23];
assign P[15][24] = x[15] & y[24];
assign P[15][25] = x[15] & y[25];
assign P[15][26] = x[15] & y[26];
assign P[15][27] = x[15] & y[27];
assign P[15][28] = x[15] & y[28];
assign P[15][29] = x[15] & y[29];
assign P[15][30] = x[15] & y[30];
assign P[15][31] = x[15] & y[31];
assign P[16][0] = x[16] & y[0];
assign P[16][1] = x[16] & y[1];
assign P[16][2] = x[16] & y[2];
assign P[16][3] = x[16] & y[3];
assign P[16][4] = x[16] & y[4];
assign P[16][5] = x[16] & y[5];
assign P[16][6] = x[16] & y[6];
assign P[16][7] = x[16] & y[7];
assign P[16][8] = x[16] & y[8];
assign P[16][9] = x[16] & y[9];
assign P[16][10] = x[16] & y[10];
assign P[16][11] = x[16] & y[11];
assign P[16][12] = x[16] & y[12];
assign P[16][13] = x[16] & y[13];
assign P[16][14] = x[16] & y[14];
assign P[16][15] = x[16] & y[15];
assign P[16][16] = x[16] & y[16];
assign P[16][17] = x[16] & y[17];
assign P[16][18] = x[16] & y[18];
assign P[16][19] = x[16] & y[19];
assign P[16][20] = x[16] & y[20];
assign P[16][21] = x[16] & y[21];
assign P[16][22] = x[16] & y[22];
assign P[16][23] = x[16] & y[23];
assign P[16][24] = x[16] & y[24];
assign P[16][25] = x[16] & y[25];
assign P[16][26] = x[16] & y[26];
assign P[16][27] = x[16] & y[27];
assign P[16][28] = x[16] & y[28];
assign P[16][29] = x[16] & y[29];
assign P[16][30] = x[16] & y[30];
assign P[16][31] = x[16] & y[31];
assign P[17][0] = x[17] & y[0];
assign P[17][1] = x[17] & y[1];
assign P[17][2] = x[17] & y[2];
assign P[17][3] = x[17] & y[3];
assign P[17][4] = x[17] & y[4];
assign P[17][5] = x[17] & y[5];
assign P[17][6] = x[17] & y[6];
assign P[17][7] = x[17] & y[7];
assign P[17][8] = x[17] & y[8];
assign P[17][9] = x[17] & y[9];
assign P[17][10] = x[17] & y[10];
assign P[17][11] = x[17] & y[11];
assign P[17][12] = x[17] & y[12];
assign P[17][13] = x[17] & y[13];
assign P[17][14] = x[17] & y[14];
assign P[17][15] = x[17] & y[15];
assign P[17][16] = x[17] & y[16];
assign P[17][17] = x[17] & y[17];
assign P[17][18] = x[17] & y[18];
assign P[17][19] = x[17] & y[19];
assign P[17][20] = x[17] & y[20];
assign P[17][21] = x[17] & y[21];
assign P[17][22] = x[17] & y[22];
assign P[17][23] = x[17] & y[23];
assign P[17][24] = x[17] & y[24];
assign P[17][25] = x[17] & y[25];
assign P[17][26] = x[17] & y[26];
assign P[17][27] = x[17] & y[27];
assign P[17][28] = x[17] & y[28];
assign P[17][29] = x[17] & y[29];
assign P[17][30] = x[17] & y[30];
assign P[17][31] = x[17] & y[31];
assign P[18][0] = x[18] & y[0];
assign P[18][1] = x[18] & y[1];
assign P[18][2] = x[18] & y[2];
assign P[18][3] = x[18] & y[3];
assign P[18][4] = x[18] & y[4];
assign P[18][5] = x[18] & y[5];
assign P[18][6] = x[18] & y[6];
assign P[18][7] = x[18] & y[7];
assign P[18][8] = x[18] & y[8];
assign P[18][9] = x[18] & y[9];
assign P[18][10] = x[18] & y[10];
assign P[18][11] = x[18] & y[11];
assign P[18][12] = x[18] & y[12];
assign P[18][13] = x[18] & y[13];
assign P[18][14] = x[18] & y[14];
assign P[18][15] = x[18] & y[15];
assign P[18][16] = x[18] & y[16];
assign P[18][17] = x[18] & y[17];
assign P[18][18] = x[18] & y[18];
assign P[18][19] = x[18] & y[19];
assign P[18][20] = x[18] & y[20];
assign P[18][21] = x[18] & y[21];
assign P[18][22] = x[18] & y[22];
assign P[18][23] = x[18] & y[23];
assign P[18][24] = x[18] & y[24];
assign P[18][25] = x[18] & y[25];
assign P[18][26] = x[18] & y[26];
assign P[18][27] = x[18] & y[27];
assign P[18][28] = x[18] & y[28];
assign P[18][29] = x[18] & y[29];
assign P[18][30] = x[18] & y[30];
assign P[18][31] = x[18] & y[31];
assign P[19][0] = x[19] & y[0];
assign P[19][1] = x[19] & y[1];
assign P[19][2] = x[19] & y[2];
assign P[19][3] = x[19] & y[3];
assign P[19][4] = x[19] & y[4];
assign P[19][5] = x[19] & y[5];
assign P[19][6] = x[19] & y[6];
assign P[19][7] = x[19] & y[7];
assign P[19][8] = x[19] & y[8];
assign P[19][9] = x[19] & y[9];
assign P[19][10] = x[19] & y[10];
assign P[19][11] = x[19] & y[11];
assign P[19][12] = x[19] & y[12];
assign P[19][13] = x[19] & y[13];
assign P[19][14] = x[19] & y[14];
assign P[19][15] = x[19] & y[15];
assign P[19][16] = x[19] & y[16];
assign P[19][17] = x[19] & y[17];
assign P[19][18] = x[19] & y[18];
assign P[19][19] = x[19] & y[19];
assign P[19][20] = x[19] & y[20];
assign P[19][21] = x[19] & y[21];
assign P[19][22] = x[19] & y[22];
assign P[19][23] = x[19] & y[23];
assign P[19][24] = x[19] & y[24];
assign P[19][25] = x[19] & y[25];
assign P[19][26] = x[19] & y[26];
assign P[19][27] = x[19] & y[27];
assign P[19][28] = x[19] & y[28];
assign P[19][29] = x[19] & y[29];
assign P[19][30] = x[19] & y[30];
assign P[19][31] = x[19] & y[31];
assign P[20][0] = x[20] & y[0];
assign P[20][1] = x[20] & y[1];
assign P[20][2] = x[20] & y[2];
assign P[20][3] = x[20] & y[3];
assign P[20][4] = x[20] & y[4];
assign P[20][5] = x[20] & y[5];
assign P[20][6] = x[20] & y[6];
assign P[20][7] = x[20] & y[7];
assign P[20][8] = x[20] & y[8];
assign P[20][9] = x[20] & y[9];
assign P[20][10] = x[20] & y[10];
assign P[20][11] = x[20] & y[11];
assign P[20][12] = x[20] & y[12];
assign P[20][13] = x[20] & y[13];
assign P[20][14] = x[20] & y[14];
assign P[20][15] = x[20] & y[15];
assign P[20][16] = x[20] & y[16];
assign P[20][17] = x[20] & y[17];
assign P[20][18] = x[20] & y[18];
assign P[20][19] = x[20] & y[19];
assign P[20][20] = x[20] & y[20];
assign P[20][21] = x[20] & y[21];
assign P[20][22] = x[20] & y[22];
assign P[20][23] = x[20] & y[23];
assign P[20][24] = x[20] & y[24];
assign P[20][25] = x[20] & y[25];
assign P[20][26] = x[20] & y[26];
assign P[20][27] = x[20] & y[27];
assign P[20][28] = x[20] & y[28];
assign P[20][29] = x[20] & y[29];
assign P[20][30] = x[20] & y[30];
assign P[20][31] = x[20] & y[31];
assign P[21][0] = x[21] & y[0];
assign P[21][1] = x[21] & y[1];
assign P[21][2] = x[21] & y[2];
assign P[21][3] = x[21] & y[3];
assign P[21][4] = x[21] & y[4];
assign P[21][5] = x[21] & y[5];
assign P[21][6] = x[21] & y[6];
assign P[21][7] = x[21] & y[7];
assign P[21][8] = x[21] & y[8];
assign P[21][9] = x[21] & y[9];
assign P[21][10] = x[21] & y[10];
assign P[21][11] = x[21] & y[11];
assign P[21][12] = x[21] & y[12];
assign P[21][13] = x[21] & y[13];
assign P[21][14] = x[21] & y[14];
assign P[21][15] = x[21] & y[15];
assign P[21][16] = x[21] & y[16];
assign P[21][17] = x[21] & y[17];
assign P[21][18] = x[21] & y[18];
assign P[21][19] = x[21] & y[19];
assign P[21][20] = x[21] & y[20];
assign P[21][21] = x[21] & y[21];
assign P[21][22] = x[21] & y[22];
assign P[21][23] = x[21] & y[23];
assign P[21][24] = x[21] & y[24];
assign P[21][25] = x[21] & y[25];
assign P[21][26] = x[21] & y[26];
assign P[21][27] = x[21] & y[27];
assign P[21][28] = x[21] & y[28];
assign P[21][29] = x[21] & y[29];
assign P[21][30] = x[21] & y[30];
assign P[21][31] = x[21] & y[31];
assign P[22][0] = x[22] & y[0];
assign P[22][1] = x[22] & y[1];
assign P[22][2] = x[22] & y[2];
assign P[22][3] = x[22] & y[3];
assign P[22][4] = x[22] & y[4];
assign P[22][5] = x[22] & y[5];
assign P[22][6] = x[22] & y[6];
assign P[22][7] = x[22] & y[7];
assign P[22][8] = x[22] & y[8];
assign P[22][9] = x[22] & y[9];
assign P[22][10] = x[22] & y[10];
assign P[22][11] = x[22] & y[11];
assign P[22][12] = x[22] & y[12];
assign P[22][13] = x[22] & y[13];
assign P[22][14] = x[22] & y[14];
assign P[22][15] = x[22] & y[15];
assign P[22][16] = x[22] & y[16];
assign P[22][17] = x[22] & y[17];
assign P[22][18] = x[22] & y[18];
assign P[22][19] = x[22] & y[19];
assign P[22][20] = x[22] & y[20];
assign P[22][21] = x[22] & y[21];
assign P[22][22] = x[22] & y[22];
assign P[22][23] = x[22] & y[23];
assign P[22][24] = x[22] & y[24];
assign P[22][25] = x[22] & y[25];
assign P[22][26] = x[22] & y[26];
assign P[22][27] = x[22] & y[27];
assign P[22][28] = x[22] & y[28];
assign P[22][29] = x[22] & y[29];
assign P[22][30] = x[22] & y[30];
assign P[22][31] = x[22] & y[31];
assign P[23][0] = x[23] & y[0];
assign P[23][1] = x[23] & y[1];
assign P[23][2] = x[23] & y[2];
assign P[23][3] = x[23] & y[3];
assign P[23][4] = x[23] & y[4];
assign P[23][5] = x[23] & y[5];
assign P[23][6] = x[23] & y[6];
assign P[23][7] = x[23] & y[7];
assign P[23][8] = x[23] & y[8];
assign P[23][9] = x[23] & y[9];
assign P[23][10] = x[23] & y[10];
assign P[23][11] = x[23] & y[11];
assign P[23][12] = x[23] & y[12];
assign P[23][13] = x[23] & y[13];
assign P[23][14] = x[23] & y[14];
assign P[23][15] = x[23] & y[15];
assign P[23][16] = x[23] & y[16];
assign P[23][17] = x[23] & y[17];
assign P[23][18] = x[23] & y[18];
assign P[23][19] = x[23] & y[19];
assign P[23][20] = x[23] & y[20];
assign P[23][21] = x[23] & y[21];
assign P[23][22] = x[23] & y[22];
assign P[23][23] = x[23] & y[23];
assign P[23][24] = x[23] & y[24];
assign P[23][25] = x[23] & y[25];
assign P[23][26] = x[23] & y[26];
assign P[23][27] = x[23] & y[27];
assign P[23][28] = x[23] & y[28];
assign P[23][29] = x[23] & y[29];
assign P[23][30] = x[23] & y[30];
assign P[23][31] = x[23] & y[31];
assign P[24][0] = x[24] & y[0];
assign P[24][1] = x[24] & y[1];
assign P[24][2] = x[24] & y[2];
assign P[24][3] = x[24] & y[3];
assign P[24][4] = x[24] & y[4];
assign P[24][5] = x[24] & y[5];
assign P[24][6] = x[24] & y[6];
assign P[24][7] = x[24] & y[7];
assign P[24][8] = x[24] & y[8];
assign P[24][9] = x[24] & y[9];
assign P[24][10] = x[24] & y[10];
assign P[24][11] = x[24] & y[11];
assign P[24][12] = x[24] & y[12];
assign P[24][13] = x[24] & y[13];
assign P[24][14] = x[24] & y[14];
assign P[24][15] = x[24] & y[15];
assign P[24][16] = x[24] & y[16];
assign P[24][17] = x[24] & y[17];
assign P[24][18] = x[24] & y[18];
assign P[24][19] = x[24] & y[19];
assign P[24][20] = x[24] & y[20];
assign P[24][21] = x[24] & y[21];
assign P[24][22] = x[24] & y[22];
assign P[24][23] = x[24] & y[23];
assign P[24][24] = x[24] & y[24];
assign P[24][25] = x[24] & y[25];
assign P[24][26] = x[24] & y[26];
assign P[24][27] = x[24] & y[27];
assign P[24][28] = x[24] & y[28];
assign P[24][29] = x[24] & y[29];
assign P[24][30] = x[24] & y[30];
assign P[24][31] = x[24] & y[31];
assign P[25][0] = x[25] & y[0];
assign P[25][1] = x[25] & y[1];
assign P[25][2] = x[25] & y[2];
assign P[25][3] = x[25] & y[3];
assign P[25][4] = x[25] & y[4];
assign P[25][5] = x[25] & y[5];
assign P[25][6] = x[25] & y[6];
assign P[25][7] = x[25] & y[7];
assign P[25][8] = x[25] & y[8];
assign P[25][9] = x[25] & y[9];
assign P[25][10] = x[25] & y[10];
assign P[25][11] = x[25] & y[11];
assign P[25][12] = x[25] & y[12];
assign P[25][13] = x[25] & y[13];
assign P[25][14] = x[25] & y[14];
assign P[25][15] = x[25] & y[15];
assign P[25][16] = x[25] & y[16];
assign P[25][17] = x[25] & y[17];
assign P[25][18] = x[25] & y[18];
assign P[25][19] = x[25] & y[19];
assign P[25][20] = x[25] & y[20];
assign P[25][21] = x[25] & y[21];
assign P[25][22] = x[25] & y[22];
assign P[25][23] = x[25] & y[23];
assign P[25][24] = x[25] & y[24];
assign P[25][25] = x[25] & y[25];
assign P[25][26] = x[25] & y[26];
assign P[25][27] = x[25] & y[27];
assign P[25][28] = x[25] & y[28];
assign P[25][29] = x[25] & y[29];
assign P[25][30] = x[25] & y[30];
assign P[25][31] = x[25] & y[31];
assign P[26][0] = x[26] & y[0];
assign P[26][1] = x[26] & y[1];
assign P[26][2] = x[26] & y[2];
assign P[26][3] = x[26] & y[3];
assign P[26][4] = x[26] & y[4];
assign P[26][5] = x[26] & y[5];
assign P[26][6] = x[26] & y[6];
assign P[26][7] = x[26] & y[7];
assign P[26][8] = x[26] & y[8];
assign P[26][9] = x[26] & y[9];
assign P[26][10] = x[26] & y[10];
assign P[26][11] = x[26] & y[11];
assign P[26][12] = x[26] & y[12];
assign P[26][13] = x[26] & y[13];
assign P[26][14] = x[26] & y[14];
assign P[26][15] = x[26] & y[15];
assign P[26][16] = x[26] & y[16];
assign P[26][17] = x[26] & y[17];
assign P[26][18] = x[26] & y[18];
assign P[26][19] = x[26] & y[19];
assign P[26][20] = x[26] & y[20];
assign P[26][21] = x[26] & y[21];
assign P[26][22] = x[26] & y[22];
assign P[26][23] = x[26] & y[23];
assign P[26][24] = x[26] & y[24];
assign P[26][25] = x[26] & y[25];
assign P[26][26] = x[26] & y[26];
assign P[26][27] = x[26] & y[27];
assign P[26][28] = x[26] & y[28];
assign P[26][29] = x[26] & y[29];
assign P[26][30] = x[26] & y[30];
assign P[26][31] = x[26] & y[31];
assign P[27][0] = x[27] & y[0];
assign P[27][1] = x[27] & y[1];
assign P[27][2] = x[27] & y[2];
assign P[27][3] = x[27] & y[3];
assign P[27][4] = x[27] & y[4];
assign P[27][5] = x[27] & y[5];
assign P[27][6] = x[27] & y[6];
assign P[27][7] = x[27] & y[7];
assign P[27][8] = x[27] & y[8];
assign P[27][9] = x[27] & y[9];
assign P[27][10] = x[27] & y[10];
assign P[27][11] = x[27] & y[11];
assign P[27][12] = x[27] & y[12];
assign P[27][13] = x[27] & y[13];
assign P[27][14] = x[27] & y[14];
assign P[27][15] = x[27] & y[15];
assign P[27][16] = x[27] & y[16];
assign P[27][17] = x[27] & y[17];
assign P[27][18] = x[27] & y[18];
assign P[27][19] = x[27] & y[19];
assign P[27][20] = x[27] & y[20];
assign P[27][21] = x[27] & y[21];
assign P[27][22] = x[27] & y[22];
assign P[27][23] = x[27] & y[23];
assign P[27][24] = x[27] & y[24];
assign P[27][25] = x[27] & y[25];
assign P[27][26] = x[27] & y[26];
assign P[27][27] = x[27] & y[27];
assign P[27][28] = x[27] & y[28];
assign P[27][29] = x[27] & y[29];
assign P[27][30] = x[27] & y[30];
assign P[27][31] = x[27] & y[31];
assign P[28][0] = x[28] & y[0];
assign P[28][1] = x[28] & y[1];
assign P[28][2] = x[28] & y[2];
assign P[28][3] = x[28] & y[3];
assign P[28][4] = x[28] & y[4];
assign P[28][5] = x[28] & y[5];
assign P[28][6] = x[28] & y[6];
assign P[28][7] = x[28] & y[7];
assign P[28][8] = x[28] & y[8];
assign P[28][9] = x[28] & y[9];
assign P[28][10] = x[28] & y[10];
assign P[28][11] = x[28] & y[11];
assign P[28][12] = x[28] & y[12];
assign P[28][13] = x[28] & y[13];
assign P[28][14] = x[28] & y[14];
assign P[28][15] = x[28] & y[15];
assign P[28][16] = x[28] & y[16];
assign P[28][17] = x[28] & y[17];
assign P[28][18] = x[28] & y[18];
assign P[28][19] = x[28] & y[19];
assign P[28][20] = x[28] & y[20];
assign P[28][21] = x[28] & y[21];
assign P[28][22] = x[28] & y[22];
assign P[28][23] = x[28] & y[23];
assign P[28][24] = x[28] & y[24];
assign P[28][25] = x[28] & y[25];
assign P[28][26] = x[28] & y[26];
assign P[28][27] = x[28] & y[27];
assign P[28][28] = x[28] & y[28];
assign P[28][29] = x[28] & y[29];
assign P[28][30] = x[28] & y[30];
assign P[28][31] = x[28] & y[31];
assign P[29][0] = x[29] & y[0];
assign P[29][1] = x[29] & y[1];
assign P[29][2] = x[29] & y[2];
assign P[29][3] = x[29] & y[3];
assign P[29][4] = x[29] & y[4];
assign P[29][5] = x[29] & y[5];
assign P[29][6] = x[29] & y[6];
assign P[29][7] = x[29] & y[7];
assign P[29][8] = x[29] & y[8];
assign P[29][9] = x[29] & y[9];
assign P[29][10] = x[29] & y[10];
assign P[29][11] = x[29] & y[11];
assign P[29][12] = x[29] & y[12];
assign P[29][13] = x[29] & y[13];
assign P[29][14] = x[29] & y[14];
assign P[29][15] = x[29] & y[15];
assign P[29][16] = x[29] & y[16];
assign P[29][17] = x[29] & y[17];
assign P[29][18] = x[29] & y[18];
assign P[29][19] = x[29] & y[19];
assign P[29][20] = x[29] & y[20];
assign P[29][21] = x[29] & y[21];
assign P[29][22] = x[29] & y[22];
assign P[29][23] = x[29] & y[23];
assign P[29][24] = x[29] & y[24];
assign P[29][25] = x[29] & y[25];
assign P[29][26] = x[29] & y[26];
assign P[29][27] = x[29] & y[27];
assign P[29][28] = x[29] & y[28];
assign P[29][29] = x[29] & y[29];
assign P[29][30] = x[29] & y[30];
assign P[29][31] = x[29] & y[31];
assign P[30][0] = x[30] & y[0];
assign P[30][1] = x[30] & y[1];
assign P[30][2] = x[30] & y[2];
assign P[30][3] = x[30] & y[3];
assign P[30][4] = x[30] & y[4];
assign P[30][5] = x[30] & y[5];
assign P[30][6] = x[30] & y[6];
assign P[30][7] = x[30] & y[7];
assign P[30][8] = x[30] & y[8];
assign P[30][9] = x[30] & y[9];
assign P[30][10] = x[30] & y[10];
assign P[30][11] = x[30] & y[11];
assign P[30][12] = x[30] & y[12];
assign P[30][13] = x[30] & y[13];
assign P[30][14] = x[30] & y[14];
assign P[30][15] = x[30] & y[15];
assign P[30][16] = x[30] & y[16];
assign P[30][17] = x[30] & y[17];
assign P[30][18] = x[30] & y[18];
assign P[30][19] = x[30] & y[19];
assign P[30][20] = x[30] & y[20];
assign P[30][21] = x[30] & y[21];
assign P[30][22] = x[30] & y[22];
assign P[30][23] = x[30] & y[23];
assign P[30][24] = x[30] & y[24];
assign P[30][25] = x[30] & y[25];
assign P[30][26] = x[30] & y[26];
assign P[30][27] = x[30] & y[27];
assign P[30][28] = x[30] & y[28];
assign P[30][29] = x[30] & y[29];
assign P[30][30] = x[30] & y[30];
assign P[30][31] = x[30] & y[31];
assign P[31][0] = x[31] & y[0];
assign P[31][1] = x[31] & y[1];
assign P[31][2] = x[31] & y[2];
assign P[31][3] = x[31] & y[3];
assign P[31][4] = x[31] & y[4];
assign P[31][5] = x[31] & y[5];
assign P[31][6] = x[31] & y[6];
assign P[31][7] = x[31] & y[7];
assign P[31][8] = x[31] & y[8];
assign P[31][9] = x[31] & y[9];
assign P[31][10] = x[31] & y[10];
assign P[31][11] = x[31] & y[11];
assign P[31][12] = x[31] & y[12];
assign P[31][13] = x[31] & y[13];
assign P[31][14] = x[31] & y[14];
assign P[31][15] = x[31] & y[15];
assign P[31][16] = x[31] & y[16];
assign P[31][17] = x[31] & y[17];
assign P[31][18] = x[31] & y[18];
assign P[31][19] = x[31] & y[19];
assign P[31][20] = x[31] & y[20];
assign P[31][21] = x[31] & y[21];
assign P[31][22] = x[31] & y[22];
assign P[31][23] = x[31] & y[23];
assign P[31][24] = x[31] & y[24];
assign P[31][25] = x[31] & y[25];
assign P[31][26] = x[31] & y[26];
assign P[31][27] = x[31] & y[27];
assign P[31][28] = x[31] & y[28];
assign P[31][29] = x[31] & y[29];
assign P[31][30] = x[31] & y[30];
assign P[31][31] = x[31] & y[31];

wire [1116:0] S;
wire [1116:0] Cout;

Half_Adder HA1 (P[0][1], P[1][0], S[0], Cout[0]);
Full_Adder FA2 (P[0][2], P[1][1], P[2][0], S[1], Cout[1]);
Full_Adder FA3 (P[0][3], P[1][2], P[2][1], S[2], Cout[2]);
Full_Adder FA4 (P[0][4], P[1][3], P[2][2], S[3], Cout[3]);
Half_Adder HA5 (P[3][1], P[4][0], S[4], Cout[4]);
Full_Adder FA6 (P[0][5], P[1][4], P[2][3], S[5], Cout[5]);
Full_Adder FA7 (P[3][2], P[4][1], P[5][0], S[6], Cout[6]);
Full_Adder FA8 (P[0][6], P[1][5], P[2][4], S[7], Cout[7]);
Full_Adder FA9 (P[3][3], P[4][2], P[5][1], S[8], Cout[8]);
Full_Adder FA10 (P[0][7], P[1][6], P[2][5], S[9], Cout[9]);
Full_Adder FA11 (P[3][4], P[4][3], P[5][2], S[10], Cout[10]);
Half_Adder HA12 (P[6][1], P[7][0], S[11], Cout[11]);
Full_Adder FA13 (P[0][8], P[1][7], P[2][6], S[12], Cout[12]);
Full_Adder FA14 (P[3][5], P[4][4], P[5][3], S[13], Cout[13]);
Full_Adder FA15 (P[6][2], P[7][1], P[8][0], S[14], Cout[14]);
Full_Adder FA16 (P[0][9], P[1][8], P[2][7], S[15], Cout[15]);
Full_Adder FA17 (P[3][6], P[4][5], P[5][4], S[16], Cout[16]);
Full_Adder FA18 (P[6][3], P[7][2], P[8][1], S[17], Cout[17]);
Full_Adder FA19 (P[0][10], P[1][9], P[2][8], S[18], Cout[18]);
Full_Adder FA20 (P[3][7], P[4][6], P[5][5], S[19], Cout[19]);
Full_Adder FA21 (P[6][4], P[7][3], P[8][2], S[20], Cout[20]);
Half_Adder HA22 (P[9][1], P[10][0], S[21], Cout[21]);
Full_Adder FA23 (P[0][11], P[1][10], P[2][9], S[22], Cout[22]);
Full_Adder FA24 (P[3][8], P[4][7], P[5][6], S[23], Cout[23]);
Full_Adder FA25 (P[6][5], P[7][4], P[8][3], S[24], Cout[24]);
Full_Adder FA26 (P[9][2], P[10][1], P[11][0], S[25], Cout[25]);
Full_Adder FA27 (P[0][12], P[1][11], P[2][10], S[26], Cout[26]);
Full_Adder FA28 (P[3][9], P[4][8], P[5][7], S[27], Cout[27]);
Full_Adder FA29 (P[6][6], P[7][5], P[8][4], S[28], Cout[28]);
Full_Adder FA30 (P[9][3], P[10][2], P[11][1], S[29], Cout[29]);
Full_Adder FA31 (P[0][13], P[1][12], P[2][11], S[30], Cout[30]);
Full_Adder FA32 (P[3][10], P[4][9], P[5][8], S[31], Cout[31]);
Full_Adder FA33 (P[6][7], P[7][6], P[8][5], S[32], Cout[32]);
Full_Adder FA34 (P[9][4], P[10][3], P[11][2], S[33], Cout[33]);
Half_Adder HA35 (P[12][1], P[13][0], S[34], Cout[34]);
Full_Adder FA36 (P[0][14], P[1][13], P[2][12], S[35], Cout[35]);
Full_Adder FA37 (P[3][11], P[4][10], P[5][9], S[36], Cout[36]);
Full_Adder FA38 (P[6][8], P[7][7], P[8][6], S[37], Cout[37]);
Full_Adder FA39 (P[9][5], P[10][4], P[11][3], S[38], Cout[38]);
Full_Adder FA40 (P[12][2], P[13][1], P[14][0], S[39], Cout[39]);
Full_Adder FA41 (P[0][15], P[1][14], P[2][13], S[40], Cout[40]);
Full_Adder FA42 (P[3][12], P[4][11], P[5][10], S[41], Cout[41]);
Full_Adder FA43 (P[6][9], P[7][8], P[8][7], S[42], Cout[42]);
Full_Adder FA44 (P[9][6], P[10][5], P[11][4], S[43], Cout[43]);
Full_Adder FA45 (P[12][3], P[13][2], P[14][1], S[44], Cout[44]);
Full_Adder FA46 (P[0][16], P[1][15], P[2][14], S[45], Cout[45]);
Full_Adder FA47 (P[3][13], P[4][12], P[5][11], S[46], Cout[46]);
Full_Adder FA48 (P[6][10], P[7][9], P[8][8], S[47], Cout[47]);
Full_Adder FA49 (P[9][7], P[10][6], P[11][5], S[48], Cout[48]);
Full_Adder FA50 (P[12][4], P[13][3], P[14][2], S[49], Cout[49]);
Half_Adder HA51 (P[15][1], P[16][0], S[50], Cout[50]);
Full_Adder FA52 (P[0][17], P[1][16], P[2][15], S[51], Cout[51]);
Full_Adder FA53 (P[3][14], P[4][13], P[5][12], S[52], Cout[52]);
Full_Adder FA54 (P[6][11], P[7][10], P[8][9], S[53], Cout[53]);
Full_Adder FA55 (P[9][8], P[10][7], P[11][6], S[54], Cout[54]);
Full_Adder FA56 (P[12][5], P[13][4], P[14][3], S[55], Cout[55]);
Full_Adder FA57 (P[15][2], P[16][1], P[17][0], S[56], Cout[56]);
Full_Adder FA58 (P[0][18], P[1][17], P[2][16], S[57], Cout[57]);
Full_Adder FA59 (P[3][15], P[4][14], P[5][13], S[58], Cout[58]);
Full_Adder FA60 (P[6][12], P[7][11], P[8][10], S[59], Cout[59]);
Full_Adder FA61 (P[9][9], P[10][8], P[11][7], S[60], Cout[60]);
Full_Adder FA62 (P[12][6], P[13][5], P[14][4], S[61], Cout[61]);
Full_Adder FA63 (P[15][3], P[16][2], P[17][1], S[62], Cout[62]);
Full_Adder FA64 (P[0][19], P[1][18], P[2][17], S[63], Cout[63]);
Full_Adder FA65 (P[3][16], P[4][15], P[5][14], S[64], Cout[64]);
Full_Adder FA66 (P[6][13], P[7][12], P[8][11], S[65], Cout[65]);
Full_Adder FA67 (P[9][10], P[10][9], P[11][8], S[66], Cout[66]);
Full_Adder FA68 (P[12][7], P[13][6], P[14][5], S[67], Cout[67]);
Full_Adder FA69 (P[15][4], P[16][3], P[17][2], S[68], Cout[68]);
Half_Adder HA70 (P[18][1], P[19][0], S[69], Cout[69]);
Full_Adder FA71 (P[0][20], P[1][19], P[2][18], S[70], Cout[70]);
Full_Adder FA72 (P[3][17], P[4][16], P[5][15], S[71], Cout[71]);
Full_Adder FA73 (P[6][14], P[7][13], P[8][12], S[72], Cout[72]);
Full_Adder FA74 (P[9][11], P[10][10], P[11][9], S[73], Cout[73]);
Full_Adder FA75 (P[12][8], P[13][7], P[14][6], S[74], Cout[74]);
Full_Adder FA76 (P[15][5], P[16][4], P[17][3], S[75], Cout[75]);
Full_Adder FA77 (P[18][2], P[19][1], P[20][0], S[76], Cout[76]);
Full_Adder FA78 (P[0][21], P[1][20], P[2][19], S[77], Cout[77]);
Full_Adder FA79 (P[3][18], P[4][17], P[5][16], S[78], Cout[78]);
Full_Adder FA80 (P[6][15], P[7][14], P[8][13], S[79], Cout[79]);
Full_Adder FA81 (P[9][12], P[10][11], P[11][10], S[80], Cout[80]);
Full_Adder FA82 (P[12][9], P[13][8], P[14][7], S[81], Cout[81]);
Full_Adder FA83 (P[15][6], P[16][5], P[17][4], S[82], Cout[82]);
Full_Adder FA84 (P[18][3], P[19][2], P[20][1], S[83], Cout[83]);
Full_Adder FA85 (P[0][22], P[1][21], P[2][20], S[84], Cout[84]);
Full_Adder FA86 (P[3][19], P[4][18], P[5][17], S[85], Cout[85]);
Full_Adder FA87 (P[6][16], P[7][15], P[8][14], S[86], Cout[86]);
Full_Adder FA88 (P[9][13], P[10][12], P[11][11], S[87], Cout[87]);
Full_Adder FA89 (P[12][10], P[13][9], P[14][8], S[88], Cout[88]);
Full_Adder FA90 (P[15][7], P[16][6], P[17][5], S[89], Cout[89]);
Full_Adder FA91 (P[18][4], P[19][3], P[20][2], S[90], Cout[90]);
Half_Adder HA92 (P[21][1], P[22][0], S[91], Cout[91]);
Full_Adder FA93 (P[0][23], P[1][22], P[2][21], S[92], Cout[92]);
Full_Adder FA94 (P[3][20], P[4][19], P[5][18], S[93], Cout[93]);
Full_Adder FA95 (P[6][17], P[7][16], P[8][15], S[94], Cout[94]);
Full_Adder FA96 (P[9][14], P[10][13], P[11][12], S[95], Cout[95]);
Full_Adder FA97 (P[12][11], P[13][10], P[14][9], S[96], Cout[96]);
Full_Adder FA98 (P[15][8], P[16][7], P[17][6], S[97], Cout[97]);
Full_Adder FA99 (P[18][5], P[19][4], P[20][3], S[98], Cout[98]);
Full_Adder FA100 (P[21][2], P[22][1], P[23][0], S[99], Cout[99]);
Full_Adder FA101 (P[0][24], P[1][23], P[2][22], S[100], Cout[100]);
Full_Adder FA102 (P[3][21], P[4][20], P[5][19], S[101], Cout[101]);
Full_Adder FA103 (P[6][18], P[7][17], P[8][16], S[102], Cout[102]);
Full_Adder FA104 (P[9][15], P[10][14], P[11][13], S[103], Cout[103]);
Full_Adder FA105 (P[12][12], P[13][11], P[14][10], S[104], Cout[104]);
Full_Adder FA106 (P[15][9], P[16][8], P[17][7], S[105], Cout[105]);
Full_Adder FA107 (P[18][6], P[19][5], P[20][4], S[106], Cout[106]);
Full_Adder FA108 (P[21][3], P[22][2], P[23][1], S[107], Cout[107]);
Full_Adder FA109 (P[0][25], P[1][24], P[2][23], S[108], Cout[108]);
Full_Adder FA110 (P[3][22], P[4][21], P[5][20], S[109], Cout[109]);
Full_Adder FA111 (P[6][19], P[7][18], P[8][17], S[110], Cout[110]);
Full_Adder FA112 (P[9][16], P[10][15], P[11][14], S[111], Cout[111]);
Full_Adder FA113 (P[12][13], P[13][12], P[14][11], S[112], Cout[112]);
Full_Adder FA114 (P[15][10], P[16][9], P[17][8], S[113], Cout[113]);
Full_Adder FA115 (P[18][7], P[19][6], P[20][5], S[114], Cout[114]);
Full_Adder FA116 (P[21][4], P[22][3], P[23][2], S[115], Cout[115]);
Half_Adder HA117 (P[24][1], P[25][0], S[116], Cout[116]);
Full_Adder FA118 (P[0][26], P[1][25], P[2][24], S[117], Cout[117]);
Full_Adder FA119 (P[3][23], P[4][22], P[5][21], S[118], Cout[118]);
Full_Adder FA120 (P[6][20], P[7][19], P[8][18], S[119], Cout[119]);
Full_Adder FA121 (P[9][17], P[10][16], P[11][15], S[120], Cout[120]);
Full_Adder FA122 (P[12][14], P[13][13], P[14][12], S[121], Cout[121]);
Full_Adder FA123 (P[15][11], P[16][10], P[17][9], S[122], Cout[122]);
Full_Adder FA124 (P[18][8], P[19][7], P[20][6], S[123], Cout[123]);
Full_Adder FA125 (P[21][5], P[22][4], P[23][3], S[124], Cout[124]);
Full_Adder FA126 (P[24][2], P[25][1], P[26][0], S[125], Cout[125]);
Full_Adder FA127 (P[0][27], P[1][26], P[2][25], S[126], Cout[126]);
Full_Adder FA128 (P[3][24], P[4][23], P[5][22], S[127], Cout[127]);
Full_Adder FA129 (P[6][21], P[7][20], P[8][19], S[128], Cout[128]);
Full_Adder FA130 (P[9][18], P[10][17], P[11][16], S[129], Cout[129]);
Full_Adder FA131 (P[12][15], P[13][14], P[14][13], S[130], Cout[130]);
Full_Adder FA132 (P[15][12], P[16][11], P[17][10], S[131], Cout[131]);
Full_Adder FA133 (P[18][9], P[19][8], P[20][7], S[132], Cout[132]);
Full_Adder FA134 (P[21][6], P[22][5], P[23][4], S[133], Cout[133]);
Full_Adder FA135 (P[24][3], P[25][2], P[26][1], S[134], Cout[134]);
Full_Adder FA136 (P[0][28], P[1][27], P[2][26], S[135], Cout[135]);
Full_Adder FA137 (P[3][25], P[4][24], P[5][23], S[136], Cout[136]);
Full_Adder FA138 (P[6][22], P[7][21], P[8][20], S[137], Cout[137]);
Full_Adder FA139 (P[9][19], P[10][18], P[11][17], S[138], Cout[138]);
Full_Adder FA140 (P[12][16], P[13][15], P[14][14], S[139], Cout[139]);
Full_Adder FA141 (P[15][13], P[16][12], P[17][11], S[140], Cout[140]);
Full_Adder FA142 (P[18][10], P[19][9], P[20][8], S[141], Cout[141]);
Full_Adder FA143 (P[21][7], P[22][6], P[23][5], S[142], Cout[142]);
Full_Adder FA144 (P[24][4], P[25][3], P[26][2], S[143], Cout[143]);
Half_Adder HA145 (P[27][1], P[28][0], S[144], Cout[144]);
Full_Adder FA146 (P[0][29], P[1][28], P[2][27], S[145], Cout[145]);
Full_Adder FA147 (P[3][26], P[4][25], P[5][24], S[146], Cout[146]);
Full_Adder FA148 (P[6][23], P[7][22], P[8][21], S[147], Cout[147]);
Full_Adder FA149 (P[9][20], P[10][19], P[11][18], S[148], Cout[148]);
Full_Adder FA150 (P[12][17], P[13][16], P[14][15], S[149], Cout[149]);
Full_Adder FA151 (P[15][14], P[16][13], P[17][12], S[150], Cout[150]);
Full_Adder FA152 (P[18][11], P[19][10], P[20][9], S[151], Cout[151]);
Full_Adder FA153 (P[21][8], P[22][7], P[23][6], S[152], Cout[152]);
Full_Adder FA154 (P[24][5], P[25][4], P[26][3], S[153], Cout[153]);
Full_Adder FA155 (P[27][2], P[28][1], P[29][0], S[154], Cout[154]);
Full_Adder FA156 (P[0][30], P[1][29], P[2][28], S[155], Cout[155]);
Full_Adder FA157 (P[3][27], P[4][26], P[5][25], S[156], Cout[156]);
Full_Adder FA158 (P[6][24], P[7][23], P[8][22], S[157], Cout[157]);
Full_Adder FA159 (P[9][21], P[10][20], P[11][19], S[158], Cout[158]);
Full_Adder FA160 (P[12][18], P[13][17], P[14][16], S[159], Cout[159]);
Full_Adder FA161 (P[15][15], P[16][14], P[17][13], S[160], Cout[160]);
Full_Adder FA162 (P[18][12], P[19][11], P[20][10], S[161], Cout[161]);
Full_Adder FA163 (P[21][9], P[22][8], P[23][7], S[162], Cout[162]);
Full_Adder FA164 (P[24][6], P[25][5], P[26][4], S[163], Cout[163]);
Full_Adder FA165 (P[27][3], P[28][2], P[29][1], S[164], Cout[164]);
Full_Adder FA166 (P[0][31], P[1][30], P[2][29], S[165], Cout[165]);
Full_Adder FA167 (P[3][28], P[4][27], P[5][26], S[166], Cout[166]);
Full_Adder FA168 (P[6][25], P[7][24], P[8][23], S[167], Cout[167]);
Full_Adder FA169 (P[9][22], P[10][21], P[11][20], S[168], Cout[168]);
Full_Adder FA170 (P[12][19], P[13][18], P[14][17], S[169], Cout[169]);
Full_Adder FA171 (P[15][16], P[16][15], P[17][14], S[170], Cout[170]);
Full_Adder FA172 (P[18][13], P[19][12], P[20][11], S[171], Cout[171]);
Full_Adder FA173 (P[21][10], P[22][9], P[23][8], S[172], Cout[172]);
Full_Adder FA174 (P[24][7], P[25][6], P[26][5], S[173], Cout[173]);
Full_Adder FA175 (P[27][4], P[28][3], P[29][2], S[174], Cout[174]);
Full_Adder FA176 (P[1][31], P[2][30], P[3][29], S[175], Cout[175]);
Full_Adder FA177 (P[4][28], P[5][27], P[6][26], S[176], Cout[176]);
Full_Adder FA178 (P[7][25], P[8][24], P[9][23], S[177], Cout[177]);
Full_Adder FA179 (P[10][22], P[11][21], P[12][20], S[178], Cout[178]);
Full_Adder FA180 (P[13][19], P[14][18], P[15][17], S[179], Cout[179]);
Full_Adder FA181 (P[16][16], P[17][15], P[18][14], S[180], Cout[180]);
Full_Adder FA182 (P[19][13], P[20][12], P[21][11], S[181], Cout[181]);
Full_Adder FA183 (P[22][10], P[23][9], P[24][8], S[182], Cout[182]);
Full_Adder FA184 (P[25][7], P[26][6], P[27][5], S[183], Cout[183]);
Half_Adder HA185 (P[28][4], P[29][3], S[184], Cout[184]);
Full_Adder FA186 (P[2][31], P[3][30], P[4][29], S[185], Cout[185]);
Full_Adder FA187 (P[5][28], P[6][27], P[7][26], S[186], Cout[186]);
Full_Adder FA188 (P[8][25], P[9][24], P[10][23], S[187], Cout[187]);
Full_Adder FA189 (P[11][22], P[12][21], P[13][20], S[188], Cout[188]);
Full_Adder FA190 (P[14][19], P[15][18], P[16][17], S[189], Cout[189]);
Full_Adder FA191 (P[17][16], P[18][15], P[19][14], S[190], Cout[190]);
Full_Adder FA192 (P[20][13], P[21][12], P[22][11], S[191], Cout[191]);
Full_Adder FA193 (P[23][10], P[24][9], P[25][8], S[192], Cout[192]);
Full_Adder FA194 (P[26][7], P[27][6], P[28][5], S[193], Cout[193]);
Full_Adder FA195 (P[3][31], P[4][30], P[5][29], S[194], Cout[194]);
Full_Adder FA196 (P[6][28], P[7][27], P[8][26], S[195], Cout[195]);
Full_Adder FA197 (P[9][25], P[10][24], P[11][23], S[196], Cout[196]);
Full_Adder FA198 (P[12][22], P[13][21], P[14][20], S[197], Cout[197]);
Full_Adder FA199 (P[15][19], P[16][18], P[17][17], S[198], Cout[198]);
Full_Adder FA200 (P[18][16], P[19][15], P[20][14], S[199], Cout[199]);
Full_Adder FA201 (P[21][13], P[22][12], P[23][11], S[200], Cout[200]);
Full_Adder FA202 (P[24][10], P[25][9], P[26][8], S[201], Cout[201]);
Full_Adder FA203 (P[27][7], P[28][6], P[29][5], S[202], Cout[202]);
Full_Adder FA204 (P[4][31], P[5][30], P[6][29], S[203], Cout[203]);
Full_Adder FA205 (P[7][28], P[8][27], P[9][26], S[204], Cout[204]);
Full_Adder FA206 (P[10][25], P[11][24], P[12][23], S[205], Cout[205]);
Full_Adder FA207 (P[13][22], P[14][21], P[15][20], S[206], Cout[206]);
Full_Adder FA208 (P[16][19], P[17][18], P[18][17], S[207], Cout[207]);
Full_Adder FA209 (P[19][16], P[20][15], P[21][14], S[208], Cout[208]);
Full_Adder FA210 (P[22][13], P[23][12], P[24][11], S[209], Cout[209]);
Full_Adder FA211 (P[25][10], P[26][9], P[27][8], S[210], Cout[210]);
Half_Adder HA212 (P[28][7], P[29][6], S[211], Cout[211]);
Full_Adder FA213 (P[5][31], P[6][30], P[7][29], S[212], Cout[212]);
Full_Adder FA214 (P[8][28], P[9][27], P[10][26], S[213], Cout[213]);
Full_Adder FA215 (P[11][25], P[12][24], P[13][23], S[214], Cout[214]);
Full_Adder FA216 (P[14][22], P[15][21], P[16][20], S[215], Cout[215]);
Full_Adder FA217 (P[17][19], P[18][18], P[19][17], S[216], Cout[216]);
Full_Adder FA218 (P[20][16], P[21][15], P[22][14], S[217], Cout[217]);
Full_Adder FA219 (P[23][13], P[24][12], P[25][11], S[218], Cout[218]);
Full_Adder FA220 (P[26][10], P[27][9], P[28][8], S[219], Cout[219]);
Full_Adder FA221 (P[6][31], P[7][30], P[8][29], S[220], Cout[220]);
Full_Adder FA222 (P[9][28], P[10][27], P[11][26], S[221], Cout[221]);
Full_Adder FA223 (P[12][25], P[13][24], P[14][23], S[222], Cout[222]);
Full_Adder FA224 (P[15][22], P[16][21], P[17][20], S[223], Cout[223]);
Full_Adder FA225 (P[18][19], P[19][18], P[20][17], S[224], Cout[224]);
Full_Adder FA226 (P[21][16], P[22][15], P[23][14], S[225], Cout[225]);
Full_Adder FA227 (P[24][13], P[25][12], P[26][11], S[226], Cout[226]);
Full_Adder FA228 (P[27][10], P[28][9], P[29][8], S[227], Cout[227]);
Full_Adder FA229 (P[7][31], P[8][30], P[9][29], S[228], Cout[228]);
Full_Adder FA230 (P[10][28], P[11][27], P[12][26], S[229], Cout[229]);
Full_Adder FA231 (P[13][25], P[14][24], P[15][23], S[230], Cout[230]);
Full_Adder FA232 (P[16][22], P[17][21], P[18][20], S[231], Cout[231]);
Full_Adder FA233 (P[19][19], P[20][18], P[21][17], S[232], Cout[232]);
Full_Adder FA234 (P[22][16], P[23][15], P[24][14], S[233], Cout[233]);
Full_Adder FA235 (P[25][13], P[26][12], P[27][11], S[234], Cout[234]);
Half_Adder HA236 (P[28][10], P[29][9], S[235], Cout[235]);
Full_Adder FA237 (P[8][31], P[9][30], P[10][29], S[236], Cout[236]);
Full_Adder FA238 (P[11][28], P[12][27], P[13][26], S[237], Cout[237]);
Full_Adder FA239 (P[14][25], P[15][24], P[16][23], S[238], Cout[238]);
Full_Adder FA240 (P[17][22], P[18][21], P[19][20], S[239], Cout[239]);
Full_Adder FA241 (P[20][19], P[21][18], P[22][17], S[240], Cout[240]);
Full_Adder FA242 (P[23][16], P[24][15], P[25][14], S[241], Cout[241]);
Full_Adder FA243 (P[26][13], P[27][12], P[28][11], S[242], Cout[242]);
Full_Adder FA244 (P[9][31], P[10][30], P[11][29], S[243], Cout[243]);
Full_Adder FA245 (P[12][28], P[13][27], P[14][26], S[244], Cout[244]);
Full_Adder FA246 (P[15][25], P[16][24], P[17][23], S[245], Cout[245]);
Full_Adder FA247 (P[18][22], P[19][21], P[20][20], S[246], Cout[246]);
Full_Adder FA248 (P[21][19], P[22][18], P[23][17], S[247], Cout[247]);
Full_Adder FA249 (P[24][16], P[25][15], P[26][14], S[248], Cout[248]);
Full_Adder FA250 (P[27][13], P[28][12], P[29][11], S[249], Cout[249]);
Full_Adder FA251 (P[10][31], P[11][30], P[12][29], S[250], Cout[250]);
Full_Adder FA252 (P[13][28], P[14][27], P[15][26], S[251], Cout[251]);
Full_Adder FA253 (P[16][25], P[17][24], P[18][23], S[252], Cout[252]);
Full_Adder FA254 (P[19][22], P[20][21], P[21][20], S[253], Cout[253]);
Full_Adder FA255 (P[22][19], P[23][18], P[24][17], S[254], Cout[254]);
Full_Adder FA256 (P[25][16], P[26][15], P[27][14], S[255], Cout[255]);
Half_Adder HA257 (P[28][13], P[29][12], S[256], Cout[256]);
Full_Adder FA258 (P[11][31], P[12][30], P[13][29], S[257], Cout[257]);
Full_Adder FA259 (P[14][28], P[15][27], P[16][26], S[258], Cout[258]);
Full_Adder FA260 (P[17][25], P[18][24], P[19][23], S[259], Cout[259]);
Full_Adder FA261 (P[20][22], P[21][21], P[22][20], S[260], Cout[260]);
Full_Adder FA262 (P[23][19], P[24][18], P[25][17], S[261], Cout[261]);
Full_Adder FA263 (P[26][16], P[27][15], P[28][14], S[262], Cout[262]);
Full_Adder FA264 (P[12][31], P[13][30], P[14][29], S[263], Cout[263]);
Full_Adder FA265 (P[15][28], P[16][27], P[17][26], S[264], Cout[264]);
Full_Adder FA266 (P[18][25], P[19][24], P[20][23], S[265], Cout[265]);
Full_Adder FA267 (P[21][22], P[22][21], P[23][20], S[266], Cout[266]);
Full_Adder FA268 (P[24][19], P[25][18], P[26][17], S[267], Cout[267]);
Full_Adder FA269 (P[27][16], P[28][15], P[29][14], S[268], Cout[268]);
Full_Adder FA270 (P[13][31], P[14][30], P[15][29], S[269], Cout[269]);
Full_Adder FA271 (P[16][28], P[17][27], P[18][26], S[270], Cout[270]);
Full_Adder FA272 (P[19][25], P[20][24], P[21][23], S[271], Cout[271]);
Full_Adder FA273 (P[22][22], P[23][21], P[24][20], S[272], Cout[272]);
Full_Adder FA274 (P[25][19], P[26][18], P[27][17], S[273], Cout[273]);
Half_Adder HA275 (P[28][16], P[29][15], S[274], Cout[274]);
Full_Adder FA276 (P[14][31], P[15][30], P[16][29], S[275], Cout[275]);
Full_Adder FA277 (P[17][28], P[18][27], P[19][26], S[276], Cout[276]);
Full_Adder FA278 (P[20][25], P[21][24], P[22][23], S[277], Cout[277]);
Full_Adder FA279 (P[23][22], P[24][21], P[25][20], S[278], Cout[278]);
Full_Adder FA280 (P[26][19], P[27][18], P[28][17], S[279], Cout[279]);
Full_Adder FA281 (P[15][31], P[16][30], P[17][29], S[280], Cout[280]);
Full_Adder FA282 (P[18][28], P[19][27], P[20][26], S[281], Cout[281]);
Full_Adder FA283 (P[21][25], P[22][24], P[23][23], S[282], Cout[282]);
Full_Adder FA284 (P[24][22], P[25][21], P[26][20], S[283], Cout[283]);
Full_Adder FA285 (P[27][19], P[28][18], P[29][17], S[284], Cout[284]);
Full_Adder FA286 (P[16][31], P[17][30], P[18][29], S[285], Cout[285]);
Full_Adder FA287 (P[19][28], P[20][27], P[21][26], S[286], Cout[286]);
Full_Adder FA288 (P[22][25], P[23][24], P[24][23], S[287], Cout[287]);
Full_Adder FA289 (P[25][22], P[26][21], P[27][20], S[288], Cout[288]);
Half_Adder HA290 (P[28][19], P[29][18], S[289], Cout[289]);
Full_Adder FA291 (P[17][31], P[18][30], P[19][29], S[290], Cout[290]);
Full_Adder FA292 (P[20][28], P[21][27], P[22][26], S[291], Cout[291]);
Full_Adder FA293 (P[23][25], P[24][24], P[25][23], S[292], Cout[292]);
Full_Adder FA294 (P[26][22], P[27][21], P[28][20], S[293], Cout[293]);
Full_Adder FA295 (P[18][31], P[19][30], P[20][29], S[294], Cout[294]);
Full_Adder FA296 (P[21][28], P[22][27], P[23][26], S[295], Cout[295]);
Full_Adder FA297 (P[24][25], P[25][24], P[26][23], S[296], Cout[296]);
Full_Adder FA298 (P[27][22], P[28][21], P[29][20], S[297], Cout[297]);
Full_Adder FA299 (P[19][31], P[20][30], P[21][29], S[298], Cout[298]);
Full_Adder FA300 (P[22][28], P[23][27], P[24][26], S[299], Cout[299]);
Full_Adder FA301 (P[25][25], P[26][24], P[27][23], S[300], Cout[300]);
Half_Adder HA302 (P[28][22], P[29][21], S[301], Cout[301]);
Full_Adder FA303 (P[20][31], P[21][30], P[22][29], S[302], Cout[302]);
Full_Adder FA304 (P[23][28], P[24][27], P[25][26], S[303], Cout[303]);
Full_Adder FA305 (P[26][25], P[27][24], P[28][23], S[304], Cout[304]);
Full_Adder FA306 (P[21][31], P[22][30], P[23][29], S[305], Cout[305]);
Full_Adder FA307 (P[24][28], P[25][27], P[26][26], S[306], Cout[306]);
Full_Adder FA308 (P[27][25], P[28][24], P[29][23], S[307], Cout[307]);
Full_Adder FA309 (P[22][31], P[23][30], P[24][29], S[308], Cout[308]);
Full_Adder FA310 (P[25][28], P[26][27], P[27][26], S[309], Cout[309]);
Half_Adder HA311 (P[28][25], P[29][24], S[310], Cout[310]);
Full_Adder FA312 (P[23][31], P[24][30], P[25][29], S[311], Cout[311]);
Full_Adder FA313 (P[26][28], P[27][27], P[28][26], S[312], Cout[312]);
Full_Adder FA314 (P[24][31], P[25][30], P[26][29], S[313], Cout[313]);
Full_Adder FA315 (P[27][28], P[28][27], P[29][26], S[314], Cout[314]);
Full_Adder FA316 (P[25][31], P[26][30], P[27][29], S[315], Cout[315]);
Half_Adder HA317 (P[28][28], P[29][27], S[316], Cout[316]);
Full_Adder FA318 (P[26][31], P[27][30], P[28][29], S[317], Cout[317]);
Full_Adder FA319 (P[27][31], P[28][30], P[29][29], S[318], Cout[318]);
Half_Adder HA320 (P[28][31], P[29][30], S[319], Cout[319]);
Half_Adder HA321 (Cout[0], S[1], S[320], Cout[320]);
Full_Adder FA322 (P[3][0], Cout[1], S[2], S[321], Cout[321]);
Full_Adder FA323 (Cout[2], S[3], S[4], S[322], Cout[322]);
Full_Adder FA324 (Cout[3], Cout[4], S[5], S[323], Cout[323]);
Full_Adder FA325 (P[6][0], Cout[5], Cout[6], S[324], Cout[324]);
Half_Adder HA326 (S[7], S[8], S[325], Cout[325]);
Full_Adder FA327 (Cout[7], Cout[8], S[9], S[326], Cout[326]);
Half_Adder HA328 (S[10], S[11], S[327], Cout[327]);
Full_Adder FA329 (Cout[9], Cout[10], Cout[11], S[328], Cout[328]);
Full_Adder FA330 (S[12], S[13], S[14], S[329], Cout[329]);
Full_Adder FA331 (P[9][0], Cout[12], Cout[13], S[330], Cout[330]);
Full_Adder FA332 (Cout[14], S[15], S[16], S[331], Cout[331]);
Full_Adder FA333 (Cout[15], Cout[16], Cout[17], S[332], Cout[332]);
Full_Adder FA334 (S[18], S[19], S[20], S[333], Cout[333]);
Full_Adder FA335 (Cout[18], Cout[19], Cout[20], S[334], Cout[334]);
Full_Adder FA336 (Cout[21], S[22], S[23], S[335], Cout[335]);
Half_Adder HA337 (S[24], S[25], S[336], Cout[336]);
Full_Adder FA338 (P[12][0], Cout[22], Cout[23], S[337], Cout[337]);
Full_Adder FA339 (Cout[24], Cout[25], S[26], S[338], Cout[338]);
Full_Adder FA340 (S[27], S[28], S[29], S[339], Cout[339]);
Full_Adder FA341 (Cout[26], Cout[27], Cout[28], S[340], Cout[340]);
Full_Adder FA342 (Cout[29], S[30], S[31], S[341], Cout[341]);
Full_Adder FA343 (S[32], S[33], S[34], S[342], Cout[342]);
Full_Adder FA344 (Cout[30], Cout[31], Cout[32], S[343], Cout[343]);
Full_Adder FA345 (Cout[33], Cout[34], S[35], S[344], Cout[344]);
Full_Adder FA346 (S[36], S[37], S[38], S[345], Cout[345]);
Full_Adder FA347 (P[15][0], Cout[35], Cout[36], S[346], Cout[346]);
Full_Adder FA348 (Cout[37], Cout[38], Cout[39], S[347], Cout[347]);
Full_Adder FA349 (S[40], S[41], S[42], S[348], Cout[348]);
Half_Adder HA350 (S[43], S[44], S[349], Cout[349]);
Full_Adder FA351 (Cout[40], Cout[41], Cout[42], S[350], Cout[350]);
Full_Adder FA352 (Cout[43], Cout[44], S[45], S[351], Cout[351]);
Full_Adder FA353 (S[46], S[47], S[48], S[352], Cout[352]);
Half_Adder HA354 (S[49], S[50], S[353], Cout[353]);
Full_Adder FA355 (Cout[45], Cout[46], Cout[47], S[354], Cout[354]);
Full_Adder FA356 (Cout[48], Cout[49], Cout[50], S[355], Cout[355]);
Full_Adder FA357 (S[51], S[52], S[53], S[356], Cout[356]);
Full_Adder FA358 (S[54], S[55], S[56], S[357], Cout[357]);
Full_Adder FA359 (P[18][0], Cout[51], Cout[52], S[358], Cout[358]);
Full_Adder FA360 (Cout[53], Cout[54], Cout[55], S[359], Cout[359]);
Full_Adder FA361 (Cout[56], S[57], S[58], S[360], Cout[360]);
Full_Adder FA362 (S[59], S[60], S[61], S[361], Cout[361]);
Full_Adder FA363 (Cout[57], Cout[58], Cout[59], S[362], Cout[362]);
Full_Adder FA364 (Cout[60], Cout[61], Cout[62], S[363], Cout[363]);
Full_Adder FA365 (S[63], S[64], S[65], S[364], Cout[364]);
Full_Adder FA366 (S[66], S[67], S[68], S[365], Cout[365]);
Full_Adder FA367 (Cout[63], Cout[64], Cout[65], S[366], Cout[366]);
Full_Adder FA368 (Cout[66], Cout[67], Cout[68], S[367], Cout[367]);
Full_Adder FA369 (Cout[69], S[70], S[71], S[368], Cout[368]);
Full_Adder FA370 (S[72], S[73], S[74], S[369], Cout[369]);
Half_Adder HA371 (S[75], S[76], S[370], Cout[370]);
Full_Adder FA372 (P[21][0], Cout[70], Cout[71], S[371], Cout[371]);
Full_Adder FA373 (Cout[72], Cout[73], Cout[74], S[372], Cout[372]);
Full_Adder FA374 (Cout[75], Cout[76], S[77], S[373], Cout[373]);
Full_Adder FA375 (S[78], S[79], S[80], S[374], Cout[374]);
Full_Adder FA376 (S[81], S[82], S[83], S[375], Cout[375]);
Full_Adder FA377 (Cout[77], Cout[78], Cout[79], S[376], Cout[376]);
Full_Adder FA378 (Cout[80], Cout[81], Cout[82], S[377], Cout[377]);
Full_Adder FA379 (Cout[83], S[84], S[85], S[378], Cout[378]);
Full_Adder FA380 (S[86], S[87], S[88], S[379], Cout[379]);
Full_Adder FA381 (S[89], S[90], S[91], S[380], Cout[380]);
Full_Adder FA382 (Cout[84], Cout[85], Cout[86], S[381], Cout[381]);
Full_Adder FA383 (Cout[87], Cout[88], Cout[89], S[382], Cout[382]);
Full_Adder FA384 (Cout[90], Cout[91], S[92], S[383], Cout[383]);
Full_Adder FA385 (S[93], S[94], S[95], S[384], Cout[384]);
Full_Adder FA386 (S[96], S[97], S[98], S[385], Cout[385]);
Full_Adder FA387 (P[24][0], Cout[92], Cout[93], S[386], Cout[386]);
Full_Adder FA388 (Cout[94], Cout[95], Cout[96], S[387], Cout[387]);
Full_Adder FA389 (Cout[97], Cout[98], Cout[99], S[388], Cout[388]);
Full_Adder FA390 (S[100], S[101], S[102], S[389], Cout[389]);
Full_Adder FA391 (S[103], S[104], S[105], S[390], Cout[390]);
Half_Adder HA392 (S[106], S[107], S[391], Cout[391]);
Full_Adder FA393 (Cout[100], Cout[101], Cout[102], S[392], Cout[392]);
Full_Adder FA394 (Cout[103], Cout[104], Cout[105], S[393], Cout[393]);
Full_Adder FA395 (Cout[106], Cout[107], S[108], S[394], Cout[394]);
Full_Adder FA396 (S[109], S[110], S[111], S[395], Cout[395]);
Full_Adder FA397 (S[112], S[113], S[114], S[396], Cout[396]);
Half_Adder HA398 (S[115], S[116], S[397], Cout[397]);
Full_Adder FA399 (Cout[108], Cout[109], Cout[110], S[398], Cout[398]);
Full_Adder FA400 (Cout[111], Cout[112], Cout[113], S[399], Cout[399]);
Full_Adder FA401 (Cout[114], Cout[115], Cout[116], S[400], Cout[400]);
Full_Adder FA402 (S[117], S[118], S[119], S[401], Cout[401]);
Full_Adder FA403 (S[120], S[121], S[122], S[402], Cout[402]);
Full_Adder FA404 (S[123], S[124], S[125], S[403], Cout[403]);
Full_Adder FA405 (P[27][0], Cout[117], Cout[118], S[404], Cout[404]);
Full_Adder FA406 (Cout[119], Cout[120], Cout[121], S[405], Cout[405]);
Full_Adder FA407 (Cout[122], Cout[123], Cout[124], S[406], Cout[406]);
Full_Adder FA408 (Cout[125], S[126], S[127], S[407], Cout[407]);
Full_Adder FA409 (S[128], S[129], S[130], S[408], Cout[408]);
Full_Adder FA410 (S[131], S[132], S[133], S[409], Cout[409]);
Full_Adder FA411 (Cout[126], Cout[127], Cout[128], S[410], Cout[410]);
Full_Adder FA412 (Cout[129], Cout[130], Cout[131], S[411], Cout[411]);
Full_Adder FA413 (Cout[132], Cout[133], Cout[134], S[412], Cout[412]);
Full_Adder FA414 (S[135], S[136], S[137], S[413], Cout[413]);
Full_Adder FA415 (S[138], S[139], S[140], S[414], Cout[414]);
Full_Adder FA416 (S[141], S[142], S[143], S[415], Cout[415]);
Full_Adder FA417 (Cout[135], Cout[136], Cout[137], S[416], Cout[416]);
Full_Adder FA418 (Cout[138], Cout[139], Cout[140], S[417], Cout[417]);
Full_Adder FA419 (Cout[141], Cout[142], Cout[143], S[418], Cout[418]);
Full_Adder FA420 (Cout[144], S[145], S[146], S[419], Cout[419]);
Full_Adder FA421 (S[147], S[148], S[149], S[420], Cout[420]);
Full_Adder FA422 (S[150], S[151], S[152], S[421], Cout[421]);
Half_Adder HA423 (S[153], S[154], S[422], Cout[422]);
Full_Adder FA424 (P[30][0], Cout[145], Cout[146], S[423], Cout[423]);
Full_Adder FA425 (Cout[147], Cout[148], Cout[149], S[424], Cout[424]);
Full_Adder FA426 (Cout[150], Cout[151], Cout[152], S[425], Cout[425]);
Full_Adder FA427 (Cout[153], Cout[154], S[155], S[426], Cout[426]);
Full_Adder FA428 (S[156], S[157], S[158], S[427], Cout[427]);
Full_Adder FA429 (S[159], S[160], S[161], S[428], Cout[428]);
Full_Adder FA430 (S[162], S[163], S[164], S[429], Cout[429]);
Full_Adder FA431 (P[30][1], P[31][0], Cout[155], S[430], Cout[430]);
Full_Adder FA432 (Cout[156], Cout[157], Cout[158], S[431], Cout[431]);
Full_Adder FA433 (Cout[159], Cout[160], Cout[161], S[432], Cout[432]);
Full_Adder FA434 (Cout[162], Cout[163], Cout[164], S[433], Cout[433]);
Full_Adder FA435 (S[165], S[166], S[167], S[434], Cout[434]);
Full_Adder FA436 (S[168], S[169], S[170], S[435], Cout[435]);
Full_Adder FA437 (S[171], S[172], S[173], S[436], Cout[436]);
Full_Adder FA438 (P[30][2], P[31][1], Cout[165], S[437], Cout[437]);
Full_Adder FA439 (Cout[166], Cout[167], Cout[168], S[438], Cout[438]);
Full_Adder FA440 (Cout[169], Cout[170], Cout[171], S[439], Cout[439]);
Full_Adder FA441 (Cout[172], Cout[173], Cout[174], S[440], Cout[440]);
Full_Adder FA442 (S[175], S[176], S[177], S[441], Cout[441]);
Full_Adder FA443 (S[178], S[179], S[180], S[442], Cout[442]);
Full_Adder FA444 (S[181], S[182], S[183], S[443], Cout[443]);
Full_Adder FA445 (P[29][4], P[30][3], P[31][2], S[444], Cout[444]);
Full_Adder FA446 (Cout[175], Cout[176], Cout[177], S[445], Cout[445]);
Full_Adder FA447 (Cout[178], Cout[179], Cout[180], S[446], Cout[446]);
Full_Adder FA448 (Cout[181], Cout[182], Cout[183], S[447], Cout[447]);
Full_Adder FA449 (Cout[184], S[185], S[186], S[448], Cout[448]);
Full_Adder FA450 (S[187], S[188], S[189], S[449], Cout[449]);
Full_Adder FA451 (S[190], S[191], S[192], S[450], Cout[450]);
Full_Adder FA452 (P[30][4], P[31][3], Cout[185], S[451], Cout[451]);
Full_Adder FA453 (Cout[186], Cout[187], Cout[188], S[452], Cout[452]);
Full_Adder FA454 (Cout[189], Cout[190], Cout[191], S[453], Cout[453]);
Full_Adder FA455 (Cout[192], Cout[193], S[194], S[454], Cout[454]);
Full_Adder FA456 (S[195], S[196], S[197], S[455], Cout[455]);
Full_Adder FA457 (S[198], S[199], S[200], S[456], Cout[456]);
Full_Adder FA458 (P[30][5], P[31][4], Cout[194], S[457], Cout[457]);
Full_Adder FA459 (Cout[195], Cout[196], Cout[197], S[458], Cout[458]);
Full_Adder FA460 (Cout[198], Cout[199], Cout[200], S[459], Cout[459]);
Full_Adder FA461 (Cout[201], Cout[202], S[203], S[460], Cout[460]);
Full_Adder FA462 (S[204], S[205], S[206], S[461], Cout[461]);
Full_Adder FA463 (S[207], S[208], S[209], S[462], Cout[462]);
Full_Adder FA464 (P[29][7], P[30][6], P[31][5], S[463], Cout[463]);
Full_Adder FA465 (Cout[203], Cout[204], Cout[205], S[464], Cout[464]);
Full_Adder FA466 (Cout[206], Cout[207], Cout[208], S[465], Cout[465]);
Full_Adder FA467 (Cout[209], Cout[210], Cout[211], S[466], Cout[466]);
Full_Adder FA468 (S[212], S[213], S[214], S[467], Cout[467]);
Full_Adder FA469 (S[215], S[216], S[217], S[468], Cout[468]);
Full_Adder FA470 (P[30][7], P[31][6], Cout[212], S[469], Cout[469]);
Full_Adder FA471 (Cout[213], Cout[214], Cout[215], S[470], Cout[470]);
Full_Adder FA472 (Cout[216], Cout[217], Cout[218], S[471], Cout[471]);
Full_Adder FA473 (Cout[219], S[220], S[221], S[472], Cout[472]);
Full_Adder FA474 (S[222], S[223], S[224], S[473], Cout[473]);
Half_Adder HA475 (S[225], S[226], S[474], Cout[474]);
Full_Adder FA476 (P[30][8], P[31][7], Cout[220], S[475], Cout[475]);
Full_Adder FA477 (Cout[221], Cout[222], Cout[223], S[476], Cout[476]);
Full_Adder FA478 (Cout[224], Cout[225], Cout[226], S[477], Cout[477]);
Full_Adder FA479 (Cout[227], S[228], S[229], S[478], Cout[478]);
Full_Adder FA480 (S[230], S[231], S[232], S[479], Cout[479]);
Half_Adder HA481 (S[233], S[234], S[480], Cout[480]);
Full_Adder FA482 (P[29][10], P[30][9], P[31][8], S[481], Cout[481]);
Full_Adder FA483 (Cout[228], Cout[229], Cout[230], S[482], Cout[482]);
Full_Adder FA484 (Cout[231], Cout[232], Cout[233], S[483], Cout[483]);
Full_Adder FA485 (Cout[234], Cout[235], S[236], S[484], Cout[484]);
Full_Adder FA486 (S[237], S[238], S[239], S[485], Cout[485]);
Half_Adder HA487 (S[240], S[241], S[486], Cout[486]);
Full_Adder FA488 (P[30][10], P[31][9], Cout[236], S[487], Cout[487]);
Full_Adder FA489 (Cout[237], Cout[238], Cout[239], S[488], Cout[488]);
Full_Adder FA490 (Cout[240], Cout[241], Cout[242], S[489], Cout[489]);
Full_Adder FA491 (S[243], S[244], S[245], S[490], Cout[490]);
Full_Adder FA492 (S[246], S[247], S[248], S[491], Cout[491]);
Full_Adder FA493 (P[30][11], P[31][10], Cout[243], S[492], Cout[492]);
Full_Adder FA494 (Cout[244], Cout[245], Cout[246], S[493], Cout[493]);
Full_Adder FA495 (Cout[247], Cout[248], Cout[249], S[494], Cout[494]);
Full_Adder FA496 (S[250], S[251], S[252], S[495], Cout[495]);
Full_Adder FA497 (S[253], S[254], S[255], S[496], Cout[496]);
Full_Adder FA498 (P[29][13], P[30][12], P[31][11], S[497], Cout[497]);
Full_Adder FA499 (Cout[250], Cout[251], Cout[252], S[498], Cout[498]);
Full_Adder FA500 (Cout[253], Cout[254], Cout[255], S[499], Cout[499]);
Full_Adder FA501 (Cout[256], S[257], S[258], S[500], Cout[500]);
Full_Adder FA502 (S[259], S[260], S[261], S[501], Cout[501]);
Full_Adder FA503 (P[30][13], P[31][12], Cout[257], S[502], Cout[502]);
Full_Adder FA504 (Cout[258], Cout[259], Cout[260], S[503], Cout[503]);
Full_Adder FA505 (Cout[261], Cout[262], S[263], S[504], Cout[504]);
Full_Adder FA506 (S[264], S[265], S[266], S[505], Cout[505]);
Full_Adder FA507 (P[30][14], P[31][13], Cout[263], S[506], Cout[506]);
Full_Adder FA508 (Cout[264], Cout[265], Cout[266], S[507], Cout[507]);
Full_Adder FA509 (Cout[267], Cout[268], S[269], S[508], Cout[508]);
Full_Adder FA510 (S[270], S[271], S[272], S[509], Cout[509]);
Full_Adder FA511 (P[29][16], P[30][15], P[31][14], S[510], Cout[510]);
Full_Adder FA512 (Cout[269], Cout[270], Cout[271], S[511], Cout[511]);
Full_Adder FA513 (Cout[272], Cout[273], Cout[274], S[512], Cout[512]);
Full_Adder FA514 (S[275], S[276], S[277], S[513], Cout[513]);
Full_Adder FA515 (P[30][16], P[31][15], Cout[275], S[514], Cout[514]);
Full_Adder FA516 (Cout[276], Cout[277], Cout[278], S[515], Cout[515]);
Full_Adder FA517 (Cout[279], S[280], S[281], S[516], Cout[516]);
Half_Adder HA518 (S[282], S[283], S[517], Cout[517]);
Full_Adder FA519 (P[30][17], P[31][16], Cout[280], S[518], Cout[518]);
Full_Adder FA520 (Cout[281], Cout[282], Cout[283], S[519], Cout[519]);
Full_Adder FA521 (Cout[284], S[285], S[286], S[520], Cout[520]);
Half_Adder HA522 (S[287], S[288], S[521], Cout[521]);
Full_Adder FA523 (P[29][19], P[30][18], P[31][17], S[522], Cout[522]);
Full_Adder FA524 (Cout[285], Cout[286], Cout[287], S[523], Cout[523]);
Full_Adder FA525 (Cout[288], Cout[289], S[290], S[524], Cout[524]);
Half_Adder HA526 (S[291], S[292], S[525], Cout[525]);
Full_Adder FA527 (P[30][19], P[31][18], Cout[290], S[526], Cout[526]);
Full_Adder FA528 (Cout[291], Cout[292], Cout[293], S[527], Cout[527]);
Full_Adder FA529 (S[294], S[295], S[296], S[528], Cout[528]);
Full_Adder FA530 (P[30][20], P[31][19], Cout[294], S[529], Cout[529]);
Full_Adder FA531 (Cout[295], Cout[296], Cout[297], S[530], Cout[530]);
Full_Adder FA532 (S[298], S[299], S[300], S[531], Cout[531]);
Full_Adder FA533 (P[29][22], P[30][21], P[31][20], S[532], Cout[532]);
Full_Adder FA534 (Cout[298], Cout[299], Cout[300], S[533], Cout[533]);
Full_Adder FA535 (Cout[301], S[302], S[303], S[534], Cout[534]);
Full_Adder FA536 (P[30][22], P[31][21], Cout[302], S[535], Cout[535]);
Full_Adder FA537 (Cout[303], Cout[304], S[305], S[536], Cout[536]);
Full_Adder FA538 (P[30][23], P[31][22], Cout[305], S[537], Cout[537]);
Full_Adder FA539 (Cout[306], Cout[307], S[308], S[538], Cout[538]);
Full_Adder FA540 (P[29][25], P[30][24], P[31][23], S[539], Cout[539]);
Full_Adder FA541 (Cout[308], Cout[309], Cout[310], S[540], Cout[540]);
Full_Adder FA542 (P[30][25], P[31][24], Cout[311], S[541], Cout[541]);
Half_Adder HA543 (Cout[312], S[313], S[542], Cout[542]);
Full_Adder FA544 (P[30][26], P[31][25], Cout[313], S[543], Cout[543]);
Half_Adder HA545 (Cout[314], S[315], S[544], Cout[544]);
Full_Adder FA546 (P[29][28], P[30][27], P[31][26], S[545], Cout[545]);
Half_Adder HA547 (Cout[315], Cout[316], S[546], Cout[546]);
Full_Adder FA548 (P[30][28], P[31][27], Cout[317], S[547], Cout[547]);
Full_Adder FA549 (P[30][29], P[31][28], Cout[318], S[548], Cout[548]);
Full_Adder FA550 (P[29][31], P[30][30], P[31][29], S[549], Cout[549]);
Half_Adder HA551 (Cout[320], S[321], S[550], Cout[550]);
Half_Adder HA552 (Cout[321], S[322], S[551], Cout[551]);
Full_Adder FA553 (S[6], Cout[322], S[323], S[552], Cout[552]);
Full_Adder FA554 (Cout[323], S[324], S[325], S[553], Cout[553]);
Full_Adder FA555 (Cout[324], Cout[325], S[326], S[554], Cout[554]);
Full_Adder FA556 (Cout[326], Cout[327], S[328], S[555], Cout[555]);
Full_Adder FA557 (S[17], Cout[328], Cout[329], S[556], Cout[556]);
Half_Adder HA558 (S[330], S[331], S[557], Cout[557]);
Full_Adder FA559 (S[21], Cout[330], Cout[331], S[558], Cout[558]);
Half_Adder HA560 (S[332], S[333], S[559], Cout[559]);
Full_Adder FA561 (Cout[332], Cout[333], S[334], S[560], Cout[560]);
Half_Adder HA562 (S[335], S[336], S[561], Cout[561]);
Full_Adder FA563 (Cout[334], Cout[335], Cout[336], S[562], Cout[562]);
Full_Adder FA564 (S[337], S[338], S[339], S[563], Cout[563]);
Full_Adder FA565 (Cout[337], Cout[338], Cout[339], S[564], Cout[564]);
Full_Adder FA566 (S[340], S[341], S[342], S[565], Cout[565]);
Full_Adder FA567 (S[39], Cout[340], Cout[341], S[566], Cout[566]);
Full_Adder FA568 (Cout[342], S[343], S[344], S[567], Cout[567]);
Full_Adder FA569 (Cout[343], Cout[344], Cout[345], S[568], Cout[568]);
Full_Adder FA570 (S[346], S[347], S[348], S[569], Cout[569]);
Full_Adder FA571 (Cout[346], Cout[347], Cout[348], S[570], Cout[570]);
Full_Adder FA572 (Cout[349], S[350], S[351], S[571], Cout[571]);
Half_Adder HA573 (S[352], S[353], S[572], Cout[572]);
Full_Adder FA574 (Cout[350], Cout[351], Cout[352], S[573], Cout[573]);
Full_Adder FA575 (Cout[353], S[354], S[355], S[574], Cout[574]);
Half_Adder HA576 (S[356], S[357], S[575], Cout[575]);
Full_Adder FA577 (S[62], Cout[354], Cout[355], S[576], Cout[576]);
Full_Adder FA578 (Cout[356], Cout[357], S[358], S[577], Cout[577]);
Full_Adder FA579 (S[359], S[360], S[361], S[578], Cout[578]);
Full_Adder FA580 (S[69], Cout[358], Cout[359], S[579], Cout[579]);
Full_Adder FA581 (Cout[360], Cout[361], S[362], S[580], Cout[580]);
Full_Adder FA582 (S[363], S[364], S[365], S[581], Cout[581]);
Full_Adder FA583 (Cout[362], Cout[363], Cout[364], S[582], Cout[582]);
Full_Adder FA584 (Cout[365], S[366], S[367], S[583], Cout[583]);
Full_Adder FA585 (S[368], S[369], S[370], S[584], Cout[584]);
Full_Adder FA586 (Cout[366], Cout[367], Cout[368], S[585], Cout[585]);
Full_Adder FA587 (Cout[369], Cout[370], S[371], S[586], Cout[586]);
Full_Adder FA588 (S[372], S[373], S[374], S[587], Cout[587]);
Full_Adder FA589 (Cout[371], Cout[372], Cout[373], S[588], Cout[588]);
Full_Adder FA590 (Cout[374], Cout[375], S[376], S[589], Cout[589]);
Full_Adder FA591 (S[377], S[378], S[379], S[590], Cout[590]);
Full_Adder FA592 (S[99], Cout[376], Cout[377], S[591], Cout[591]);
Full_Adder FA593 (Cout[378], Cout[379], Cout[380], S[592], Cout[592]);
Full_Adder FA594 (S[381], S[382], S[383], S[593], Cout[593]);
Half_Adder HA595 (S[384], S[385], S[594], Cout[594]);
Full_Adder FA596 (Cout[381], Cout[382], Cout[383], S[595], Cout[595]);
Full_Adder FA597 (Cout[384], Cout[385], S[386], S[596], Cout[596]);
Full_Adder FA598 (S[387], S[388], S[389], S[597], Cout[597]);
Half_Adder HA599 (S[390], S[391], S[598], Cout[598]);
Full_Adder FA600 (Cout[386], Cout[387], Cout[388], S[599], Cout[599]);
Full_Adder FA601 (Cout[389], Cout[390], Cout[391], S[600], Cout[600]);
Full_Adder FA602 (S[392], S[393], S[394], S[601], Cout[601]);
Full_Adder FA603 (S[395], S[396], S[397], S[602], Cout[602]);
Full_Adder FA604 (Cout[392], Cout[393], Cout[394], S[603], Cout[603]);
Full_Adder FA605 (Cout[395], Cout[396], Cout[397], S[604], Cout[604]);
Full_Adder FA606 (S[398], S[399], S[400], S[605], Cout[605]);
Full_Adder FA607 (S[401], S[402], S[403], S[606], Cout[606]);
Full_Adder FA608 (S[134], Cout[398], Cout[399], S[607], Cout[607]);
Full_Adder FA609 (Cout[400], Cout[401], Cout[402], S[608], Cout[608]);
Full_Adder FA610 (Cout[403], S[404], S[405], S[609], Cout[609]);
Full_Adder FA611 (S[406], S[407], S[408], S[610], Cout[610]);
Full_Adder FA612 (S[144], Cout[404], Cout[405], S[611], Cout[611]);
Full_Adder FA613 (Cout[406], Cout[407], Cout[408], S[612], Cout[612]);
Full_Adder FA614 (Cout[409], S[410], S[411], S[613], Cout[613]);
Full_Adder FA615 (S[412], S[413], S[414], S[614], Cout[614]);
Full_Adder FA616 (Cout[410], Cout[411], Cout[412], S[615], Cout[615]);
Full_Adder FA617 (Cout[413], Cout[414], Cout[415], S[616], Cout[616]);
Full_Adder FA618 (S[416], S[417], S[418], S[617], Cout[617]);
Full_Adder FA619 (S[419], S[420], S[421], S[618], Cout[618]);
Full_Adder FA620 (Cout[416], Cout[417], Cout[418], S[619], Cout[619]);
Full_Adder FA621 (Cout[419], Cout[420], Cout[421], S[620], Cout[620]);
Full_Adder FA622 (Cout[422], S[423], S[424], S[621], Cout[621]);
Full_Adder FA623 (S[425], S[426], S[427], S[622], Cout[622]);
Half_Adder HA624 (S[428], S[429], S[623], Cout[623]);
Full_Adder FA625 (S[174], Cout[423], Cout[424], S[624], Cout[624]);
Full_Adder FA626 (Cout[425], Cout[426], Cout[427], S[625], Cout[625]);
Full_Adder FA627 (Cout[428], Cout[429], S[430], S[626], Cout[626]);
Full_Adder FA628 (S[431], S[432], S[433], S[627], Cout[627]);
Full_Adder FA629 (S[434], S[435], S[436], S[628], Cout[628]);
Full_Adder FA630 (S[184], Cout[430], Cout[431], S[629], Cout[629]);
Full_Adder FA631 (Cout[432], Cout[433], Cout[434], S[630], Cout[630]);
Full_Adder FA632 (Cout[435], Cout[436], S[437], S[631], Cout[631]);
Full_Adder FA633 (S[438], S[439], S[440], S[632], Cout[632]);
Full_Adder FA634 (S[441], S[442], S[443], S[633], Cout[633]);
Full_Adder FA635 (S[193], Cout[437], Cout[438], S[634], Cout[634]);
Full_Adder FA636 (Cout[439], Cout[440], Cout[441], S[635], Cout[635]);
Full_Adder FA637 (Cout[442], Cout[443], S[444], S[636], Cout[636]);
Full_Adder FA638 (S[445], S[446], S[447], S[637], Cout[637]);
Full_Adder FA639 (S[448], S[449], S[450], S[638], Cout[638]);
Full_Adder FA640 (S[201], S[202], Cout[444], S[639], Cout[639]);
Full_Adder FA641 (Cout[445], Cout[446], Cout[447], S[640], Cout[640]);
Full_Adder FA642 (Cout[448], Cout[449], Cout[450], S[641], Cout[641]);
Full_Adder FA643 (S[451], S[452], S[453], S[642], Cout[642]);
Full_Adder FA644 (S[454], S[455], S[456], S[643], Cout[643]);
Full_Adder FA645 (S[210], S[211], Cout[451], S[644], Cout[644]);
Full_Adder FA646 (Cout[452], Cout[453], Cout[454], S[645], Cout[645]);
Full_Adder FA647 (Cout[455], Cout[456], S[457], S[646], Cout[646]);
Full_Adder FA648 (S[458], S[459], S[460], S[647], Cout[647]);
Half_Adder HA649 (S[461], S[462], S[648], Cout[648]);
Full_Adder FA650 (S[218], S[219], Cout[457], S[649], Cout[649]);
Full_Adder FA651 (Cout[458], Cout[459], Cout[460], S[650], Cout[650]);
Full_Adder FA652 (Cout[461], Cout[462], S[463], S[651], Cout[651]);
Full_Adder FA653 (S[464], S[465], S[466], S[652], Cout[652]);
Half_Adder HA654 (S[467], S[468], S[653], Cout[653]);
Full_Adder FA655 (S[227], Cout[463], Cout[464], S[654], Cout[654]);
Full_Adder FA656 (Cout[465], Cout[466], Cout[467], S[655], Cout[655]);
Full_Adder FA657 (Cout[468], S[469], S[470], S[656], Cout[656]);
Full_Adder FA658 (S[471], S[472], S[473], S[657], Cout[657]);
Full_Adder FA659 (S[235], Cout[469], Cout[470], S[658], Cout[658]);
Full_Adder FA660 (Cout[471], Cout[472], Cout[473], S[659], Cout[659]);
Full_Adder FA661 (Cout[474], S[475], S[476], S[660], Cout[660]);
Full_Adder FA662 (S[477], S[478], S[479], S[661], Cout[661]);
Full_Adder FA663 (S[242], Cout[475], Cout[476], S[662], Cout[662]);
Full_Adder FA664 (Cout[477], Cout[478], Cout[479], S[663], Cout[663]);
Full_Adder FA665 (Cout[480], S[481], S[482], S[664], Cout[664]);
Full_Adder FA666 (S[483], S[484], S[485], S[665], Cout[665]);
Full_Adder FA667 (S[249], Cout[481], Cout[482], S[666], Cout[666]);
Full_Adder FA668 (Cout[483], Cout[484], Cout[485], S[667], Cout[667]);
Full_Adder FA669 (Cout[486], S[487], S[488], S[668], Cout[668]);
Full_Adder FA670 (S[489], S[490], S[491], S[669], Cout[669]);
Full_Adder FA671 (S[256], Cout[487], Cout[488], S[670], Cout[670]);
Full_Adder FA672 (Cout[489], Cout[490], Cout[491], S[671], Cout[671]);
Full_Adder FA673 (S[492], S[493], S[494], S[672], Cout[672]);
Half_Adder HA674 (S[495], S[496], S[673], Cout[673]);
Full_Adder FA675 (S[262], Cout[492], Cout[493], S[674], Cout[674]);
Full_Adder FA676 (Cout[494], Cout[495], Cout[496], S[675], Cout[675]);
Full_Adder FA677 (S[497], S[498], S[499], S[676], Cout[676]);
Half_Adder HA678 (S[500], S[501], S[677], Cout[677]);
Full_Adder FA679 (S[267], S[268], Cout[497], S[678], Cout[678]);
Full_Adder FA680 (Cout[498], Cout[499], Cout[500], S[679], Cout[679]);
Full_Adder FA681 (Cout[501], S[502], S[503], S[680], Cout[680]);
Half_Adder HA682 (S[504], S[505], S[681], Cout[681]);
Full_Adder FA683 (S[273], S[274], Cout[502], S[682], Cout[682]);
Full_Adder FA684 (Cout[503], Cout[504], Cout[505], S[683], Cout[683]);
Full_Adder FA685 (S[506], S[507], S[508], S[684], Cout[684]);
Full_Adder FA686 (S[278], S[279], Cout[506], S[685], Cout[685]);
Full_Adder FA687 (Cout[507], Cout[508], Cout[509], S[686], Cout[686]);
Full_Adder FA688 (S[510], S[511], S[512], S[687], Cout[687]);
Full_Adder FA689 (S[284], Cout[510], Cout[511], S[688], Cout[688]);
Full_Adder FA690 (Cout[512], Cout[513], S[514], S[689], Cout[689]);
Full_Adder FA691 (S[515], S[516], S[517], S[690], Cout[690]);
Full_Adder FA692 (S[289], Cout[514], Cout[515], S[691], Cout[691]);
Full_Adder FA693 (Cout[516], Cout[517], S[518], S[692], Cout[692]);
Full_Adder FA694 (S[519], S[520], S[521], S[693], Cout[693]);
Full_Adder FA695 (S[293], Cout[518], Cout[519], S[694], Cout[694]);
Full_Adder FA696 (Cout[520], Cout[521], S[522], S[695], Cout[695]);
Full_Adder FA697 (S[523], S[524], S[525], S[696], Cout[696]);
Full_Adder FA698 (S[297], Cout[522], Cout[523], S[697], Cout[697]);
Full_Adder FA699 (Cout[524], Cout[525], S[526], S[698], Cout[698]);
Half_Adder HA700 (S[527], S[528], S[699], Cout[699]);
Full_Adder FA701 (S[301], Cout[526], Cout[527], S[700], Cout[700]);
Full_Adder FA702 (Cout[528], S[529], S[530], S[701], Cout[701]);
Full_Adder FA703 (S[304], Cout[529], Cout[530], S[702], Cout[702]);
Full_Adder FA704 (Cout[531], S[532], S[533], S[703], Cout[703]);
Full_Adder FA705 (S[306], S[307], Cout[532], S[704], Cout[704]);
Full_Adder FA706 (Cout[533], Cout[534], S[535], S[705], Cout[705]);
Full_Adder FA707 (S[309], S[310], Cout[535], S[706], Cout[706]);
Full_Adder FA708 (Cout[536], S[537], S[538], S[707], Cout[707]);
Full_Adder FA709 (S[311], S[312], Cout[537], S[708], Cout[708]);
Full_Adder FA710 (Cout[538], S[539], S[540], S[709], Cout[709]);
Full_Adder FA711 (S[314], Cout[539], Cout[540], S[710], Cout[710]);
Half_Adder HA712 (S[541], S[542], S[711], Cout[711]);
Full_Adder FA713 (S[316], Cout[541], Cout[542], S[712], Cout[712]);
Half_Adder HA714 (S[543], S[544], S[713], Cout[713]);
Full_Adder FA715 (S[317], Cout[543], Cout[544], S[714], Cout[714]);
Half_Adder HA716 (S[545], S[546], S[715], Cout[715]);
Full_Adder FA717 (S[318], Cout[545], Cout[546], S[716], Cout[716]);
Full_Adder FA718 (S[319], Cout[547], S[548], S[717], Cout[717]);
Full_Adder FA719 (Cout[319], Cout[548], S[549], S[718], Cout[718]);
Full_Adder FA720 (P[30][31], P[31][30], Cout[549], S[719], Cout[719]);
Half_Adder HA721 (Cout[550], S[551], S[720], Cout[720]);
Half_Adder HA722 (Cout[551], S[552], S[721], Cout[721]);
Half_Adder HA723 (Cout[552], S[553], S[722], Cout[722]);
Full_Adder FA724 (S[327], Cout[553], S[554], S[723], Cout[723]);
Full_Adder FA725 (S[329], Cout[554], S[555], S[724], Cout[724]);
Full_Adder FA726 (Cout[555], S[556], S[557], S[725], Cout[725]);
Full_Adder FA727 (Cout[556], Cout[557], S[558], S[726], Cout[726]);
Full_Adder FA728 (Cout[558], Cout[559], S[560], S[727], Cout[727]);
Full_Adder FA729 (Cout[560], Cout[561], S[562], S[728], Cout[728]);
Full_Adder FA730 (Cout[562], Cout[563], S[564], S[729], Cout[729]);
Full_Adder FA731 (S[345], Cout[564], Cout[565], S[730], Cout[730]);
Half_Adder HA732 (S[566], S[567], S[731], Cout[731]);
Full_Adder FA733 (S[349], Cout[566], Cout[567], S[732], Cout[732]);
Half_Adder HA734 (S[568], S[569], S[733], Cout[733]);
Full_Adder FA735 (Cout[568], Cout[569], S[570], S[734], Cout[734]);
Half_Adder HA736 (S[571], S[572], S[735], Cout[735]);
Full_Adder FA737 (Cout[570], Cout[571], Cout[572], S[736], Cout[736]);
Full_Adder FA738 (S[573], S[574], S[575], S[737], Cout[737]);
Full_Adder FA739 (Cout[573], Cout[574], Cout[575], S[738], Cout[738]);
Full_Adder FA740 (S[576], S[577], S[578], S[739], Cout[739]);
Full_Adder FA741 (Cout[576], Cout[577], Cout[578], S[740], Cout[740]);
Full_Adder FA742 (S[579], S[580], S[581], S[741], Cout[741]);
Full_Adder FA743 (Cout[579], Cout[580], Cout[581], S[742], Cout[742]);
Full_Adder FA744 (S[582], S[583], S[584], S[743], Cout[743]);
Full_Adder FA745 (S[375], Cout[582], Cout[583], S[744], Cout[744]);
Full_Adder FA746 (Cout[584], S[585], S[586], S[745], Cout[745]);
Full_Adder FA747 (S[380], Cout[585], Cout[586], S[746], Cout[746]);
Full_Adder FA748 (Cout[587], S[588], S[589], S[747], Cout[747]);
Full_Adder FA749 (Cout[588], Cout[589], Cout[590], S[748], Cout[748]);
Full_Adder FA750 (S[591], S[592], S[593], S[749], Cout[749]);
Full_Adder FA751 (Cout[591], Cout[592], Cout[593], S[750], Cout[750]);
Full_Adder FA752 (Cout[594], S[595], S[596], S[751], Cout[751]);
Half_Adder HA753 (S[597], S[598], S[752], Cout[752]);
Full_Adder FA754 (Cout[595], Cout[596], Cout[597], S[753], Cout[753]);
Full_Adder FA755 (Cout[598], S[599], S[600], S[754], Cout[754]);
Half_Adder HA756 (S[601], S[602], S[755], Cout[755]);
Full_Adder FA757 (Cout[599], Cout[600], Cout[601], S[756], Cout[756]);
Full_Adder FA758 (Cout[602], S[603], S[604], S[757], Cout[757]);
Half_Adder HA759 (S[605], S[606], S[758], Cout[758]);
Full_Adder FA760 (S[409], Cout[603], Cout[604], S[759], Cout[759]);
Full_Adder FA761 (Cout[605], Cout[606], S[607], S[760], Cout[760]);
Full_Adder FA762 (S[608], S[609], S[610], S[761], Cout[761]);
Full_Adder FA763 (S[415], Cout[607], Cout[608], S[762], Cout[762]);
Full_Adder FA764 (Cout[609], Cout[610], S[611], S[763], Cout[763]);
Full_Adder FA765 (S[612], S[613], S[614], S[764], Cout[764]);
Full_Adder FA766 (S[422], Cout[611], Cout[612], S[765], Cout[765]);
Full_Adder FA767 (Cout[613], Cout[614], S[615], S[766], Cout[766]);
Full_Adder FA768 (S[616], S[617], S[618], S[767], Cout[767]);
Full_Adder FA769 (Cout[615], Cout[616], Cout[617], S[768], Cout[768]);
Full_Adder FA770 (Cout[618], S[619], S[620], S[769], Cout[769]);
Full_Adder FA771 (S[621], S[622], S[623], S[770], Cout[770]);
Full_Adder FA772 (Cout[619], Cout[620], Cout[621], S[771], Cout[771]);
Full_Adder FA773 (Cout[622], Cout[623], S[624], S[772], Cout[772]);
Full_Adder FA774 (S[625], S[626], S[627], S[773], Cout[773]);
Full_Adder FA775 (Cout[624], Cout[625], Cout[626], S[774], Cout[774]);
Full_Adder FA776 (Cout[627], Cout[628], S[629], S[775], Cout[775]);
Full_Adder FA777 (S[630], S[631], S[632], S[776], Cout[776]);
Full_Adder FA778 (Cout[629], Cout[630], Cout[631], S[777], Cout[777]);
Full_Adder FA779 (Cout[632], Cout[633], S[634], S[778], Cout[778]);
Full_Adder FA780 (S[635], S[636], S[637], S[779], Cout[779]);
Full_Adder FA781 (Cout[634], Cout[635], Cout[636], S[780], Cout[780]);
Full_Adder FA782 (Cout[637], Cout[638], S[639], S[781], Cout[781]);
Full_Adder FA783 (S[640], S[641], S[642], S[782], Cout[782]);
Full_Adder FA784 (Cout[639], Cout[640], Cout[641], S[783], Cout[783]);
Full_Adder FA785 (Cout[642], Cout[643], S[644], S[784], Cout[784]);
Full_Adder FA786 (S[645], S[646], S[647], S[785], Cout[785]);
Full_Adder FA787 (Cout[644], Cout[645], Cout[646], S[786], Cout[786]);
Full_Adder FA788 (Cout[647], Cout[648], S[649], S[787], Cout[787]);
Full_Adder FA789 (S[650], S[651], S[652], S[788], Cout[788]);
Full_Adder FA790 (S[474], Cout[649], Cout[650], S[789], Cout[789]);
Full_Adder FA791 (Cout[651], Cout[652], Cout[653], S[790], Cout[790]);
Full_Adder FA792 (S[654], S[655], S[656], S[791], Cout[791]);
Full_Adder FA793 (S[480], Cout[654], Cout[655], S[792], Cout[792]);
Full_Adder FA794 (Cout[656], Cout[657], S[658], S[793], Cout[793]);
Half_Adder HA795 (S[659], S[660], S[794], Cout[794]);
Full_Adder FA796 (S[486], Cout[658], Cout[659], S[795], Cout[795]);
Full_Adder FA797 (Cout[660], Cout[661], S[662], S[796], Cout[796]);
Half_Adder HA798 (S[663], S[664], S[797], Cout[797]);
Full_Adder FA799 (Cout[662], Cout[663], Cout[664], S[798], Cout[798]);
Full_Adder FA800 (Cout[665], S[666], S[667], S[799], Cout[799]);
Full_Adder FA801 (Cout[666], Cout[667], Cout[668], S[800], Cout[800]);
Full_Adder FA802 (Cout[669], S[670], S[671], S[801], Cout[801]);
Full_Adder FA803 (Cout[670], Cout[671], Cout[672], S[802], Cout[802]);
Full_Adder FA804 (Cout[673], S[674], S[675], S[803], Cout[803]);
Full_Adder FA805 (Cout[674], Cout[675], Cout[676], S[804], Cout[804]);
Full_Adder FA806 (Cout[677], S[678], S[679], S[805], Cout[805]);
Full_Adder FA807 (S[509], Cout[678], Cout[679], S[806], Cout[806]);
Full_Adder FA808 (Cout[680], Cout[681], S[682], S[807], Cout[807]);
Full_Adder FA809 (S[513], Cout[682], Cout[683], S[808], Cout[808]);
Full_Adder FA810 (Cout[684], S[685], S[686], S[809], Cout[809]);
Full_Adder FA811 (Cout[685], Cout[686], Cout[687], S[810], Cout[810]);
Half_Adder HA812 (S[688], S[689], S[811], Cout[811]);
Full_Adder FA813 (Cout[688], Cout[689], Cout[690], S[812], Cout[812]);
Half_Adder HA814 (S[691], S[692], S[813], Cout[813]);
Full_Adder FA815 (Cout[691], Cout[692], Cout[693], S[814], Cout[814]);
Half_Adder HA816 (S[694], S[695], S[815], Cout[815]);
Full_Adder FA817 (Cout[694], Cout[695], Cout[696], S[816], Cout[816]);
Half_Adder HA818 (S[697], S[698], S[817], Cout[817]);
Full_Adder FA819 (S[531], Cout[697], Cout[698], S[818], Cout[818]);
Half_Adder HA820 (Cout[699], S[700], S[819], Cout[819]);
Full_Adder FA821 (S[534], Cout[700], Cout[701], S[820], Cout[820]);
Full_Adder FA822 (S[536], Cout[702], Cout[703], S[821], Cout[821]);
Full_Adder FA823 (Cout[704], Cout[705], S[706], S[822], Cout[822]);
Full_Adder FA824 (Cout[706], Cout[707], S[708], S[823], Cout[823]);
Full_Adder FA825 (Cout[708], Cout[709], S[710], S[824], Cout[824]);
Full_Adder FA826 (Cout[710], Cout[711], S[712], S[825], Cout[825]);
Full_Adder FA827 (Cout[712], Cout[713], S[714], S[826], Cout[826]);
Full_Adder FA828 (S[547], Cout[714], Cout[715], S[827], Cout[827]);
Half_Adder HA829 (Cout[720], S[721], S[828], Cout[828]);
Half_Adder HA830 (Cout[721], S[722], S[829], Cout[829]);
Half_Adder HA831 (Cout[722], S[723], S[830], Cout[830]);
Half_Adder HA832 (Cout[723], S[724], S[831], Cout[831]);
Half_Adder HA833 (Cout[724], S[725], S[832], Cout[832]);
Full_Adder FA834 (S[559], Cout[725], S[726], S[833], Cout[833]);
Full_Adder FA835 (S[561], Cout[726], S[727], S[834], Cout[834]);
Full_Adder FA836 (S[563], Cout[727], S[728], S[835], Cout[835]);
Full_Adder FA837 (S[565], Cout[728], S[729], S[836], Cout[836]);
Full_Adder FA838 (Cout[729], S[730], S[731], S[837], Cout[837]);
Full_Adder FA839 (Cout[730], Cout[731], S[732], S[838], Cout[838]);
Full_Adder FA840 (Cout[732], Cout[733], S[734], S[839], Cout[839]);
Full_Adder FA841 (Cout[734], Cout[735], S[736], S[840], Cout[840]);
Full_Adder FA842 (Cout[736], Cout[737], S[738], S[841], Cout[841]);
Full_Adder FA843 (Cout[738], Cout[739], S[740], S[842], Cout[842]);
Full_Adder FA844 (Cout[740], Cout[741], S[742], S[843], Cout[843]);
Full_Adder FA845 (S[587], Cout[742], Cout[743], S[844], Cout[844]);
Half_Adder HA846 (S[744], S[745], S[845], Cout[845]);
Full_Adder FA847 (S[590], Cout[744], Cout[745], S[846], Cout[846]);
Half_Adder HA848 (S[746], S[747], S[847], Cout[847]);
Full_Adder FA849 (S[594], Cout[746], Cout[747], S[848], Cout[848]);
Half_Adder HA850 (S[748], S[749], S[849], Cout[849]);
Full_Adder FA851 (Cout[748], Cout[749], S[750], S[850], Cout[850]);
Half_Adder HA852 (S[751], S[752], S[851], Cout[851]);
Full_Adder FA853 (Cout[750], Cout[751], Cout[752], S[852], Cout[852]);
Full_Adder FA854 (S[753], S[754], S[755], S[853], Cout[853]);
Full_Adder FA855 (Cout[753], Cout[754], Cout[755], S[854], Cout[854]);
Full_Adder FA856 (S[756], S[757], S[758], S[855], Cout[855]);
Full_Adder FA857 (Cout[756], Cout[757], Cout[758], S[856], Cout[856]);
Full_Adder FA858 (S[759], S[760], S[761], S[857], Cout[857]);
Full_Adder FA859 (Cout[759], Cout[760], Cout[761], S[858], Cout[858]);
Full_Adder FA860 (S[762], S[763], S[764], S[859], Cout[859]);
Full_Adder FA861 (Cout[762], Cout[763], Cout[764], S[860], Cout[860]);
Full_Adder FA862 (S[765], S[766], S[767], S[861], Cout[861]);
Full_Adder FA863 (Cout[765], Cout[766], Cout[767], S[862], Cout[862]);
Full_Adder FA864 (S[768], S[769], S[770], S[863], Cout[863]);
Full_Adder FA865 (S[628], Cout[768], Cout[769], S[864], Cout[864]);
Full_Adder FA866 (Cout[770], S[771], S[772], S[865], Cout[865]);
Full_Adder FA867 (S[633], Cout[771], Cout[772], S[866], Cout[866]);
Full_Adder FA868 (Cout[773], S[774], S[775], S[867], Cout[867]);
Full_Adder FA869 (S[638], Cout[774], Cout[775], S[868], Cout[868]);
Full_Adder FA870 (Cout[776], S[777], S[778], S[869], Cout[869]);
Full_Adder FA871 (S[643], Cout[777], Cout[778], S[870], Cout[870]);
Full_Adder FA872 (Cout[779], S[780], S[781], S[871], Cout[871]);
Full_Adder FA873 (S[648], Cout[780], Cout[781], S[872], Cout[872]);
Full_Adder FA874 (Cout[782], S[783], S[784], S[873], Cout[873]);
Full_Adder FA875 (S[653], Cout[783], Cout[784], S[874], Cout[874]);
Full_Adder FA876 (Cout[785], S[786], S[787], S[875], Cout[875]);
Full_Adder FA877 (S[657], Cout[786], Cout[787], S[876], Cout[876]);
Full_Adder FA878 (Cout[788], S[789], S[790], S[877], Cout[877]);
Full_Adder FA879 (S[661], Cout[789], Cout[790], S[878], Cout[878]);
Full_Adder FA880 (Cout[791], S[792], S[793], S[879], Cout[879]);
Full_Adder FA881 (S[665], Cout[792], Cout[793], S[880], Cout[880]);
Full_Adder FA882 (Cout[794], S[795], S[796], S[881], Cout[881]);
Full_Adder FA883 (S[668], S[669], Cout[795], S[882], Cout[882]);
Full_Adder FA884 (Cout[796], Cout[797], S[798], S[883], Cout[883]);
Full_Adder FA885 (S[672], S[673], Cout[798], S[884], Cout[884]);
Half_Adder HA886 (Cout[799], S[800], S[885], Cout[885]);
Full_Adder FA887 (S[676], S[677], Cout[800], S[886], Cout[886]);
Half_Adder HA888 (Cout[801], S[802], S[887], Cout[887]);
Full_Adder FA889 (S[680], S[681], Cout[802], S[888], Cout[888]);
Half_Adder HA890 (Cout[803], S[804], S[889], Cout[889]);
Full_Adder FA891 (S[683], S[684], Cout[804], S[890], Cout[890]);
Half_Adder HA892 (Cout[805], S[806], S[891], Cout[891]);
Full_Adder FA893 (S[687], Cout[806], Cout[807], S[892], Cout[892]);
Full_Adder FA894 (S[690], Cout[808], Cout[809], S[893], Cout[893]);
Full_Adder FA895 (S[693], Cout[810], Cout[811], S[894], Cout[894]);
Full_Adder FA896 (S[696], Cout[812], Cout[813], S[895], Cout[895]);
Full_Adder FA897 (S[699], Cout[814], Cout[815], S[896], Cout[896]);
Full_Adder FA898 (S[701], Cout[816], Cout[817], S[897], Cout[897]);
Full_Adder FA899 (S[702], S[703], Cout[818], S[898], Cout[898]);
Full_Adder FA900 (S[704], S[705], Cout[820], S[899], Cout[899]);
Half_Adder HA901 (S[707], Cout[821], S[900], Cout[900]);
Half_Adder HA902 (S[709], Cout[822], S[901], Cout[901]);
Half_Adder HA903 (S[711], Cout[823], S[902], Cout[902]);
Half_Adder HA904 (S[713], Cout[824], S[903], Cout[903]);
Half_Adder HA905 (S[715], Cout[825], S[904], Cout[904]);
Half_Adder HA906 (S[716], Cout[826], S[905], Cout[905]);
Half_Adder HA907 (Cout[716], S[717], S[906], Cout[906]);
Half_Adder HA908 (Cout[828], S[829], S[907], Cout[907]);
Half_Adder HA909 (Cout[829], S[830], S[908], Cout[908]);
Half_Adder HA910 (Cout[830], S[831], S[909], Cout[909]);
Half_Adder HA911 (Cout[831], S[832], S[910], Cout[910]);
Half_Adder HA912 (Cout[832], S[833], S[911], Cout[911]);
Half_Adder HA913 (Cout[833], S[834], S[912], Cout[912]);
Half_Adder HA914 (Cout[834], S[835], S[913], Cout[913]);
Half_Adder HA915 (Cout[835], S[836], S[914], Cout[914]);
Half_Adder HA916 (Cout[836], S[837], S[915], Cout[915]);
Full_Adder FA917 (S[733], Cout[837], S[838], S[916], Cout[916]);
Full_Adder FA918 (S[735], Cout[838], S[839], S[917], Cout[917]);
Full_Adder FA919 (S[737], Cout[839], S[840], S[918], Cout[918]);
Full_Adder FA920 (S[739], Cout[840], S[841], S[919], Cout[919]);
Full_Adder FA921 (S[741], Cout[841], S[842], S[920], Cout[920]);
Full_Adder FA922 (S[743], Cout[842], S[843], S[921], Cout[921]);
Full_Adder FA923 (Cout[843], S[844], S[845], S[922], Cout[922]);
Full_Adder FA924 (Cout[844], Cout[845], S[846], S[923], Cout[923]);
Full_Adder FA925 (Cout[846], Cout[847], S[848], S[924], Cout[924]);
Full_Adder FA926 (Cout[848], Cout[849], S[850], S[925], Cout[925]);
Full_Adder FA927 (Cout[850], Cout[851], S[852], S[926], Cout[926]);
Full_Adder FA928 (Cout[852], Cout[853], S[854], S[927], Cout[927]);
Full_Adder FA929 (Cout[854], Cout[855], S[856], S[928], Cout[928]);
Full_Adder FA930 (Cout[856], Cout[857], S[858], S[929], Cout[929]);
Full_Adder FA931 (Cout[858], Cout[859], S[860], S[930], Cout[930]);
Full_Adder FA932 (Cout[860], Cout[861], S[862], S[931], Cout[931]);
Full_Adder FA933 (S[773], Cout[862], Cout[863], S[932], Cout[932]);
Full_Adder FA934 (S[776], Cout[864], Cout[865], S[933], Cout[933]);
Full_Adder FA935 (S[779], Cout[866], Cout[867], S[934], Cout[934]);
Full_Adder FA936 (S[782], Cout[868], Cout[869], S[935], Cout[935]);
Full_Adder FA937 (S[785], Cout[870], Cout[871], S[936], Cout[936]);
Full_Adder FA938 (S[788], Cout[872], Cout[873], S[937], Cout[937]);
Full_Adder FA939 (S[791], Cout[874], Cout[875], S[938], Cout[938]);
Full_Adder FA940 (S[794], Cout[876], Cout[877], S[939], Cout[939]);
Full_Adder FA941 (S[797], Cout[878], Cout[879], S[940], Cout[940]);
Full_Adder FA942 (S[799], Cout[880], Cout[881], S[941], Cout[941]);
Full_Adder FA943 (S[801], Cout[882], Cout[883], S[942], Cout[942]);
Full_Adder FA944 (S[803], Cout[884], Cout[885], S[943], Cout[943]);
Full_Adder FA945 (S[805], Cout[886], Cout[887], S[944], Cout[944]);
Full_Adder FA946 (S[807], Cout[888], Cout[889], S[945], Cout[945]);
Full_Adder FA947 (S[808], S[809], Cout[890], S[946], Cout[946]);
Half_Adder HA948 (S[810], S[811], S[947], Cout[947]);
Half_Adder HA949 (S[812], S[813], S[948], Cout[948]);
Half_Adder HA950 (S[814], S[815], S[949], Cout[949]);
Half_Adder HA951 (S[816], S[817], S[950], Cout[950]);
Half_Adder HA952 (S[818], S[819], S[951], Cout[951]);
Half_Adder HA953 (Cout[819], S[820], S[952], Cout[952]);
Half_Adder HA954 (Cout[907], S[908], S[953], Cout[953]);
Half_Adder HA955 (Cout[908], S[909], S[954], Cout[954]);
Half_Adder HA956 (Cout[909], S[910], S[955], Cout[955]);
Half_Adder HA957 (Cout[910], S[911], S[956], Cout[956]);
Half_Adder HA958 (Cout[911], S[912], S[957], Cout[957]);
Half_Adder HA959 (Cout[912], S[913], S[958], Cout[958]);
Half_Adder HA960 (Cout[913], S[914], S[959], Cout[959]);
Half_Adder HA961 (Cout[914], S[915], S[960], Cout[960]);
Half_Adder HA962 (Cout[915], S[916], S[961], Cout[961]);
Half_Adder HA963 (Cout[916], S[917], S[962], Cout[962]);
Half_Adder HA964 (Cout[917], S[918], S[963], Cout[963]);
Half_Adder HA965 (Cout[918], S[919], S[964], Cout[964]);
Half_Adder HA966 (Cout[919], S[920], S[965], Cout[965]);
Half_Adder HA967 (Cout[920], S[921], S[966], Cout[966]);
Half_Adder HA968 (Cout[921], S[922], S[967], Cout[967]);
Full_Adder FA969 (S[847], Cout[922], S[923], S[968], Cout[968]);
Full_Adder FA970 (S[849], Cout[923], S[924], S[969], Cout[969]);
Full_Adder FA971 (S[851], Cout[924], S[925], S[970], Cout[970]);
Full_Adder FA972 (S[853], Cout[925], S[926], S[971], Cout[971]);
Full_Adder FA973 (S[855], Cout[926], S[927], S[972], Cout[972]);
Full_Adder FA974 (S[857], Cout[927], S[928], S[973], Cout[973]);
Full_Adder FA975 (S[859], Cout[928], S[929], S[974], Cout[974]);
Full_Adder FA976 (S[861], Cout[929], S[930], S[975], Cout[975]);
Full_Adder FA977 (S[863], Cout[930], S[931], S[976], Cout[976]);
Full_Adder FA978 (S[864], S[865], Cout[931], S[977], Cout[977]);
Full_Adder FA979 (S[866], S[867], Cout[932], S[978], Cout[978]);
Full_Adder FA980 (S[868], S[869], Cout[933], S[979], Cout[979]);
Full_Adder FA981 (S[870], S[871], Cout[934], S[980], Cout[980]);
Full_Adder FA982 (S[872], S[873], Cout[935], S[981], Cout[981]);
Full_Adder FA983 (S[874], S[875], Cout[936], S[982], Cout[982]);
Full_Adder FA984 (S[876], S[877], Cout[937], S[983], Cout[983]);
Full_Adder FA985 (S[878], S[879], Cout[938], S[984], Cout[984]);
Full_Adder FA986 (S[880], S[881], Cout[939], S[985], Cout[985]);
Full_Adder FA987 (S[882], S[883], Cout[940], S[986], Cout[986]);
Full_Adder FA988 (S[884], S[885], Cout[941], S[987], Cout[987]);
Full_Adder FA989 (S[886], S[887], Cout[942], S[988], Cout[988]);
Full_Adder FA990 (S[888], S[889], Cout[943], S[989], Cout[989]);
Full_Adder FA991 (S[890], S[891], Cout[944], S[990], Cout[990]);
Full_Adder FA992 (Cout[891], S[892], Cout[945], S[991], Cout[991]);
Full_Adder FA993 (Cout[892], S[893], Cout[946], S[992], Cout[992]);
Full_Adder FA994 (Cout[893], S[894], Cout[947], S[993], Cout[993]);
Full_Adder FA995 (Cout[894], S[895], Cout[948], S[994], Cout[994]);
Full_Adder FA996 (Cout[895], S[896], Cout[949], S[995], Cout[995]);
Full_Adder FA997 (Cout[896], S[897], Cout[950], S[996], Cout[996]);
Full_Adder FA998 (Cout[897], S[898], Cout[951], S[997], Cout[997]);
Full_Adder FA999 (S[821], Cout[898], S[899], S[998], Cout[998]);
Half_Adder HA1000 (S[822], Cout[899], S[999], Cout[999]);
Half_Adder HA1001 (S[823], Cout[900], S[1000], Cout[1000]);
Half_Adder HA1002 (S[824], Cout[901], S[1001], Cout[1001]);
Half_Adder HA1003 (S[825], Cout[902], S[1002], Cout[1002]);
Half_Adder HA1004 (S[826], Cout[903], S[1003], Cout[1003]);
Half_Adder HA1005 (S[827], Cout[904], S[1004], Cout[1004]);
Half_Adder HA1006 (Cout[827], Cout[905], S[1005], Cout[1005]);
Half_Adder HA1007 (Cout[717], S[718], S[1006], Cout[1006]);
Half_Adder HA1008 (Cout[953], S[954], S[1007], Cout[1007]);
Half_Adder HA1009 (Cout[954], S[955], S[1008], Cout[1008]);
Half_Adder HA1010 (Cout[955], S[956], S[1009], Cout[1009]);
Half_Adder HA1011 (Cout[956], S[957], S[1010], Cout[1010]);
Half_Adder HA1012 (Cout[957], S[958], S[1011], Cout[1011]);
Half_Adder HA1013 (Cout[958], S[959], S[1012], Cout[1012]);
Half_Adder HA1014 (Cout[959], S[960], S[1013], Cout[1013]);
Half_Adder HA1015 (Cout[960], S[961], S[1014], Cout[1014]);
Half_Adder HA1016 (Cout[961], S[962], S[1015], Cout[1015]);
Half_Adder HA1017 (Cout[962], S[963], S[1016], Cout[1016]);
Half_Adder HA1018 (Cout[963], S[964], S[1017], Cout[1017]);
Half_Adder HA1019 (Cout[964], S[965], S[1018], Cout[1018]);
Half_Adder HA1020 (Cout[965], S[966], S[1019], Cout[1019]);
Half_Adder HA1021 (Cout[966], S[967], S[1020], Cout[1020]);
Half_Adder HA1022 (Cout[967], S[968], S[1021], Cout[1021]);
Half_Adder HA1023 (Cout[968], S[969], S[1022], Cout[1022]);
Half_Adder HA1024 (Cout[969], S[970], S[1023], Cout[1023]);
Half_Adder HA1025 (Cout[970], S[971], S[1024], Cout[1024]);
Half_Adder HA1026 (Cout[971], S[972], S[1025], Cout[1025]);
Half_Adder HA1027 (Cout[972], S[973], S[1026], Cout[1026]);
Half_Adder HA1028 (Cout[973], S[974], S[1027], Cout[1027]);
Half_Adder HA1029 (Cout[974], S[975], S[1028], Cout[1028]);
Half_Adder HA1030 (Cout[975], S[976], S[1029], Cout[1029]);
Full_Adder FA1031 (S[932], Cout[976], S[977], S[1030], Cout[1030]);
Full_Adder FA1032 (S[933], Cout[977], S[978], S[1031], Cout[1031]);
Full_Adder FA1033 (S[934], Cout[978], S[979], S[1032], Cout[1032]);
Full_Adder FA1034 (S[935], Cout[979], S[980], S[1033], Cout[1033]);
Full_Adder FA1035 (S[936], Cout[980], S[981], S[1034], Cout[1034]);
Full_Adder FA1036 (S[937], Cout[981], S[982], S[1035], Cout[1035]);
Full_Adder FA1037 (S[938], Cout[982], S[983], S[1036], Cout[1036]);
Full_Adder FA1038 (S[939], Cout[983], S[984], S[1037], Cout[1037]);
Full_Adder FA1039 (S[940], Cout[984], S[985], S[1038], Cout[1038]);
Full_Adder FA1040 (S[941], Cout[985], S[986], S[1039], Cout[1039]);
Full_Adder FA1041 (S[942], Cout[986], S[987], S[1040], Cout[1040]);
Full_Adder FA1042 (S[943], Cout[987], S[988], S[1041], Cout[1041]);
Full_Adder FA1043 (S[944], Cout[988], S[989], S[1042], Cout[1042]);
Full_Adder FA1044 (S[945], Cout[989], S[990], S[1043], Cout[1043]);
Full_Adder FA1045 (S[946], Cout[990], S[991], S[1044], Cout[1044]);
Full_Adder FA1046 (S[947], Cout[991], S[992], S[1045], Cout[1045]);
Full_Adder FA1047 (S[948], Cout[992], S[993], S[1046], Cout[1046]);
Full_Adder FA1048 (S[949], Cout[993], S[994], S[1047], Cout[1047]);
Full_Adder FA1049 (S[950], Cout[994], S[995], S[1048], Cout[1048]);
Full_Adder FA1050 (S[951], Cout[995], S[996], S[1049], Cout[1049]);
Full_Adder FA1051 (S[952], Cout[996], S[997], S[1050], Cout[1050]);
Full_Adder FA1052 (Cout[952], Cout[997], S[998], S[1051], Cout[1051]);
Full_Adder FA1053 (S[900], Cout[998], S[999], S[1052], Cout[1052]);
Full_Adder FA1054 (S[901], Cout[999], S[1000], S[1053], Cout[1053]);
Full_Adder FA1055 (S[902], Cout[1000], S[1001], S[1054], Cout[1054]);
Full_Adder FA1056 (S[903], Cout[1001], S[1002], S[1055], Cout[1055]);
Full_Adder FA1057 (S[904], Cout[1002], S[1003], S[1056], Cout[1056]);
Full_Adder FA1058 (S[905], Cout[1003], S[1004], S[1057], Cout[1057]);
Full_Adder FA1059 (S[906], Cout[1004], S[1005], S[1058], Cout[1058]);
Full_Adder FA1060 (Cout[906], Cout[1005], S[1006], S[1059], Cout[1059]);
Full_Adder FA1061 (Cout[718], S[719], Cout[1006], S[1060], Cout[1060]);
Half_Adder HA1062 (P[31][31], Cout[719], S[1061], Cout[1061]);
Half_Adder HA1063 (Cout[1007], S[1008], S[1062], Cout[1062]);
Full_Adder FA1064 (Cout[1008], S[1009], Cout[1062], S[1063], Cout[1063]);
Full_Adder FA1065 (Cout[1009], S[1010], Cout[1063], S[1064], Cout[1064]);
Full_Adder FA1066 (Cout[1010], S[1011], Cout[1064], S[1065], Cout[1065]);
Full_Adder FA1067 (Cout[1011], S[1012], Cout[1065], S[1066], Cout[1066]);
Full_Adder FA1068 (Cout[1012], S[1013], Cout[1066], S[1067], Cout[1067]);
Full_Adder FA1069 (Cout[1013], S[1014], Cout[1067], S[1068], Cout[1068]);
Full_Adder FA1070 (Cout[1014], S[1015], Cout[1068], S[1069], Cout[1069]);
Full_Adder FA1071 (Cout[1015], S[1016], Cout[1069], S[1070], Cout[1070]);
Full_Adder FA1072 (Cout[1016], S[1017], Cout[1070], S[1071], Cout[1071]);
Full_Adder FA1073 (Cout[1017], S[1018], Cout[1071], S[1072], Cout[1072]);
Full_Adder FA1074 (Cout[1018], S[1019], Cout[1072], S[1073], Cout[1073]);
Full_Adder FA1075 (Cout[1019], S[1020], Cout[1073], S[1074], Cout[1074]);
Full_Adder FA1076 (Cout[1020], S[1021], Cout[1074], S[1075], Cout[1075]);
Full_Adder FA1077 (Cout[1021], S[1022], Cout[1075], S[1076], Cout[1076]);
Full_Adder FA1078 (Cout[1022], S[1023], Cout[1076], S[1077], Cout[1077]);
Full_Adder FA1079 (Cout[1023], S[1024], Cout[1077], S[1078], Cout[1078]);
Full_Adder FA1080 (Cout[1024], S[1025], Cout[1078], S[1079], Cout[1079]);
Full_Adder FA1081 (Cout[1025], S[1026], Cout[1079], S[1080], Cout[1080]);
Full_Adder FA1082 (Cout[1026], S[1027], Cout[1080], S[1081], Cout[1081]);
Full_Adder FA1083 (Cout[1027], S[1028], Cout[1081], S[1082], Cout[1082]);
Full_Adder FA1084 (Cout[1028], S[1029], Cout[1082], S[1083], Cout[1083]);
Full_Adder FA1085 (Cout[1029], S[1030], Cout[1083], S[1084], Cout[1084]);
Full_Adder FA1086 (Cout[1030], S[1031], Cout[1084], S[1085], Cout[1085]);
Full_Adder FA1087 (Cout[1031], S[1032], Cout[1085], S[1086], Cout[1086]);
Full_Adder FA1088 (Cout[1032], S[1033], Cout[1086], S[1087], Cout[1087]);
Full_Adder FA1089 (Cout[1033], S[1034], Cout[1087], S[1088], Cout[1088]);
Full_Adder FA1090 (Cout[1034], S[1035], Cout[1088], S[1089], Cout[1089]);
Full_Adder FA1091 (Cout[1035], S[1036], Cout[1089], S[1090], Cout[1090]);
Full_Adder FA1092 (Cout[1036], S[1037], Cout[1090], S[1091], Cout[1091]);
Full_Adder FA1093 (Cout[1037], S[1038], Cout[1091], S[1092], Cout[1092]);
Full_Adder FA1094 (Cout[1038], S[1039], Cout[1092], S[1093], Cout[1093]);
Full_Adder FA1095 (Cout[1039], S[1040], Cout[1093], S[1094], Cout[1094]);
Full_Adder FA1096 (Cout[1040], S[1041], Cout[1094], S[1095], Cout[1095]);
Full_Adder FA1097 (Cout[1041], S[1042], Cout[1095], S[1096], Cout[1096]);
Full_Adder FA1098 (Cout[1042], S[1043], Cout[1096], S[1097], Cout[1097]);
Full_Adder FA1099 (Cout[1043], S[1044], Cout[1097], S[1098], Cout[1098]);
Full_Adder FA1100 (Cout[1044], S[1045], Cout[1098], S[1099], Cout[1099]);
Full_Adder FA1101 (Cout[1045], S[1046], Cout[1099], S[1100], Cout[1100]);
Full_Adder FA1102 (Cout[1046], S[1047], Cout[1100], S[1101], Cout[1101]);
Full_Adder FA1103 (Cout[1047], S[1048], Cout[1101], S[1102], Cout[1102]);
Full_Adder FA1104 (Cout[1048], S[1049], Cout[1102], S[1103], Cout[1103]);
Full_Adder FA1105 (Cout[1049], S[1050], Cout[1103], S[1104], Cout[1104]);
Full_Adder FA1106 (Cout[1050], S[1051], Cout[1104], S[1105], Cout[1105]);
Full_Adder FA1107 (Cout[1051], S[1052], Cout[1105], S[1106], Cout[1106]);
Full_Adder FA1108 (Cout[1052], S[1053], Cout[1106], S[1107], Cout[1107]);
Full_Adder FA1109 (Cout[1053], S[1054], Cout[1107], S[1108], Cout[1108]);
Full_Adder FA1110 (Cout[1054], S[1055], Cout[1108], S[1109], Cout[1109]);
Full_Adder FA1111 (Cout[1055], S[1056], Cout[1109], S[1110], Cout[1110]);
Full_Adder FA1112 (Cout[1056], S[1057], Cout[1110], S[1111], Cout[1111]);
Full_Adder FA1113 (Cout[1057], S[1058], Cout[1111], S[1112], Cout[1112]);
Full_Adder FA1114 (Cout[1058], S[1059], Cout[1112], S[1113], Cout[1113]);
Full_Adder FA1115 (Cout[1059], S[1060], Cout[1113], S[1114], Cout[1114]);
Full_Adder FA1116 (Cout[1060], S[1061], Cout[1114], S[1115], Cout[1115]);
Half_Adder HA1117 (Cout[1061], Cout[1115], S[1116], Cout[1116]);

assign z[63] = S[1116];
assign z[62] = S[1115];
assign z[61] = S[1114];
assign z[60] = S[1113];
assign z[59] = S[1112];
assign z[58] = S[1111];
assign z[57] = S[1110];
assign z[56] = S[1109];
assign z[55] = S[1108];
assign z[54] = S[1107];
assign z[53] = S[1106];
assign z[52] = S[1105];
assign z[51] = S[1104];
assign z[50] = S[1103];
assign z[49] = S[1102];
assign z[48] = S[1101];
assign z[47] = S[1100];
assign z[46] = S[1099];
assign z[45] = S[1098];
assign z[44] = S[1097];
assign z[43] = S[1096];
assign z[42] = S[1095];
assign z[41] = S[1094];
assign z[40] = S[1093];
assign z[39] = S[1092];
assign z[38] = S[1091];
assign z[37] = S[1090];
assign z[36] = S[1089];
assign z[35] = S[1088];
assign z[34] = S[1087];
assign z[33] = S[1086];
assign z[32] = S[1085];
assign z[31] = S[1084];
assign z[30] = S[1083];
assign z[29] = S[1082];
assign z[28] = S[1081];
assign z[27] = S[1080];
assign z[26] = S[1079];
assign z[25] = S[1078];
assign z[24] = S[1077];
assign z[23] = S[1076];
assign z[22] = S[1075];
assign z[21] = S[1074];
assign z[20] = S[1073];
assign z[19] = S[1072];
assign z[18] = S[1071];
assign z[17] = S[1070];
assign z[16] = S[1069];
assign z[15] = S[1068];
assign z[14] = S[1067];
assign z[13] = S[1066];
assign z[12] = S[1065];
assign z[11] = S[1064];
assign z[10] = S[1063];
assign z[9] = S[1062];
assign z[8] = S[1007];
assign z[7] = S[953];
assign z[6] = S[907];
assign z[5] = S[828];
assign z[4] = S[720];
assign z[3] = S[550];
assign z[2] = S[320];
assign z[1] = S[0];
assign z[0] = P[0][0];

endmodule
